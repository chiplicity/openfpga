magic
tech sky130A
magscale 1 2
timestamp 1605122071
<< locali >>
rect 22845 12155 22879 12325
rect 18061 5627 18095 5865
rect 9873 3043 9907 3145
<< viali >>
rect 23489 24361 23523 24395
rect 24593 24225 24627 24259
rect 24777 24089 24811 24123
rect 24777 23817 24811 23851
rect 24409 23681 24443 23715
rect 24593 23613 24627 23647
rect 25237 23477 25271 23511
rect 24777 23273 24811 23307
rect 12817 23205 12851 23239
rect 12541 23137 12575 23171
rect 24593 23137 24627 23171
rect 24777 22729 24811 22763
rect 24593 22525 24627 22559
rect 25145 22525 25179 22559
rect 12633 22389 12667 22423
rect 24409 22389 24443 22423
rect 23857 22117 23891 22151
rect 23581 22049 23615 22083
rect 24869 22049 24903 22083
rect 25053 21913 25087 21947
rect 24869 21641 24903 21675
rect 25145 21641 25179 21675
rect 14565 21505 14599 21539
rect 23949 21505 23983 21539
rect 14289 21437 14323 21471
rect 15025 21437 15059 21471
rect 23489 21437 23523 21471
rect 23673 21437 23707 21471
rect 24961 21437 24995 21471
rect 25513 21437 25547 21471
rect 24409 21369 24443 21403
rect 25053 21097 25087 21131
rect 23581 20961 23615 20995
rect 24869 20961 24903 20995
rect 23765 20893 23799 20927
rect 16865 20553 16899 20587
rect 24777 20553 24811 20587
rect 16681 20349 16715 20383
rect 17233 20349 17267 20383
rect 24593 20349 24627 20383
rect 25145 20349 25179 20383
rect 23857 20213 23891 20247
rect 25513 20213 25547 20247
rect 17316 19941 17350 19975
rect 23765 19941 23799 19975
rect 23489 19873 23523 19907
rect 17049 19805 17083 19839
rect 18429 19669 18463 19703
rect 17141 19465 17175 19499
rect 17417 19397 17451 19431
rect 23949 19329 23983 19363
rect 15669 19261 15703 19295
rect 15945 19261 15979 19295
rect 23673 19261 23707 19295
rect 24409 19261 24443 19295
rect 24961 19261 24995 19295
rect 25513 19261 25547 19295
rect 16405 19193 16439 19227
rect 23489 19125 23523 19159
rect 25145 19125 25179 19159
rect 24777 18921 24811 18955
rect 24593 18785 24627 18819
rect 15025 18377 15059 18411
rect 24685 18377 24719 18411
rect 13553 18173 13587 18207
rect 14289 18173 14323 18207
rect 14841 18173 14875 18207
rect 13829 18105 13863 18139
rect 15393 18105 15427 18139
rect 24777 17833 24811 17867
rect 11621 17765 11655 17799
rect 11345 17697 11379 17731
rect 24593 17697 24627 17731
rect 24777 17289 24811 17323
rect 13461 17153 13495 17187
rect 13185 17085 13219 17119
rect 13921 17085 13955 17119
rect 24593 17085 24627 17119
rect 11437 16949 11471 16983
rect 24409 16949 24443 16983
rect 25145 16949 25179 16983
rect 22937 16745 22971 16779
rect 16313 16609 16347 16643
rect 16589 16609 16623 16643
rect 22753 16609 22787 16643
rect 25145 16201 25179 16235
rect 23949 16065 23983 16099
rect 23673 15997 23707 16031
rect 24409 15997 24443 16031
rect 24961 15997 24995 16031
rect 25513 15997 25547 16031
rect 16405 15861 16439 15895
rect 22753 15861 22787 15895
rect 23397 15657 23431 15691
rect 22201 15589 22235 15623
rect 21925 15521 21959 15555
rect 23213 15521 23247 15555
rect 25881 15113 25915 15147
rect 24225 14977 24259 15011
rect 23949 14909 23983 14943
rect 24685 14909 24719 14943
rect 25237 14909 25271 14943
rect 21925 14773 21959 14807
rect 23213 14773 23247 14807
rect 25421 14773 25455 14807
rect 24777 14569 24811 14603
rect 22477 14501 22511 14535
rect 22201 14433 22235 14467
rect 24593 14433 24627 14467
rect 18889 14025 18923 14059
rect 24685 14025 24719 14059
rect 25605 14025 25639 14059
rect 25145 13957 25179 13991
rect 23949 13889 23983 13923
rect 22661 13821 22695 13855
rect 23489 13821 23523 13855
rect 23673 13821 23707 13855
rect 24961 13821 24995 13855
rect 19257 13685 19291 13719
rect 19625 13685 19659 13719
rect 21097 13685 21131 13719
rect 22109 13685 22143 13719
rect 19257 13481 19291 13515
rect 24777 13481 24811 13515
rect 19625 13345 19659 13379
rect 23489 13345 23523 13379
rect 24593 13345 24627 13379
rect 19717 13277 19751 13311
rect 19809 13277 19843 13311
rect 21465 13277 21499 13311
rect 22477 13277 22511 13311
rect 18705 13209 18739 13243
rect 23673 13209 23707 13243
rect 19073 13141 19107 13175
rect 21189 13141 21223 13175
rect 24041 13141 24075 13175
rect 18521 12937 18555 12971
rect 18981 12937 19015 12971
rect 20269 12937 20303 12971
rect 23489 12937 23523 12971
rect 24685 12937 24719 12971
rect 25145 12937 25179 12971
rect 22661 12869 22695 12903
rect 19533 12801 19567 12835
rect 21281 12801 21315 12835
rect 23949 12801 23983 12835
rect 19441 12733 19475 12767
rect 22477 12733 22511 12767
rect 23673 12733 23707 12767
rect 24961 12733 24995 12767
rect 25513 12733 25547 12767
rect 18797 12665 18831 12699
rect 19349 12665 19383 12699
rect 20637 12665 20671 12699
rect 21097 12665 21131 12699
rect 16773 12597 16807 12631
rect 20729 12597 20763 12631
rect 21189 12597 21223 12631
rect 21741 12597 21775 12631
rect 23121 12597 23155 12631
rect 17141 12393 17175 12427
rect 18245 12393 18279 12427
rect 19073 12393 19107 12427
rect 23121 12393 23155 12427
rect 18981 12325 19015 12359
rect 21180 12325 21214 12359
rect 22845 12325 22879 12359
rect 23489 12325 23523 12359
rect 24961 12325 24995 12359
rect 17509 12257 17543 12291
rect 17601 12257 17635 12291
rect 19441 12257 19475 12291
rect 17693 12189 17727 12223
rect 19533 12189 19567 12223
rect 19625 12189 19659 12223
rect 20085 12189 20119 12223
rect 20913 12189 20947 12223
rect 24685 12257 24719 12291
rect 23581 12189 23615 12223
rect 23673 12189 23707 12223
rect 22569 12121 22603 12155
rect 22845 12121 22879 12155
rect 18613 12053 18647 12087
rect 20453 12053 20487 12087
rect 22293 12053 22327 12087
rect 22937 12053 22971 12087
rect 24225 12053 24259 12087
rect 16865 11849 16899 11883
rect 17785 11849 17819 11883
rect 20913 11849 20947 11883
rect 21833 11849 21867 11883
rect 25329 11849 25363 11883
rect 16957 11713 16991 11747
rect 19073 11713 19107 11747
rect 22661 11713 22695 11747
rect 15209 11645 15243 11679
rect 19533 11645 19567 11679
rect 23673 11645 23707 11679
rect 15485 11577 15519 11611
rect 18521 11577 18555 11611
rect 19778 11577 19812 11611
rect 21557 11577 21591 11611
rect 23121 11577 23155 11611
rect 23489 11577 23523 11611
rect 23918 11577 23952 11611
rect 16037 11509 16071 11543
rect 16313 11509 16347 11543
rect 17417 11509 17451 11543
rect 18429 11509 18463 11543
rect 22017 11509 22051 11543
rect 22385 11509 22419 11543
rect 22477 11509 22511 11543
rect 25053 11509 25087 11543
rect 15301 11305 15335 11339
rect 20269 11305 20303 11339
rect 20545 11305 20579 11339
rect 21189 11305 21223 11339
rect 22661 11305 22695 11339
rect 23213 11305 23247 11339
rect 15669 11169 15703 11203
rect 17049 11169 17083 11203
rect 18889 11169 18923 11203
rect 19156 11169 19190 11203
rect 21537 11169 21571 11203
rect 23489 11169 23523 11203
rect 23756 11169 23790 11203
rect 14197 11101 14231 11135
rect 15761 11101 15795 11135
rect 15853 11101 15887 11135
rect 21281 11101 21315 11135
rect 14841 11033 14875 11067
rect 16589 10965 16623 10999
rect 16957 10965 16991 10999
rect 18337 10965 18371 10999
rect 24869 10965 24903 10999
rect 15945 10761 15979 10795
rect 16865 10761 16899 10795
rect 19441 10761 19475 10795
rect 19809 10761 19843 10795
rect 21281 10761 21315 10795
rect 21925 10761 21959 10795
rect 24777 10761 24811 10795
rect 25421 10761 25455 10795
rect 14381 10693 14415 10727
rect 16037 10693 16071 10727
rect 20085 10693 20119 10727
rect 22017 10693 22051 10727
rect 14933 10625 14967 10659
rect 16681 10625 16715 10659
rect 17417 10625 17451 10659
rect 20729 10625 20763 10659
rect 20821 10625 20855 10659
rect 22477 10625 22511 10659
rect 22661 10625 22695 10659
rect 24225 10625 24259 10659
rect 25053 10625 25087 10659
rect 13001 10557 13035 10591
rect 13093 10557 13127 10591
rect 16405 10557 16439 10591
rect 17325 10557 17359 10591
rect 18061 10557 18095 10591
rect 22385 10557 22419 10591
rect 23121 10557 23155 10591
rect 24133 10557 24167 10591
rect 25237 10557 25271 10591
rect 25789 10557 25823 10591
rect 13369 10489 13403 10523
rect 14841 10489 14875 10523
rect 18328 10489 18362 10523
rect 20637 10489 20671 10523
rect 23489 10489 23523 10523
rect 13829 10421 13863 10455
rect 14289 10421 14323 10455
rect 14749 10421 14783 10455
rect 15393 10421 15427 10455
rect 16497 10421 16531 10455
rect 17233 10421 17267 10455
rect 20269 10421 20303 10455
rect 23673 10421 23707 10455
rect 24041 10421 24075 10455
rect 12909 10217 12943 10251
rect 14749 10217 14783 10251
rect 15117 10217 15151 10251
rect 15577 10217 15611 10251
rect 17785 10217 17819 10251
rect 18153 10217 18187 10251
rect 18337 10217 18371 10251
rect 18613 10217 18647 10251
rect 19625 10217 19659 10251
rect 20177 10217 20211 10251
rect 21281 10217 21315 10251
rect 21649 10217 21683 10251
rect 22661 10217 22695 10251
rect 13829 10149 13863 10183
rect 21741 10149 21775 10183
rect 22385 10149 22419 10183
rect 23550 10149 23584 10183
rect 13921 10081 13955 10115
rect 14197 10081 14231 10115
rect 16129 10081 16163 10115
rect 16396 10081 16430 10115
rect 18521 10081 18555 10115
rect 18981 10081 19015 10115
rect 19073 10081 19107 10115
rect 20361 10081 20395 10115
rect 23121 10081 23155 10115
rect 23305 10081 23339 10115
rect 19165 10013 19199 10047
rect 19993 10013 20027 10047
rect 21925 10013 21959 10047
rect 17509 9945 17543 9979
rect 21189 9945 21223 9979
rect 16037 9877 16071 9911
rect 20729 9877 20763 9911
rect 24685 9877 24719 9911
rect 24961 9877 24995 9911
rect 14289 9673 14323 9707
rect 16957 9673 16991 9707
rect 19717 9673 19751 9707
rect 13277 9605 13311 9639
rect 19441 9605 19475 9639
rect 20085 9605 20119 9639
rect 23121 9605 23155 9639
rect 13921 9537 13955 9571
rect 17877 9537 17911 9571
rect 23765 9537 23799 9571
rect 13185 9469 13219 9503
rect 13645 9469 13679 9503
rect 14841 9469 14875 9503
rect 17233 9469 17267 9503
rect 18061 9469 18095 9503
rect 20269 9469 20303 9503
rect 20525 9469 20559 9503
rect 22293 9469 22327 9503
rect 22477 9469 22511 9503
rect 25421 9469 25455 9503
rect 14749 9401 14783 9435
rect 15086 9401 15120 9435
rect 18306 9401 18340 9435
rect 23489 9401 23523 9435
rect 24032 9401 24066 9435
rect 12817 9333 12851 9367
rect 13737 9333 13771 9367
rect 16221 9333 16255 9367
rect 16589 9333 16623 9367
rect 17049 9333 17083 9367
rect 21649 9333 21683 9367
rect 21925 9333 21959 9367
rect 22661 9333 22695 9367
rect 25145 9333 25179 9367
rect 11989 9129 12023 9163
rect 13369 9129 13403 9163
rect 13553 9129 13587 9163
rect 18061 9129 18095 9163
rect 20269 9129 20303 9163
rect 21189 9129 21223 9163
rect 23305 9129 23339 9163
rect 16948 9061 16982 9095
rect 19349 9061 19383 9095
rect 12357 8993 12391 9027
rect 13921 8993 13955 9027
rect 14013 8993 14047 9027
rect 15577 8993 15611 9027
rect 16681 8993 16715 9027
rect 19257 8993 19291 9027
rect 20729 8993 20763 9027
rect 21557 8993 21591 9027
rect 22293 8993 22327 9027
rect 22937 8993 22971 9027
rect 23664 8993 23698 9027
rect 12449 8925 12483 8959
rect 12541 8925 12575 8959
rect 14105 8925 14139 8959
rect 19533 8925 19567 8959
rect 21649 8925 21683 8959
rect 21833 8925 21867 8959
rect 23397 8925 23431 8959
rect 15761 8857 15795 8891
rect 14565 8789 14599 8823
rect 15117 8789 15151 8823
rect 16129 8789 16163 8823
rect 16589 8789 16623 8823
rect 18613 8789 18647 8823
rect 18889 8789 18923 8823
rect 19901 8789 19935 8823
rect 24777 8789 24811 8823
rect 11253 8585 11287 8619
rect 12081 8585 12115 8619
rect 13185 8585 13219 8619
rect 15025 8585 15059 8619
rect 16129 8585 16163 8619
rect 17141 8585 17175 8619
rect 18613 8585 18647 8619
rect 20453 8585 20487 8619
rect 20729 8585 20763 8619
rect 21281 8585 21315 8619
rect 23489 8585 23523 8619
rect 23121 8517 23155 8551
rect 23673 8517 23707 8551
rect 24685 8517 24719 8551
rect 12449 8449 12483 8483
rect 13645 8449 13679 8483
rect 16773 8449 16807 8483
rect 17509 8449 17543 8483
rect 21925 8449 21959 8483
rect 22293 8449 22327 8483
rect 24133 8449 24167 8483
rect 24225 8449 24259 8483
rect 13461 8381 13495 8415
rect 16037 8381 16071 8415
rect 16497 8381 16531 8415
rect 19073 8381 19107 8415
rect 21649 8381 21683 8415
rect 25237 8381 25271 8415
rect 25973 8381 26007 8415
rect 11345 8313 11379 8347
rect 13912 8313 13946 8347
rect 15669 8313 15703 8347
rect 18981 8313 19015 8347
rect 19340 8313 19374 8347
rect 21189 8313 21223 8347
rect 22661 8313 22695 8347
rect 24041 8313 24075 8347
rect 25513 8313 25547 8347
rect 15853 8245 15887 8279
rect 16589 8245 16623 8279
rect 18061 8245 18095 8279
rect 21741 8245 21775 8279
rect 25145 8245 25179 8279
rect 9965 8041 9999 8075
rect 10977 8041 11011 8075
rect 14841 8041 14875 8075
rect 16957 8041 16991 8075
rect 17233 8041 17267 8075
rect 17693 8041 17727 8075
rect 18521 8041 18555 8075
rect 19533 8041 19567 8075
rect 21281 8041 21315 8075
rect 22017 8041 22051 8075
rect 23029 8041 23063 8075
rect 24133 8041 24167 8075
rect 25145 8041 25179 8075
rect 12081 7973 12115 8007
rect 12786 7973 12820 8007
rect 15844 7973 15878 8007
rect 20729 7973 20763 8007
rect 22937 7973 22971 8007
rect 23765 7973 23799 8007
rect 11345 7905 11379 7939
rect 15025 7905 15059 7939
rect 18889 7905 18923 7939
rect 20269 7905 20303 7939
rect 24501 7905 24535 7939
rect 24593 7905 24627 7939
rect 11437 7837 11471 7871
rect 11621 7837 11655 7871
rect 12541 7837 12575 7871
rect 15577 7837 15611 7871
rect 18981 7837 19015 7871
rect 19073 7837 19107 7871
rect 21373 7837 21407 7871
rect 21557 7837 21591 7871
rect 23121 7837 23155 7871
rect 24777 7837 24811 7871
rect 19993 7769 20027 7803
rect 20085 7769 20119 7803
rect 12357 7701 12391 7735
rect 13921 7701 13955 7735
rect 14197 7701 14231 7735
rect 14565 7701 14599 7735
rect 17969 7701 18003 7735
rect 18429 7701 18463 7735
rect 20913 7701 20947 7735
rect 22385 7701 22419 7735
rect 22569 7701 22603 7735
rect 12265 7497 12299 7531
rect 13001 7497 13035 7531
rect 14013 7497 14047 7531
rect 15945 7497 15979 7531
rect 16221 7497 16255 7531
rect 17417 7497 17451 7531
rect 18337 7497 18371 7531
rect 19809 7497 19843 7531
rect 20637 7497 20671 7531
rect 22109 7497 22143 7531
rect 23029 7497 23063 7531
rect 25421 7497 25455 7531
rect 20453 7429 20487 7463
rect 12817 7361 12851 7395
rect 13645 7361 13679 7395
rect 14473 7361 14507 7395
rect 21189 7361 21223 7395
rect 22385 7361 22419 7395
rect 23673 7361 23707 7395
rect 10149 7293 10183 7327
rect 13369 7293 13403 7327
rect 14565 7293 14599 7327
rect 14832 7293 14866 7327
rect 16773 7293 16807 7327
rect 18429 7293 18463 7327
rect 21097 7293 21131 7327
rect 22201 7293 22235 7327
rect 10057 7225 10091 7259
rect 10416 7225 10450 7259
rect 18674 7225 18708 7259
rect 23918 7225 23952 7259
rect 9689 7157 9723 7191
rect 11529 7157 11563 7191
rect 11805 7157 11839 7191
rect 13461 7157 13495 7191
rect 16589 7157 16623 7191
rect 16957 7157 16991 7191
rect 17785 7157 17819 7191
rect 20177 7157 20211 7191
rect 21005 7157 21039 7191
rect 21741 7157 21775 7191
rect 23489 7157 23523 7191
rect 25053 7157 25087 7191
rect 12909 6953 12943 6987
rect 13277 6953 13311 6987
rect 14013 6953 14047 6987
rect 14841 6953 14875 6987
rect 16589 6953 16623 6987
rect 19993 6953 20027 6987
rect 20361 6953 20395 6987
rect 22385 6953 22419 6987
rect 22753 6953 22787 6987
rect 24869 6953 24903 6987
rect 23458 6885 23492 6919
rect 10333 6817 10367 6851
rect 11437 6817 11471 6851
rect 11796 6817 11830 6851
rect 14105 6817 14139 6851
rect 16037 6817 16071 6851
rect 16497 6817 16531 6851
rect 17693 6817 17727 6851
rect 17960 6817 17994 6851
rect 21005 6817 21039 6851
rect 21272 6817 21306 6851
rect 23213 6817 23247 6851
rect 10425 6749 10459 6783
rect 10609 6749 10643 6783
rect 11529 6749 11563 6783
rect 16681 6749 16715 6783
rect 25421 6749 25455 6783
rect 9965 6681 9999 6715
rect 15577 6681 15611 6715
rect 16129 6681 16163 6715
rect 9505 6613 9539 6647
rect 11069 6613 11103 6647
rect 14289 6613 14323 6647
rect 17601 6613 17635 6647
rect 19073 6613 19107 6647
rect 19349 6613 19383 6647
rect 20729 6613 20763 6647
rect 23121 6613 23155 6647
rect 24593 6613 24627 6647
rect 10057 6409 10091 6443
rect 11529 6409 11563 6443
rect 12173 6409 12207 6443
rect 13277 6409 13311 6443
rect 14841 6409 14875 6443
rect 16221 6409 16255 6443
rect 16405 6409 16439 6443
rect 17785 6409 17819 6443
rect 18245 6409 18279 6443
rect 19717 6409 19751 6443
rect 21281 6409 21315 6443
rect 21557 6409 21591 6443
rect 22017 6409 22051 6443
rect 23489 6409 23523 6443
rect 25513 6409 25547 6443
rect 15209 6341 15243 6375
rect 19257 6341 19291 6375
rect 23121 6341 23155 6375
rect 9137 6273 9171 6307
rect 9689 6273 9723 6307
rect 15945 6273 15979 6307
rect 16957 6273 16991 6307
rect 18797 6273 18831 6307
rect 23857 6273 23891 6307
rect 10149 6205 10183 6239
rect 13461 6205 13495 6239
rect 13717 6205 13751 6239
rect 16773 6205 16807 6239
rect 18613 6205 18647 6239
rect 18705 6205 18739 6239
rect 19901 6205 19935 6239
rect 20157 6205 20191 6239
rect 22477 6205 22511 6239
rect 24124 6205 24158 6239
rect 9045 6137 9079 6171
rect 10416 6137 10450 6171
rect 12449 6137 12483 6171
rect 11805 6069 11839 6103
rect 13001 6069 13035 6103
rect 15577 6069 15611 6103
rect 16865 6069 16899 6103
rect 22661 6069 22695 6103
rect 25237 6069 25271 6103
rect 8585 5865 8619 5899
rect 10241 5865 10275 5899
rect 13645 5865 13679 5899
rect 14105 5865 14139 5899
rect 15853 5865 15887 5899
rect 17417 5865 17451 5899
rect 18061 5865 18095 5899
rect 18153 5865 18187 5899
rect 18337 5865 18371 5899
rect 20361 5865 20395 5899
rect 23305 5865 23339 5899
rect 23673 5865 23707 5899
rect 12510 5797 12544 5831
rect 17877 5797 17911 5831
rect 10609 5729 10643 5763
rect 16221 5729 16255 5763
rect 10057 5661 10091 5695
rect 10701 5661 10735 5695
rect 10885 5661 10919 5695
rect 12265 5661 12299 5695
rect 16313 5661 16347 5695
rect 16405 5661 16439 5695
rect 24124 5797 24158 5831
rect 18705 5729 18739 5763
rect 20913 5729 20947 5763
rect 22661 5729 22695 5763
rect 23857 5729 23891 5763
rect 25513 5729 25547 5763
rect 18797 5661 18831 5695
rect 18889 5661 18923 5695
rect 22753 5661 22787 5695
rect 22937 5661 22971 5695
rect 18061 5593 18095 5627
rect 22293 5593 22327 5627
rect 9505 5525 9539 5559
rect 11529 5525 11563 5559
rect 15669 5525 15703 5559
rect 16957 5525 16991 5559
rect 19993 5525 20027 5559
rect 21097 5525 21131 5559
rect 22109 5525 22143 5559
rect 25237 5525 25271 5559
rect 9505 5321 9539 5355
rect 11345 5321 11379 5355
rect 14657 5321 14691 5355
rect 15761 5321 15795 5355
rect 18337 5321 18371 5355
rect 19901 5321 19935 5355
rect 20913 5321 20947 5355
rect 22017 5321 22051 5355
rect 23121 5321 23155 5355
rect 23489 5321 23523 5355
rect 24041 5321 24075 5355
rect 15577 5253 15611 5287
rect 16865 5253 16899 5287
rect 23949 5253 23983 5287
rect 13277 5185 13311 5219
rect 16405 5185 16439 5219
rect 18889 5185 18923 5219
rect 20453 5185 20487 5219
rect 21557 5185 21591 5219
rect 22661 5185 22695 5219
rect 24501 5185 24535 5219
rect 24685 5185 24719 5219
rect 9965 5117 9999 5151
rect 10232 5117 10266 5151
rect 12173 5117 12207 5151
rect 16129 5117 16163 5151
rect 17785 5117 17819 5151
rect 18705 5117 18739 5151
rect 18797 5117 18831 5151
rect 19441 5117 19475 5151
rect 22385 5117 22419 5151
rect 25053 5117 25087 5151
rect 11713 5049 11747 5083
rect 13185 5049 13219 5083
rect 13522 5049 13556 5083
rect 19809 5049 19843 5083
rect 20269 5049 20303 5083
rect 21833 5049 21867 5083
rect 24409 5049 24443 5083
rect 25421 5049 25455 5083
rect 7941 4981 7975 5015
rect 8861 4981 8895 5015
rect 8953 4981 8987 5015
rect 9781 4981 9815 5015
rect 12633 4981 12667 5015
rect 15301 4981 15335 5015
rect 16221 4981 16255 5015
rect 17417 4981 17451 5015
rect 20361 4981 20395 5015
rect 22477 4981 22511 5015
rect 25605 4981 25639 5015
rect 8677 4777 8711 4811
rect 9873 4777 9907 4811
rect 10977 4777 11011 4811
rect 11437 4777 11471 4811
rect 12817 4777 12851 4811
rect 14381 4777 14415 4811
rect 15117 4777 15151 4811
rect 17141 4777 17175 4811
rect 18337 4777 18371 4811
rect 21557 4777 21591 4811
rect 22017 4777 22051 4811
rect 22109 4777 22143 4811
rect 24133 4777 24167 4811
rect 25053 4777 25087 4811
rect 25421 4777 25455 4811
rect 10333 4709 10367 4743
rect 15669 4709 15703 4743
rect 17969 4709 18003 4743
rect 20085 4709 20119 4743
rect 23121 4709 23155 4743
rect 23581 4709 23615 4743
rect 24041 4709 24075 4743
rect 8493 4641 8527 4675
rect 10241 4641 10275 4675
rect 11805 4641 11839 4675
rect 13257 4641 13291 4675
rect 16028 4641 16062 4675
rect 18696 4641 18730 4675
rect 21005 4641 21039 4675
rect 22477 4641 22511 4675
rect 24777 4641 24811 4675
rect 25237 4641 25271 4675
rect 7481 4573 7515 4607
rect 10517 4573 10551 4607
rect 11897 4573 11931 4607
rect 12081 4573 12115 4607
rect 13001 4573 13035 4607
rect 15761 4573 15795 4607
rect 18429 4573 18463 4607
rect 22569 4573 22603 4607
rect 22661 4573 22695 4607
rect 24225 4573 24259 4607
rect 9505 4505 9539 4539
rect 23673 4505 23707 4539
rect 8401 4437 8435 4471
rect 9137 4437 9171 4471
rect 11253 4437 11287 4471
rect 12541 4437 12575 4471
rect 19809 4437 19843 4471
rect 21189 4437 21223 4471
rect 8677 4233 8711 4267
rect 12817 4233 12851 4267
rect 14381 4233 14415 4267
rect 15669 4233 15703 4267
rect 18613 4233 18647 4267
rect 21005 4233 21039 4267
rect 23489 4233 23523 4267
rect 24409 4233 24443 4267
rect 25421 4233 25455 4267
rect 18337 4165 18371 4199
rect 22753 4165 22787 4199
rect 23121 4165 23155 4199
rect 8309 4097 8343 4131
rect 9229 4097 9263 4131
rect 9321 4097 9355 4131
rect 10977 4097 11011 4131
rect 13093 4097 13127 4131
rect 13921 4097 13955 4131
rect 14657 4097 14691 4131
rect 15301 4097 15335 4131
rect 17877 4097 17911 4131
rect 19349 4097 19383 4131
rect 19901 4097 19935 4131
rect 21833 4097 21867 4131
rect 25053 4097 25087 4131
rect 7665 4029 7699 4063
rect 9137 4029 9171 4063
rect 13645 4029 13679 4063
rect 15761 4029 15795 4063
rect 16028 4029 16062 4063
rect 19257 4029 19291 4063
rect 23949 4029 23983 4063
rect 24869 4029 24903 4063
rect 9965 3961 9999 3995
rect 19165 3961 19199 3995
rect 20177 3961 20211 3995
rect 20729 3961 20763 3995
rect 21649 3961 21683 3995
rect 7849 3893 7883 3927
rect 8769 3893 8803 3927
rect 10333 3893 10367 3927
rect 10701 3893 10735 3927
rect 10793 3893 10827 3927
rect 11437 3893 11471 3927
rect 11713 3893 11747 3927
rect 12081 3893 12115 3927
rect 13277 3893 13311 3927
rect 13737 3893 13771 3927
rect 17141 3893 17175 3927
rect 17417 3893 17451 3927
rect 18797 3893 18831 3927
rect 21281 3893 21315 3927
rect 21741 3893 21775 3927
rect 22293 3893 22327 3927
rect 24225 3893 24259 3927
rect 24777 3893 24811 3927
rect 8033 3689 8067 3723
rect 9505 3689 9539 3723
rect 12449 3689 12483 3723
rect 13001 3689 13035 3723
rect 14013 3689 14047 3723
rect 15025 3689 15059 3723
rect 15669 3689 15703 3723
rect 17693 3689 17727 3723
rect 18429 3689 18463 3723
rect 18797 3689 18831 3723
rect 23765 3689 23799 3723
rect 9045 3621 9079 3655
rect 13369 3621 13403 3655
rect 13921 3621 13955 3655
rect 16037 3621 16071 3655
rect 17601 3621 17635 3655
rect 19901 3621 19935 3655
rect 20729 3621 20763 3655
rect 24308 3621 24342 3655
rect 6929 3553 6963 3587
rect 8401 3553 8435 3587
rect 9965 3553 9999 3587
rect 11336 3553 11370 3587
rect 16681 3553 16715 3587
rect 19165 3553 19199 3587
rect 21649 3553 21683 3587
rect 21833 3553 21867 3587
rect 22089 3553 22123 3587
rect 8493 3485 8527 3519
rect 8677 3485 8711 3519
rect 11069 3485 11103 3519
rect 14197 3485 14231 3519
rect 16129 3485 16163 3519
rect 16313 3485 16347 3519
rect 17877 3485 17911 3519
rect 19257 3485 19291 3519
rect 19441 3485 19475 3519
rect 24041 3485 24075 3519
rect 7941 3417 7975 3451
rect 10517 3417 10551 3451
rect 13553 3417 13587 3451
rect 15577 3417 15611 3451
rect 17233 3417 17267 3451
rect 7113 3349 7147 3383
rect 7573 3349 7607 3383
rect 10149 3349 10183 3383
rect 10977 3349 11011 3383
rect 21373 3349 21407 3383
rect 23213 3349 23247 3383
rect 25421 3349 25455 3383
rect 5825 3145 5859 3179
rect 6285 3145 6319 3179
rect 6653 3145 6687 3179
rect 7021 3145 7055 3179
rect 9873 3145 9907 3179
rect 11529 3145 11563 3179
rect 11805 3145 11839 3179
rect 14105 3145 14139 3179
rect 15393 3145 15427 3179
rect 16865 3145 16899 3179
rect 17693 3145 17727 3179
rect 20085 3145 20119 3179
rect 20545 3145 20579 3179
rect 21097 3145 21131 3179
rect 25053 3145 25087 3179
rect 7665 3077 7699 3111
rect 8585 3077 8619 3111
rect 15025 3077 15059 3111
rect 17325 3077 17359 3111
rect 19717 3077 19751 3111
rect 23489 3077 23523 3111
rect 24777 3077 24811 3111
rect 8125 3009 8159 3043
rect 9229 3009 9263 3043
rect 9873 3009 9907 3043
rect 9965 3009 9999 3043
rect 10149 3009 10183 3043
rect 12449 3009 12483 3043
rect 15485 3009 15519 3043
rect 18061 3009 18095 3043
rect 21189 3009 21223 3043
rect 23121 3009 23155 3043
rect 24317 3009 24351 3043
rect 5641 2941 5675 2975
rect 7481 2941 7515 2975
rect 8493 2941 8527 2975
rect 8953 2941 8987 2975
rect 9045 2941 9079 2975
rect 24133 2941 24167 2975
rect 9597 2873 9631 2907
rect 10416 2873 10450 2907
rect 12265 2873 12299 2907
rect 12716 2873 12750 2907
rect 14657 2873 14691 2907
rect 15752 2873 15786 2907
rect 18306 2873 18340 2907
rect 21456 2873 21490 2907
rect 24041 2873 24075 2907
rect 13829 2805 13863 2839
rect 19441 2805 19475 2839
rect 22569 2805 22603 2839
rect 23673 2805 23707 2839
rect 25421 2805 25455 2839
rect 5641 2601 5675 2635
rect 6377 2601 6411 2635
rect 8125 2601 8159 2635
rect 11529 2601 11563 2635
rect 11897 2601 11931 2635
rect 14013 2601 14047 2635
rect 14749 2601 14783 2635
rect 16865 2601 16899 2635
rect 17233 2601 17267 2635
rect 17601 2601 17635 2635
rect 18153 2601 18187 2635
rect 20269 2601 20303 2635
rect 21005 2601 21039 2635
rect 22201 2601 22235 2635
rect 22937 2601 22971 2635
rect 25605 2601 25639 2635
rect 8033 2533 8067 2567
rect 8493 2533 8527 2567
rect 9597 2533 9631 2567
rect 15301 2533 15335 2567
rect 15752 2533 15786 2567
rect 18797 2533 18831 2567
rect 19156 2533 19190 2567
rect 24409 2533 24443 2567
rect 5733 2465 5767 2499
rect 6745 2465 6779 2499
rect 7021 2465 7055 2499
rect 10057 2465 10091 2499
rect 10416 2465 10450 2499
rect 12633 2465 12667 2499
rect 12900 2465 12934 2499
rect 14381 2465 14415 2499
rect 15485 2465 15519 2499
rect 18889 2465 18923 2499
rect 20637 2465 20671 2499
rect 22293 2465 22327 2499
rect 23489 2465 23523 2499
rect 24501 2465 24535 2499
rect 4721 2397 4755 2431
rect 7665 2397 7699 2431
rect 8585 2397 8619 2431
rect 8769 2397 8803 2431
rect 10149 2397 10183 2431
rect 12449 2397 12483 2431
rect 21649 2397 21683 2431
rect 22385 2397 22419 2431
rect 23857 2397 23891 2431
rect 24593 2397 24627 2431
rect 25053 2397 25087 2431
rect 21833 2329 21867 2363
rect 24041 2329 24075 2363
rect 5917 2261 5951 2295
rect 7205 2261 7239 2295
rect 9229 2261 9263 2295
<< metal1 >>
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 23477 24395 23535 24401
rect 23477 24361 23489 24395
rect 23523 24392 23535 24395
rect 24762 24392 24768 24404
rect 23523 24364 24768 24392
rect 23523 24361 23535 24364
rect 23477 24355 23535 24361
rect 24762 24352 24768 24364
rect 24820 24352 24826 24404
rect 24581 24259 24639 24265
rect 24581 24225 24593 24259
rect 24627 24256 24639 24259
rect 25222 24256 25228 24268
rect 24627 24228 25228 24256
rect 24627 24225 24639 24228
rect 24581 24219 24639 24225
rect 25222 24216 25228 24228
rect 25280 24216 25286 24268
rect 24762 24120 24768 24132
rect 24723 24092 24768 24120
rect 24762 24080 24768 24092
rect 24820 24080 24826 24132
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 24670 23808 24676 23860
rect 24728 23848 24734 23860
rect 24765 23851 24823 23857
rect 24765 23848 24777 23851
rect 24728 23820 24777 23848
rect 24728 23808 24734 23820
rect 24765 23817 24777 23820
rect 24811 23817 24823 23851
rect 24765 23811 24823 23817
rect 24394 23712 24400 23724
rect 24355 23684 24400 23712
rect 24394 23672 24400 23684
rect 24452 23712 24458 23724
rect 24452 23684 24624 23712
rect 24452 23672 24458 23684
rect 24596 23653 24624 23684
rect 24581 23647 24639 23653
rect 24581 23613 24593 23647
rect 24627 23613 24639 23647
rect 24581 23607 24639 23613
rect 25222 23508 25228 23520
rect 25183 23480 25228 23508
rect 25222 23468 25228 23480
rect 25280 23468 25286 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 24118 23264 24124 23316
rect 24176 23304 24182 23316
rect 24765 23307 24823 23313
rect 24765 23304 24777 23307
rect 24176 23276 24777 23304
rect 24176 23264 24182 23276
rect 24765 23273 24777 23276
rect 24811 23273 24823 23307
rect 24765 23267 24823 23273
rect 12802 23236 12808 23248
rect 12763 23208 12808 23236
rect 12802 23196 12808 23208
rect 12860 23196 12866 23248
rect 12526 23168 12532 23180
rect 12487 23140 12532 23168
rect 12526 23128 12532 23140
rect 12584 23128 12590 23180
rect 23842 23128 23848 23180
rect 23900 23168 23906 23180
rect 24581 23171 24639 23177
rect 24581 23168 24593 23171
rect 23900 23140 24593 23168
rect 23900 23128 23906 23140
rect 24581 23137 24593 23140
rect 24627 23137 24639 23171
rect 24581 23131 24639 23137
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 24762 22760 24768 22772
rect 24723 22732 24768 22760
rect 24762 22720 24768 22732
rect 24820 22720 24826 22772
rect 25222 22584 25228 22636
rect 25280 22624 25286 22636
rect 26234 22624 26240 22636
rect 25280 22596 26240 22624
rect 25280 22584 25286 22596
rect 26234 22584 26240 22596
rect 26292 22584 26298 22636
rect 24578 22556 24584 22568
rect 24539 22528 24584 22556
rect 24578 22516 24584 22528
rect 24636 22556 24642 22568
rect 25133 22559 25191 22565
rect 25133 22556 25145 22559
rect 24636 22528 25145 22556
rect 24636 22516 24642 22528
rect 25133 22525 25145 22528
rect 25179 22525 25191 22559
rect 25133 22519 25191 22525
rect 11974 22380 11980 22432
rect 12032 22420 12038 22432
rect 12526 22420 12532 22432
rect 12032 22392 12532 22420
rect 12032 22380 12038 22392
rect 12526 22380 12532 22392
rect 12584 22420 12590 22432
rect 12621 22423 12679 22429
rect 12621 22420 12633 22423
rect 12584 22392 12633 22420
rect 12584 22380 12590 22392
rect 12621 22389 12633 22392
rect 12667 22389 12679 22423
rect 12621 22383 12679 22389
rect 23842 22380 23848 22432
rect 23900 22420 23906 22432
rect 24397 22423 24455 22429
rect 24397 22420 24409 22423
rect 23900 22392 24409 22420
rect 23900 22380 23906 22392
rect 24397 22389 24409 22392
rect 24443 22389 24455 22423
rect 24397 22383 24455 22389
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 23842 22148 23848 22160
rect 23803 22120 23848 22148
rect 23842 22108 23848 22120
rect 23900 22108 23906 22160
rect 23474 22040 23480 22092
rect 23532 22080 23538 22092
rect 23569 22083 23627 22089
rect 23569 22080 23581 22083
rect 23532 22052 23581 22080
rect 23532 22040 23538 22052
rect 23569 22049 23581 22052
rect 23615 22049 23627 22083
rect 24854 22080 24860 22092
rect 24815 22052 24860 22080
rect 23569 22043 23627 22049
rect 24854 22040 24860 22052
rect 24912 22040 24918 22092
rect 23382 21972 23388 22024
rect 23440 22012 23446 22024
rect 24210 22012 24216 22024
rect 23440 21984 24216 22012
rect 23440 21972 23446 21984
rect 24210 21972 24216 21984
rect 24268 21972 24274 22024
rect 25038 21944 25044 21956
rect 24999 21916 25044 21944
rect 25038 21904 25044 21916
rect 25096 21904 25102 21956
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 24854 21672 24860 21684
rect 24815 21644 24860 21672
rect 24854 21632 24860 21644
rect 24912 21632 24918 21684
rect 25130 21672 25136 21684
rect 25091 21644 25136 21672
rect 25130 21632 25136 21644
rect 25188 21632 25194 21684
rect 14550 21536 14556 21548
rect 14511 21508 14556 21536
rect 14550 21496 14556 21508
rect 14608 21496 14614 21548
rect 23937 21539 23995 21545
rect 23937 21505 23949 21539
rect 23983 21536 23995 21539
rect 24872 21536 24900 21632
rect 23983 21508 24900 21536
rect 23983 21505 23995 21508
rect 23937 21499 23995 21505
rect 13998 21428 14004 21480
rect 14056 21468 14062 21480
rect 14277 21471 14335 21477
rect 14277 21468 14289 21471
rect 14056 21440 14289 21468
rect 14056 21428 14062 21440
rect 14277 21437 14289 21440
rect 14323 21468 14335 21471
rect 15013 21471 15071 21477
rect 15013 21468 15025 21471
rect 14323 21440 15025 21468
rect 14323 21437 14335 21440
rect 14277 21431 14335 21437
rect 15013 21437 15025 21440
rect 15059 21437 15071 21471
rect 23474 21468 23480 21480
rect 23435 21440 23480 21468
rect 15013 21431 15071 21437
rect 23474 21428 23480 21440
rect 23532 21428 23538 21480
rect 23566 21428 23572 21480
rect 23624 21468 23630 21480
rect 23661 21471 23719 21477
rect 23661 21468 23673 21471
rect 23624 21440 23673 21468
rect 23624 21428 23630 21440
rect 23661 21437 23673 21440
rect 23707 21437 23719 21471
rect 23661 21431 23719 21437
rect 23676 21400 23704 21431
rect 23750 21428 23756 21480
rect 23808 21468 23814 21480
rect 24949 21471 25007 21477
rect 24949 21468 24961 21471
rect 23808 21440 24961 21468
rect 23808 21428 23814 21440
rect 24949 21437 24961 21440
rect 24995 21468 25007 21471
rect 25501 21471 25559 21477
rect 25501 21468 25513 21471
rect 24995 21440 25513 21468
rect 24995 21437 25007 21440
rect 24949 21431 25007 21437
rect 25501 21437 25513 21440
rect 25547 21437 25559 21471
rect 25501 21431 25559 21437
rect 24397 21403 24455 21409
rect 24397 21400 24409 21403
rect 23676 21372 24409 21400
rect 24397 21369 24409 21372
rect 24443 21369 24455 21403
rect 24397 21363 24455 21369
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 25041 21131 25099 21137
rect 25041 21097 25053 21131
rect 25087 21128 25099 21131
rect 25222 21128 25228 21140
rect 25087 21100 25228 21128
rect 25087 21097 25099 21100
rect 25041 21091 25099 21097
rect 25222 21088 25228 21100
rect 25280 21088 25286 21140
rect 23569 20995 23627 21001
rect 23569 20961 23581 20995
rect 23615 20992 23627 20995
rect 23842 20992 23848 21004
rect 23615 20964 23848 20992
rect 23615 20961 23627 20964
rect 23569 20955 23627 20961
rect 23842 20952 23848 20964
rect 23900 20952 23906 21004
rect 24854 20992 24860 21004
rect 24815 20964 24860 20992
rect 24854 20952 24860 20964
rect 24912 20952 24918 21004
rect 23750 20924 23756 20936
rect 23711 20896 23756 20924
rect 23750 20884 23756 20896
rect 23808 20884 23814 20936
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 16850 20584 16856 20596
rect 16811 20556 16856 20584
rect 16850 20544 16856 20556
rect 16908 20544 16914 20596
rect 24670 20544 24676 20596
rect 24728 20584 24734 20596
rect 24765 20587 24823 20593
rect 24765 20584 24777 20587
rect 24728 20556 24777 20584
rect 24728 20544 24734 20556
rect 24765 20553 24777 20556
rect 24811 20553 24823 20587
rect 24765 20547 24823 20553
rect 16574 20340 16580 20392
rect 16632 20380 16638 20392
rect 16669 20383 16727 20389
rect 16669 20380 16681 20383
rect 16632 20352 16681 20380
rect 16632 20340 16638 20352
rect 16669 20349 16681 20352
rect 16715 20380 16727 20383
rect 17221 20383 17279 20389
rect 17221 20380 17233 20383
rect 16715 20352 17233 20380
rect 16715 20349 16727 20352
rect 16669 20343 16727 20349
rect 17221 20349 17233 20352
rect 17267 20349 17279 20383
rect 17221 20343 17279 20349
rect 23934 20340 23940 20392
rect 23992 20380 23998 20392
rect 24581 20383 24639 20389
rect 24581 20380 24593 20383
rect 23992 20352 24593 20380
rect 23992 20340 23998 20352
rect 24581 20349 24593 20352
rect 24627 20380 24639 20383
rect 25133 20383 25191 20389
rect 25133 20380 25145 20383
rect 24627 20352 25145 20380
rect 24627 20349 24639 20352
rect 24581 20343 24639 20349
rect 25133 20349 25145 20352
rect 25179 20349 25191 20383
rect 25133 20343 25191 20349
rect 23842 20244 23848 20256
rect 23803 20216 23848 20244
rect 23842 20204 23848 20216
rect 23900 20204 23906 20256
rect 25498 20244 25504 20256
rect 25459 20216 25504 20244
rect 25498 20204 25504 20216
rect 25556 20204 25562 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 17304 19975 17362 19981
rect 17304 19941 17316 19975
rect 17350 19972 17362 19975
rect 17494 19972 17500 19984
rect 17350 19944 17500 19972
rect 17350 19941 17362 19944
rect 17304 19935 17362 19941
rect 17494 19932 17500 19944
rect 17552 19932 17558 19984
rect 23753 19975 23811 19981
rect 23753 19941 23765 19975
rect 23799 19972 23811 19975
rect 24854 19972 24860 19984
rect 23799 19944 24860 19972
rect 23799 19941 23811 19944
rect 23753 19935 23811 19941
rect 24854 19932 24860 19944
rect 24912 19972 24918 19984
rect 25498 19972 25504 19984
rect 24912 19944 25504 19972
rect 24912 19932 24918 19944
rect 25498 19932 25504 19944
rect 25556 19932 25562 19984
rect 23474 19904 23480 19916
rect 23435 19876 23480 19904
rect 23474 19864 23480 19876
rect 23532 19864 23538 19916
rect 17034 19836 17040 19848
rect 16995 19808 17040 19836
rect 17034 19796 17040 19808
rect 17092 19796 17098 19848
rect 18230 19660 18236 19712
rect 18288 19700 18294 19712
rect 18417 19703 18475 19709
rect 18417 19700 18429 19703
rect 18288 19672 18429 19700
rect 18288 19660 18294 19672
rect 18417 19669 18429 19672
rect 18463 19669 18475 19703
rect 18417 19663 18475 19669
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 17129 19499 17187 19505
rect 17129 19465 17141 19499
rect 17175 19496 17187 19499
rect 17494 19496 17500 19508
rect 17175 19468 17500 19496
rect 17175 19465 17187 19468
rect 17129 19459 17187 19465
rect 17494 19456 17500 19468
rect 17552 19456 17558 19508
rect 17034 19388 17040 19440
rect 17092 19428 17098 19440
rect 17405 19431 17463 19437
rect 17405 19428 17417 19431
rect 17092 19400 17417 19428
rect 17092 19388 17098 19400
rect 17405 19397 17417 19400
rect 17451 19428 17463 19431
rect 17862 19428 17868 19440
rect 17451 19400 17868 19428
rect 17451 19397 17463 19400
rect 17405 19391 17463 19397
rect 17862 19388 17868 19400
rect 17920 19388 17926 19440
rect 23934 19360 23940 19372
rect 23895 19332 23940 19360
rect 23934 19320 23940 19332
rect 23992 19320 23998 19372
rect 15286 19252 15292 19304
rect 15344 19292 15350 19304
rect 15657 19295 15715 19301
rect 15657 19292 15669 19295
rect 15344 19264 15669 19292
rect 15344 19252 15350 19264
rect 15657 19261 15669 19264
rect 15703 19261 15715 19295
rect 15657 19255 15715 19261
rect 15933 19295 15991 19301
rect 15933 19261 15945 19295
rect 15979 19292 15991 19295
rect 16482 19292 16488 19304
rect 15979 19264 16488 19292
rect 15979 19261 15991 19264
rect 15933 19255 15991 19261
rect 15672 19224 15700 19255
rect 16482 19252 16488 19264
rect 16540 19252 16546 19304
rect 23658 19292 23664 19304
rect 23619 19264 23664 19292
rect 23658 19252 23664 19264
rect 23716 19292 23722 19304
rect 24397 19295 24455 19301
rect 24397 19292 24409 19295
rect 23716 19264 24409 19292
rect 23716 19252 23722 19264
rect 24397 19261 24409 19264
rect 24443 19261 24455 19295
rect 24946 19292 24952 19304
rect 24907 19264 24952 19292
rect 24397 19255 24455 19261
rect 24946 19252 24952 19264
rect 25004 19292 25010 19304
rect 25501 19295 25559 19301
rect 25501 19292 25513 19295
rect 25004 19264 25513 19292
rect 25004 19252 25010 19264
rect 25501 19261 25513 19264
rect 25547 19261 25559 19295
rect 25501 19255 25559 19261
rect 26234 19252 26240 19304
rect 26292 19292 26298 19304
rect 26878 19292 26884 19304
rect 26292 19264 26884 19292
rect 26292 19252 26298 19264
rect 26878 19252 26884 19264
rect 26936 19252 26942 19304
rect 16393 19227 16451 19233
rect 16393 19224 16405 19227
rect 15672 19196 16405 19224
rect 16393 19193 16405 19196
rect 16439 19193 16451 19227
rect 16393 19187 16451 19193
rect 23474 19156 23480 19168
rect 23435 19128 23480 19156
rect 23474 19116 23480 19128
rect 23532 19116 23538 19168
rect 24854 19116 24860 19168
rect 24912 19156 24918 19168
rect 25133 19159 25191 19165
rect 25133 19156 25145 19159
rect 24912 19128 25145 19156
rect 24912 19116 24918 19128
rect 25133 19125 25145 19128
rect 25179 19125 25191 19159
rect 25133 19119 25191 19125
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 24670 18912 24676 18964
rect 24728 18952 24734 18964
rect 24765 18955 24823 18961
rect 24765 18952 24777 18955
rect 24728 18924 24777 18952
rect 24728 18912 24734 18924
rect 24765 18921 24777 18924
rect 24811 18921 24823 18955
rect 24765 18915 24823 18921
rect 24578 18816 24584 18828
rect 24539 18788 24584 18816
rect 24578 18776 24584 18788
rect 24636 18776 24642 18828
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 14826 18368 14832 18420
rect 14884 18408 14890 18420
rect 15013 18411 15071 18417
rect 15013 18408 15025 18411
rect 14884 18380 15025 18408
rect 14884 18368 14890 18380
rect 15013 18377 15025 18380
rect 15059 18377 15071 18411
rect 24670 18408 24676 18420
rect 24631 18380 24676 18408
rect 15013 18371 15071 18377
rect 24670 18368 24676 18380
rect 24728 18368 24734 18420
rect 13538 18204 13544 18216
rect 13499 18176 13544 18204
rect 13538 18164 13544 18176
rect 13596 18204 13602 18216
rect 14277 18207 14335 18213
rect 14277 18204 14289 18207
rect 13596 18176 14289 18204
rect 13596 18164 13602 18176
rect 14277 18173 14289 18176
rect 14323 18173 14335 18207
rect 14277 18167 14335 18173
rect 14829 18207 14887 18213
rect 14829 18173 14841 18207
rect 14875 18173 14887 18207
rect 14829 18167 14887 18173
rect 13814 18136 13820 18148
rect 13775 18108 13820 18136
rect 13814 18096 13820 18108
rect 13872 18096 13878 18148
rect 13906 18096 13912 18148
rect 13964 18136 13970 18148
rect 14844 18136 14872 18167
rect 15381 18139 15439 18145
rect 15381 18136 15393 18139
rect 13964 18108 15393 18136
rect 13964 18096 13970 18108
rect 15381 18105 15393 18108
rect 15427 18105 15439 18139
rect 15381 18099 15439 18105
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 24762 17864 24768 17876
rect 24723 17836 24768 17864
rect 24762 17824 24768 17836
rect 24820 17824 24826 17876
rect 11606 17796 11612 17808
rect 11567 17768 11612 17796
rect 11606 17756 11612 17768
rect 11664 17756 11670 17808
rect 11333 17731 11391 17737
rect 11333 17697 11345 17731
rect 11379 17728 11391 17731
rect 11422 17728 11428 17740
rect 11379 17700 11428 17728
rect 11379 17697 11391 17700
rect 11333 17691 11391 17697
rect 11422 17688 11428 17700
rect 11480 17688 11486 17740
rect 24581 17731 24639 17737
rect 24581 17697 24593 17731
rect 24627 17728 24639 17731
rect 25038 17728 25044 17740
rect 24627 17700 25044 17728
rect 24627 17697 24639 17700
rect 24581 17691 24639 17697
rect 25038 17688 25044 17700
rect 25096 17688 25102 17740
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 24670 17280 24676 17332
rect 24728 17320 24734 17332
rect 24765 17323 24823 17329
rect 24765 17320 24777 17323
rect 24728 17292 24777 17320
rect 24728 17280 24734 17292
rect 24765 17289 24777 17292
rect 24811 17289 24823 17323
rect 24765 17283 24823 17289
rect 13449 17187 13507 17193
rect 13449 17153 13461 17187
rect 13495 17184 13507 17187
rect 13722 17184 13728 17196
rect 13495 17156 13728 17184
rect 13495 17153 13507 17156
rect 13449 17147 13507 17153
rect 13722 17144 13728 17156
rect 13780 17144 13786 17196
rect 13170 17116 13176 17128
rect 13131 17088 13176 17116
rect 13170 17076 13176 17088
rect 13228 17116 13234 17128
rect 13909 17119 13967 17125
rect 13909 17116 13921 17119
rect 13228 17088 13921 17116
rect 13228 17076 13234 17088
rect 13909 17085 13921 17088
rect 13955 17085 13967 17119
rect 24581 17119 24639 17125
rect 24581 17116 24593 17119
rect 13909 17079 13967 17085
rect 24412 17088 24593 17116
rect 11425 16983 11483 16989
rect 11425 16949 11437 16983
rect 11471 16980 11483 16983
rect 11514 16980 11520 16992
rect 11471 16952 11520 16980
rect 11471 16949 11483 16952
rect 11425 16943 11483 16949
rect 11514 16940 11520 16952
rect 11572 16940 11578 16992
rect 23934 16940 23940 16992
rect 23992 16980 23998 16992
rect 24412 16989 24440 17088
rect 24581 17085 24593 17088
rect 24627 17085 24639 17119
rect 24581 17079 24639 17085
rect 24397 16983 24455 16989
rect 24397 16980 24409 16983
rect 23992 16952 24409 16980
rect 23992 16940 23998 16952
rect 24397 16949 24409 16952
rect 24443 16949 24455 16983
rect 24397 16943 24455 16949
rect 25038 16940 25044 16992
rect 25096 16980 25102 16992
rect 25133 16983 25191 16989
rect 25133 16980 25145 16983
rect 25096 16952 25145 16980
rect 25096 16940 25102 16952
rect 25133 16949 25145 16952
rect 25179 16949 25191 16983
rect 25133 16943 25191 16949
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 22922 16776 22928 16788
rect 22883 16748 22928 16776
rect 22922 16736 22928 16748
rect 22980 16736 22986 16788
rect 16301 16643 16359 16649
rect 16301 16609 16313 16643
rect 16347 16609 16359 16643
rect 16574 16640 16580 16652
rect 16535 16612 16580 16640
rect 16301 16603 16359 16609
rect 16316 16572 16344 16603
rect 16574 16600 16580 16612
rect 16632 16600 16638 16652
rect 22738 16640 22744 16652
rect 22699 16612 22744 16640
rect 22738 16600 22744 16612
rect 22796 16600 22802 16652
rect 16482 16572 16488 16584
rect 16316 16544 16488 16572
rect 16482 16532 16488 16544
rect 16540 16532 16546 16584
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 25130 16232 25136 16244
rect 25091 16204 25136 16232
rect 25130 16192 25136 16204
rect 25188 16192 25194 16244
rect 23934 16096 23940 16108
rect 23895 16068 23940 16096
rect 23934 16056 23940 16068
rect 23992 16056 23998 16108
rect 23658 16028 23664 16040
rect 23619 16000 23664 16028
rect 23658 15988 23664 16000
rect 23716 16028 23722 16040
rect 24397 16031 24455 16037
rect 24397 16028 24409 16031
rect 23716 16000 24409 16028
rect 23716 15988 23722 16000
rect 24397 15997 24409 16000
rect 24443 15997 24455 16031
rect 24397 15991 24455 15997
rect 24854 15988 24860 16040
rect 24912 16028 24918 16040
rect 24949 16031 25007 16037
rect 24949 16028 24961 16031
rect 24912 16000 24961 16028
rect 24912 15988 24918 16000
rect 24949 15997 24961 16000
rect 24995 16028 25007 16031
rect 25501 16031 25559 16037
rect 25501 16028 25513 16031
rect 24995 16000 25513 16028
rect 24995 15997 25007 16000
rect 24949 15991 25007 15997
rect 25501 15997 25513 16000
rect 25547 15997 25559 16031
rect 25501 15991 25559 15997
rect 16393 15895 16451 15901
rect 16393 15861 16405 15895
rect 16439 15892 16451 15895
rect 16482 15892 16488 15904
rect 16439 15864 16488 15892
rect 16439 15861 16451 15864
rect 16393 15855 16451 15861
rect 16482 15852 16488 15864
rect 16540 15852 16546 15904
rect 22186 15852 22192 15904
rect 22244 15892 22250 15904
rect 22738 15892 22744 15904
rect 22244 15864 22744 15892
rect 22244 15852 22250 15864
rect 22738 15852 22744 15864
rect 22796 15852 22802 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 23382 15688 23388 15700
rect 23343 15660 23388 15688
rect 23382 15648 23388 15660
rect 23440 15648 23446 15700
rect 22186 15620 22192 15632
rect 22147 15592 22192 15620
rect 22186 15580 22192 15592
rect 22244 15580 22250 15632
rect 21910 15552 21916 15564
rect 21871 15524 21916 15552
rect 21910 15512 21916 15524
rect 21968 15512 21974 15564
rect 23198 15552 23204 15564
rect 23159 15524 23204 15552
rect 23198 15512 23204 15524
rect 23256 15512 23262 15564
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 25866 15144 25872 15156
rect 25827 15116 25872 15144
rect 25866 15104 25872 15116
rect 25924 15104 25930 15156
rect 24213 15011 24271 15017
rect 24213 14977 24225 15011
rect 24259 15008 24271 15011
rect 24762 15008 24768 15020
rect 24259 14980 24768 15008
rect 24259 14977 24271 14980
rect 24213 14971 24271 14977
rect 24762 14968 24768 14980
rect 24820 14968 24826 15020
rect 23842 14900 23848 14952
rect 23900 14940 23906 14952
rect 23937 14943 23995 14949
rect 23937 14940 23949 14943
rect 23900 14912 23949 14940
rect 23900 14900 23906 14912
rect 23937 14909 23949 14912
rect 23983 14940 23995 14943
rect 24673 14943 24731 14949
rect 24673 14940 24685 14943
rect 23983 14912 24685 14940
rect 23983 14909 23995 14912
rect 23937 14903 23995 14909
rect 24673 14909 24685 14912
rect 24719 14909 24731 14943
rect 24673 14903 24731 14909
rect 25225 14943 25283 14949
rect 25225 14909 25237 14943
rect 25271 14940 25283 14943
rect 25866 14940 25872 14952
rect 25271 14912 25872 14940
rect 25271 14909 25283 14912
rect 25225 14903 25283 14909
rect 25866 14900 25872 14912
rect 25924 14900 25930 14952
rect 21910 14804 21916 14816
rect 21871 14776 21916 14804
rect 21910 14764 21916 14776
rect 21968 14764 21974 14816
rect 22462 14764 22468 14816
rect 22520 14804 22526 14816
rect 23198 14804 23204 14816
rect 22520 14776 23204 14804
rect 22520 14764 22526 14776
rect 23198 14764 23204 14776
rect 23256 14764 23262 14816
rect 25409 14807 25467 14813
rect 25409 14773 25421 14807
rect 25455 14804 25467 14807
rect 25682 14804 25688 14816
rect 25455 14776 25688 14804
rect 25455 14773 25467 14776
rect 25409 14767 25467 14773
rect 25682 14764 25688 14776
rect 25740 14764 25746 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 24670 14560 24676 14612
rect 24728 14600 24734 14612
rect 24765 14603 24823 14609
rect 24765 14600 24777 14603
rect 24728 14572 24777 14600
rect 24728 14560 24734 14572
rect 24765 14569 24777 14572
rect 24811 14569 24823 14603
rect 24765 14563 24823 14569
rect 22462 14532 22468 14544
rect 22423 14504 22468 14532
rect 22462 14492 22468 14504
rect 22520 14492 22526 14544
rect 22189 14467 22247 14473
rect 22189 14433 22201 14467
rect 22235 14464 22247 14467
rect 22738 14464 22744 14476
rect 22235 14436 22744 14464
rect 22235 14433 22247 14436
rect 22189 14427 22247 14433
rect 22738 14424 22744 14436
rect 22796 14424 22802 14476
rect 24581 14467 24639 14473
rect 24581 14433 24593 14467
rect 24627 14464 24639 14467
rect 24670 14464 24676 14476
rect 24627 14436 24676 14464
rect 24627 14433 24639 14436
rect 24581 14427 24639 14433
rect 24670 14424 24676 14436
rect 24728 14424 24734 14476
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 17862 14016 17868 14068
rect 17920 14056 17926 14068
rect 18322 14056 18328 14068
rect 17920 14028 18328 14056
rect 17920 14016 17926 14028
rect 18322 14016 18328 14028
rect 18380 14056 18386 14068
rect 18877 14059 18935 14065
rect 18877 14056 18889 14059
rect 18380 14028 18889 14056
rect 18380 14016 18386 14028
rect 18877 14025 18889 14028
rect 18923 14025 18935 14059
rect 24670 14056 24676 14068
rect 18877 14019 18935 14025
rect 23952 14028 24676 14056
rect 23952 13929 23980 14028
rect 24670 14016 24676 14028
rect 24728 14016 24734 14068
rect 25590 14056 25596 14068
rect 25551 14028 25596 14056
rect 25590 14016 25596 14028
rect 25648 14016 25654 14068
rect 25130 13988 25136 14000
rect 25091 13960 25136 13988
rect 25130 13948 25136 13960
rect 25188 13948 25194 14000
rect 23937 13923 23995 13929
rect 23937 13889 23949 13923
rect 23983 13889 23995 13923
rect 23937 13883 23995 13889
rect 22649 13855 22707 13861
rect 22649 13821 22661 13855
rect 22695 13852 22707 13855
rect 22738 13852 22744 13864
rect 22695 13824 22744 13852
rect 22695 13821 22707 13824
rect 22649 13815 22707 13821
rect 22738 13812 22744 13824
rect 22796 13812 22802 13864
rect 23477 13855 23535 13861
rect 23477 13821 23489 13855
rect 23523 13852 23535 13855
rect 23661 13855 23719 13861
rect 23661 13852 23673 13855
rect 23523 13824 23673 13852
rect 23523 13821 23535 13824
rect 23477 13815 23535 13821
rect 23661 13821 23673 13824
rect 23707 13852 23719 13855
rect 24026 13852 24032 13864
rect 23707 13824 24032 13852
rect 23707 13821 23719 13824
rect 23661 13815 23719 13821
rect 24026 13812 24032 13824
rect 24084 13812 24090 13864
rect 24949 13855 25007 13861
rect 24949 13821 24961 13855
rect 24995 13852 25007 13855
rect 25590 13852 25596 13864
rect 24995 13824 25596 13852
rect 24995 13821 25007 13824
rect 24949 13815 25007 13821
rect 25590 13812 25596 13824
rect 25648 13812 25654 13864
rect 19242 13716 19248 13728
rect 19203 13688 19248 13716
rect 19242 13676 19248 13688
rect 19300 13676 19306 13728
rect 19518 13676 19524 13728
rect 19576 13716 19582 13728
rect 19613 13719 19671 13725
rect 19613 13716 19625 13719
rect 19576 13688 19625 13716
rect 19576 13676 19582 13688
rect 19613 13685 19625 13688
rect 19659 13685 19671 13719
rect 19613 13679 19671 13685
rect 21085 13719 21143 13725
rect 21085 13685 21097 13719
rect 21131 13716 21143 13719
rect 21634 13716 21640 13728
rect 21131 13688 21640 13716
rect 21131 13685 21143 13688
rect 21085 13679 21143 13685
rect 21634 13676 21640 13688
rect 21692 13676 21698 13728
rect 22094 13676 22100 13728
rect 22152 13716 22158 13728
rect 22152 13688 22197 13716
rect 22152 13676 22158 13688
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 19150 13472 19156 13524
rect 19208 13512 19214 13524
rect 19245 13515 19303 13521
rect 19245 13512 19257 13515
rect 19208 13484 19257 13512
rect 19208 13472 19214 13484
rect 19245 13481 19257 13484
rect 19291 13481 19303 13515
rect 19245 13475 19303 13481
rect 24210 13472 24216 13524
rect 24268 13512 24274 13524
rect 24765 13515 24823 13521
rect 24765 13512 24777 13515
rect 24268 13484 24777 13512
rect 24268 13472 24274 13484
rect 24765 13481 24777 13484
rect 24811 13481 24823 13515
rect 24765 13475 24823 13481
rect 18506 13336 18512 13388
rect 18564 13376 18570 13388
rect 19518 13376 19524 13388
rect 18564 13348 19524 13376
rect 18564 13336 18570 13348
rect 19518 13336 19524 13348
rect 19576 13376 19582 13388
rect 19613 13379 19671 13385
rect 19613 13376 19625 13379
rect 19576 13348 19625 13376
rect 19576 13336 19582 13348
rect 19613 13345 19625 13348
rect 19659 13345 19671 13379
rect 23474 13376 23480 13388
rect 23435 13348 23480 13376
rect 19613 13339 19671 13345
rect 23474 13336 23480 13348
rect 23532 13336 23538 13388
rect 24581 13379 24639 13385
rect 24581 13345 24593 13379
rect 24627 13376 24639 13379
rect 24670 13376 24676 13388
rect 24627 13348 24676 13376
rect 24627 13345 24639 13348
rect 24581 13339 24639 13345
rect 24670 13336 24676 13348
rect 24728 13336 24734 13388
rect 19242 13268 19248 13320
rect 19300 13308 19306 13320
rect 19705 13311 19763 13317
rect 19705 13308 19717 13311
rect 19300 13280 19717 13308
rect 19300 13268 19306 13280
rect 19705 13277 19717 13280
rect 19751 13277 19763 13311
rect 19705 13271 19763 13277
rect 19797 13311 19855 13317
rect 19797 13277 19809 13311
rect 19843 13308 19855 13311
rect 20070 13308 20076 13320
rect 19843 13280 20076 13308
rect 19843 13277 19855 13280
rect 19797 13271 19855 13277
rect 20070 13268 20076 13280
rect 20128 13268 20134 13320
rect 21453 13311 21511 13317
rect 21453 13277 21465 13311
rect 21499 13308 21511 13311
rect 21542 13308 21548 13320
rect 21499 13280 21548 13308
rect 21499 13277 21511 13280
rect 21453 13271 21511 13277
rect 21542 13268 21548 13280
rect 21600 13268 21606 13320
rect 22465 13311 22523 13317
rect 22465 13277 22477 13311
rect 22511 13308 22523 13311
rect 22554 13308 22560 13320
rect 22511 13280 22560 13308
rect 22511 13277 22523 13280
rect 22465 13271 22523 13277
rect 22554 13268 22560 13280
rect 22612 13268 22618 13320
rect 18693 13243 18751 13249
rect 18693 13209 18705 13243
rect 18739 13240 18751 13243
rect 19518 13240 19524 13252
rect 18739 13212 19524 13240
rect 18739 13209 18751 13212
rect 18693 13203 18751 13209
rect 19518 13200 19524 13212
rect 19576 13200 19582 13252
rect 23658 13240 23664 13252
rect 23619 13212 23664 13240
rect 23658 13200 23664 13212
rect 23716 13200 23722 13252
rect 19061 13175 19119 13181
rect 19061 13141 19073 13175
rect 19107 13172 19119 13175
rect 19426 13172 19432 13184
rect 19107 13144 19432 13172
rect 19107 13141 19119 13144
rect 19061 13135 19119 13141
rect 19426 13132 19432 13144
rect 19484 13132 19490 13184
rect 21174 13172 21180 13184
rect 21135 13144 21180 13172
rect 21174 13132 21180 13144
rect 21232 13132 21238 13184
rect 23934 13132 23940 13184
rect 23992 13172 23998 13184
rect 24029 13175 24087 13181
rect 24029 13172 24041 13175
rect 23992 13144 24041 13172
rect 23992 13132 23998 13144
rect 24029 13141 24041 13144
rect 24075 13141 24087 13175
rect 24029 13135 24087 13141
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 18506 12968 18512 12980
rect 18467 12940 18512 12968
rect 18506 12928 18512 12940
rect 18564 12928 18570 12980
rect 18969 12971 19027 12977
rect 18969 12937 18981 12971
rect 19015 12968 19027 12971
rect 19242 12968 19248 12980
rect 19015 12940 19248 12968
rect 19015 12937 19027 12940
rect 18969 12931 19027 12937
rect 19242 12928 19248 12940
rect 19300 12928 19306 12980
rect 20257 12971 20315 12977
rect 20257 12937 20269 12971
rect 20303 12968 20315 12971
rect 21266 12968 21272 12980
rect 20303 12940 21272 12968
rect 20303 12937 20315 12940
rect 20257 12931 20315 12937
rect 21266 12928 21272 12940
rect 21324 12928 21330 12980
rect 23474 12968 23480 12980
rect 23435 12940 23480 12968
rect 23474 12928 23480 12940
rect 23532 12928 23538 12980
rect 23934 12968 23940 12980
rect 23676 12940 23940 12968
rect 19334 12860 19340 12912
rect 19392 12900 19398 12912
rect 22646 12900 22652 12912
rect 19392 12872 22508 12900
rect 22607 12872 22652 12900
rect 19392 12860 19398 12872
rect 19518 12832 19524 12844
rect 19479 12804 19524 12832
rect 19518 12792 19524 12804
rect 19576 12792 19582 12844
rect 21174 12792 21180 12844
rect 21232 12832 21238 12844
rect 21269 12835 21327 12841
rect 21269 12832 21281 12835
rect 21232 12804 21281 12832
rect 21232 12792 21238 12804
rect 21269 12801 21281 12804
rect 21315 12801 21327 12835
rect 22480 12832 22508 12872
rect 22646 12860 22652 12872
rect 22704 12860 22710 12912
rect 23676 12832 23704 12940
rect 23934 12928 23940 12940
rect 23992 12928 23998 12980
rect 24670 12968 24676 12980
rect 24631 12940 24676 12968
rect 24670 12928 24676 12940
rect 24728 12928 24734 12980
rect 24946 12928 24952 12980
rect 25004 12968 25010 12980
rect 25133 12971 25191 12977
rect 25133 12968 25145 12971
rect 25004 12940 25145 12968
rect 25004 12928 25010 12940
rect 25133 12937 25145 12940
rect 25179 12937 25191 12971
rect 25133 12931 25191 12937
rect 22480 12804 23704 12832
rect 21269 12795 21327 12801
rect 19150 12724 19156 12776
rect 19208 12764 19214 12776
rect 19426 12764 19432 12776
rect 19208 12736 19432 12764
rect 19208 12724 19214 12736
rect 19426 12724 19432 12736
rect 19484 12724 19490 12776
rect 23676 12773 23704 12804
rect 23937 12835 23995 12841
rect 23937 12801 23949 12835
rect 23983 12832 23995 12835
rect 24688 12832 24716 12928
rect 23983 12804 24716 12832
rect 23983 12801 23995 12804
rect 23937 12795 23995 12801
rect 22465 12767 22523 12773
rect 22465 12733 22477 12767
rect 22511 12764 22523 12767
rect 23661 12767 23719 12773
rect 22511 12736 23152 12764
rect 22511 12733 22523 12736
rect 22465 12727 22523 12733
rect 18782 12696 18788 12708
rect 18743 12668 18788 12696
rect 18782 12656 18788 12668
rect 18840 12696 18846 12708
rect 19337 12699 19395 12705
rect 19337 12696 19349 12699
rect 18840 12668 19349 12696
rect 18840 12656 18846 12668
rect 19337 12665 19349 12668
rect 19383 12665 19395 12699
rect 19337 12659 19395 12665
rect 20625 12699 20683 12705
rect 20625 12665 20637 12699
rect 20671 12696 20683 12699
rect 21085 12699 21143 12705
rect 21085 12696 21097 12699
rect 20671 12668 21097 12696
rect 20671 12665 20683 12668
rect 20625 12659 20683 12665
rect 21085 12665 21097 12668
rect 21131 12696 21143 12699
rect 21358 12696 21364 12708
rect 21131 12668 21364 12696
rect 21131 12665 21143 12668
rect 21085 12659 21143 12665
rect 21358 12656 21364 12668
rect 21416 12656 21422 12708
rect 16206 12588 16212 12640
rect 16264 12628 16270 12640
rect 16761 12631 16819 12637
rect 16761 12628 16773 12631
rect 16264 12600 16773 12628
rect 16264 12588 16270 12600
rect 16761 12597 16773 12600
rect 16807 12597 16819 12631
rect 16761 12591 16819 12597
rect 20530 12588 20536 12640
rect 20588 12628 20594 12640
rect 20717 12631 20775 12637
rect 20717 12628 20729 12631
rect 20588 12600 20729 12628
rect 20588 12588 20594 12600
rect 20717 12597 20729 12600
rect 20763 12597 20775 12631
rect 20717 12591 20775 12597
rect 21177 12631 21235 12637
rect 21177 12597 21189 12631
rect 21223 12628 21235 12631
rect 21266 12628 21272 12640
rect 21223 12600 21272 12628
rect 21223 12597 21235 12600
rect 21177 12591 21235 12597
rect 21266 12588 21272 12600
rect 21324 12588 21330 12640
rect 21726 12628 21732 12640
rect 21687 12600 21732 12628
rect 21726 12588 21732 12600
rect 21784 12588 21790 12640
rect 23124 12637 23152 12736
rect 23661 12733 23673 12767
rect 23707 12733 23719 12767
rect 24946 12764 24952 12776
rect 24859 12736 24952 12764
rect 23661 12727 23719 12733
rect 24946 12724 24952 12736
rect 25004 12764 25010 12776
rect 25501 12767 25559 12773
rect 25501 12764 25513 12767
rect 25004 12736 25513 12764
rect 25004 12724 25010 12736
rect 25501 12733 25513 12736
rect 25547 12733 25559 12767
rect 25501 12727 25559 12733
rect 23109 12631 23167 12637
rect 23109 12597 23121 12631
rect 23155 12628 23167 12631
rect 23382 12628 23388 12640
rect 23155 12600 23388 12628
rect 23155 12597 23167 12600
rect 23109 12591 23167 12597
rect 23382 12588 23388 12600
rect 23440 12588 23446 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 17126 12424 17132 12436
rect 17087 12396 17132 12424
rect 17126 12384 17132 12396
rect 17184 12384 17190 12436
rect 18233 12427 18291 12433
rect 18233 12393 18245 12427
rect 18279 12424 18291 12427
rect 18322 12424 18328 12436
rect 18279 12396 18328 12424
rect 18279 12393 18291 12396
rect 18233 12387 18291 12393
rect 18322 12384 18328 12396
rect 18380 12384 18386 12436
rect 19058 12424 19064 12436
rect 19019 12396 19064 12424
rect 19058 12384 19064 12396
rect 19116 12384 19122 12436
rect 22738 12384 22744 12436
rect 22796 12424 22802 12436
rect 23109 12427 23167 12433
rect 23109 12424 23121 12427
rect 22796 12396 23121 12424
rect 22796 12384 22802 12396
rect 23109 12393 23121 12396
rect 23155 12393 23167 12427
rect 23109 12387 23167 12393
rect 18969 12359 19027 12365
rect 18969 12325 18981 12359
rect 19015 12356 19027 12359
rect 19242 12356 19248 12368
rect 19015 12328 19248 12356
rect 19015 12325 19027 12328
rect 18969 12319 19027 12325
rect 19242 12316 19248 12328
rect 19300 12316 19306 12368
rect 19334 12316 19340 12368
rect 19392 12356 19398 12368
rect 20070 12356 20076 12368
rect 19392 12328 20076 12356
rect 19392 12316 19398 12328
rect 20070 12316 20076 12328
rect 20128 12316 20134 12368
rect 21174 12365 21180 12368
rect 21168 12356 21180 12365
rect 21135 12328 21180 12356
rect 21168 12319 21180 12328
rect 21174 12316 21180 12319
rect 21232 12316 21238 12368
rect 22833 12359 22891 12365
rect 22833 12325 22845 12359
rect 22879 12356 22891 12359
rect 23477 12359 23535 12365
rect 23477 12356 23489 12359
rect 22879 12328 23489 12356
rect 22879 12325 22891 12328
rect 22833 12319 22891 12325
rect 23477 12325 23489 12328
rect 23523 12325 23535 12359
rect 24946 12356 24952 12368
rect 24907 12328 24952 12356
rect 23477 12319 23535 12325
rect 24946 12316 24952 12328
rect 25004 12316 25010 12368
rect 17402 12248 17408 12300
rect 17460 12288 17466 12300
rect 17497 12291 17555 12297
rect 17497 12288 17509 12291
rect 17460 12260 17509 12288
rect 17460 12248 17466 12260
rect 17497 12257 17509 12260
rect 17543 12257 17555 12291
rect 17497 12251 17555 12257
rect 17586 12248 17592 12300
rect 17644 12288 17650 12300
rect 19426 12288 19432 12300
rect 17644 12260 17689 12288
rect 19387 12260 19432 12288
rect 17644 12248 17650 12260
rect 19426 12248 19432 12260
rect 19484 12248 19490 12300
rect 21726 12288 21732 12300
rect 20916 12260 21732 12288
rect 17678 12220 17684 12232
rect 17639 12192 17684 12220
rect 17678 12180 17684 12192
rect 17736 12180 17742 12232
rect 19521 12223 19579 12229
rect 19521 12220 19533 12223
rect 18616 12192 19533 12220
rect 18616 12096 18644 12192
rect 19521 12189 19533 12192
rect 19567 12189 19579 12223
rect 19521 12183 19579 12189
rect 19610 12180 19616 12232
rect 19668 12220 19674 12232
rect 20916 12229 20944 12260
rect 21726 12248 21732 12260
rect 21784 12248 21790 12300
rect 24670 12288 24676 12300
rect 24631 12260 24676 12288
rect 24670 12248 24676 12260
rect 24728 12248 24734 12300
rect 20073 12223 20131 12229
rect 20073 12220 20085 12223
rect 19668 12192 20085 12220
rect 19668 12180 19674 12192
rect 20073 12189 20085 12192
rect 20119 12189 20131 12223
rect 20901 12223 20959 12229
rect 20901 12220 20913 12223
rect 20073 12183 20131 12189
rect 20456 12192 20913 12220
rect 18598 12084 18604 12096
rect 18559 12056 18604 12084
rect 18598 12044 18604 12056
rect 18656 12044 18662 12096
rect 20162 12044 20168 12096
rect 20220 12084 20226 12096
rect 20456 12093 20484 12192
rect 20901 12189 20913 12192
rect 20947 12189 20959 12223
rect 20901 12183 20959 12189
rect 23569 12223 23627 12229
rect 23569 12189 23581 12223
rect 23615 12189 23627 12223
rect 23569 12183 23627 12189
rect 22557 12155 22615 12161
rect 22557 12152 22569 12155
rect 22112 12124 22569 12152
rect 20441 12087 20499 12093
rect 20441 12084 20453 12087
rect 20220 12056 20453 12084
rect 20220 12044 20226 12056
rect 20441 12053 20453 12056
rect 20487 12053 20499 12087
rect 20441 12047 20499 12053
rect 21266 12044 21272 12096
rect 21324 12084 21330 12096
rect 22112 12084 22140 12124
rect 22557 12121 22569 12124
rect 22603 12152 22615 12155
rect 22833 12155 22891 12161
rect 22833 12152 22845 12155
rect 22603 12124 22845 12152
rect 22603 12121 22615 12124
rect 22557 12115 22615 12121
rect 22833 12121 22845 12124
rect 22879 12121 22891 12155
rect 22833 12115 22891 12121
rect 22278 12084 22284 12096
rect 21324 12056 22140 12084
rect 22239 12056 22284 12084
rect 21324 12044 21330 12056
rect 22278 12044 22284 12056
rect 22336 12044 22342 12096
rect 22922 12084 22928 12096
rect 22883 12056 22928 12084
rect 22922 12044 22928 12056
rect 22980 12084 22986 12096
rect 23584 12084 23612 12183
rect 23658 12180 23664 12232
rect 23716 12220 23722 12232
rect 23716 12192 23761 12220
rect 23716 12180 23722 12192
rect 24210 12084 24216 12096
rect 22980 12056 23612 12084
rect 24171 12056 24216 12084
rect 22980 12044 22986 12056
rect 24210 12044 24216 12056
rect 24268 12044 24274 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 16850 11880 16856 11892
rect 16763 11852 16856 11880
rect 16850 11840 16856 11852
rect 16908 11880 16914 11892
rect 17586 11880 17592 11892
rect 16908 11852 17592 11880
rect 16908 11840 16914 11852
rect 17586 11840 17592 11852
rect 17644 11840 17650 11892
rect 17678 11840 17684 11892
rect 17736 11880 17742 11892
rect 17773 11883 17831 11889
rect 17773 11880 17785 11883
rect 17736 11852 17785 11880
rect 17736 11840 17742 11852
rect 17773 11849 17785 11852
rect 17819 11880 17831 11883
rect 17954 11880 17960 11892
rect 17819 11852 17960 11880
rect 17819 11849 17831 11852
rect 17773 11843 17831 11849
rect 17954 11840 17960 11852
rect 18012 11840 18018 11892
rect 20901 11883 20959 11889
rect 20901 11849 20913 11883
rect 20947 11880 20959 11883
rect 21174 11880 21180 11892
rect 20947 11852 21180 11880
rect 20947 11849 20959 11852
rect 20901 11843 20959 11849
rect 21174 11840 21180 11852
rect 21232 11840 21238 11892
rect 21358 11840 21364 11892
rect 21416 11880 21422 11892
rect 21821 11883 21879 11889
rect 21821 11880 21833 11883
rect 21416 11852 21833 11880
rect 21416 11840 21422 11852
rect 21821 11849 21833 11852
rect 21867 11880 21879 11883
rect 22370 11880 22376 11892
rect 21867 11852 22376 11880
rect 21867 11849 21879 11852
rect 21821 11843 21879 11849
rect 22370 11840 22376 11852
rect 22428 11840 22434 11892
rect 24670 11840 24676 11892
rect 24728 11880 24734 11892
rect 25317 11883 25375 11889
rect 25317 11880 25329 11883
rect 24728 11852 25329 11880
rect 24728 11840 24734 11852
rect 25317 11849 25329 11852
rect 25363 11849 25375 11883
rect 25317 11843 25375 11849
rect 16945 11747 17003 11753
rect 16945 11713 16957 11747
rect 16991 11744 17003 11747
rect 19061 11747 19119 11753
rect 19061 11744 19073 11747
rect 16991 11716 19073 11744
rect 16991 11713 17003 11716
rect 16945 11707 17003 11713
rect 19061 11713 19073 11716
rect 19107 11744 19119 11747
rect 19426 11744 19432 11756
rect 19107 11716 19432 11744
rect 19107 11713 19119 11716
rect 19061 11707 19119 11713
rect 19426 11704 19432 11716
rect 19484 11704 19490 11756
rect 22646 11744 22652 11756
rect 22559 11716 22652 11744
rect 22646 11704 22652 11716
rect 22704 11744 22710 11756
rect 22704 11716 23152 11744
rect 22704 11704 22710 11716
rect 15197 11679 15255 11685
rect 15197 11645 15209 11679
rect 15243 11645 15255 11679
rect 15197 11639 15255 11645
rect 15212 11540 15240 11639
rect 15654 11636 15660 11688
rect 15712 11676 15718 11688
rect 16114 11676 16120 11688
rect 15712 11648 16120 11676
rect 15712 11636 15718 11648
rect 16114 11636 16120 11648
rect 16172 11636 16178 11688
rect 18322 11636 18328 11688
rect 18380 11676 18386 11688
rect 18874 11676 18880 11688
rect 18380 11648 18880 11676
rect 18380 11636 18386 11648
rect 18874 11636 18880 11648
rect 18932 11676 18938 11688
rect 19521 11679 19579 11685
rect 19521 11676 19533 11679
rect 18932 11648 19533 11676
rect 18932 11636 18938 11648
rect 19521 11645 19533 11648
rect 19567 11676 19579 11679
rect 20162 11676 20168 11688
rect 19567 11648 20168 11676
rect 19567 11645 19579 11648
rect 19521 11639 19579 11645
rect 20162 11636 20168 11648
rect 20220 11636 20226 11688
rect 15470 11608 15476 11620
rect 15431 11580 15476 11608
rect 15470 11568 15476 11580
rect 15528 11568 15534 11620
rect 18509 11611 18567 11617
rect 18509 11577 18521 11611
rect 18555 11608 18567 11611
rect 19334 11608 19340 11620
rect 18555 11580 19340 11608
rect 18555 11577 18567 11580
rect 18509 11571 18567 11577
rect 19334 11568 19340 11580
rect 19392 11568 19398 11620
rect 19610 11608 19616 11620
rect 19523 11580 19616 11608
rect 19610 11568 19616 11580
rect 19668 11608 19674 11620
rect 19766 11611 19824 11617
rect 19766 11608 19778 11611
rect 19668 11580 19778 11608
rect 19668 11568 19674 11580
rect 19766 11577 19778 11580
rect 19812 11608 19824 11611
rect 20254 11608 20260 11620
rect 19812 11580 20260 11608
rect 19812 11577 19824 11580
rect 19766 11571 19824 11577
rect 20254 11568 20260 11580
rect 20312 11568 20318 11620
rect 23124 11617 23152 11716
rect 23661 11679 23719 11685
rect 23661 11645 23673 11679
rect 23707 11676 23719 11679
rect 24210 11676 24216 11688
rect 23707 11648 24216 11676
rect 23707 11645 23719 11648
rect 23661 11639 23719 11645
rect 24210 11636 24216 11648
rect 24268 11636 24274 11688
rect 21545 11611 21603 11617
rect 21545 11577 21557 11611
rect 21591 11608 21603 11611
rect 23109 11611 23167 11617
rect 21591 11580 22508 11608
rect 21591 11577 21603 11580
rect 21545 11571 21603 11577
rect 16022 11540 16028 11552
rect 15212 11512 16028 11540
rect 16022 11500 16028 11512
rect 16080 11500 16086 11552
rect 16114 11500 16120 11552
rect 16172 11540 16178 11552
rect 16301 11543 16359 11549
rect 16301 11540 16313 11543
rect 16172 11512 16313 11540
rect 16172 11500 16178 11512
rect 16301 11509 16313 11512
rect 16347 11509 16359 11543
rect 17402 11540 17408 11552
rect 17363 11512 17408 11540
rect 16301 11503 16359 11509
rect 17402 11500 17408 11512
rect 17460 11500 17466 11552
rect 18417 11543 18475 11549
rect 18417 11509 18429 11543
rect 18463 11540 18475 11543
rect 19628 11540 19656 11568
rect 18463 11512 19656 11540
rect 22005 11543 22063 11549
rect 18463 11509 18475 11512
rect 18417 11503 18475 11509
rect 22005 11509 22017 11543
rect 22051 11540 22063 11543
rect 22186 11540 22192 11552
rect 22051 11512 22192 11540
rect 22051 11509 22063 11512
rect 22005 11503 22063 11509
rect 22186 11500 22192 11512
rect 22244 11500 22250 11552
rect 22370 11540 22376 11552
rect 22331 11512 22376 11540
rect 22370 11500 22376 11512
rect 22428 11500 22434 11552
rect 22480 11549 22508 11580
rect 23109 11577 23121 11611
rect 23155 11608 23167 11611
rect 23477 11611 23535 11617
rect 23477 11608 23489 11611
rect 23155 11580 23489 11608
rect 23155 11577 23167 11580
rect 23109 11571 23167 11577
rect 23477 11577 23489 11580
rect 23523 11608 23535 11611
rect 23906 11611 23964 11617
rect 23906 11608 23918 11611
rect 23523 11580 23918 11608
rect 23523 11577 23535 11580
rect 23477 11571 23535 11577
rect 23906 11577 23918 11580
rect 23952 11577 23964 11611
rect 23906 11571 23964 11577
rect 22465 11543 22523 11549
rect 22465 11509 22477 11543
rect 22511 11540 22523 11543
rect 23382 11540 23388 11552
rect 22511 11512 23388 11540
rect 22511 11509 22523 11512
rect 22465 11503 22523 11509
rect 23382 11500 23388 11512
rect 23440 11500 23446 11552
rect 24762 11500 24768 11552
rect 24820 11540 24826 11552
rect 25041 11543 25099 11549
rect 25041 11540 25053 11543
rect 24820 11512 25053 11540
rect 24820 11500 24826 11512
rect 25041 11509 25053 11512
rect 25087 11509 25099 11543
rect 25041 11503 25099 11509
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 15286 11336 15292 11348
rect 15247 11308 15292 11336
rect 15286 11296 15292 11308
rect 15344 11296 15350 11348
rect 20254 11336 20260 11348
rect 20215 11308 20260 11336
rect 20254 11296 20260 11308
rect 20312 11296 20318 11348
rect 20530 11336 20536 11348
rect 20491 11308 20536 11336
rect 20530 11296 20536 11308
rect 20588 11296 20594 11348
rect 21174 11336 21180 11348
rect 21135 11308 21180 11336
rect 21174 11296 21180 11308
rect 21232 11296 21238 11348
rect 22646 11336 22652 11348
rect 22607 11308 22652 11336
rect 22646 11296 22652 11308
rect 22704 11296 22710 11348
rect 23201 11339 23259 11345
rect 23201 11305 23213 11339
rect 23247 11336 23259 11339
rect 23658 11336 23664 11348
rect 23247 11308 23664 11336
rect 23247 11305 23259 11308
rect 23201 11299 23259 11305
rect 23658 11296 23664 11308
rect 23716 11296 23722 11348
rect 24210 11268 24216 11280
rect 23492 11240 24216 11268
rect 23492 11212 23520 11240
rect 24210 11228 24216 11240
rect 24268 11228 24274 11280
rect 15378 11160 15384 11212
rect 15436 11200 15442 11212
rect 15657 11203 15715 11209
rect 15657 11200 15669 11203
rect 15436 11172 15669 11200
rect 15436 11160 15442 11172
rect 15657 11169 15669 11172
rect 15703 11169 15715 11203
rect 17034 11200 17040 11212
rect 16995 11172 17040 11200
rect 15657 11163 15715 11169
rect 17034 11160 17040 11172
rect 17092 11160 17098 11212
rect 18874 11200 18880 11212
rect 18835 11172 18880 11200
rect 18874 11160 18880 11172
rect 18932 11160 18938 11212
rect 19150 11209 19156 11212
rect 19144 11163 19156 11209
rect 19208 11200 19214 11212
rect 19208 11172 19244 11200
rect 19150 11160 19156 11163
rect 19208 11160 19214 11172
rect 21358 11160 21364 11212
rect 21416 11200 21422 11212
rect 21525 11203 21583 11209
rect 21525 11200 21537 11203
rect 21416 11172 21537 11200
rect 21416 11160 21422 11172
rect 21525 11169 21537 11172
rect 21571 11200 21583 11203
rect 22278 11200 22284 11212
rect 21571 11172 22284 11200
rect 21571 11169 21583 11172
rect 21525 11163 21583 11169
rect 22278 11160 22284 11172
rect 22336 11160 22342 11212
rect 23474 11200 23480 11212
rect 23387 11172 23480 11200
rect 23474 11160 23480 11172
rect 23532 11160 23538 11212
rect 23566 11160 23572 11212
rect 23624 11200 23630 11212
rect 23744 11203 23802 11209
rect 23744 11200 23756 11203
rect 23624 11172 23756 11200
rect 23624 11160 23630 11172
rect 23744 11169 23756 11172
rect 23790 11200 23802 11203
rect 24762 11200 24768 11212
rect 23790 11172 24768 11200
rect 23790 11169 23802 11172
rect 23744 11163 23802 11169
rect 24762 11160 24768 11172
rect 24820 11160 24826 11212
rect 13722 11092 13728 11144
rect 13780 11132 13786 11144
rect 14185 11135 14243 11141
rect 14185 11132 14197 11135
rect 13780 11104 14197 11132
rect 13780 11092 13786 11104
rect 14185 11101 14197 11104
rect 14231 11101 14243 11135
rect 14185 11095 14243 11101
rect 15286 11092 15292 11144
rect 15344 11132 15350 11144
rect 15749 11135 15807 11141
rect 15749 11132 15761 11135
rect 15344 11104 15761 11132
rect 15344 11092 15350 11104
rect 15749 11101 15761 11104
rect 15795 11101 15807 11135
rect 15749 11095 15807 11101
rect 15838 11092 15844 11144
rect 15896 11132 15902 11144
rect 15896 11104 15941 11132
rect 15896 11092 15902 11104
rect 20162 11092 20168 11144
rect 20220 11132 20226 11144
rect 21269 11135 21327 11141
rect 21269 11132 21281 11135
rect 20220 11104 21281 11132
rect 20220 11092 20226 11104
rect 21269 11101 21281 11104
rect 21315 11101 21327 11135
rect 21269 11095 21327 11101
rect 14734 11024 14740 11076
rect 14792 11064 14798 11076
rect 14829 11067 14887 11073
rect 14829 11064 14841 11067
rect 14792 11036 14841 11064
rect 14792 11024 14798 11036
rect 14829 11033 14841 11036
rect 14875 11033 14887 11067
rect 14829 11027 14887 11033
rect 22370 11024 22376 11076
rect 22428 11064 22434 11076
rect 22428 11036 23428 11064
rect 22428 11024 22434 11036
rect 16577 10999 16635 11005
rect 16577 10965 16589 10999
rect 16623 10996 16635 10999
rect 16666 10996 16672 11008
rect 16623 10968 16672 10996
rect 16623 10965 16635 10968
rect 16577 10959 16635 10965
rect 16666 10956 16672 10968
rect 16724 10956 16730 11008
rect 16945 10999 17003 11005
rect 16945 10965 16957 10999
rect 16991 10996 17003 10999
rect 17126 10996 17132 11008
rect 16991 10968 17132 10996
rect 16991 10965 17003 10968
rect 16945 10959 17003 10965
rect 17126 10956 17132 10968
rect 17184 10956 17190 11008
rect 18046 10956 18052 11008
rect 18104 10996 18110 11008
rect 18325 10999 18383 11005
rect 18325 10996 18337 10999
rect 18104 10968 18337 10996
rect 18104 10956 18110 10968
rect 18325 10965 18337 10968
rect 18371 10965 18383 10999
rect 23400 10996 23428 11036
rect 24210 10996 24216 11008
rect 23400 10968 24216 10996
rect 18325 10959 18383 10965
rect 24210 10956 24216 10968
rect 24268 10956 24274 11008
rect 24854 10996 24860 11008
rect 24815 10968 24860 10996
rect 24854 10956 24860 10968
rect 24912 10956 24918 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 15933 10795 15991 10801
rect 15933 10761 15945 10795
rect 15979 10792 15991 10795
rect 16206 10792 16212 10804
rect 15979 10764 16212 10792
rect 15979 10761 15991 10764
rect 15933 10755 15991 10761
rect 16206 10752 16212 10764
rect 16264 10752 16270 10804
rect 16666 10752 16672 10804
rect 16724 10752 16730 10804
rect 16850 10792 16856 10804
rect 16811 10764 16856 10792
rect 16850 10752 16856 10764
rect 16908 10752 16914 10804
rect 19150 10752 19156 10804
rect 19208 10792 19214 10804
rect 19429 10795 19487 10801
rect 19429 10792 19441 10795
rect 19208 10764 19441 10792
rect 19208 10752 19214 10764
rect 19429 10761 19441 10764
rect 19475 10761 19487 10795
rect 19429 10755 19487 10761
rect 19797 10795 19855 10801
rect 19797 10761 19809 10795
rect 19843 10792 19855 10795
rect 21269 10795 21327 10801
rect 21269 10792 21281 10795
rect 19843 10764 21281 10792
rect 19843 10761 19855 10764
rect 19797 10755 19855 10761
rect 14369 10727 14427 10733
rect 14369 10693 14381 10727
rect 14415 10724 14427 10727
rect 15286 10724 15292 10736
rect 14415 10696 15292 10724
rect 14415 10693 14427 10696
rect 14369 10687 14427 10693
rect 15286 10684 15292 10696
rect 15344 10684 15350 10736
rect 16025 10727 16083 10733
rect 16025 10693 16037 10727
rect 16071 10724 16083 10727
rect 16390 10724 16396 10736
rect 16071 10696 16396 10724
rect 16071 10693 16083 10696
rect 16025 10687 16083 10693
rect 16390 10684 16396 10696
rect 16448 10684 16454 10736
rect 16684 10724 16712 10752
rect 16684 10696 17540 10724
rect 14918 10656 14924 10668
rect 14879 10628 14924 10656
rect 14918 10616 14924 10628
rect 14976 10616 14982 10668
rect 16669 10659 16727 10665
rect 16669 10625 16681 10659
rect 16715 10656 16727 10659
rect 17402 10656 17408 10668
rect 16715 10628 17264 10656
rect 17363 10628 17408 10656
rect 16715 10625 16727 10628
rect 16669 10619 16727 10625
rect 12989 10591 13047 10597
rect 12989 10557 13001 10591
rect 13035 10588 13047 10591
rect 13078 10588 13084 10600
rect 13035 10560 13084 10588
rect 13035 10557 13047 10560
rect 12989 10551 13047 10557
rect 13078 10548 13084 10560
rect 13136 10548 13142 10600
rect 16206 10548 16212 10600
rect 16264 10588 16270 10600
rect 16393 10591 16451 10597
rect 16393 10588 16405 10591
rect 16264 10560 16405 10588
rect 16264 10548 16270 10560
rect 16393 10557 16405 10560
rect 16439 10557 16451 10591
rect 16393 10551 16451 10557
rect 12618 10480 12624 10532
rect 12676 10520 12682 10532
rect 13357 10523 13415 10529
rect 13357 10520 13369 10523
rect 12676 10492 13369 10520
rect 12676 10480 12682 10492
rect 13357 10489 13369 10492
rect 13403 10489 13415 10523
rect 14829 10523 14887 10529
rect 14829 10520 14841 10523
rect 13357 10483 13415 10489
rect 13832 10492 14841 10520
rect 13832 10464 13860 10492
rect 14829 10489 14841 10492
rect 14875 10489 14887 10523
rect 17236 10520 17264 10628
rect 17402 10616 17408 10628
rect 17460 10616 17466 10668
rect 17313 10591 17371 10597
rect 17313 10557 17325 10591
rect 17359 10588 17371 10591
rect 17512 10588 17540 10696
rect 19334 10684 19340 10736
rect 19392 10724 19398 10736
rect 20073 10727 20131 10733
rect 20073 10724 20085 10727
rect 19392 10696 20085 10724
rect 19392 10684 19398 10696
rect 20073 10693 20085 10696
rect 20119 10693 20131 10727
rect 20073 10687 20131 10693
rect 17359 10560 17540 10588
rect 17359 10557 17371 10560
rect 17313 10551 17371 10557
rect 17586 10548 17592 10600
rect 17644 10588 17650 10600
rect 18049 10591 18107 10597
rect 18049 10588 18061 10591
rect 17644 10560 18061 10588
rect 17644 10548 17650 10560
rect 18049 10557 18061 10560
rect 18095 10588 18107 10591
rect 18874 10588 18880 10600
rect 18095 10560 18880 10588
rect 18095 10557 18107 10560
rect 18049 10551 18107 10557
rect 18874 10548 18880 10560
rect 18932 10548 18938 10600
rect 18316 10523 18374 10529
rect 18316 10520 18328 10523
rect 17236 10492 18328 10520
rect 14829 10483 14887 10489
rect 18316 10489 18328 10492
rect 18362 10520 18374 10523
rect 18690 10520 18696 10532
rect 18362 10492 18696 10520
rect 18362 10489 18374 10492
rect 18316 10483 18374 10489
rect 18690 10480 18696 10492
rect 18748 10480 18754 10532
rect 20088 10520 20116 10687
rect 20530 10616 20536 10668
rect 20588 10656 20594 10668
rect 20824 10665 20852 10764
rect 21269 10761 21281 10764
rect 21315 10792 21327 10795
rect 21358 10792 21364 10804
rect 21315 10764 21364 10792
rect 21315 10761 21327 10764
rect 21269 10755 21327 10761
rect 21358 10752 21364 10764
rect 21416 10752 21422 10804
rect 21913 10795 21971 10801
rect 21913 10761 21925 10795
rect 21959 10792 21971 10795
rect 22094 10792 22100 10804
rect 21959 10764 22100 10792
rect 21959 10761 21971 10764
rect 21913 10755 21971 10761
rect 22094 10752 22100 10764
rect 22152 10752 22158 10804
rect 24762 10792 24768 10804
rect 24723 10764 24768 10792
rect 24762 10752 24768 10764
rect 24820 10752 24826 10804
rect 25406 10792 25412 10804
rect 25367 10764 25412 10792
rect 25406 10752 25412 10764
rect 25464 10752 25470 10804
rect 20898 10684 20904 10736
rect 20956 10724 20962 10736
rect 22005 10727 22063 10733
rect 22005 10724 22017 10727
rect 20956 10696 22017 10724
rect 20956 10684 20962 10696
rect 22005 10693 22017 10696
rect 22051 10693 22063 10727
rect 23566 10724 23572 10736
rect 22005 10687 22063 10693
rect 22664 10696 23572 10724
rect 20717 10659 20775 10665
rect 20717 10656 20729 10659
rect 20588 10628 20729 10656
rect 20588 10616 20594 10628
rect 20717 10625 20729 10628
rect 20763 10625 20775 10659
rect 20717 10619 20775 10625
rect 20809 10659 20867 10665
rect 20809 10625 20821 10659
rect 20855 10625 20867 10659
rect 20809 10619 20867 10625
rect 22186 10616 22192 10668
rect 22244 10656 22250 10668
rect 22465 10659 22523 10665
rect 22465 10656 22477 10659
rect 22244 10628 22477 10656
rect 22244 10616 22250 10628
rect 22465 10625 22477 10628
rect 22511 10625 22523 10659
rect 22465 10619 22523 10625
rect 22554 10616 22560 10668
rect 22612 10656 22618 10668
rect 22664 10665 22692 10696
rect 23566 10684 23572 10696
rect 23624 10684 23630 10736
rect 22649 10659 22707 10665
rect 22649 10656 22661 10659
rect 22612 10628 22661 10656
rect 22612 10616 22618 10628
rect 22649 10625 22661 10628
rect 22695 10625 22707 10659
rect 22649 10619 22707 10625
rect 23474 10616 23480 10668
rect 23532 10656 23538 10668
rect 24213 10659 24271 10665
rect 24213 10656 24225 10659
rect 23532 10628 24225 10656
rect 23532 10616 23538 10628
rect 24213 10625 24225 10628
rect 24259 10656 24271 10659
rect 24854 10656 24860 10668
rect 24259 10628 24860 10656
rect 24259 10625 24271 10628
rect 24213 10619 24271 10625
rect 24854 10616 24860 10628
rect 24912 10656 24918 10668
rect 25041 10659 25099 10665
rect 25041 10656 25053 10659
rect 24912 10628 25053 10656
rect 24912 10616 24918 10628
rect 25041 10625 25053 10628
rect 25087 10625 25099 10659
rect 25041 10619 25099 10625
rect 22094 10548 22100 10600
rect 22152 10588 22158 10600
rect 22373 10591 22431 10597
rect 22373 10588 22385 10591
rect 22152 10560 22385 10588
rect 22152 10548 22158 10560
rect 22373 10557 22385 10560
rect 22419 10557 22431 10591
rect 22373 10551 22431 10557
rect 23109 10591 23167 10597
rect 23109 10557 23121 10591
rect 23155 10588 23167 10591
rect 24118 10588 24124 10600
rect 23155 10560 24124 10588
rect 23155 10557 23167 10560
rect 23109 10551 23167 10557
rect 24118 10548 24124 10560
rect 24176 10548 24182 10600
rect 25222 10588 25228 10600
rect 25183 10560 25228 10588
rect 25222 10548 25228 10560
rect 25280 10588 25286 10600
rect 25777 10591 25835 10597
rect 25777 10588 25789 10591
rect 25280 10560 25789 10588
rect 25280 10548 25286 10560
rect 25777 10557 25789 10560
rect 25823 10557 25835 10591
rect 25777 10551 25835 10557
rect 20625 10523 20683 10529
rect 20625 10520 20637 10523
rect 20088 10492 20637 10520
rect 20625 10489 20637 10492
rect 20671 10489 20683 10523
rect 20625 10483 20683 10489
rect 23477 10523 23535 10529
rect 23477 10489 23489 10523
rect 23523 10520 23535 10523
rect 23523 10492 24072 10520
rect 23523 10489 23535 10492
rect 23477 10483 23535 10489
rect 13814 10452 13820 10464
rect 13775 10424 13820 10452
rect 13814 10412 13820 10424
rect 13872 10412 13878 10464
rect 14274 10452 14280 10464
rect 14235 10424 14280 10452
rect 14274 10412 14280 10424
rect 14332 10452 14338 10464
rect 14737 10455 14795 10461
rect 14737 10452 14749 10455
rect 14332 10424 14749 10452
rect 14332 10412 14338 10424
rect 14737 10421 14749 10424
rect 14783 10421 14795 10455
rect 15378 10452 15384 10464
rect 15339 10424 15384 10452
rect 14737 10415 14795 10421
rect 15378 10412 15384 10424
rect 15436 10412 15442 10464
rect 16114 10412 16120 10464
rect 16172 10452 16178 10464
rect 16485 10455 16543 10461
rect 16485 10452 16497 10455
rect 16172 10424 16497 10452
rect 16172 10412 16178 10424
rect 16485 10421 16497 10424
rect 16531 10421 16543 10455
rect 16485 10415 16543 10421
rect 17126 10412 17132 10464
rect 17184 10452 17190 10464
rect 17221 10455 17279 10461
rect 17221 10452 17233 10455
rect 17184 10424 17233 10452
rect 17184 10412 17190 10424
rect 17221 10421 17233 10424
rect 17267 10421 17279 10455
rect 20254 10452 20260 10464
rect 20215 10424 20260 10452
rect 17221 10415 17279 10421
rect 20254 10412 20260 10424
rect 20312 10412 20318 10464
rect 23661 10455 23719 10461
rect 23661 10421 23673 10455
rect 23707 10452 23719 10455
rect 23934 10452 23940 10464
rect 23707 10424 23940 10452
rect 23707 10421 23719 10424
rect 23661 10415 23719 10421
rect 23934 10412 23940 10424
rect 23992 10412 23998 10464
rect 24044 10461 24072 10492
rect 24029 10455 24087 10461
rect 24029 10421 24041 10455
rect 24075 10452 24087 10455
rect 24118 10452 24124 10464
rect 24075 10424 24124 10452
rect 24075 10421 24087 10424
rect 24029 10415 24087 10421
rect 24118 10412 24124 10424
rect 24176 10412 24182 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 12894 10248 12900 10260
rect 12855 10220 12900 10248
rect 12894 10208 12900 10220
rect 12952 10208 12958 10260
rect 14737 10251 14795 10257
rect 14737 10217 14749 10251
rect 14783 10248 14795 10251
rect 14918 10248 14924 10260
rect 14783 10220 14924 10248
rect 14783 10217 14795 10220
rect 14737 10211 14795 10217
rect 14918 10208 14924 10220
rect 14976 10208 14982 10260
rect 15105 10251 15163 10257
rect 15105 10217 15117 10251
rect 15151 10248 15163 10251
rect 15286 10248 15292 10260
rect 15151 10220 15292 10248
rect 15151 10217 15163 10220
rect 15105 10211 15163 10217
rect 15286 10208 15292 10220
rect 15344 10208 15350 10260
rect 15565 10251 15623 10257
rect 15565 10217 15577 10251
rect 15611 10248 15623 10251
rect 15838 10248 15844 10260
rect 15611 10220 15844 10248
rect 15611 10217 15623 10220
rect 15565 10211 15623 10217
rect 15838 10208 15844 10220
rect 15896 10208 15902 10260
rect 17034 10208 17040 10260
rect 17092 10248 17098 10260
rect 17773 10251 17831 10257
rect 17773 10248 17785 10251
rect 17092 10220 17785 10248
rect 17092 10208 17098 10220
rect 17773 10217 17785 10220
rect 17819 10217 17831 10251
rect 17773 10211 17831 10217
rect 17954 10208 17960 10260
rect 18012 10248 18018 10260
rect 18141 10251 18199 10257
rect 18141 10248 18153 10251
rect 18012 10220 18153 10248
rect 18012 10208 18018 10220
rect 18141 10217 18153 10220
rect 18187 10217 18199 10251
rect 18141 10211 18199 10217
rect 18325 10251 18383 10257
rect 18325 10217 18337 10251
rect 18371 10217 18383 10251
rect 18598 10248 18604 10260
rect 18559 10220 18604 10248
rect 18325 10211 18383 10217
rect 13817 10183 13875 10189
rect 13817 10149 13829 10183
rect 13863 10180 13875 10183
rect 17586 10180 17592 10192
rect 13863 10152 17592 10180
rect 13863 10149 13875 10152
rect 13817 10143 13875 10149
rect 13906 10112 13912 10124
rect 13867 10084 13912 10112
rect 13906 10072 13912 10084
rect 13964 10072 13970 10124
rect 14182 10112 14188 10124
rect 14143 10084 14188 10112
rect 14182 10072 14188 10084
rect 14240 10072 14246 10124
rect 16132 10121 16160 10152
rect 17586 10140 17592 10152
rect 17644 10140 17650 10192
rect 18340 10180 18368 10211
rect 18598 10208 18604 10220
rect 18656 10208 18662 10260
rect 18690 10208 18696 10260
rect 18748 10248 18754 10260
rect 19613 10251 19671 10257
rect 19613 10248 19625 10251
rect 18748 10220 19625 10248
rect 18748 10208 18754 10220
rect 19613 10217 19625 10220
rect 19659 10217 19671 10251
rect 20162 10248 20168 10260
rect 20123 10220 20168 10248
rect 19613 10211 19671 10217
rect 20162 10208 20168 10220
rect 20220 10208 20226 10260
rect 21266 10248 21272 10260
rect 21227 10220 21272 10248
rect 21266 10208 21272 10220
rect 21324 10208 21330 10260
rect 21634 10248 21640 10260
rect 21595 10220 21640 10248
rect 21634 10208 21640 10220
rect 21692 10208 21698 10260
rect 22186 10208 22192 10260
rect 22244 10248 22250 10260
rect 22649 10251 22707 10257
rect 22649 10248 22661 10251
rect 22244 10220 22661 10248
rect 22244 10208 22250 10220
rect 22649 10217 22661 10220
rect 22695 10217 22707 10251
rect 22649 10211 22707 10217
rect 20254 10180 20260 10192
rect 18340 10152 20260 10180
rect 20254 10140 20260 10152
rect 20312 10180 20318 10192
rect 21729 10183 21787 10189
rect 20312 10152 20392 10180
rect 20312 10140 20318 10152
rect 16390 10121 16396 10124
rect 16117 10115 16175 10121
rect 16117 10081 16129 10115
rect 16163 10081 16175 10115
rect 16384 10112 16396 10121
rect 16351 10084 16396 10112
rect 16117 10075 16175 10081
rect 16384 10075 16396 10084
rect 16390 10072 16396 10075
rect 16448 10072 16454 10124
rect 18046 10072 18052 10124
rect 18104 10112 18110 10124
rect 18509 10115 18567 10121
rect 18509 10112 18521 10115
rect 18104 10084 18521 10112
rect 18104 10072 18110 10084
rect 18509 10081 18521 10084
rect 18555 10081 18567 10115
rect 18509 10075 18567 10081
rect 18598 10072 18604 10124
rect 18656 10112 18662 10124
rect 18969 10115 19027 10121
rect 18969 10112 18981 10115
rect 18656 10084 18981 10112
rect 18656 10072 18662 10084
rect 18969 10081 18981 10084
rect 19015 10081 19027 10115
rect 18969 10075 19027 10081
rect 19058 10072 19064 10124
rect 19116 10112 19122 10124
rect 20364 10121 20392 10152
rect 21729 10149 21741 10183
rect 21775 10180 21787 10183
rect 21910 10180 21916 10192
rect 21775 10152 21916 10180
rect 21775 10149 21787 10152
rect 21729 10143 21787 10149
rect 21910 10140 21916 10152
rect 21968 10140 21974 10192
rect 22373 10183 22431 10189
rect 22373 10149 22385 10183
rect 22419 10180 22431 10183
rect 22554 10180 22560 10192
rect 22419 10152 22560 10180
rect 22419 10149 22431 10152
rect 22373 10143 22431 10149
rect 22554 10140 22560 10152
rect 22612 10140 22618 10192
rect 23474 10140 23480 10192
rect 23532 10189 23538 10192
rect 23532 10183 23596 10189
rect 23532 10149 23550 10183
rect 23584 10149 23596 10183
rect 23532 10143 23596 10149
rect 23532 10140 23538 10143
rect 20349 10115 20407 10121
rect 19116 10084 19161 10112
rect 19116 10072 19122 10084
rect 20349 10081 20361 10115
rect 20395 10081 20407 10115
rect 20349 10075 20407 10081
rect 23109 10115 23167 10121
rect 23109 10081 23121 10115
rect 23155 10112 23167 10115
rect 23290 10112 23296 10124
rect 23155 10084 23296 10112
rect 23155 10081 23167 10084
rect 23109 10075 23167 10081
rect 23290 10072 23296 10084
rect 23348 10072 23354 10124
rect 19150 10004 19156 10056
rect 19208 10044 19214 10056
rect 19702 10044 19708 10056
rect 19208 10016 19708 10044
rect 19208 10004 19214 10016
rect 19702 10004 19708 10016
rect 19760 10044 19766 10056
rect 19981 10047 20039 10053
rect 19981 10044 19993 10047
rect 19760 10016 19993 10044
rect 19760 10004 19766 10016
rect 19981 10013 19993 10016
rect 20027 10013 20039 10047
rect 19981 10007 20039 10013
rect 21913 10047 21971 10053
rect 21913 10013 21925 10047
rect 21959 10044 21971 10047
rect 22002 10044 22008 10056
rect 21959 10016 22008 10044
rect 21959 10013 21971 10016
rect 21913 10007 21971 10013
rect 17497 9979 17555 9985
rect 17497 9945 17509 9979
rect 17543 9976 17555 9979
rect 18690 9976 18696 9988
rect 17543 9948 18696 9976
rect 17543 9945 17555 9948
rect 17497 9939 17555 9945
rect 16025 9911 16083 9917
rect 16025 9877 16037 9911
rect 16071 9908 16083 9911
rect 17512 9908 17540 9939
rect 18690 9936 18696 9948
rect 18748 9936 18754 9988
rect 21177 9979 21235 9985
rect 21177 9945 21189 9979
rect 21223 9976 21235 9979
rect 21928 9976 21956 10007
rect 22002 10004 22008 10016
rect 22060 10004 22066 10056
rect 21223 9948 21956 9976
rect 21223 9945 21235 9948
rect 21177 9939 21235 9945
rect 16071 9880 17540 9908
rect 16071 9877 16083 9880
rect 16025 9871 16083 9877
rect 19150 9868 19156 9920
rect 19208 9908 19214 9920
rect 20717 9911 20775 9917
rect 20717 9908 20729 9911
rect 19208 9880 20729 9908
rect 19208 9868 19214 9880
rect 20717 9877 20729 9880
rect 20763 9877 20775 9911
rect 20717 9871 20775 9877
rect 24210 9868 24216 9920
rect 24268 9908 24274 9920
rect 24673 9911 24731 9917
rect 24673 9908 24685 9911
rect 24268 9880 24685 9908
rect 24268 9868 24274 9880
rect 24673 9877 24685 9880
rect 24719 9877 24731 9911
rect 24946 9908 24952 9920
rect 24907 9880 24952 9908
rect 24673 9871 24731 9877
rect 24946 9868 24952 9880
rect 25004 9868 25010 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 13906 9664 13912 9716
rect 13964 9704 13970 9716
rect 14277 9707 14335 9713
rect 14277 9704 14289 9707
rect 13964 9676 14289 9704
rect 13964 9664 13970 9676
rect 14277 9673 14289 9676
rect 14323 9673 14335 9707
rect 16942 9704 16948 9716
rect 16855 9676 16948 9704
rect 14277 9667 14335 9673
rect 16942 9664 16948 9676
rect 17000 9704 17006 9716
rect 17402 9704 17408 9716
rect 17000 9676 17408 9704
rect 17000 9664 17006 9676
rect 17402 9664 17408 9676
rect 17460 9664 17466 9716
rect 19242 9704 19248 9716
rect 18064 9676 19248 9704
rect 13265 9639 13323 9645
rect 13265 9605 13277 9639
rect 13311 9636 13323 9639
rect 13924 9636 13952 9664
rect 18064 9648 18092 9676
rect 19242 9664 19248 9676
rect 19300 9664 19306 9716
rect 19702 9704 19708 9716
rect 19663 9676 19708 9704
rect 19702 9664 19708 9676
rect 19760 9664 19766 9716
rect 13311 9608 13952 9636
rect 13311 9605 13323 9608
rect 13265 9599 13323 9605
rect 14734 9596 14740 9648
rect 14792 9636 14798 9648
rect 18046 9636 18052 9648
rect 14792 9608 14872 9636
rect 14792 9596 14798 9608
rect 13354 9528 13360 9580
rect 13412 9568 13418 9580
rect 13909 9571 13967 9577
rect 13909 9568 13921 9571
rect 13412 9540 13921 9568
rect 13412 9528 13418 9540
rect 13909 9537 13921 9540
rect 13955 9568 13967 9571
rect 13955 9540 14780 9568
rect 13955 9537 13967 9540
rect 13909 9531 13967 9537
rect 13173 9503 13231 9509
rect 13173 9469 13185 9503
rect 13219 9500 13231 9503
rect 13633 9503 13691 9509
rect 13633 9500 13645 9503
rect 13219 9472 13645 9500
rect 13219 9469 13231 9472
rect 13173 9463 13231 9469
rect 13633 9469 13645 9472
rect 13679 9500 13691 9503
rect 13722 9500 13728 9512
rect 13679 9472 13728 9500
rect 13679 9469 13691 9472
rect 13633 9463 13691 9469
rect 13722 9460 13728 9472
rect 13780 9460 13786 9512
rect 14752 9444 14780 9540
rect 14844 9509 14872 9608
rect 17236 9608 18052 9636
rect 17236 9512 17264 9608
rect 18046 9596 18052 9608
rect 18104 9596 18110 9648
rect 19429 9639 19487 9645
rect 19429 9605 19441 9639
rect 19475 9636 19487 9639
rect 19518 9636 19524 9648
rect 19475 9608 19524 9636
rect 19475 9605 19487 9608
rect 19429 9599 19487 9605
rect 19518 9596 19524 9608
rect 19576 9596 19582 9648
rect 20070 9636 20076 9648
rect 20031 9608 20076 9636
rect 20070 9596 20076 9608
rect 20128 9596 20134 9648
rect 23106 9636 23112 9648
rect 23067 9608 23112 9636
rect 23106 9596 23112 9608
rect 23164 9596 23170 9648
rect 17862 9568 17868 9580
rect 17823 9540 17868 9568
rect 17862 9528 17868 9540
rect 17920 9528 17926 9580
rect 20088 9568 20116 9596
rect 20088 9540 20392 9568
rect 20364 9512 20392 9540
rect 14829 9503 14887 9509
rect 14829 9469 14841 9503
rect 14875 9500 14887 9503
rect 14918 9500 14924 9512
rect 14875 9472 14924 9500
rect 14875 9469 14887 9472
rect 14829 9463 14887 9469
rect 14918 9460 14924 9472
rect 14976 9460 14982 9512
rect 17218 9500 17224 9512
rect 17179 9472 17224 9500
rect 17218 9460 17224 9472
rect 17276 9460 17282 9512
rect 17678 9460 17684 9512
rect 17736 9500 17742 9512
rect 18049 9503 18107 9509
rect 18049 9500 18061 9503
rect 17736 9472 18061 9500
rect 17736 9460 17742 9472
rect 18049 9469 18061 9472
rect 18095 9500 18107 9503
rect 19150 9500 19156 9512
rect 18095 9472 19156 9500
rect 18095 9469 18107 9472
rect 18049 9463 18107 9469
rect 19150 9460 19156 9472
rect 19208 9460 19214 9512
rect 20162 9460 20168 9512
rect 20220 9500 20226 9512
rect 20257 9503 20315 9509
rect 20257 9500 20269 9503
rect 20220 9472 20269 9500
rect 20220 9460 20226 9472
rect 20257 9469 20269 9472
rect 20303 9469 20315 9503
rect 20257 9463 20315 9469
rect 20346 9460 20352 9512
rect 20404 9500 20410 9512
rect 20513 9503 20571 9509
rect 20513 9500 20525 9503
rect 20404 9472 20525 9500
rect 20404 9460 20410 9472
rect 20513 9469 20525 9472
rect 20559 9469 20571 9503
rect 20513 9463 20571 9469
rect 21634 9460 21640 9512
rect 21692 9500 21698 9512
rect 22281 9503 22339 9509
rect 22281 9500 22293 9503
rect 21692 9472 22293 9500
rect 21692 9460 21698 9472
rect 22281 9469 22293 9472
rect 22327 9469 22339 9503
rect 22281 9463 22339 9469
rect 22465 9503 22523 9509
rect 22465 9469 22477 9503
rect 22511 9500 22523 9503
rect 23124 9500 23152 9596
rect 23290 9528 23296 9580
rect 23348 9568 23354 9580
rect 23753 9571 23811 9577
rect 23753 9568 23765 9571
rect 23348 9540 23765 9568
rect 23348 9528 23354 9540
rect 23753 9537 23765 9540
rect 23799 9537 23811 9571
rect 23753 9531 23811 9537
rect 22511 9472 23152 9500
rect 23768 9500 23796 9531
rect 24946 9500 24952 9512
rect 23768 9472 24952 9500
rect 22511 9469 22523 9472
rect 22465 9463 22523 9469
rect 24946 9460 24952 9472
rect 25004 9500 25010 9512
rect 25409 9503 25467 9509
rect 25409 9500 25421 9503
rect 25004 9472 25421 9500
rect 25004 9460 25010 9472
rect 25409 9469 25421 9472
rect 25455 9469 25467 9503
rect 25409 9463 25467 9469
rect 14734 9432 14740 9444
rect 14695 9404 14740 9432
rect 14734 9392 14740 9404
rect 14792 9432 14798 9444
rect 15074 9435 15132 9441
rect 15074 9432 15086 9435
rect 14792 9404 15086 9432
rect 14792 9392 14798 9404
rect 15074 9401 15086 9404
rect 15120 9401 15132 9435
rect 15074 9395 15132 9401
rect 17954 9392 17960 9444
rect 18012 9432 18018 9444
rect 18294 9435 18352 9441
rect 18294 9432 18306 9435
rect 18012 9404 18306 9432
rect 18012 9392 18018 9404
rect 18294 9401 18306 9404
rect 18340 9401 18352 9435
rect 18294 9395 18352 9401
rect 23477 9435 23535 9441
rect 23477 9401 23489 9435
rect 23523 9432 23535 9435
rect 24020 9435 24078 9441
rect 24020 9432 24032 9435
rect 23523 9404 24032 9432
rect 23523 9401 23535 9404
rect 23477 9395 23535 9401
rect 24020 9401 24032 9404
rect 24066 9432 24078 9435
rect 24762 9432 24768 9444
rect 24066 9404 24768 9432
rect 24066 9401 24078 9404
rect 24020 9395 24078 9401
rect 24762 9392 24768 9404
rect 24820 9392 24826 9444
rect 12805 9367 12863 9373
rect 12805 9333 12817 9367
rect 12851 9364 12863 9367
rect 12986 9364 12992 9376
rect 12851 9336 12992 9364
rect 12851 9333 12863 9336
rect 12805 9327 12863 9333
rect 12986 9324 12992 9336
rect 13044 9364 13050 9376
rect 13725 9367 13783 9373
rect 13725 9364 13737 9367
rect 13044 9336 13737 9364
rect 13044 9324 13050 9336
rect 13725 9333 13737 9336
rect 13771 9333 13783 9367
rect 13725 9327 13783 9333
rect 16209 9367 16267 9373
rect 16209 9333 16221 9367
rect 16255 9364 16267 9367
rect 16390 9364 16396 9376
rect 16255 9336 16396 9364
rect 16255 9333 16267 9336
rect 16209 9327 16267 9333
rect 16390 9324 16396 9336
rect 16448 9364 16454 9376
rect 16574 9364 16580 9376
rect 16448 9336 16580 9364
rect 16448 9324 16454 9336
rect 16574 9324 16580 9336
rect 16632 9324 16638 9376
rect 17034 9364 17040 9376
rect 16995 9336 17040 9364
rect 17034 9324 17040 9336
rect 17092 9324 17098 9376
rect 21634 9364 21640 9376
rect 21595 9336 21640 9364
rect 21634 9324 21640 9336
rect 21692 9324 21698 9376
rect 21910 9364 21916 9376
rect 21871 9336 21916 9364
rect 21910 9324 21916 9336
rect 21968 9324 21974 9376
rect 22646 9364 22652 9376
rect 22607 9336 22652 9364
rect 22646 9324 22652 9336
rect 22704 9324 22710 9376
rect 23198 9324 23204 9376
rect 23256 9364 23262 9376
rect 23750 9364 23756 9376
rect 23256 9336 23756 9364
rect 23256 9324 23262 9336
rect 23750 9324 23756 9336
rect 23808 9324 23814 9376
rect 25130 9364 25136 9376
rect 25091 9336 25136 9364
rect 25130 9324 25136 9336
rect 25188 9324 25194 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 11974 9160 11980 9172
rect 11935 9132 11980 9160
rect 11974 9120 11980 9132
rect 12032 9120 12038 9172
rect 13354 9160 13360 9172
rect 13315 9132 13360 9160
rect 13354 9120 13360 9132
rect 13412 9120 13418 9172
rect 13538 9160 13544 9172
rect 13499 9132 13544 9160
rect 13538 9120 13544 9132
rect 13596 9120 13602 9172
rect 17954 9120 17960 9172
rect 18012 9160 18018 9172
rect 18049 9163 18107 9169
rect 18049 9160 18061 9163
rect 18012 9132 18061 9160
rect 18012 9120 18018 9132
rect 18049 9129 18061 9132
rect 18095 9129 18107 9163
rect 20254 9160 20260 9172
rect 20215 9132 20260 9160
rect 18049 9123 18107 9129
rect 20254 9120 20260 9132
rect 20312 9120 20318 9172
rect 21174 9160 21180 9172
rect 21135 9132 21180 9160
rect 21174 9120 21180 9132
rect 21232 9120 21238 9172
rect 23293 9163 23351 9169
rect 23293 9129 23305 9163
rect 23339 9160 23351 9163
rect 23382 9160 23388 9172
rect 23339 9132 23388 9160
rect 23339 9129 23351 9132
rect 23293 9123 23351 9129
rect 23382 9120 23388 9132
rect 23440 9120 23446 9172
rect 16942 9101 16948 9104
rect 16936 9092 16948 9101
rect 16903 9064 16948 9092
rect 16936 9055 16948 9064
rect 16942 9052 16948 9055
rect 17000 9052 17006 9104
rect 19337 9095 19395 9101
rect 19337 9061 19349 9095
rect 19383 9092 19395 9095
rect 19426 9092 19432 9104
rect 19383 9064 19432 9092
rect 19383 9061 19395 9064
rect 19337 9055 19395 9061
rect 19426 9052 19432 9064
rect 19484 9052 19490 9104
rect 22462 9052 22468 9104
rect 22520 9092 22526 9104
rect 24670 9092 24676 9104
rect 22520 9064 24676 9092
rect 22520 9052 22526 9064
rect 24670 9052 24676 9064
rect 24728 9052 24734 9104
rect 12342 9024 12348 9036
rect 12303 8996 12348 9024
rect 12342 8984 12348 8996
rect 12400 8984 12406 9036
rect 13446 8984 13452 9036
rect 13504 9024 13510 9036
rect 13909 9027 13967 9033
rect 13909 9024 13921 9027
rect 13504 8996 13921 9024
rect 13504 8984 13510 8996
rect 13909 8993 13921 8996
rect 13955 8993 13967 9027
rect 13909 8987 13967 8993
rect 14001 9027 14059 9033
rect 14001 8993 14013 9027
rect 14047 9024 14059 9027
rect 14550 9024 14556 9036
rect 14047 8996 14556 9024
rect 14047 8993 14059 8996
rect 14001 8987 14059 8993
rect 14550 8984 14556 8996
rect 14608 8984 14614 9036
rect 15470 8984 15476 9036
rect 15528 9024 15534 9036
rect 15565 9027 15623 9033
rect 15565 9024 15577 9027
rect 15528 8996 15577 9024
rect 15528 8984 15534 8996
rect 15565 8993 15577 8996
rect 15611 8993 15623 9027
rect 15565 8987 15623 8993
rect 16669 9027 16727 9033
rect 16669 8993 16681 9027
rect 16715 9024 16727 9027
rect 17678 9024 17684 9036
rect 16715 8996 17684 9024
rect 16715 8993 16727 8996
rect 16669 8987 16727 8993
rect 17678 8984 17684 8996
rect 17736 8984 17742 9036
rect 18966 8984 18972 9036
rect 19024 9024 19030 9036
rect 19245 9027 19303 9033
rect 19245 9024 19257 9027
rect 19024 8996 19257 9024
rect 19024 8984 19030 8996
rect 19245 8993 19257 8996
rect 19291 8993 19303 9027
rect 19245 8987 19303 8993
rect 20717 9027 20775 9033
rect 20717 8993 20729 9027
rect 20763 9024 20775 9027
rect 21266 9024 21272 9036
rect 20763 8996 21272 9024
rect 20763 8993 20775 8996
rect 20717 8987 20775 8993
rect 21266 8984 21272 8996
rect 21324 9024 21330 9036
rect 21545 9027 21603 9033
rect 21545 9024 21557 9027
rect 21324 8996 21557 9024
rect 21324 8984 21330 8996
rect 21545 8993 21557 8996
rect 21591 8993 21603 9027
rect 21545 8987 21603 8993
rect 22281 9027 22339 9033
rect 22281 8993 22293 9027
rect 22327 9024 22339 9027
rect 22925 9027 22983 9033
rect 22925 9024 22937 9027
rect 22327 8996 22937 9024
rect 22327 8993 22339 8996
rect 22281 8987 22339 8993
rect 22925 8993 22937 8996
rect 22971 9024 22983 9027
rect 23290 9024 23296 9036
rect 22971 8996 23296 9024
rect 22971 8993 22983 8996
rect 22925 8987 22983 8993
rect 23290 8984 23296 8996
rect 23348 8984 23354 9036
rect 23652 9027 23710 9033
rect 23652 8993 23664 9027
rect 23698 9024 23710 9027
rect 24210 9024 24216 9036
rect 23698 8996 24216 9024
rect 23698 8993 23710 8996
rect 23652 8987 23710 8993
rect 24210 8984 24216 8996
rect 24268 8984 24274 9036
rect 11238 8916 11244 8968
rect 11296 8956 11302 8968
rect 12437 8959 12495 8965
rect 12437 8956 12449 8959
rect 11296 8928 12449 8956
rect 11296 8916 11302 8928
rect 12437 8925 12449 8928
rect 12483 8925 12495 8959
rect 12437 8919 12495 8925
rect 12529 8959 12587 8965
rect 12529 8925 12541 8959
rect 12575 8925 12587 8959
rect 12529 8919 12587 8925
rect 14093 8959 14151 8965
rect 14093 8925 14105 8959
rect 14139 8925 14151 8959
rect 14093 8919 14151 8925
rect 19521 8959 19579 8965
rect 19521 8925 19533 8959
rect 19567 8925 19579 8959
rect 19521 8919 19579 8925
rect 12250 8848 12256 8900
rect 12308 8888 12314 8900
rect 12544 8888 12572 8919
rect 12308 8860 12572 8888
rect 12308 8848 12314 8860
rect 13170 8848 13176 8900
rect 13228 8888 13234 8900
rect 14108 8888 14136 8919
rect 13228 8860 14136 8888
rect 13228 8848 13234 8860
rect 14918 8848 14924 8900
rect 14976 8848 14982 8900
rect 15746 8888 15752 8900
rect 15707 8860 15752 8888
rect 15746 8848 15752 8860
rect 15804 8848 15810 8900
rect 19242 8848 19248 8900
rect 19300 8888 19306 8900
rect 19536 8888 19564 8919
rect 21450 8916 21456 8968
rect 21508 8956 21514 8968
rect 21637 8959 21695 8965
rect 21637 8956 21649 8959
rect 21508 8928 21649 8956
rect 21508 8916 21514 8928
rect 21637 8925 21649 8928
rect 21683 8925 21695 8959
rect 21637 8919 21695 8925
rect 21821 8959 21879 8965
rect 21821 8925 21833 8959
rect 21867 8956 21879 8959
rect 22002 8956 22008 8968
rect 21867 8928 22008 8956
rect 21867 8925 21879 8928
rect 21821 8919 21879 8925
rect 22002 8916 22008 8928
rect 22060 8916 22066 8968
rect 23385 8959 23443 8965
rect 23385 8925 23397 8959
rect 23431 8925 23443 8959
rect 23385 8919 23443 8925
rect 19300 8860 19564 8888
rect 19300 8848 19306 8860
rect 13538 8780 13544 8832
rect 13596 8820 13602 8832
rect 14553 8823 14611 8829
rect 14553 8820 14565 8823
rect 13596 8792 14565 8820
rect 13596 8780 13602 8792
rect 14553 8789 14565 8792
rect 14599 8820 14611 8823
rect 14936 8820 14964 8848
rect 14599 8792 14964 8820
rect 15105 8823 15163 8829
rect 14599 8789 14611 8792
rect 14553 8783 14611 8789
rect 15105 8789 15117 8823
rect 15151 8820 15163 8823
rect 15286 8820 15292 8832
rect 15151 8792 15292 8820
rect 15151 8789 15163 8792
rect 15105 8783 15163 8789
rect 15286 8780 15292 8792
rect 15344 8780 15350 8832
rect 16022 8780 16028 8832
rect 16080 8820 16086 8832
rect 16117 8823 16175 8829
rect 16117 8820 16129 8823
rect 16080 8792 16129 8820
rect 16080 8780 16086 8792
rect 16117 8789 16129 8792
rect 16163 8789 16175 8823
rect 16117 8783 16175 8789
rect 16577 8823 16635 8829
rect 16577 8789 16589 8823
rect 16623 8820 16635 8823
rect 16666 8820 16672 8832
rect 16623 8792 16672 8820
rect 16623 8789 16635 8792
rect 16577 8783 16635 8789
rect 16666 8780 16672 8792
rect 16724 8820 16730 8832
rect 17862 8820 17868 8832
rect 16724 8792 17868 8820
rect 16724 8780 16730 8792
rect 17862 8780 17868 8792
rect 17920 8780 17926 8832
rect 18598 8820 18604 8832
rect 18559 8792 18604 8820
rect 18598 8780 18604 8792
rect 18656 8780 18662 8832
rect 18874 8820 18880 8832
rect 18835 8792 18880 8820
rect 18874 8780 18880 8792
rect 18932 8780 18938 8832
rect 19334 8780 19340 8832
rect 19392 8820 19398 8832
rect 19889 8823 19947 8829
rect 19889 8820 19901 8823
rect 19392 8792 19901 8820
rect 19392 8780 19398 8792
rect 19889 8789 19901 8792
rect 19935 8789 19947 8823
rect 23400 8820 23428 8919
rect 25130 8888 25136 8900
rect 24311 8860 25136 8888
rect 23566 8820 23572 8832
rect 23400 8792 23572 8820
rect 19889 8783 19947 8789
rect 23566 8780 23572 8792
rect 23624 8820 23630 8832
rect 24311 8820 24339 8860
rect 25130 8848 25136 8860
rect 25188 8848 25194 8900
rect 24762 8820 24768 8832
rect 23624 8792 24339 8820
rect 24723 8792 24768 8820
rect 23624 8780 23630 8792
rect 24762 8780 24768 8792
rect 24820 8780 24826 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 10962 8576 10968 8628
rect 11020 8616 11026 8628
rect 11238 8616 11244 8628
rect 11020 8588 11244 8616
rect 11020 8576 11026 8588
rect 11238 8576 11244 8588
rect 11296 8576 11302 8628
rect 12069 8619 12127 8625
rect 12069 8585 12081 8619
rect 12115 8616 12127 8619
rect 12342 8616 12348 8628
rect 12115 8588 12348 8616
rect 12115 8585 12127 8588
rect 12069 8579 12127 8585
rect 12342 8576 12348 8588
rect 12400 8576 12406 8628
rect 13170 8616 13176 8628
rect 13131 8588 13176 8616
rect 13170 8576 13176 8588
rect 13228 8576 13234 8628
rect 14734 8576 14740 8628
rect 14792 8616 14798 8628
rect 15013 8619 15071 8625
rect 15013 8616 15025 8619
rect 14792 8588 15025 8616
rect 14792 8576 14798 8588
rect 15013 8585 15025 8588
rect 15059 8585 15071 8619
rect 16114 8616 16120 8628
rect 16075 8588 16120 8616
rect 15013 8579 15071 8585
rect 16114 8576 16120 8588
rect 16172 8576 16178 8628
rect 16942 8576 16948 8628
rect 17000 8616 17006 8628
rect 17129 8619 17187 8625
rect 17129 8616 17141 8619
rect 17000 8588 17141 8616
rect 17000 8576 17006 8588
rect 17129 8585 17141 8588
rect 17175 8585 17187 8619
rect 17129 8579 17187 8585
rect 18601 8619 18659 8625
rect 18601 8585 18613 8619
rect 18647 8616 18659 8619
rect 19426 8616 19432 8628
rect 18647 8588 19432 8616
rect 18647 8585 18659 8588
rect 18601 8579 18659 8585
rect 19426 8576 19432 8588
rect 19484 8616 19490 8628
rect 19484 8588 20300 8616
rect 19484 8576 19490 8588
rect 12360 8480 12388 8576
rect 20272 8548 20300 8588
rect 20346 8576 20352 8628
rect 20404 8616 20410 8628
rect 20441 8619 20499 8625
rect 20441 8616 20453 8619
rect 20404 8588 20453 8616
rect 20404 8576 20410 8588
rect 20441 8585 20453 8588
rect 20487 8585 20499 8619
rect 20714 8616 20720 8628
rect 20675 8588 20720 8616
rect 20441 8579 20499 8585
rect 20714 8576 20720 8588
rect 20772 8576 20778 8628
rect 21266 8616 21272 8628
rect 21227 8588 21272 8616
rect 21266 8576 21272 8588
rect 21324 8576 21330 8628
rect 23474 8616 23480 8628
rect 23435 8588 23480 8616
rect 23474 8576 23480 8588
rect 23532 8576 23538 8628
rect 24210 8616 24216 8628
rect 23584 8588 24216 8616
rect 23109 8551 23167 8557
rect 20272 8520 20392 8548
rect 20364 8492 20392 8520
rect 23109 8517 23121 8551
rect 23155 8548 23167 8551
rect 23584 8548 23612 8588
rect 24210 8576 24216 8588
rect 24268 8576 24274 8628
rect 23155 8520 23612 8548
rect 23661 8551 23719 8557
rect 23155 8517 23167 8520
rect 23109 8511 23167 8517
rect 23661 8517 23673 8551
rect 23707 8517 23719 8551
rect 24673 8551 24731 8557
rect 24673 8548 24685 8551
rect 23661 8511 23719 8517
rect 24136 8520 24685 8548
rect 12437 8483 12495 8489
rect 12437 8480 12449 8483
rect 12360 8452 12449 8480
rect 12437 8449 12449 8452
rect 12483 8449 12495 8483
rect 12437 8443 12495 8449
rect 12526 8440 12532 8492
rect 12584 8480 12590 8492
rect 13538 8480 13544 8492
rect 12584 8452 13544 8480
rect 12584 8440 12590 8452
rect 13538 8440 13544 8452
rect 13596 8480 13602 8492
rect 13633 8483 13691 8489
rect 13633 8480 13645 8483
rect 13596 8452 13645 8480
rect 13596 8440 13602 8452
rect 13633 8449 13645 8452
rect 13679 8449 13691 8483
rect 13633 8443 13691 8449
rect 16574 8440 16580 8492
rect 16632 8480 16638 8492
rect 16761 8483 16819 8489
rect 16761 8480 16773 8483
rect 16632 8452 16773 8480
rect 16632 8440 16638 8452
rect 16761 8449 16773 8452
rect 16807 8480 16819 8483
rect 17497 8483 17555 8489
rect 17497 8480 17509 8483
rect 16807 8452 17509 8480
rect 16807 8449 16819 8452
rect 16761 8443 16819 8449
rect 17497 8449 17509 8452
rect 17543 8449 17555 8483
rect 17497 8443 17555 8449
rect 20346 8440 20352 8492
rect 20404 8440 20410 8492
rect 21266 8440 21272 8492
rect 21324 8480 21330 8492
rect 21913 8483 21971 8489
rect 21913 8480 21925 8483
rect 21324 8452 21925 8480
rect 21324 8440 21330 8452
rect 21913 8449 21925 8452
rect 21959 8480 21971 8483
rect 22281 8483 22339 8489
rect 22281 8480 22293 8483
rect 21959 8452 22293 8480
rect 21959 8449 21971 8452
rect 21913 8443 21971 8449
rect 22281 8449 22293 8452
rect 22327 8449 22339 8483
rect 22281 8443 22339 8449
rect 13446 8412 13452 8424
rect 13407 8384 13452 8412
rect 13446 8372 13452 8384
rect 13504 8372 13510 8424
rect 15010 8372 15016 8424
rect 15068 8412 15074 8424
rect 15286 8412 15292 8424
rect 15068 8384 15292 8412
rect 15068 8372 15074 8384
rect 15286 8372 15292 8384
rect 15344 8412 15350 8424
rect 16025 8415 16083 8421
rect 16025 8412 16037 8415
rect 15344 8384 16037 8412
rect 15344 8372 15350 8384
rect 16025 8381 16037 8384
rect 16071 8381 16083 8415
rect 16025 8375 16083 8381
rect 11333 8347 11391 8353
rect 11333 8313 11345 8347
rect 11379 8344 11391 8347
rect 11974 8344 11980 8356
rect 11379 8316 11980 8344
rect 11379 8313 11391 8316
rect 11333 8307 11391 8313
rect 11974 8304 11980 8316
rect 12032 8304 12038 8356
rect 13900 8347 13958 8353
rect 13900 8313 13912 8347
rect 13946 8344 13958 8347
rect 13998 8344 14004 8356
rect 13946 8316 14004 8344
rect 13946 8313 13958 8316
rect 13900 8307 13958 8313
rect 13998 8304 14004 8316
rect 14056 8304 14062 8356
rect 15470 8304 15476 8356
rect 15528 8344 15534 8356
rect 15657 8347 15715 8353
rect 15657 8344 15669 8347
rect 15528 8316 15669 8344
rect 15528 8304 15534 8316
rect 15657 8313 15669 8316
rect 15703 8344 15715 8347
rect 15746 8344 15752 8356
rect 15703 8316 15752 8344
rect 15703 8313 15715 8316
rect 15657 8307 15715 8313
rect 15746 8304 15752 8316
rect 15804 8304 15810 8356
rect 16040 8344 16068 8375
rect 16114 8372 16120 8424
rect 16172 8412 16178 8424
rect 16485 8415 16543 8421
rect 16485 8412 16497 8415
rect 16172 8384 16497 8412
rect 16172 8372 16178 8384
rect 16485 8381 16497 8384
rect 16531 8381 16543 8415
rect 16485 8375 16543 8381
rect 19061 8415 19119 8421
rect 19061 8381 19073 8415
rect 19107 8412 19119 8415
rect 19150 8412 19156 8424
rect 19107 8384 19156 8412
rect 19107 8381 19119 8384
rect 19061 8375 19119 8381
rect 19150 8372 19156 8384
rect 19208 8372 19214 8424
rect 20714 8372 20720 8424
rect 20772 8412 20778 8424
rect 21637 8415 21695 8421
rect 21637 8412 21649 8415
rect 20772 8384 21649 8412
rect 20772 8372 20778 8384
rect 21637 8381 21649 8384
rect 21683 8412 21695 8415
rect 21726 8412 21732 8424
rect 21683 8384 21732 8412
rect 21683 8381 21695 8384
rect 21637 8375 21695 8381
rect 21726 8372 21732 8384
rect 21784 8372 21790 8424
rect 23676 8412 23704 8511
rect 23934 8440 23940 8492
rect 23992 8480 23998 8492
rect 24136 8489 24164 8520
rect 24673 8517 24685 8520
rect 24719 8517 24731 8551
rect 24673 8511 24731 8517
rect 24121 8483 24179 8489
rect 24121 8480 24133 8483
rect 23992 8452 24133 8480
rect 23992 8440 23998 8452
rect 24121 8449 24133 8452
rect 24167 8449 24179 8483
rect 24121 8443 24179 8449
rect 24210 8440 24216 8492
rect 24268 8480 24274 8492
rect 24268 8452 24313 8480
rect 24268 8440 24274 8452
rect 25225 8415 25283 8421
rect 25225 8412 25237 8415
rect 23676 8384 25237 8412
rect 25225 8381 25237 8384
rect 25271 8412 25283 8415
rect 25961 8415 26019 8421
rect 25961 8412 25973 8415
rect 25271 8384 25973 8412
rect 25271 8381 25283 8384
rect 25225 8375 25283 8381
rect 25961 8381 25973 8384
rect 26007 8381 26019 8415
rect 25961 8375 26019 8381
rect 17034 8344 17040 8356
rect 16040 8316 17040 8344
rect 17034 8304 17040 8316
rect 17092 8304 17098 8356
rect 18966 8344 18972 8356
rect 18927 8316 18972 8344
rect 18966 8304 18972 8316
rect 19024 8304 19030 8356
rect 19328 8347 19386 8353
rect 19328 8313 19340 8347
rect 19374 8344 19386 8347
rect 19518 8344 19524 8356
rect 19374 8316 19524 8344
rect 19374 8313 19386 8316
rect 19328 8307 19386 8313
rect 19518 8304 19524 8316
rect 19576 8304 19582 8356
rect 21177 8347 21235 8353
rect 21177 8313 21189 8347
rect 21223 8344 21235 8347
rect 21223 8316 21404 8344
rect 21223 8313 21235 8316
rect 21177 8307 21235 8313
rect 15286 8236 15292 8288
rect 15344 8276 15350 8288
rect 15841 8279 15899 8285
rect 15841 8276 15853 8279
rect 15344 8248 15853 8276
rect 15344 8236 15350 8248
rect 15841 8245 15853 8248
rect 15887 8245 15899 8279
rect 15841 8239 15899 8245
rect 16577 8279 16635 8285
rect 16577 8245 16589 8279
rect 16623 8276 16635 8279
rect 16666 8276 16672 8288
rect 16623 8248 16672 8276
rect 16623 8245 16635 8248
rect 16577 8239 16635 8245
rect 16666 8236 16672 8248
rect 16724 8236 16730 8288
rect 18046 8276 18052 8288
rect 18007 8248 18052 8276
rect 18046 8236 18052 8248
rect 18104 8236 18110 8288
rect 21376 8276 21404 8316
rect 21450 8304 21456 8356
rect 21508 8344 21514 8356
rect 22649 8347 22707 8353
rect 22649 8344 22661 8347
rect 21508 8316 22661 8344
rect 21508 8304 21514 8316
rect 22649 8313 22661 8316
rect 22695 8313 22707 8347
rect 22649 8307 22707 8313
rect 23474 8304 23480 8356
rect 23532 8344 23538 8356
rect 24029 8347 24087 8353
rect 24029 8344 24041 8347
rect 23532 8316 24041 8344
rect 23532 8304 23538 8316
rect 24029 8313 24041 8316
rect 24075 8313 24087 8347
rect 25498 8344 25504 8356
rect 25459 8316 25504 8344
rect 24029 8307 24087 8313
rect 25498 8304 25504 8316
rect 25556 8304 25562 8356
rect 21729 8279 21787 8285
rect 21729 8276 21741 8279
rect 21376 8248 21741 8276
rect 21729 8245 21741 8248
rect 21775 8276 21787 8279
rect 21910 8276 21916 8288
rect 21775 8248 21916 8276
rect 21775 8245 21787 8248
rect 21729 8239 21787 8245
rect 21910 8236 21916 8248
rect 21968 8236 21974 8288
rect 25130 8276 25136 8288
rect 25091 8248 25136 8276
rect 25130 8236 25136 8248
rect 25188 8236 25194 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 9953 8075 10011 8081
rect 9953 8041 9965 8075
rect 9999 8072 10011 8075
rect 10686 8072 10692 8084
rect 9999 8044 10692 8072
rect 9999 8041 10011 8044
rect 9953 8035 10011 8041
rect 10686 8032 10692 8044
rect 10744 8032 10750 8084
rect 10962 8072 10968 8084
rect 10923 8044 10968 8072
rect 10962 8032 10968 8044
rect 11020 8032 11026 8084
rect 14366 8032 14372 8084
rect 14424 8072 14430 8084
rect 14829 8075 14887 8081
rect 14829 8072 14841 8075
rect 14424 8044 14841 8072
rect 14424 8032 14430 8044
rect 14829 8041 14841 8044
rect 14875 8072 14887 8075
rect 16942 8072 16948 8084
rect 14875 8044 16712 8072
rect 16903 8044 16948 8072
rect 14875 8041 14887 8044
rect 14829 8035 14887 8041
rect 12069 8007 12127 8013
rect 12069 7973 12081 8007
rect 12115 8004 12127 8007
rect 12250 8004 12256 8016
rect 12115 7976 12256 8004
rect 12115 7973 12127 7976
rect 12069 7967 12127 7973
rect 12250 7964 12256 7976
rect 12308 8004 12314 8016
rect 15838 8013 15844 8016
rect 12774 8007 12832 8013
rect 12774 8004 12786 8007
rect 12308 7976 12786 8004
rect 12308 7964 12314 7976
rect 12774 7973 12786 7976
rect 12820 7973 12832 8007
rect 15832 8004 15844 8013
rect 15799 7976 15844 8004
rect 12774 7967 12832 7973
rect 15832 7967 15844 7976
rect 15838 7964 15844 7967
rect 15896 7964 15902 8016
rect 16684 8004 16712 8044
rect 16942 8032 16948 8044
rect 17000 8032 17006 8084
rect 17218 8072 17224 8084
rect 17179 8044 17224 8072
rect 17218 8032 17224 8044
rect 17276 8032 17282 8084
rect 17678 8072 17684 8084
rect 17639 8044 17684 8072
rect 17678 8032 17684 8044
rect 17736 8032 17742 8084
rect 18506 8072 18512 8084
rect 18467 8044 18512 8072
rect 18506 8032 18512 8044
rect 18564 8032 18570 8084
rect 19518 8072 19524 8084
rect 19479 8044 19524 8072
rect 19518 8032 19524 8044
rect 19576 8032 19582 8084
rect 21269 8075 21327 8081
rect 21269 8041 21281 8075
rect 21315 8072 21327 8075
rect 21726 8072 21732 8084
rect 21315 8044 21732 8072
rect 21315 8041 21327 8044
rect 21269 8035 21327 8041
rect 21726 8032 21732 8044
rect 21784 8032 21790 8084
rect 22002 8072 22008 8084
rect 21963 8044 22008 8072
rect 22002 8032 22008 8044
rect 22060 8032 22066 8084
rect 22738 8032 22744 8084
rect 22796 8072 22802 8084
rect 23017 8075 23075 8081
rect 23017 8072 23029 8075
rect 22796 8044 23029 8072
rect 22796 8032 22802 8044
rect 23017 8041 23029 8044
rect 23063 8072 23075 8075
rect 24121 8075 24179 8081
rect 24121 8072 24133 8075
rect 23063 8044 24133 8072
rect 23063 8041 23075 8044
rect 23017 8035 23075 8041
rect 24121 8041 24133 8044
rect 24167 8041 24179 8075
rect 25130 8072 25136 8084
rect 25091 8044 25136 8072
rect 24121 8035 24179 8041
rect 25130 8032 25136 8044
rect 25188 8032 25194 8084
rect 17696 8004 17724 8032
rect 16684 7976 17724 8004
rect 20717 8007 20775 8013
rect 20717 7973 20729 8007
rect 20763 8004 20775 8007
rect 20806 8004 20812 8016
rect 20763 7976 20812 8004
rect 20763 7973 20775 7976
rect 20717 7967 20775 7973
rect 20806 7964 20812 7976
rect 20864 8004 20870 8016
rect 21634 8004 21640 8016
rect 20864 7976 21640 8004
rect 20864 7964 20870 7976
rect 21634 7964 21640 7976
rect 21692 7964 21698 8016
rect 22830 7964 22836 8016
rect 22888 8004 22894 8016
rect 22925 8007 22983 8013
rect 22925 8004 22937 8007
rect 22888 7976 22937 8004
rect 22888 7964 22894 7976
rect 22925 7973 22937 7976
rect 22971 7973 22983 8007
rect 22925 7967 22983 7973
rect 23753 8007 23811 8013
rect 23753 7973 23765 8007
rect 23799 8004 23811 8007
rect 24210 8004 24216 8016
rect 23799 7976 24216 8004
rect 23799 7973 23811 7976
rect 23753 7967 23811 7973
rect 24210 7964 24216 7976
rect 24268 7964 24274 8016
rect 11333 7939 11391 7945
rect 11333 7905 11345 7939
rect 11379 7936 11391 7939
rect 11790 7936 11796 7948
rect 11379 7908 11796 7936
rect 11379 7905 11391 7908
rect 11333 7899 11391 7905
rect 11790 7896 11796 7908
rect 11848 7896 11854 7948
rect 14642 7896 14648 7948
rect 14700 7936 14706 7948
rect 15010 7936 15016 7948
rect 14700 7908 15016 7936
rect 14700 7896 14706 7908
rect 15010 7896 15016 7908
rect 15068 7896 15074 7948
rect 17954 7896 17960 7948
rect 18012 7936 18018 7948
rect 18877 7939 18935 7945
rect 18877 7936 18889 7939
rect 18012 7908 18889 7936
rect 18012 7896 18018 7908
rect 18877 7905 18889 7908
rect 18923 7905 18935 7939
rect 20254 7936 20260 7948
rect 20215 7908 20260 7936
rect 18877 7899 18935 7905
rect 20254 7896 20260 7908
rect 20312 7896 20318 7948
rect 23198 7936 23204 7948
rect 21376 7908 23204 7936
rect 11054 7828 11060 7880
rect 11112 7868 11118 7880
rect 11425 7871 11483 7877
rect 11425 7868 11437 7871
rect 11112 7840 11437 7868
rect 11112 7828 11118 7840
rect 11425 7837 11437 7840
rect 11471 7837 11483 7871
rect 11606 7868 11612 7880
rect 11567 7840 11612 7868
rect 11425 7831 11483 7837
rect 11606 7828 11612 7840
rect 11664 7828 11670 7880
rect 12526 7868 12532 7880
rect 12360 7840 12532 7868
rect 11330 7692 11336 7744
rect 11388 7732 11394 7744
rect 12360 7741 12388 7840
rect 12526 7828 12532 7840
rect 12584 7828 12590 7880
rect 15470 7828 15476 7880
rect 15528 7868 15534 7880
rect 15565 7871 15623 7877
rect 15565 7868 15577 7871
rect 15528 7840 15577 7868
rect 15528 7828 15534 7840
rect 15565 7837 15577 7840
rect 15611 7837 15623 7871
rect 18966 7868 18972 7880
rect 18927 7840 18972 7868
rect 15565 7831 15623 7837
rect 18966 7828 18972 7840
rect 19024 7828 19030 7880
rect 19058 7828 19064 7880
rect 19116 7868 19122 7880
rect 19116 7840 19161 7868
rect 19116 7828 19122 7840
rect 20346 7828 20352 7880
rect 20404 7868 20410 7880
rect 21376 7877 21404 7908
rect 23198 7896 23204 7908
rect 23256 7896 23262 7948
rect 23474 7896 23480 7948
rect 23532 7936 23538 7948
rect 24118 7936 24124 7948
rect 23532 7908 24124 7936
rect 23532 7896 23538 7908
rect 24118 7896 24124 7908
rect 24176 7936 24182 7948
rect 24489 7939 24547 7945
rect 24489 7936 24501 7939
rect 24176 7908 24501 7936
rect 24176 7896 24182 7908
rect 24489 7905 24501 7908
rect 24535 7905 24547 7939
rect 24489 7899 24547 7905
rect 24581 7939 24639 7945
rect 24581 7905 24593 7939
rect 24627 7936 24639 7939
rect 25406 7936 25412 7948
rect 24627 7908 25412 7936
rect 24627 7905 24639 7908
rect 24581 7899 24639 7905
rect 25406 7896 25412 7908
rect 25464 7896 25470 7948
rect 21361 7871 21419 7877
rect 21361 7868 21373 7871
rect 20404 7840 21373 7868
rect 20404 7828 20410 7840
rect 21361 7837 21373 7840
rect 21407 7837 21419 7871
rect 21361 7831 21419 7837
rect 21545 7871 21603 7877
rect 21545 7837 21557 7871
rect 21591 7868 21603 7871
rect 21634 7868 21640 7880
rect 21591 7840 21640 7868
rect 21591 7837 21603 7840
rect 21545 7831 21603 7837
rect 21634 7828 21640 7840
rect 21692 7828 21698 7880
rect 23014 7828 23020 7880
rect 23072 7868 23078 7880
rect 23109 7871 23167 7877
rect 23109 7868 23121 7871
rect 23072 7840 23121 7868
rect 23072 7828 23078 7840
rect 23109 7837 23121 7840
rect 23155 7837 23167 7871
rect 24762 7868 24768 7880
rect 24723 7840 24768 7868
rect 23109 7831 23167 7837
rect 24762 7828 24768 7840
rect 24820 7828 24826 7880
rect 19978 7800 19984 7812
rect 19891 7772 19984 7800
rect 19978 7760 19984 7772
rect 20036 7800 20042 7812
rect 20073 7803 20131 7809
rect 20073 7800 20085 7803
rect 20036 7772 20085 7800
rect 20036 7760 20042 7772
rect 20073 7769 20085 7772
rect 20119 7800 20131 7803
rect 21082 7800 21088 7812
rect 20119 7772 21088 7800
rect 20119 7769 20131 7772
rect 20073 7763 20131 7769
rect 21082 7760 21088 7772
rect 21140 7760 21146 7812
rect 12345 7735 12403 7741
rect 12345 7732 12357 7735
rect 11388 7704 12357 7732
rect 11388 7692 11394 7704
rect 12345 7701 12357 7704
rect 12391 7701 12403 7735
rect 12345 7695 12403 7701
rect 13909 7735 13967 7741
rect 13909 7701 13921 7735
rect 13955 7732 13967 7735
rect 13998 7732 14004 7744
rect 13955 7704 14004 7732
rect 13955 7701 13967 7704
rect 13909 7695 13967 7701
rect 13998 7692 14004 7704
rect 14056 7732 14062 7744
rect 14185 7735 14243 7741
rect 14185 7732 14197 7735
rect 14056 7704 14197 7732
rect 14056 7692 14062 7704
rect 14185 7701 14197 7704
rect 14231 7701 14243 7735
rect 14550 7732 14556 7744
rect 14511 7704 14556 7732
rect 14185 7695 14243 7701
rect 14550 7692 14556 7704
rect 14608 7692 14614 7744
rect 17954 7732 17960 7744
rect 17915 7704 17960 7732
rect 17954 7692 17960 7704
rect 18012 7692 18018 7744
rect 18417 7735 18475 7741
rect 18417 7701 18429 7735
rect 18463 7732 18475 7735
rect 19242 7732 19248 7744
rect 18463 7704 19248 7732
rect 18463 7701 18475 7704
rect 18417 7695 18475 7701
rect 19242 7692 19248 7704
rect 19300 7692 19306 7744
rect 20714 7692 20720 7744
rect 20772 7732 20778 7744
rect 20901 7735 20959 7741
rect 20901 7732 20913 7735
rect 20772 7704 20913 7732
rect 20772 7692 20778 7704
rect 20901 7701 20913 7704
rect 20947 7701 20959 7735
rect 20901 7695 20959 7701
rect 22186 7692 22192 7744
rect 22244 7732 22250 7744
rect 22373 7735 22431 7741
rect 22373 7732 22385 7735
rect 22244 7704 22385 7732
rect 22244 7692 22250 7704
rect 22373 7701 22385 7704
rect 22419 7732 22431 7735
rect 22557 7735 22615 7741
rect 22557 7732 22569 7735
rect 22419 7704 22569 7732
rect 22419 7701 22431 7704
rect 22373 7695 22431 7701
rect 22557 7701 22569 7704
rect 22603 7701 22615 7735
rect 22557 7695 22615 7701
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 4154 7488 4160 7540
rect 4212 7528 4218 7540
rect 5442 7528 5448 7540
rect 4212 7500 5448 7528
rect 4212 7488 4218 7500
rect 5442 7488 5448 7500
rect 5500 7488 5506 7540
rect 12250 7528 12256 7540
rect 12211 7500 12256 7528
rect 12250 7488 12256 7500
rect 12308 7488 12314 7540
rect 12986 7528 12992 7540
rect 12947 7500 12992 7528
rect 12986 7488 12992 7500
rect 13044 7488 13050 7540
rect 13998 7528 14004 7540
rect 13959 7500 14004 7528
rect 13998 7488 14004 7500
rect 14056 7488 14062 7540
rect 15838 7488 15844 7540
rect 15896 7528 15902 7540
rect 15933 7531 15991 7537
rect 15933 7528 15945 7531
rect 15896 7500 15945 7528
rect 15896 7488 15902 7500
rect 15933 7497 15945 7500
rect 15979 7528 15991 7531
rect 16209 7531 16267 7537
rect 16209 7528 16221 7531
rect 15979 7500 16221 7528
rect 15979 7497 15991 7500
rect 15933 7491 15991 7497
rect 16209 7497 16221 7500
rect 16255 7497 16267 7531
rect 17402 7528 17408 7540
rect 17363 7500 17408 7528
rect 16209 7491 16267 7497
rect 17402 7488 17408 7500
rect 17460 7488 17466 7540
rect 18325 7531 18383 7537
rect 18325 7497 18337 7531
rect 18371 7528 18383 7531
rect 19058 7528 19064 7540
rect 18371 7500 19064 7528
rect 18371 7497 18383 7500
rect 18325 7491 18383 7497
rect 19058 7488 19064 7500
rect 19116 7528 19122 7540
rect 19518 7528 19524 7540
rect 19116 7500 19524 7528
rect 19116 7488 19122 7500
rect 19518 7488 19524 7500
rect 19576 7528 19582 7540
rect 19797 7531 19855 7537
rect 19797 7528 19809 7531
rect 19576 7500 19809 7528
rect 19576 7488 19582 7500
rect 19797 7497 19809 7500
rect 19843 7497 19855 7531
rect 20622 7528 20628 7540
rect 20583 7500 20628 7528
rect 19797 7491 19855 7497
rect 20622 7488 20628 7500
rect 20680 7488 20686 7540
rect 22097 7531 22155 7537
rect 22097 7497 22109 7531
rect 22143 7528 22155 7531
rect 22830 7528 22836 7540
rect 22143 7500 22836 7528
rect 22143 7497 22155 7500
rect 22097 7491 22155 7497
rect 22830 7488 22836 7500
rect 22888 7488 22894 7540
rect 23014 7528 23020 7540
rect 22975 7500 23020 7528
rect 23014 7488 23020 7500
rect 23072 7488 23078 7540
rect 25406 7528 25412 7540
rect 25367 7500 25412 7528
rect 25406 7488 25412 7500
rect 25464 7488 25470 7540
rect 12802 7392 12808 7404
rect 12763 7364 12808 7392
rect 12802 7352 12808 7364
rect 12860 7392 12866 7404
rect 13633 7395 13691 7401
rect 12860 7364 13400 7392
rect 12860 7352 12866 7364
rect 13372 7333 13400 7364
rect 13633 7361 13645 7395
rect 13679 7392 13691 7395
rect 14016 7392 14044 7488
rect 19426 7420 19432 7472
rect 19484 7460 19490 7472
rect 20441 7463 20499 7469
rect 20441 7460 20453 7463
rect 19484 7432 20453 7460
rect 19484 7420 19490 7432
rect 20441 7429 20453 7432
rect 20487 7429 20499 7463
rect 20441 7423 20499 7429
rect 13679 7364 14044 7392
rect 14461 7395 14519 7401
rect 13679 7361 13691 7364
rect 13633 7355 13691 7361
rect 14461 7361 14473 7395
rect 14507 7392 14519 7395
rect 14507 7364 14688 7392
rect 14507 7361 14519 7364
rect 14461 7355 14519 7361
rect 10137 7327 10195 7333
rect 10137 7324 10149 7327
rect 9968 7296 10149 7324
rect 9677 7191 9735 7197
rect 9677 7157 9689 7191
rect 9723 7188 9735 7191
rect 9968 7188 9996 7296
rect 10137 7293 10149 7296
rect 10183 7293 10195 7327
rect 10137 7287 10195 7293
rect 13357 7327 13415 7333
rect 13357 7293 13369 7327
rect 13403 7293 13415 7327
rect 13357 7287 13415 7293
rect 14366 7284 14372 7336
rect 14424 7324 14430 7336
rect 14553 7327 14611 7333
rect 14553 7324 14565 7327
rect 14424 7296 14565 7324
rect 14424 7284 14430 7296
rect 14553 7293 14565 7296
rect 14599 7293 14611 7327
rect 14660 7324 14688 7364
rect 14826 7333 14832 7336
rect 14820 7324 14832 7333
rect 14660 7296 14832 7324
rect 14553 7287 14611 7293
rect 14820 7287 14832 7296
rect 14826 7284 14832 7287
rect 14884 7284 14890 7336
rect 16761 7327 16819 7333
rect 16761 7293 16773 7327
rect 16807 7324 16819 7327
rect 17402 7324 17408 7336
rect 16807 7296 17408 7324
rect 16807 7293 16819 7296
rect 16761 7287 16819 7293
rect 17402 7284 17408 7296
rect 17460 7284 17466 7336
rect 17586 7284 17592 7336
rect 17644 7324 17650 7336
rect 18417 7327 18475 7333
rect 18417 7324 18429 7327
rect 17644 7296 18429 7324
rect 17644 7284 17650 7296
rect 18417 7293 18429 7296
rect 18463 7324 18475 7327
rect 19150 7324 19156 7336
rect 18463 7296 19156 7324
rect 18463 7293 18475 7296
rect 18417 7287 18475 7293
rect 19150 7284 19156 7296
rect 19208 7324 19214 7336
rect 19978 7324 19984 7336
rect 19208 7296 19984 7324
rect 19208 7284 19214 7296
rect 19978 7284 19984 7296
rect 20036 7284 20042 7336
rect 20456 7324 20484 7423
rect 21174 7392 21180 7404
rect 21135 7364 21180 7392
rect 21174 7352 21180 7364
rect 21232 7352 21238 7404
rect 22370 7392 22376 7404
rect 22331 7364 22376 7392
rect 22370 7352 22376 7364
rect 22428 7352 22434 7404
rect 23198 7352 23204 7404
rect 23256 7392 23262 7404
rect 23566 7392 23572 7404
rect 23256 7364 23572 7392
rect 23256 7352 23262 7364
rect 23566 7352 23572 7364
rect 23624 7392 23630 7404
rect 23661 7395 23719 7401
rect 23661 7392 23673 7395
rect 23624 7364 23673 7392
rect 23624 7352 23630 7364
rect 23661 7361 23673 7364
rect 23707 7361 23719 7395
rect 23661 7355 23719 7361
rect 21085 7327 21143 7333
rect 21085 7324 21097 7327
rect 20456 7296 21097 7324
rect 21085 7293 21097 7296
rect 21131 7293 21143 7327
rect 22186 7324 22192 7336
rect 22147 7296 22192 7324
rect 21085 7287 21143 7293
rect 22186 7284 22192 7296
rect 22244 7284 22250 7336
rect 10045 7259 10103 7265
rect 10045 7225 10057 7259
rect 10091 7256 10103 7259
rect 10404 7259 10462 7265
rect 10404 7256 10416 7259
rect 10091 7228 10416 7256
rect 10091 7225 10103 7228
rect 10045 7219 10103 7225
rect 10404 7225 10416 7228
rect 10450 7256 10462 7259
rect 10778 7256 10784 7268
rect 10450 7228 10784 7256
rect 10450 7225 10462 7228
rect 10404 7219 10462 7225
rect 10778 7216 10784 7228
rect 10836 7216 10842 7268
rect 18662 7259 18720 7265
rect 18662 7256 18674 7259
rect 17788 7228 18674 7256
rect 11330 7188 11336 7200
rect 9723 7160 11336 7188
rect 9723 7157 9735 7160
rect 9677 7151 9735 7157
rect 11330 7148 11336 7160
rect 11388 7148 11394 7200
rect 11517 7191 11575 7197
rect 11517 7157 11529 7191
rect 11563 7188 11575 7191
rect 11606 7188 11612 7200
rect 11563 7160 11612 7188
rect 11563 7157 11575 7160
rect 11517 7151 11575 7157
rect 11606 7148 11612 7160
rect 11664 7148 11670 7200
rect 11790 7188 11796 7200
rect 11751 7160 11796 7188
rect 11790 7148 11796 7160
rect 11848 7148 11854 7200
rect 13446 7188 13452 7200
rect 13407 7160 13452 7188
rect 13446 7148 13452 7160
rect 13504 7148 13510 7200
rect 16574 7188 16580 7200
rect 16535 7160 16580 7188
rect 16574 7148 16580 7160
rect 16632 7148 16638 7200
rect 16666 7148 16672 7200
rect 16724 7188 16730 7200
rect 16945 7191 17003 7197
rect 16945 7188 16957 7191
rect 16724 7160 16957 7188
rect 16724 7148 16730 7160
rect 16945 7157 16957 7160
rect 16991 7157 17003 7191
rect 16945 7151 17003 7157
rect 17678 7148 17684 7200
rect 17736 7188 17742 7200
rect 17788 7197 17816 7228
rect 18662 7225 18674 7228
rect 18708 7225 18720 7259
rect 18662 7219 18720 7225
rect 23658 7216 23664 7268
rect 23716 7256 23722 7268
rect 23906 7259 23964 7265
rect 23906 7256 23918 7259
rect 23716 7228 23918 7256
rect 23716 7216 23722 7228
rect 23906 7225 23918 7228
rect 23952 7225 23964 7259
rect 23906 7219 23964 7225
rect 17773 7191 17831 7197
rect 17773 7188 17785 7191
rect 17736 7160 17785 7188
rect 17736 7148 17742 7160
rect 17773 7157 17785 7160
rect 17819 7157 17831 7191
rect 17773 7151 17831 7157
rect 20165 7191 20223 7197
rect 20165 7157 20177 7191
rect 20211 7188 20223 7191
rect 20346 7188 20352 7200
rect 20211 7160 20352 7188
rect 20211 7157 20223 7160
rect 20165 7151 20223 7157
rect 20346 7148 20352 7160
rect 20404 7148 20410 7200
rect 20990 7188 20996 7200
rect 20951 7160 20996 7188
rect 20990 7148 20996 7160
rect 21048 7148 21054 7200
rect 21726 7188 21732 7200
rect 21687 7160 21732 7188
rect 21726 7148 21732 7160
rect 21784 7148 21790 7200
rect 23474 7188 23480 7200
rect 23435 7160 23480 7188
rect 23474 7148 23480 7160
rect 23532 7148 23538 7200
rect 25038 7188 25044 7200
rect 24999 7160 25044 7188
rect 25038 7148 25044 7160
rect 25096 7148 25102 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 12250 6944 12256 6996
rect 12308 6984 12314 6996
rect 12897 6987 12955 6993
rect 12897 6984 12909 6987
rect 12308 6956 12909 6984
rect 12308 6944 12314 6956
rect 12897 6953 12909 6956
rect 12943 6953 12955 6987
rect 12897 6947 12955 6953
rect 13265 6987 13323 6993
rect 13265 6953 13277 6987
rect 13311 6984 13323 6987
rect 13446 6984 13452 6996
rect 13311 6956 13452 6984
rect 13311 6953 13323 6956
rect 13265 6947 13323 6953
rect 13446 6944 13452 6956
rect 13504 6944 13510 6996
rect 14001 6987 14059 6993
rect 14001 6953 14013 6987
rect 14047 6984 14059 6987
rect 14366 6984 14372 6996
rect 14047 6956 14372 6984
rect 14047 6953 14059 6956
rect 14001 6947 14059 6953
rect 14366 6944 14372 6956
rect 14424 6984 14430 6996
rect 14550 6984 14556 6996
rect 14424 6956 14556 6984
rect 14424 6944 14430 6956
rect 14550 6944 14556 6956
rect 14608 6944 14614 6996
rect 14642 6944 14648 6996
rect 14700 6984 14706 6996
rect 14829 6987 14887 6993
rect 14829 6984 14841 6987
rect 14700 6956 14841 6984
rect 14700 6944 14706 6956
rect 14829 6953 14841 6956
rect 14875 6953 14887 6987
rect 14829 6947 14887 6953
rect 16482 6944 16488 6996
rect 16540 6984 16546 6996
rect 16577 6987 16635 6993
rect 16577 6984 16589 6987
rect 16540 6956 16589 6984
rect 16540 6944 16546 6956
rect 16577 6953 16589 6956
rect 16623 6953 16635 6987
rect 16577 6947 16635 6953
rect 19981 6987 20039 6993
rect 19981 6953 19993 6987
rect 20027 6984 20039 6987
rect 20162 6984 20168 6996
rect 20027 6956 20168 6984
rect 20027 6953 20039 6956
rect 19981 6947 20039 6953
rect 20162 6944 20168 6956
rect 20220 6944 20226 6996
rect 20349 6987 20407 6993
rect 20349 6953 20361 6987
rect 20395 6984 20407 6987
rect 21174 6984 21180 6996
rect 20395 6956 21180 6984
rect 20395 6953 20407 6956
rect 20349 6947 20407 6953
rect 16500 6916 16528 6944
rect 16408 6888 16528 6916
rect 10318 6848 10324 6860
rect 10279 6820 10324 6848
rect 10318 6808 10324 6820
rect 10376 6808 10382 6860
rect 11425 6851 11483 6857
rect 11425 6817 11437 6851
rect 11471 6848 11483 6851
rect 11606 6848 11612 6860
rect 11471 6820 11612 6848
rect 11471 6817 11483 6820
rect 11425 6811 11483 6817
rect 11606 6808 11612 6820
rect 11664 6848 11670 6860
rect 11784 6851 11842 6857
rect 11784 6848 11796 6851
rect 11664 6820 11796 6848
rect 11664 6808 11670 6820
rect 11784 6817 11796 6820
rect 11830 6848 11842 6851
rect 12158 6848 12164 6860
rect 11830 6820 12164 6848
rect 11830 6817 11842 6820
rect 11784 6811 11842 6817
rect 12158 6808 12164 6820
rect 12216 6808 12222 6860
rect 14090 6848 14096 6860
rect 14051 6820 14096 6848
rect 14090 6808 14096 6820
rect 14148 6808 14154 6860
rect 16025 6851 16083 6857
rect 16025 6817 16037 6851
rect 16071 6848 16083 6851
rect 16408 6848 16436 6888
rect 19334 6876 19340 6928
rect 19392 6916 19398 6928
rect 20364 6916 20392 6947
rect 21174 6944 21180 6956
rect 21232 6944 21238 6996
rect 22002 6944 22008 6996
rect 22060 6984 22066 6996
rect 22373 6987 22431 6993
rect 22373 6984 22385 6987
rect 22060 6956 22385 6984
rect 22060 6944 22066 6956
rect 22373 6953 22385 6956
rect 22419 6953 22431 6987
rect 22738 6984 22744 6996
rect 22699 6956 22744 6984
rect 22373 6947 22431 6953
rect 19392 6888 20392 6916
rect 22388 6916 22416 6947
rect 22738 6944 22744 6956
rect 22796 6944 22802 6996
rect 24762 6944 24768 6996
rect 24820 6984 24826 6996
rect 24857 6987 24915 6993
rect 24857 6984 24869 6987
rect 24820 6956 24869 6984
rect 24820 6944 24826 6956
rect 24857 6953 24869 6956
rect 24903 6953 24915 6987
rect 24857 6947 24915 6953
rect 23474 6925 23480 6928
rect 23446 6919 23480 6925
rect 23446 6916 23458 6919
rect 22388 6888 23458 6916
rect 19392 6876 19398 6888
rect 23446 6885 23458 6888
rect 23532 6916 23538 6928
rect 23532 6888 23594 6916
rect 23446 6879 23480 6885
rect 23474 6876 23480 6879
rect 23532 6876 23538 6888
rect 16071 6820 16436 6848
rect 16485 6851 16543 6857
rect 16071 6817 16083 6820
rect 16025 6811 16083 6817
rect 16485 6817 16497 6851
rect 16531 6817 16543 6851
rect 16485 6811 16543 6817
rect 10134 6740 10140 6792
rect 10192 6780 10198 6792
rect 10413 6783 10471 6789
rect 10413 6780 10425 6783
rect 10192 6752 10425 6780
rect 10192 6740 10198 6752
rect 10413 6749 10425 6752
rect 10459 6749 10471 6783
rect 10413 6743 10471 6749
rect 10597 6783 10655 6789
rect 10597 6749 10609 6783
rect 10643 6780 10655 6783
rect 10778 6780 10784 6792
rect 10643 6752 10784 6780
rect 10643 6749 10655 6752
rect 10597 6743 10655 6749
rect 10778 6740 10784 6752
rect 10836 6740 10842 6792
rect 11330 6740 11336 6792
rect 11388 6780 11394 6792
rect 11517 6783 11575 6789
rect 11517 6780 11529 6783
rect 11388 6752 11529 6780
rect 11388 6740 11394 6752
rect 11517 6749 11529 6752
rect 11563 6749 11575 6783
rect 11517 6743 11575 6749
rect 15930 6740 15936 6792
rect 15988 6780 15994 6792
rect 15988 6752 16160 6780
rect 15988 6740 15994 6752
rect 9953 6715 10011 6721
rect 9953 6681 9965 6715
rect 9999 6712 10011 6715
rect 10042 6712 10048 6724
rect 9999 6684 10048 6712
rect 9999 6681 10011 6684
rect 9953 6675 10011 6681
rect 10042 6672 10048 6684
rect 10100 6672 10106 6724
rect 13262 6672 13268 6724
rect 13320 6712 13326 6724
rect 15470 6712 15476 6724
rect 13320 6684 15476 6712
rect 13320 6672 13326 6684
rect 15470 6672 15476 6684
rect 15528 6712 15534 6724
rect 16132 6721 16160 6752
rect 16298 6740 16304 6792
rect 16356 6780 16362 6792
rect 16500 6780 16528 6811
rect 16574 6808 16580 6860
rect 16632 6848 16638 6860
rect 17402 6848 17408 6860
rect 16632 6820 17408 6848
rect 16632 6808 16638 6820
rect 17402 6808 17408 6820
rect 17460 6848 17466 6860
rect 17586 6848 17592 6860
rect 17460 6820 17592 6848
rect 17460 6808 17466 6820
rect 17586 6808 17592 6820
rect 17644 6848 17650 6860
rect 17954 6857 17960 6860
rect 17681 6851 17739 6857
rect 17681 6848 17693 6851
rect 17644 6820 17693 6848
rect 17644 6808 17650 6820
rect 17681 6817 17693 6820
rect 17727 6817 17739 6851
rect 17948 6848 17960 6857
rect 17867 6820 17960 6848
rect 17681 6811 17739 6817
rect 17948 6811 17960 6820
rect 18012 6848 18018 6860
rect 18230 6848 18236 6860
rect 18012 6820 18236 6848
rect 17954 6808 17960 6811
rect 18012 6808 18018 6820
rect 18230 6808 18236 6820
rect 18288 6808 18294 6860
rect 20993 6851 21051 6857
rect 20993 6817 21005 6851
rect 21039 6848 21051 6851
rect 21082 6848 21088 6860
rect 21039 6820 21088 6848
rect 21039 6817 21051 6820
rect 20993 6811 21051 6817
rect 21082 6808 21088 6820
rect 21140 6808 21146 6860
rect 21266 6857 21272 6860
rect 21260 6848 21272 6857
rect 21227 6820 21272 6848
rect 21260 6811 21272 6820
rect 21266 6808 21272 6811
rect 21324 6808 21330 6860
rect 23198 6848 23204 6860
rect 23159 6820 23204 6848
rect 23198 6808 23204 6820
rect 23256 6808 23262 6860
rect 16356 6752 16528 6780
rect 16669 6783 16727 6789
rect 16356 6740 16362 6752
rect 16669 6749 16681 6783
rect 16715 6749 16727 6783
rect 16669 6743 16727 6749
rect 15565 6715 15623 6721
rect 15565 6712 15577 6715
rect 15528 6684 15577 6712
rect 15528 6672 15534 6684
rect 15565 6681 15577 6684
rect 15611 6681 15623 6715
rect 15565 6675 15623 6681
rect 16117 6715 16175 6721
rect 16117 6681 16129 6715
rect 16163 6681 16175 6715
rect 16684 6712 16712 6743
rect 24946 6740 24952 6792
rect 25004 6780 25010 6792
rect 25409 6783 25467 6789
rect 25409 6780 25421 6783
rect 25004 6752 25421 6780
rect 25004 6740 25010 6752
rect 25409 6749 25421 6752
rect 25455 6749 25467 6783
rect 25409 6743 25467 6749
rect 16117 6675 16175 6681
rect 16408 6684 16712 6712
rect 9493 6647 9551 6653
rect 9493 6613 9505 6647
rect 9539 6644 9551 6647
rect 9858 6644 9864 6656
rect 9539 6616 9864 6644
rect 9539 6613 9551 6616
rect 9493 6607 9551 6613
rect 9858 6604 9864 6616
rect 9916 6604 9922 6656
rect 11054 6644 11060 6656
rect 11015 6616 11060 6644
rect 11054 6604 11060 6616
rect 11112 6604 11118 6656
rect 14274 6644 14280 6656
rect 14235 6616 14280 6644
rect 14274 6604 14280 6616
rect 14332 6604 14338 6656
rect 15930 6604 15936 6656
rect 15988 6644 15994 6656
rect 16408 6644 16436 6684
rect 17586 6644 17592 6656
rect 15988 6616 16436 6644
rect 17547 6616 17592 6644
rect 15988 6604 15994 6616
rect 17586 6604 17592 6616
rect 17644 6604 17650 6656
rect 19058 6644 19064 6656
rect 19019 6616 19064 6644
rect 19058 6604 19064 6616
rect 19116 6604 19122 6656
rect 19334 6644 19340 6656
rect 19295 6616 19340 6644
rect 19334 6604 19340 6616
rect 19392 6604 19398 6656
rect 20717 6647 20775 6653
rect 20717 6613 20729 6647
rect 20763 6644 20775 6647
rect 20990 6644 20996 6656
rect 20763 6616 20996 6644
rect 20763 6613 20775 6616
rect 20717 6607 20775 6613
rect 20990 6604 20996 6616
rect 21048 6644 21054 6656
rect 21358 6644 21364 6656
rect 21048 6616 21364 6644
rect 21048 6604 21054 6616
rect 21358 6604 21364 6616
rect 21416 6604 21422 6656
rect 23109 6647 23167 6653
rect 23109 6613 23121 6647
rect 23155 6644 23167 6647
rect 23566 6644 23572 6656
rect 23155 6616 23572 6644
rect 23155 6613 23167 6616
rect 23109 6607 23167 6613
rect 23566 6604 23572 6616
rect 23624 6644 23630 6656
rect 24581 6647 24639 6653
rect 24581 6644 24593 6647
rect 23624 6616 24593 6644
rect 23624 6604 23630 6616
rect 24581 6613 24593 6616
rect 24627 6613 24639 6647
rect 24581 6607 24639 6613
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 10045 6443 10103 6449
rect 10045 6440 10057 6443
rect 9140 6412 10057 6440
rect 9140 6313 9168 6412
rect 10045 6409 10057 6412
rect 10091 6440 10103 6443
rect 10318 6440 10324 6452
rect 10091 6412 10324 6440
rect 10091 6409 10103 6412
rect 10045 6403 10103 6409
rect 10318 6400 10324 6412
rect 10376 6400 10382 6452
rect 10778 6400 10784 6452
rect 10836 6440 10842 6452
rect 11517 6443 11575 6449
rect 11517 6440 11529 6443
rect 10836 6412 11529 6440
rect 10836 6400 10842 6412
rect 11517 6409 11529 6412
rect 11563 6409 11575 6443
rect 12158 6440 12164 6452
rect 12119 6412 12164 6440
rect 11517 6403 11575 6409
rect 12158 6400 12164 6412
rect 12216 6400 12222 6452
rect 13170 6400 13176 6452
rect 13228 6440 13234 6452
rect 13265 6443 13323 6449
rect 13265 6440 13277 6443
rect 13228 6412 13277 6440
rect 13228 6400 13234 6412
rect 13265 6409 13277 6412
rect 13311 6409 13323 6443
rect 14826 6440 14832 6452
rect 14787 6412 14832 6440
rect 13265 6403 13323 6409
rect 9125 6307 9183 6313
rect 9125 6273 9137 6307
rect 9171 6273 9183 6307
rect 9125 6267 9183 6273
rect 9677 6307 9735 6313
rect 9677 6273 9689 6307
rect 9723 6304 9735 6307
rect 13280 6304 13308 6403
rect 14826 6400 14832 6412
rect 14884 6400 14890 6452
rect 16206 6440 16212 6452
rect 16167 6412 16212 6440
rect 16206 6400 16212 6412
rect 16264 6400 16270 6452
rect 16390 6440 16396 6452
rect 16351 6412 16396 6440
rect 16390 6400 16396 6412
rect 16448 6400 16454 6452
rect 17773 6443 17831 6449
rect 17773 6409 17785 6443
rect 17819 6440 17831 6443
rect 17954 6440 17960 6452
rect 17819 6412 17960 6440
rect 17819 6409 17831 6412
rect 17773 6403 17831 6409
rect 17954 6400 17960 6412
rect 18012 6400 18018 6452
rect 18233 6443 18291 6449
rect 18233 6409 18245 6443
rect 18279 6440 18291 6443
rect 18966 6440 18972 6452
rect 18279 6412 18972 6440
rect 18279 6409 18291 6412
rect 18233 6403 18291 6409
rect 18966 6400 18972 6412
rect 19024 6440 19030 6452
rect 19334 6440 19340 6452
rect 19024 6412 19340 6440
rect 19024 6400 19030 6412
rect 19334 6400 19340 6412
rect 19392 6400 19398 6452
rect 19518 6400 19524 6452
rect 19576 6440 19582 6452
rect 19705 6443 19763 6449
rect 19705 6440 19717 6443
rect 19576 6412 19717 6440
rect 19576 6400 19582 6412
rect 19705 6409 19717 6412
rect 19751 6409 19763 6443
rect 21266 6440 21272 6452
rect 21227 6412 21272 6440
rect 19705 6403 19763 6409
rect 15197 6375 15255 6381
rect 15197 6341 15209 6375
rect 15243 6372 15255 6375
rect 16298 6372 16304 6384
rect 15243 6344 16304 6372
rect 15243 6341 15255 6344
rect 15197 6335 15255 6341
rect 16298 6332 16304 6344
rect 16356 6332 16362 6384
rect 19245 6375 19303 6381
rect 19245 6341 19257 6375
rect 19291 6341 19303 6375
rect 19245 6335 19303 6341
rect 15933 6307 15991 6313
rect 9723 6276 10272 6304
rect 13280 6276 13584 6304
rect 9723 6273 9735 6276
rect 9677 6267 9735 6273
rect 9950 6196 9956 6248
rect 10008 6236 10014 6248
rect 10137 6239 10195 6245
rect 10137 6236 10149 6239
rect 10008 6208 10149 6236
rect 10008 6196 10014 6208
rect 10137 6205 10149 6208
rect 10183 6205 10195 6239
rect 10244 6236 10272 6276
rect 13556 6248 13584 6276
rect 15933 6273 15945 6307
rect 15979 6304 15991 6307
rect 16945 6307 17003 6313
rect 16945 6304 16957 6307
rect 15979 6276 16957 6304
rect 15979 6273 15991 6276
rect 15933 6267 15991 6273
rect 16945 6273 16957 6276
rect 16991 6304 17003 6307
rect 17678 6304 17684 6316
rect 16991 6276 17684 6304
rect 16991 6273 17003 6276
rect 16945 6267 17003 6273
rect 17678 6264 17684 6276
rect 17736 6304 17742 6316
rect 18785 6307 18843 6313
rect 18785 6304 18797 6307
rect 17736 6276 18797 6304
rect 17736 6264 17742 6276
rect 18785 6273 18797 6276
rect 18831 6304 18843 6307
rect 19058 6304 19064 6316
rect 18831 6276 19064 6304
rect 18831 6273 18843 6276
rect 18785 6267 18843 6273
rect 19058 6264 19064 6276
rect 19116 6304 19122 6316
rect 19260 6304 19288 6335
rect 19116 6276 19288 6304
rect 19720 6304 19748 6403
rect 21266 6400 21272 6412
rect 21324 6440 21330 6452
rect 21545 6443 21603 6449
rect 21545 6440 21557 6443
rect 21324 6412 21557 6440
rect 21324 6400 21330 6412
rect 21545 6409 21557 6412
rect 21591 6409 21603 6443
rect 21545 6403 21603 6409
rect 22005 6443 22063 6449
rect 22005 6409 22017 6443
rect 22051 6440 22063 6443
rect 23198 6440 23204 6452
rect 22051 6412 23204 6440
rect 22051 6409 22063 6412
rect 22005 6403 22063 6409
rect 21082 6332 21088 6384
rect 21140 6372 21146 6384
rect 22020 6372 22048 6403
rect 23198 6400 23204 6412
rect 23256 6400 23262 6452
rect 23474 6440 23480 6452
rect 23435 6412 23480 6440
rect 23474 6400 23480 6412
rect 23532 6400 23538 6452
rect 25038 6400 25044 6452
rect 25096 6440 25102 6452
rect 25501 6443 25559 6449
rect 25501 6440 25513 6443
rect 25096 6412 25513 6440
rect 25096 6400 25102 6412
rect 25501 6409 25513 6412
rect 25547 6409 25559 6443
rect 25501 6403 25559 6409
rect 21140 6344 22048 6372
rect 23109 6375 23167 6381
rect 21140 6332 21146 6344
rect 23109 6341 23121 6375
rect 23155 6372 23167 6375
rect 23382 6372 23388 6384
rect 23155 6344 23388 6372
rect 23155 6341 23167 6344
rect 23109 6335 23167 6341
rect 19720 6276 20024 6304
rect 19116 6264 19122 6276
rect 10778 6236 10784 6248
rect 10244 6208 10784 6236
rect 10137 6199 10195 6205
rect 10778 6196 10784 6208
rect 10836 6196 10842 6248
rect 13262 6196 13268 6248
rect 13320 6236 13326 6248
rect 13449 6239 13507 6245
rect 13449 6236 13461 6239
rect 13320 6208 13461 6236
rect 13320 6196 13326 6208
rect 13449 6205 13461 6208
rect 13495 6205 13507 6239
rect 13449 6199 13507 6205
rect 13538 6196 13544 6248
rect 13596 6236 13602 6248
rect 13705 6239 13763 6245
rect 13705 6236 13717 6239
rect 13596 6208 13717 6236
rect 13596 6196 13602 6208
rect 13705 6205 13717 6208
rect 13751 6205 13763 6239
rect 13705 6199 13763 6205
rect 16206 6196 16212 6248
rect 16264 6236 16270 6248
rect 16761 6239 16819 6245
rect 16761 6236 16773 6239
rect 16264 6208 16773 6236
rect 16264 6196 16270 6208
rect 16761 6205 16773 6208
rect 16807 6205 16819 6239
rect 16761 6199 16819 6205
rect 17586 6196 17592 6248
rect 17644 6236 17650 6248
rect 18322 6236 18328 6248
rect 17644 6208 18328 6236
rect 17644 6196 17650 6208
rect 18322 6196 18328 6208
rect 18380 6236 18386 6248
rect 18601 6239 18659 6245
rect 18601 6236 18613 6239
rect 18380 6208 18613 6236
rect 18380 6196 18386 6208
rect 18601 6205 18613 6208
rect 18647 6205 18659 6239
rect 18601 6199 18659 6205
rect 18693 6239 18751 6245
rect 18693 6205 18705 6239
rect 18739 6236 18751 6239
rect 19242 6236 19248 6248
rect 18739 6208 19248 6236
rect 18739 6205 18751 6208
rect 18693 6199 18751 6205
rect 19242 6196 19248 6208
rect 19300 6196 19306 6248
rect 19889 6239 19947 6245
rect 19889 6205 19901 6239
rect 19935 6205 19947 6239
rect 19996 6236 20024 6276
rect 20145 6239 20203 6245
rect 20145 6236 20157 6239
rect 19996 6208 20157 6236
rect 19889 6199 19947 6205
rect 20145 6205 20157 6208
rect 20191 6205 20203 6239
rect 20145 6199 20203 6205
rect 22465 6239 22523 6245
rect 22465 6205 22477 6239
rect 22511 6236 22523 6239
rect 23124 6236 23152 6335
rect 23382 6332 23388 6344
rect 23440 6332 23446 6384
rect 23198 6264 23204 6316
rect 23256 6304 23262 6316
rect 23845 6307 23903 6313
rect 23845 6304 23857 6307
rect 23256 6276 23857 6304
rect 23256 6264 23262 6276
rect 23845 6273 23857 6276
rect 23891 6273 23903 6307
rect 23845 6267 23903 6273
rect 22511 6208 23152 6236
rect 24112 6239 24170 6245
rect 22511 6205 22523 6208
rect 22465 6199 22523 6205
rect 24112 6205 24124 6239
rect 24158 6236 24170 6239
rect 25038 6236 25044 6248
rect 24158 6208 25044 6236
rect 24158 6205 24170 6208
rect 24112 6199 24170 6205
rect 9033 6171 9091 6177
rect 9033 6137 9045 6171
rect 9079 6168 9091 6171
rect 10404 6171 10462 6177
rect 9079 6140 10180 6168
rect 9079 6137 9091 6140
rect 9033 6131 9091 6137
rect 10152 6112 10180 6140
rect 10404 6137 10416 6171
rect 10450 6168 10462 6171
rect 12437 6171 12495 6177
rect 10450 6140 11836 6168
rect 10450 6137 10462 6140
rect 10404 6131 10462 6137
rect 11808 6112 11836 6140
rect 12437 6137 12449 6171
rect 12483 6168 12495 6171
rect 19904 6168 19932 6199
rect 25038 6196 25044 6208
rect 25096 6196 25102 6248
rect 19978 6168 19984 6180
rect 12483 6140 13676 6168
rect 19904 6140 19984 6168
rect 12483 6137 12495 6140
rect 12437 6131 12495 6137
rect 10134 6060 10140 6112
rect 10192 6060 10198 6112
rect 11790 6100 11796 6112
rect 11751 6072 11796 6100
rect 11790 6060 11796 6072
rect 11848 6060 11854 6112
rect 12989 6103 13047 6109
rect 12989 6069 13001 6103
rect 13035 6100 13047 6103
rect 13262 6100 13268 6112
rect 13035 6072 13268 6100
rect 13035 6069 13047 6072
rect 12989 6063 13047 6069
rect 13262 6060 13268 6072
rect 13320 6060 13326 6112
rect 13648 6100 13676 6140
rect 19978 6128 19984 6140
rect 20036 6128 20042 6180
rect 13722 6100 13728 6112
rect 13648 6072 13728 6100
rect 13722 6060 13728 6072
rect 13780 6060 13786 6112
rect 15565 6103 15623 6109
rect 15565 6069 15577 6103
rect 15611 6100 15623 6103
rect 15930 6100 15936 6112
rect 15611 6072 15936 6100
rect 15611 6069 15623 6072
rect 15565 6063 15623 6069
rect 15930 6060 15936 6072
rect 15988 6060 15994 6112
rect 16850 6100 16856 6112
rect 16811 6072 16856 6100
rect 16850 6060 16856 6072
rect 16908 6060 16914 6112
rect 22646 6100 22652 6112
rect 22607 6072 22652 6100
rect 22646 6060 22652 6072
rect 22704 6060 22710 6112
rect 25222 6100 25228 6112
rect 25183 6072 25228 6100
rect 25222 6060 25228 6072
rect 25280 6060 25286 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 8570 5896 8576 5908
rect 8531 5868 8576 5896
rect 8570 5856 8576 5868
rect 8628 5856 8634 5908
rect 10134 5856 10140 5908
rect 10192 5896 10198 5908
rect 10229 5899 10287 5905
rect 10229 5896 10241 5899
rect 10192 5868 10241 5896
rect 10192 5856 10198 5868
rect 10229 5865 10241 5868
rect 10275 5865 10287 5899
rect 10229 5859 10287 5865
rect 13538 5856 13544 5908
rect 13596 5896 13602 5908
rect 13633 5899 13691 5905
rect 13633 5896 13645 5899
rect 13596 5868 13645 5896
rect 13596 5856 13602 5868
rect 13633 5865 13645 5868
rect 13679 5865 13691 5899
rect 14090 5896 14096 5908
rect 14051 5868 14096 5896
rect 13633 5859 13691 5865
rect 14090 5856 14096 5868
rect 14148 5856 14154 5908
rect 15562 5856 15568 5908
rect 15620 5896 15626 5908
rect 15841 5899 15899 5905
rect 15841 5896 15853 5899
rect 15620 5868 15853 5896
rect 15620 5856 15626 5868
rect 15841 5865 15853 5868
rect 15887 5865 15899 5899
rect 17402 5896 17408 5908
rect 17363 5868 17408 5896
rect 15841 5859 15899 5865
rect 17402 5856 17408 5868
rect 17460 5856 17466 5908
rect 17954 5856 17960 5908
rect 18012 5896 18018 5908
rect 18049 5899 18107 5905
rect 18049 5896 18061 5899
rect 18012 5868 18061 5896
rect 18012 5856 18018 5868
rect 18049 5865 18061 5868
rect 18095 5896 18107 5899
rect 18141 5899 18199 5905
rect 18141 5896 18153 5899
rect 18095 5868 18153 5896
rect 18095 5865 18107 5868
rect 18049 5859 18107 5865
rect 18141 5865 18153 5868
rect 18187 5865 18199 5899
rect 18322 5896 18328 5908
rect 18283 5868 18328 5896
rect 18141 5859 18199 5865
rect 18322 5856 18328 5868
rect 18380 5856 18386 5908
rect 19978 5856 19984 5908
rect 20036 5896 20042 5908
rect 20349 5899 20407 5905
rect 20349 5896 20361 5899
rect 20036 5868 20361 5896
rect 20036 5856 20042 5868
rect 20349 5865 20361 5868
rect 20395 5896 20407 5899
rect 21082 5896 21088 5908
rect 20395 5868 21088 5896
rect 20395 5865 20407 5868
rect 20349 5859 20407 5865
rect 21082 5856 21088 5868
rect 21140 5856 21146 5908
rect 23198 5856 23204 5908
rect 23256 5896 23262 5908
rect 23293 5899 23351 5905
rect 23293 5896 23305 5899
rect 23256 5868 23305 5896
rect 23256 5856 23262 5868
rect 23293 5865 23305 5868
rect 23339 5896 23351 5899
rect 23661 5899 23719 5905
rect 23661 5896 23673 5899
rect 23339 5868 23673 5896
rect 23339 5865 23351 5868
rect 23293 5859 23351 5865
rect 12434 5788 12440 5840
rect 12492 5837 12498 5840
rect 12492 5831 12556 5837
rect 12492 5797 12510 5831
rect 12544 5797 12556 5831
rect 12492 5791 12556 5797
rect 17865 5831 17923 5837
rect 17865 5797 17877 5831
rect 17911 5828 17923 5831
rect 19242 5828 19248 5840
rect 17911 5800 19248 5828
rect 17911 5797 17923 5800
rect 17865 5791 17923 5797
rect 12492 5788 12498 5791
rect 19242 5788 19248 5800
rect 19300 5788 19306 5840
rect 9766 5720 9772 5772
rect 9824 5760 9830 5772
rect 10597 5763 10655 5769
rect 10597 5760 10609 5763
rect 9824 5732 10609 5760
rect 9824 5720 9830 5732
rect 10597 5729 10609 5732
rect 10643 5729 10655 5763
rect 16206 5760 16212 5772
rect 16167 5732 16212 5760
rect 10597 5723 10655 5729
rect 16206 5720 16212 5732
rect 16264 5720 16270 5772
rect 18230 5720 18236 5772
rect 18288 5760 18294 5772
rect 18693 5763 18751 5769
rect 18693 5760 18705 5763
rect 18288 5732 18705 5760
rect 18288 5720 18294 5732
rect 18693 5729 18705 5732
rect 18739 5760 18751 5763
rect 19518 5760 19524 5772
rect 18739 5732 19524 5760
rect 18739 5729 18751 5732
rect 18693 5723 18751 5729
rect 19518 5720 19524 5732
rect 19576 5720 19582 5772
rect 20898 5760 20904 5772
rect 20859 5732 20904 5760
rect 20898 5720 20904 5732
rect 20956 5720 20962 5772
rect 22002 5720 22008 5772
rect 22060 5760 22066 5772
rect 22649 5763 22707 5769
rect 22649 5760 22661 5763
rect 22060 5732 22661 5760
rect 22060 5720 22066 5732
rect 22649 5729 22661 5732
rect 22695 5729 22707 5763
rect 23400 5760 23428 5868
rect 23661 5865 23673 5868
rect 23707 5865 23719 5899
rect 23661 5859 23719 5865
rect 23474 5788 23480 5840
rect 23532 5828 23538 5840
rect 24112 5831 24170 5837
rect 24112 5828 24124 5831
rect 23532 5800 24124 5828
rect 23532 5788 23538 5800
rect 24112 5797 24124 5800
rect 24158 5828 24170 5831
rect 25222 5828 25228 5840
rect 24158 5800 25228 5828
rect 24158 5797 24170 5800
rect 24112 5791 24170 5797
rect 25222 5788 25228 5800
rect 25280 5788 25286 5840
rect 23845 5763 23903 5769
rect 23845 5760 23857 5763
rect 23400 5732 23857 5760
rect 22649 5723 22707 5729
rect 23845 5729 23857 5732
rect 23891 5760 23903 5763
rect 25501 5763 25559 5769
rect 25501 5760 25513 5763
rect 23891 5732 25513 5760
rect 23891 5729 23903 5732
rect 23845 5723 23903 5729
rect 25501 5729 25513 5732
rect 25547 5729 25559 5763
rect 25501 5723 25559 5729
rect 10045 5695 10103 5701
rect 10045 5661 10057 5695
rect 10091 5692 10103 5695
rect 10226 5692 10232 5704
rect 10091 5664 10232 5692
rect 10091 5661 10103 5664
rect 10045 5655 10103 5661
rect 10226 5652 10232 5664
rect 10284 5652 10290 5704
rect 10689 5695 10747 5701
rect 10689 5661 10701 5695
rect 10735 5692 10747 5695
rect 10778 5692 10784 5704
rect 10735 5664 10784 5692
rect 10735 5661 10747 5664
rect 10689 5655 10747 5661
rect 9674 5584 9680 5636
rect 9732 5624 9738 5636
rect 10704 5624 10732 5655
rect 10778 5652 10784 5664
rect 10836 5652 10842 5704
rect 10873 5695 10931 5701
rect 10873 5661 10885 5695
rect 10919 5692 10931 5695
rect 10962 5692 10968 5704
rect 10919 5664 10968 5692
rect 10919 5661 10931 5664
rect 10873 5655 10931 5661
rect 10962 5652 10968 5664
rect 11020 5692 11026 5704
rect 11790 5692 11796 5704
rect 11020 5664 11796 5692
rect 11020 5652 11026 5664
rect 11790 5652 11796 5664
rect 11848 5652 11854 5704
rect 12253 5695 12311 5701
rect 12253 5661 12265 5695
rect 12299 5661 12311 5695
rect 12253 5655 12311 5661
rect 12268 5624 12296 5655
rect 15746 5652 15752 5704
rect 15804 5692 15810 5704
rect 16301 5695 16359 5701
rect 16301 5692 16313 5695
rect 15804 5664 16313 5692
rect 15804 5652 15810 5664
rect 16301 5661 16313 5664
rect 16347 5661 16359 5695
rect 16301 5655 16359 5661
rect 16393 5695 16451 5701
rect 16393 5661 16405 5695
rect 16439 5661 16451 5695
rect 16393 5655 16451 5661
rect 16408 5624 16436 5655
rect 18138 5652 18144 5704
rect 18196 5692 18202 5704
rect 18785 5695 18843 5701
rect 18785 5692 18797 5695
rect 18196 5664 18797 5692
rect 18196 5652 18202 5664
rect 18785 5661 18797 5664
rect 18831 5661 18843 5695
rect 18785 5655 18843 5661
rect 18877 5695 18935 5701
rect 18877 5661 18889 5695
rect 18923 5661 18935 5695
rect 22738 5692 22744 5704
rect 22699 5664 22744 5692
rect 18877 5655 18935 5661
rect 9732 5596 10732 5624
rect 11532 5596 12296 5624
rect 15672 5596 16436 5624
rect 18049 5627 18107 5633
rect 9732 5584 9738 5596
rect 9493 5559 9551 5565
rect 9493 5525 9505 5559
rect 9539 5556 9551 5559
rect 9950 5556 9956 5568
rect 9539 5528 9956 5556
rect 9539 5525 9551 5528
rect 9493 5519 9551 5525
rect 9950 5516 9956 5528
rect 10008 5516 10014 5568
rect 11330 5516 11336 5568
rect 11388 5556 11394 5568
rect 11532 5565 11560 5596
rect 11517 5559 11575 5565
rect 11517 5556 11529 5559
rect 11388 5528 11529 5556
rect 11388 5516 11394 5528
rect 11517 5525 11529 5528
rect 11563 5525 11575 5559
rect 11517 5519 11575 5525
rect 15562 5516 15568 5568
rect 15620 5556 15626 5568
rect 15672 5565 15700 5596
rect 18049 5593 18061 5627
rect 18095 5624 18107 5627
rect 18598 5624 18604 5636
rect 18095 5596 18604 5624
rect 18095 5593 18107 5596
rect 18049 5587 18107 5593
rect 18598 5584 18604 5596
rect 18656 5624 18662 5636
rect 18892 5624 18920 5655
rect 22738 5652 22744 5664
rect 22796 5652 22802 5704
rect 22925 5695 22983 5701
rect 22925 5661 22937 5695
rect 22971 5692 22983 5695
rect 23474 5692 23480 5704
rect 22971 5664 23480 5692
rect 22971 5661 22983 5664
rect 22925 5655 22983 5661
rect 23474 5652 23480 5664
rect 23532 5652 23538 5704
rect 18656 5596 18920 5624
rect 22281 5627 22339 5633
rect 18656 5584 18662 5596
rect 22281 5593 22293 5627
rect 22327 5624 22339 5627
rect 23382 5624 23388 5636
rect 22327 5596 23388 5624
rect 22327 5593 22339 5596
rect 22281 5587 22339 5593
rect 23382 5584 23388 5596
rect 23440 5584 23446 5636
rect 15657 5559 15715 5565
rect 15657 5556 15669 5559
rect 15620 5528 15669 5556
rect 15620 5516 15626 5528
rect 15657 5525 15669 5528
rect 15703 5525 15715 5559
rect 15657 5519 15715 5525
rect 16850 5516 16856 5568
rect 16908 5556 16914 5568
rect 16945 5559 17003 5565
rect 16945 5556 16957 5559
rect 16908 5528 16957 5556
rect 16908 5516 16914 5528
rect 16945 5525 16957 5528
rect 16991 5556 17003 5559
rect 17862 5556 17868 5568
rect 16991 5528 17868 5556
rect 16991 5525 17003 5528
rect 16945 5519 17003 5525
rect 17862 5516 17868 5528
rect 17920 5516 17926 5568
rect 19981 5559 20039 5565
rect 19981 5525 19993 5559
rect 20027 5556 20039 5559
rect 20346 5556 20352 5568
rect 20027 5528 20352 5556
rect 20027 5525 20039 5528
rect 19981 5519 20039 5525
rect 20346 5516 20352 5528
rect 20404 5516 20410 5568
rect 21082 5556 21088 5568
rect 21043 5528 21088 5556
rect 21082 5516 21088 5528
rect 21140 5516 21146 5568
rect 22094 5516 22100 5568
rect 22152 5556 22158 5568
rect 22152 5528 22197 5556
rect 22152 5516 22158 5528
rect 24854 5516 24860 5568
rect 24912 5556 24918 5568
rect 25225 5559 25283 5565
rect 25225 5556 25237 5559
rect 24912 5528 25237 5556
rect 24912 5516 24918 5528
rect 25225 5525 25237 5528
rect 25271 5525 25283 5559
rect 25225 5519 25283 5525
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 9493 5355 9551 5361
rect 9493 5321 9505 5355
rect 9539 5352 9551 5355
rect 9582 5352 9588 5364
rect 9539 5324 9588 5352
rect 9539 5321 9551 5324
rect 9493 5315 9551 5321
rect 9582 5312 9588 5324
rect 9640 5312 9646 5364
rect 11333 5355 11391 5361
rect 11333 5321 11345 5355
rect 11379 5352 11391 5355
rect 11790 5352 11796 5364
rect 11379 5324 11796 5352
rect 11379 5321 11391 5324
rect 11333 5315 11391 5321
rect 11790 5312 11796 5324
rect 11848 5312 11854 5364
rect 14642 5352 14648 5364
rect 14603 5324 14648 5352
rect 14642 5312 14648 5324
rect 14700 5312 14706 5364
rect 15746 5352 15752 5364
rect 15707 5324 15752 5352
rect 15746 5312 15752 5324
rect 15804 5312 15810 5364
rect 17954 5312 17960 5364
rect 18012 5352 18018 5364
rect 18325 5355 18383 5361
rect 18325 5352 18337 5355
rect 18012 5324 18337 5352
rect 18012 5312 18018 5324
rect 18325 5321 18337 5324
rect 18371 5321 18383 5355
rect 18325 5315 18383 5321
rect 19334 5312 19340 5364
rect 19392 5352 19398 5364
rect 19889 5355 19947 5361
rect 19889 5352 19901 5355
rect 19392 5324 19901 5352
rect 19392 5312 19398 5324
rect 19889 5321 19901 5324
rect 19935 5321 19947 5355
rect 20898 5352 20904 5364
rect 20859 5324 20904 5352
rect 19889 5315 19947 5321
rect 20898 5312 20904 5324
rect 20956 5312 20962 5364
rect 22002 5352 22008 5364
rect 21963 5324 22008 5352
rect 22002 5312 22008 5324
rect 22060 5312 22066 5364
rect 23109 5355 23167 5361
rect 23109 5321 23121 5355
rect 23155 5352 23167 5355
rect 23474 5352 23480 5364
rect 23155 5324 23480 5352
rect 23155 5321 23167 5324
rect 23109 5315 23167 5321
rect 23474 5312 23480 5324
rect 23532 5312 23538 5364
rect 23842 5312 23848 5364
rect 23900 5352 23906 5364
rect 24029 5355 24087 5361
rect 24029 5352 24041 5355
rect 23900 5324 24041 5352
rect 23900 5312 23906 5324
rect 24029 5321 24041 5324
rect 24075 5321 24087 5355
rect 24029 5315 24087 5321
rect 14458 5244 14464 5296
rect 14516 5284 14522 5296
rect 15565 5287 15623 5293
rect 15565 5284 15577 5287
rect 14516 5256 15577 5284
rect 14516 5244 14522 5256
rect 15565 5253 15577 5256
rect 15611 5284 15623 5287
rect 15611 5256 16160 5284
rect 15611 5253 15623 5256
rect 15565 5247 15623 5253
rect 13262 5216 13268 5228
rect 13223 5188 13268 5216
rect 13262 5176 13268 5188
rect 13320 5176 13326 5228
rect 14366 5176 14372 5228
rect 14424 5176 14430 5228
rect 9950 5148 9956 5160
rect 9863 5120 9956 5148
rect 9950 5108 9956 5120
rect 10008 5108 10014 5160
rect 10226 5157 10232 5160
rect 10220 5148 10232 5157
rect 10187 5120 10232 5148
rect 10220 5111 10232 5120
rect 10226 5108 10232 5111
rect 10284 5108 10290 5160
rect 11330 5108 11336 5160
rect 11388 5148 11394 5160
rect 12161 5151 12219 5157
rect 12161 5148 12173 5151
rect 11388 5120 12173 5148
rect 11388 5108 11394 5120
rect 12161 5117 12173 5120
rect 12207 5148 12219 5151
rect 12342 5148 12348 5160
rect 12207 5120 12348 5148
rect 12207 5117 12219 5120
rect 12161 5111 12219 5117
rect 12342 5108 12348 5120
rect 12400 5108 12406 5160
rect 14384 5148 14412 5176
rect 14458 5148 14464 5160
rect 14384 5120 14464 5148
rect 14458 5108 14464 5120
rect 14516 5108 14522 5160
rect 16132 5157 16160 5256
rect 16206 5244 16212 5296
rect 16264 5284 16270 5296
rect 16853 5287 16911 5293
rect 16853 5284 16865 5287
rect 16264 5256 16865 5284
rect 16264 5244 16270 5256
rect 16853 5253 16865 5256
rect 16899 5284 16911 5287
rect 18046 5284 18052 5296
rect 16899 5256 18052 5284
rect 16899 5253 16911 5256
rect 16853 5247 16911 5253
rect 18046 5244 18052 5256
rect 18104 5244 18110 5296
rect 23937 5287 23995 5293
rect 23937 5253 23949 5287
rect 23983 5284 23995 5287
rect 23983 5256 24716 5284
rect 23983 5253 23995 5256
rect 23937 5247 23995 5253
rect 16390 5216 16396 5228
rect 16351 5188 16396 5216
rect 16390 5176 16396 5188
rect 16448 5176 16454 5228
rect 18598 5176 18604 5228
rect 18656 5216 18662 5228
rect 18877 5219 18935 5225
rect 18877 5216 18889 5219
rect 18656 5188 18889 5216
rect 18656 5176 18662 5188
rect 18877 5185 18889 5188
rect 18923 5216 18935 5219
rect 20441 5219 20499 5225
rect 20441 5216 20453 5219
rect 18923 5188 20453 5216
rect 18923 5185 18935 5188
rect 18877 5179 18935 5185
rect 20441 5185 20453 5188
rect 20487 5185 20499 5219
rect 20441 5179 20499 5185
rect 21545 5219 21603 5225
rect 21545 5185 21557 5219
rect 21591 5216 21603 5219
rect 22646 5216 22652 5228
rect 21591 5188 22652 5216
rect 21591 5185 21603 5188
rect 21545 5179 21603 5185
rect 22646 5176 22652 5188
rect 22704 5176 22710 5228
rect 23474 5176 23480 5228
rect 23532 5216 23538 5228
rect 24688 5225 24716 5256
rect 24489 5219 24547 5225
rect 24489 5216 24501 5219
rect 23532 5188 24501 5216
rect 23532 5176 23538 5188
rect 24489 5185 24501 5188
rect 24535 5185 24547 5219
rect 24489 5179 24547 5185
rect 24673 5219 24731 5225
rect 24673 5185 24685 5219
rect 24719 5216 24731 5219
rect 24762 5216 24768 5228
rect 24719 5188 24768 5216
rect 24719 5185 24731 5188
rect 24673 5179 24731 5185
rect 16117 5151 16175 5157
rect 16117 5117 16129 5151
rect 16163 5117 16175 5151
rect 16117 5111 16175 5117
rect 17678 5108 17684 5160
rect 17736 5148 17742 5160
rect 17773 5151 17831 5157
rect 17773 5148 17785 5151
rect 17736 5120 17785 5148
rect 17736 5108 17742 5120
rect 17773 5117 17785 5120
rect 17819 5148 17831 5151
rect 18693 5151 18751 5157
rect 18693 5148 18705 5151
rect 17819 5120 18705 5148
rect 17819 5117 17831 5120
rect 17773 5111 17831 5117
rect 18693 5117 18705 5120
rect 18739 5117 18751 5151
rect 18693 5111 18751 5117
rect 18785 5151 18843 5157
rect 18785 5117 18797 5151
rect 18831 5148 18843 5151
rect 18966 5148 18972 5160
rect 18831 5120 18972 5148
rect 18831 5117 18843 5120
rect 18785 5111 18843 5117
rect 18966 5108 18972 5120
rect 19024 5108 19030 5160
rect 19429 5151 19487 5157
rect 19429 5117 19441 5151
rect 19475 5148 19487 5151
rect 19518 5148 19524 5160
rect 19475 5120 19524 5148
rect 19475 5117 19487 5120
rect 19429 5111 19487 5117
rect 19518 5108 19524 5120
rect 19576 5148 19582 5160
rect 22094 5148 22100 5160
rect 19576 5120 22100 5148
rect 19576 5108 19582 5120
rect 22094 5108 22100 5120
rect 22152 5148 22158 5160
rect 22373 5151 22431 5157
rect 22373 5148 22385 5151
rect 22152 5120 22385 5148
rect 22152 5108 22158 5120
rect 22373 5117 22385 5120
rect 22419 5148 22431 5151
rect 23382 5148 23388 5160
rect 22419 5120 23388 5148
rect 22419 5117 22431 5120
rect 22373 5111 22431 5117
rect 23382 5108 23388 5120
rect 23440 5108 23446 5160
rect 24504 5148 24532 5179
rect 24762 5176 24768 5188
rect 24820 5176 24826 5228
rect 25041 5151 25099 5157
rect 25041 5148 25053 5151
rect 24504 5120 25053 5148
rect 25041 5117 25053 5120
rect 25087 5117 25099 5151
rect 25041 5111 25099 5117
rect 9968 5080 9996 5108
rect 11701 5083 11759 5089
rect 11701 5080 11713 5083
rect 9968 5052 11713 5080
rect 11701 5049 11713 5052
rect 11747 5080 11759 5083
rect 12526 5080 12532 5092
rect 11747 5052 12532 5080
rect 11747 5049 11759 5052
rect 11701 5043 11759 5049
rect 12526 5040 12532 5052
rect 12584 5040 12590 5092
rect 13173 5083 13231 5089
rect 13173 5049 13185 5083
rect 13219 5080 13231 5083
rect 13510 5083 13568 5089
rect 13510 5080 13522 5083
rect 13219 5052 13522 5080
rect 13219 5049 13231 5052
rect 13173 5043 13231 5049
rect 13510 5049 13522 5052
rect 13556 5080 13568 5083
rect 14366 5080 14372 5092
rect 13556 5052 14372 5080
rect 13556 5049 13568 5052
rect 13510 5043 13568 5049
rect 14366 5040 14372 5052
rect 14424 5040 14430 5092
rect 18138 5080 18144 5092
rect 17420 5052 18144 5080
rect 7929 5015 7987 5021
rect 7929 4981 7941 5015
rect 7975 5012 7987 5015
rect 8478 5012 8484 5024
rect 7975 4984 8484 5012
rect 7975 4981 7987 4984
rect 7929 4975 7987 4981
rect 8478 4972 8484 4984
rect 8536 4972 8542 5024
rect 8846 5012 8852 5024
rect 8807 4984 8852 5012
rect 8846 4972 8852 4984
rect 8904 4972 8910 5024
rect 8941 5015 8999 5021
rect 8941 4981 8953 5015
rect 8987 5012 8999 5015
rect 9582 5012 9588 5024
rect 8987 4984 9588 5012
rect 8987 4981 8999 4984
rect 8941 4975 8999 4981
rect 9582 4972 9588 4984
rect 9640 4972 9646 5024
rect 9766 5012 9772 5024
rect 9727 4984 9772 5012
rect 9766 4972 9772 4984
rect 9824 4972 9830 5024
rect 12434 4972 12440 5024
rect 12492 5012 12498 5024
rect 12621 5015 12679 5021
rect 12621 5012 12633 5015
rect 12492 4984 12633 5012
rect 12492 4972 12498 4984
rect 12621 4981 12633 4984
rect 12667 4981 12679 5015
rect 12621 4975 12679 4981
rect 15289 5015 15347 5021
rect 15289 4981 15301 5015
rect 15335 5012 15347 5015
rect 16114 5012 16120 5024
rect 15335 4984 16120 5012
rect 15335 4981 15347 4984
rect 15289 4975 15347 4981
rect 16114 4972 16120 4984
rect 16172 5012 16178 5024
rect 16209 5015 16267 5021
rect 16209 5012 16221 5015
rect 16172 4984 16221 5012
rect 16172 4972 16178 4984
rect 16209 4981 16221 4984
rect 16255 4981 16267 5015
rect 16209 4975 16267 4981
rect 16942 4972 16948 5024
rect 17000 5012 17006 5024
rect 17420 5021 17448 5052
rect 18138 5040 18144 5052
rect 18196 5040 18202 5092
rect 19797 5083 19855 5089
rect 19797 5049 19809 5083
rect 19843 5080 19855 5083
rect 20257 5083 20315 5089
rect 20257 5080 20269 5083
rect 19843 5052 20269 5080
rect 19843 5049 19855 5052
rect 19797 5043 19855 5049
rect 20257 5049 20269 5052
rect 20303 5080 20315 5083
rect 20438 5080 20444 5092
rect 20303 5052 20444 5080
rect 20303 5049 20315 5052
rect 20257 5043 20315 5049
rect 20438 5040 20444 5052
rect 20496 5040 20502 5092
rect 21818 5080 21824 5092
rect 21779 5052 21824 5080
rect 21818 5040 21824 5052
rect 21876 5040 21882 5092
rect 23658 5040 23664 5092
rect 23716 5080 23722 5092
rect 24397 5083 24455 5089
rect 24397 5080 24409 5083
rect 23716 5052 24409 5080
rect 23716 5040 23722 5052
rect 24397 5049 24409 5052
rect 24443 5080 24455 5083
rect 25409 5083 25467 5089
rect 25409 5080 25421 5083
rect 24443 5052 25421 5080
rect 24443 5049 24455 5052
rect 24397 5043 24455 5049
rect 25409 5049 25421 5052
rect 25455 5049 25467 5083
rect 25409 5043 25467 5049
rect 17405 5015 17463 5021
rect 17405 5012 17417 5015
rect 17000 4984 17417 5012
rect 17000 4972 17006 4984
rect 17405 4981 17417 4984
rect 17451 4981 17463 5015
rect 20346 5012 20352 5024
rect 20307 4984 20352 5012
rect 17405 4975 17463 4981
rect 20346 4972 20352 4984
rect 20404 4972 20410 5024
rect 21836 5012 21864 5040
rect 22465 5015 22523 5021
rect 22465 5012 22477 5015
rect 21836 4984 22477 5012
rect 22465 4981 22477 4984
rect 22511 5012 22523 5015
rect 22922 5012 22928 5024
rect 22511 4984 22928 5012
rect 22511 4981 22523 4984
rect 22465 4975 22523 4981
rect 22922 4972 22928 4984
rect 22980 4972 22986 5024
rect 25590 5012 25596 5024
rect 25551 4984 25596 5012
rect 25590 4972 25596 4984
rect 25648 4972 25654 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 8662 4808 8668 4820
rect 8623 4780 8668 4808
rect 8662 4768 8668 4780
rect 8720 4768 8726 4820
rect 9861 4811 9919 4817
rect 9861 4777 9873 4811
rect 9907 4808 9919 4811
rect 10686 4808 10692 4820
rect 9907 4780 10692 4808
rect 9907 4777 9919 4780
rect 9861 4771 9919 4777
rect 10686 4768 10692 4780
rect 10744 4768 10750 4820
rect 10962 4808 10968 4820
rect 10923 4780 10968 4808
rect 10962 4768 10968 4780
rect 11020 4768 11026 4820
rect 11422 4808 11428 4820
rect 11383 4780 11428 4808
rect 11422 4768 11428 4780
rect 11480 4768 11486 4820
rect 12342 4768 12348 4820
rect 12400 4808 12406 4820
rect 12805 4811 12863 4817
rect 12805 4808 12817 4811
rect 12400 4780 12817 4808
rect 12400 4768 12406 4780
rect 12805 4777 12817 4780
rect 12851 4808 12863 4811
rect 13262 4808 13268 4820
rect 12851 4780 13268 4808
rect 12851 4777 12863 4780
rect 12805 4771 12863 4777
rect 13262 4768 13268 4780
rect 13320 4808 13326 4820
rect 14182 4808 14188 4820
rect 13320 4780 14188 4808
rect 13320 4768 13326 4780
rect 14182 4768 14188 4780
rect 14240 4768 14246 4820
rect 14366 4808 14372 4820
rect 14327 4780 14372 4808
rect 14366 4768 14372 4780
rect 14424 4768 14430 4820
rect 15105 4811 15163 4817
rect 15105 4777 15117 4811
rect 15151 4808 15163 4811
rect 15746 4808 15752 4820
rect 15151 4780 15752 4808
rect 15151 4777 15163 4780
rect 15105 4771 15163 4777
rect 15746 4768 15752 4780
rect 15804 4768 15810 4820
rect 16390 4768 16396 4820
rect 16448 4808 16454 4820
rect 17129 4811 17187 4817
rect 17129 4808 17141 4811
rect 16448 4780 17141 4808
rect 16448 4768 16454 4780
rect 17129 4777 17141 4780
rect 17175 4777 17187 4811
rect 17129 4771 17187 4777
rect 18325 4811 18383 4817
rect 18325 4777 18337 4811
rect 18371 4808 18383 4811
rect 18966 4808 18972 4820
rect 18371 4780 18972 4808
rect 18371 4777 18383 4780
rect 18325 4771 18383 4777
rect 18966 4768 18972 4780
rect 19024 4768 19030 4820
rect 21266 4768 21272 4820
rect 21324 4808 21330 4820
rect 21545 4811 21603 4817
rect 21545 4808 21557 4811
rect 21324 4780 21557 4808
rect 21324 4768 21330 4780
rect 21545 4777 21557 4780
rect 21591 4777 21603 4811
rect 22002 4808 22008 4820
rect 21963 4780 22008 4808
rect 21545 4771 21603 4777
rect 22002 4768 22008 4780
rect 22060 4768 22066 4820
rect 22097 4811 22155 4817
rect 22097 4777 22109 4811
rect 22143 4808 22155 4811
rect 24121 4811 24179 4817
rect 24121 4808 24133 4811
rect 22143 4780 24133 4808
rect 22143 4777 22155 4780
rect 22097 4771 22155 4777
rect 24121 4777 24133 4780
rect 24167 4808 24179 4811
rect 25041 4811 25099 4817
rect 25041 4808 25053 4811
rect 24167 4780 25053 4808
rect 24167 4777 24179 4780
rect 24121 4771 24179 4777
rect 25041 4777 25053 4780
rect 25087 4777 25099 4811
rect 25406 4808 25412 4820
rect 25367 4780 25412 4808
rect 25041 4771 25099 4777
rect 25406 4768 25412 4780
rect 25464 4768 25470 4820
rect 9490 4700 9496 4752
rect 9548 4740 9554 4752
rect 10321 4743 10379 4749
rect 10321 4740 10333 4743
rect 9548 4712 10333 4740
rect 9548 4700 9554 4712
rect 10321 4709 10333 4712
rect 10367 4740 10379 4743
rect 11054 4740 11060 4752
rect 10367 4712 11060 4740
rect 10367 4709 10379 4712
rect 10321 4703 10379 4709
rect 11054 4700 11060 4712
rect 11112 4700 11118 4752
rect 15657 4743 15715 4749
rect 15657 4709 15669 4743
rect 15703 4740 15715 4743
rect 16408 4740 16436 4768
rect 15703 4712 16436 4740
rect 17957 4743 18015 4749
rect 15703 4709 15715 4712
rect 15657 4703 15715 4709
rect 17957 4709 17969 4743
rect 18003 4740 18015 4743
rect 18598 4740 18604 4752
rect 18003 4712 18604 4740
rect 18003 4709 18015 4712
rect 17957 4703 18015 4709
rect 18598 4700 18604 4712
rect 18656 4740 18662 4752
rect 20073 4743 20131 4749
rect 20073 4740 20085 4743
rect 18656 4712 20085 4740
rect 18656 4700 18662 4712
rect 20073 4709 20085 4712
rect 20119 4709 20131 4743
rect 22370 4740 22376 4752
rect 20073 4703 20131 4709
rect 21008 4712 22376 4740
rect 21008 4684 21036 4712
rect 22370 4700 22376 4712
rect 22428 4700 22434 4752
rect 22738 4700 22744 4752
rect 22796 4740 22802 4752
rect 23109 4743 23167 4749
rect 23109 4740 23121 4743
rect 22796 4712 23121 4740
rect 22796 4700 22802 4712
rect 23109 4709 23121 4712
rect 23155 4740 23167 4743
rect 23290 4740 23296 4752
rect 23155 4712 23296 4740
rect 23155 4709 23167 4712
rect 23109 4703 23167 4709
rect 23290 4700 23296 4712
rect 23348 4700 23354 4752
rect 23566 4700 23572 4752
rect 23624 4740 23630 4752
rect 23624 4712 23669 4740
rect 23624 4700 23630 4712
rect 23750 4700 23756 4752
rect 23808 4740 23814 4752
rect 24029 4743 24087 4749
rect 24029 4740 24041 4743
rect 23808 4712 24041 4740
rect 23808 4700 23814 4712
rect 24029 4709 24041 4712
rect 24075 4740 24087 4743
rect 24946 4740 24952 4752
rect 24075 4712 24952 4740
rect 24075 4709 24087 4712
rect 24029 4703 24087 4709
rect 24946 4700 24952 4712
rect 25004 4700 25010 4752
rect 8481 4675 8539 4681
rect 8481 4641 8493 4675
rect 8527 4672 8539 4675
rect 8754 4672 8760 4684
rect 8527 4644 8760 4672
rect 8527 4641 8539 4644
rect 8481 4635 8539 4641
rect 8754 4632 8760 4644
rect 8812 4632 8818 4684
rect 10134 4632 10140 4684
rect 10192 4672 10198 4684
rect 10229 4675 10287 4681
rect 10229 4672 10241 4675
rect 10192 4644 10241 4672
rect 10192 4632 10198 4644
rect 10229 4641 10241 4644
rect 10275 4641 10287 4675
rect 10229 4635 10287 4641
rect 11698 4632 11704 4684
rect 11756 4672 11762 4684
rect 11793 4675 11851 4681
rect 11793 4672 11805 4675
rect 11756 4644 11805 4672
rect 11756 4632 11762 4644
rect 11793 4641 11805 4644
rect 11839 4641 11851 4675
rect 11793 4635 11851 4641
rect 12802 4632 12808 4684
rect 12860 4672 12866 4684
rect 13245 4675 13303 4681
rect 13245 4672 13257 4675
rect 12860 4644 13257 4672
rect 12860 4632 12866 4644
rect 13245 4641 13257 4644
rect 13291 4672 13303 4675
rect 13538 4672 13544 4684
rect 13291 4644 13544 4672
rect 13291 4641 13303 4644
rect 13245 4635 13303 4641
rect 13538 4632 13544 4644
rect 13596 4632 13602 4684
rect 16022 4681 16028 4684
rect 16016 4672 16028 4681
rect 15983 4644 16028 4672
rect 16016 4635 16028 4644
rect 16022 4632 16028 4635
rect 16080 4632 16086 4684
rect 18322 4632 18328 4684
rect 18380 4672 18386 4684
rect 18684 4675 18742 4681
rect 18684 4672 18696 4675
rect 18380 4644 18696 4672
rect 18380 4632 18386 4644
rect 18684 4641 18696 4644
rect 18730 4672 18742 4675
rect 19242 4672 19248 4684
rect 18730 4644 19248 4672
rect 18730 4641 18742 4644
rect 18684 4635 18742 4641
rect 19242 4632 19248 4644
rect 19300 4632 19306 4684
rect 20990 4672 20996 4684
rect 20903 4644 20996 4672
rect 20990 4632 20996 4644
rect 21048 4632 21054 4684
rect 22278 4632 22284 4684
rect 22336 4672 22342 4684
rect 22465 4675 22523 4681
rect 22465 4672 22477 4675
rect 22336 4644 22477 4672
rect 22336 4632 22342 4644
rect 22465 4641 22477 4644
rect 22511 4641 22523 4675
rect 22465 4635 22523 4641
rect 7466 4604 7472 4616
rect 7427 4576 7472 4604
rect 7466 4564 7472 4576
rect 7524 4564 7530 4616
rect 10502 4604 10508 4616
rect 10463 4576 10508 4604
rect 10502 4564 10508 4576
rect 10560 4564 10566 4616
rect 11885 4607 11943 4613
rect 11885 4573 11897 4607
rect 11931 4573 11943 4607
rect 12066 4604 12072 4616
rect 12027 4576 12072 4604
rect 11885 4567 11943 4573
rect 9493 4539 9551 4545
rect 9493 4505 9505 4539
rect 9539 4536 9551 4539
rect 10520 4536 10548 4564
rect 9539 4508 10548 4536
rect 9539 4505 9551 4508
rect 9493 4499 9551 4505
rect 8386 4468 8392 4480
rect 8347 4440 8392 4468
rect 8386 4428 8392 4440
rect 8444 4428 8450 4480
rect 9125 4471 9183 4477
rect 9125 4437 9137 4471
rect 9171 4468 9183 4471
rect 9306 4468 9312 4480
rect 9171 4440 9312 4468
rect 9171 4437 9183 4440
rect 9125 4431 9183 4437
rect 9306 4428 9312 4440
rect 9364 4428 9370 4480
rect 11238 4468 11244 4480
rect 11199 4440 11244 4468
rect 11238 4428 11244 4440
rect 11296 4468 11302 4480
rect 11900 4468 11928 4567
rect 12066 4564 12072 4576
rect 12124 4564 12130 4616
rect 12989 4607 13047 4613
rect 12989 4604 13001 4607
rect 12544 4576 13001 4604
rect 12544 4480 12572 4576
rect 12989 4573 13001 4576
rect 13035 4573 13047 4607
rect 12989 4567 13047 4573
rect 15470 4564 15476 4616
rect 15528 4604 15534 4616
rect 15749 4607 15807 4613
rect 15749 4604 15761 4607
rect 15528 4576 15761 4604
rect 15528 4564 15534 4576
rect 15749 4573 15761 4576
rect 15795 4573 15807 4607
rect 15749 4567 15807 4573
rect 17402 4564 17408 4616
rect 17460 4604 17466 4616
rect 17862 4604 17868 4616
rect 17460 4576 17868 4604
rect 17460 4564 17466 4576
rect 17862 4564 17868 4576
rect 17920 4604 17926 4616
rect 18417 4607 18475 4613
rect 18417 4604 18429 4607
rect 17920 4576 18429 4604
rect 17920 4564 17926 4576
rect 18417 4573 18429 4576
rect 18463 4573 18475 4607
rect 22554 4604 22560 4616
rect 22467 4576 22560 4604
rect 18417 4567 18475 4573
rect 22554 4564 22560 4576
rect 22612 4564 22618 4616
rect 22646 4564 22652 4616
rect 22704 4604 22710 4616
rect 23106 4604 23112 4616
rect 22704 4576 23112 4604
rect 22704 4564 22710 4576
rect 23106 4564 23112 4576
rect 23164 4564 23170 4616
rect 23584 4604 23612 4700
rect 24765 4675 24823 4681
rect 24765 4641 24777 4675
rect 24811 4672 24823 4675
rect 25038 4672 25044 4684
rect 24811 4644 25044 4672
rect 24811 4641 24823 4644
rect 24765 4635 24823 4641
rect 25038 4632 25044 4644
rect 25096 4632 25102 4684
rect 25222 4672 25228 4684
rect 25183 4644 25228 4672
rect 25222 4632 25228 4644
rect 25280 4632 25286 4684
rect 24213 4607 24271 4613
rect 24213 4604 24225 4607
rect 23584 4576 24225 4604
rect 24213 4573 24225 4576
rect 24259 4573 24271 4607
rect 24213 4567 24271 4573
rect 22572 4536 22600 4564
rect 22738 4536 22744 4548
rect 22572 4508 22744 4536
rect 22738 4496 22744 4508
rect 22796 4496 22802 4548
rect 23658 4536 23664 4548
rect 23619 4508 23664 4536
rect 23658 4496 23664 4508
rect 23716 4496 23722 4548
rect 12526 4468 12532 4480
rect 11296 4440 11928 4468
rect 12487 4440 12532 4468
rect 11296 4428 11302 4440
rect 12526 4428 12532 4440
rect 12584 4428 12590 4480
rect 19794 4468 19800 4480
rect 19755 4440 19800 4468
rect 19794 4428 19800 4440
rect 19852 4428 19858 4480
rect 21174 4468 21180 4480
rect 21135 4440 21180 4468
rect 21174 4428 21180 4440
rect 21232 4428 21238 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 8665 4267 8723 4273
rect 8665 4233 8677 4267
rect 8711 4264 8723 4267
rect 8754 4264 8760 4276
rect 8711 4236 8760 4264
rect 8711 4233 8723 4236
rect 8665 4227 8723 4233
rect 8754 4224 8760 4236
rect 8812 4224 8818 4276
rect 9674 4224 9680 4276
rect 9732 4264 9738 4276
rect 11330 4264 11336 4276
rect 9732 4236 11336 4264
rect 9732 4224 9738 4236
rect 11330 4224 11336 4236
rect 11388 4224 11394 4276
rect 12802 4264 12808 4276
rect 12763 4236 12808 4264
rect 12802 4224 12808 4236
rect 12860 4224 12866 4276
rect 14366 4264 14372 4276
rect 14327 4236 14372 4264
rect 14366 4224 14372 4236
rect 14424 4224 14430 4276
rect 15657 4267 15715 4273
rect 15657 4233 15669 4267
rect 15703 4264 15715 4267
rect 16022 4264 16028 4276
rect 15703 4236 16028 4264
rect 15703 4233 15715 4236
rect 15657 4227 15715 4233
rect 16022 4224 16028 4236
rect 16080 4264 16086 4276
rect 18601 4267 18659 4273
rect 18601 4264 18613 4267
rect 16080 4236 18613 4264
rect 16080 4224 16086 4236
rect 18601 4233 18613 4236
rect 18647 4233 18659 4267
rect 20990 4264 20996 4276
rect 20951 4236 20996 4264
rect 18601 4227 18659 4233
rect 8294 4128 8300 4140
rect 7668 4100 8300 4128
rect 7668 4069 7696 4100
rect 8294 4088 8300 4100
rect 8352 4088 8358 4140
rect 8386 4088 8392 4140
rect 8444 4128 8450 4140
rect 9217 4131 9275 4137
rect 9217 4128 9229 4131
rect 8444 4100 9229 4128
rect 8444 4088 8450 4100
rect 9217 4097 9229 4100
rect 9263 4097 9275 4131
rect 9217 4091 9275 4097
rect 7653 4063 7711 4069
rect 7653 4029 7665 4063
rect 7699 4029 7711 4063
rect 7653 4023 7711 4029
rect 8846 4020 8852 4072
rect 8904 4060 8910 4072
rect 9125 4063 9183 4069
rect 9125 4060 9137 4063
rect 8904 4032 9137 4060
rect 8904 4020 8910 4032
rect 9125 4029 9137 4032
rect 9171 4029 9183 4063
rect 9232 4060 9260 4091
rect 9306 4088 9312 4140
rect 9364 4128 9370 4140
rect 10962 4128 10968 4140
rect 9364 4100 9409 4128
rect 10923 4100 10968 4128
rect 9364 4088 9370 4100
rect 10962 4088 10968 4100
rect 11020 4088 11026 4140
rect 13078 4128 13084 4140
rect 13039 4100 13084 4128
rect 13078 4088 13084 4100
rect 13136 4128 13142 4140
rect 13909 4131 13967 4137
rect 13136 4100 13676 4128
rect 13136 4088 13142 4100
rect 9398 4060 9404 4072
rect 9232 4032 9404 4060
rect 9125 4023 9183 4029
rect 9398 4020 9404 4032
rect 9456 4020 9462 4072
rect 13648 4069 13676 4100
rect 13909 4097 13921 4131
rect 13955 4128 13967 4131
rect 14384 4128 14412 4224
rect 18322 4196 18328 4208
rect 18283 4168 18328 4196
rect 18322 4156 18328 4168
rect 18380 4156 18386 4208
rect 18616 4196 18644 4227
rect 20990 4224 20996 4236
rect 21048 4224 21054 4276
rect 23477 4267 23535 4273
rect 23477 4233 23489 4267
rect 23523 4264 23535 4267
rect 23750 4264 23756 4276
rect 23523 4236 23756 4264
rect 23523 4233 23535 4236
rect 23477 4227 23535 4233
rect 23750 4224 23756 4236
rect 23808 4224 23814 4276
rect 24026 4224 24032 4276
rect 24084 4264 24090 4276
rect 24397 4267 24455 4273
rect 24397 4264 24409 4267
rect 24084 4236 24409 4264
rect 24084 4224 24090 4236
rect 24397 4233 24409 4236
rect 24443 4233 24455 4267
rect 24397 4227 24455 4233
rect 25222 4224 25228 4276
rect 25280 4264 25286 4276
rect 25409 4267 25467 4273
rect 25409 4264 25421 4267
rect 25280 4236 25421 4264
rect 25280 4224 25286 4236
rect 25409 4233 25421 4236
rect 25455 4233 25467 4267
rect 25409 4227 25467 4233
rect 19794 4196 19800 4208
rect 18616 4168 19800 4196
rect 13955 4100 14412 4128
rect 13955 4097 13967 4100
rect 13909 4091 13967 4097
rect 14550 4088 14556 4140
rect 14608 4128 14614 4140
rect 14645 4131 14703 4137
rect 14645 4128 14657 4131
rect 14608 4100 14657 4128
rect 14608 4088 14614 4100
rect 14645 4097 14657 4100
rect 14691 4128 14703 4131
rect 14734 4128 14740 4140
rect 14691 4100 14740 4128
rect 14691 4097 14703 4100
rect 14645 4091 14703 4097
rect 14734 4088 14740 4100
rect 14792 4088 14798 4140
rect 15289 4131 15347 4137
rect 15289 4097 15301 4131
rect 15335 4128 15347 4131
rect 17862 4128 17868 4140
rect 15335 4100 15884 4128
rect 17823 4100 17868 4128
rect 15335 4097 15347 4100
rect 15289 4091 15347 4097
rect 13633 4063 13691 4069
rect 13633 4029 13645 4063
rect 13679 4029 13691 4063
rect 13633 4023 13691 4029
rect 15470 4020 15476 4072
rect 15528 4060 15534 4072
rect 15749 4063 15807 4069
rect 15749 4060 15761 4063
rect 15528 4032 15761 4060
rect 15528 4020 15534 4032
rect 15749 4029 15761 4032
rect 15795 4029 15807 4063
rect 15856 4060 15884 4100
rect 17862 4088 17868 4100
rect 17920 4088 17926 4140
rect 19352 4137 19380 4168
rect 19794 4156 19800 4168
rect 19852 4156 19858 4208
rect 21266 4156 21272 4208
rect 21324 4196 21330 4208
rect 22738 4196 22744 4208
rect 21324 4168 21864 4196
rect 22699 4168 22744 4196
rect 21324 4156 21330 4168
rect 19337 4131 19395 4137
rect 19337 4097 19349 4131
rect 19383 4097 19395 4131
rect 19337 4091 19395 4097
rect 19889 4131 19947 4137
rect 19889 4097 19901 4131
rect 19935 4128 19947 4131
rect 20622 4128 20628 4140
rect 19935 4100 20628 4128
rect 19935 4097 19947 4100
rect 19889 4091 19947 4097
rect 16016 4063 16074 4069
rect 16016 4060 16028 4063
rect 15856 4032 16028 4060
rect 15749 4023 15807 4029
rect 16016 4029 16028 4032
rect 16062 4060 16074 4063
rect 16390 4060 16396 4072
rect 16062 4032 16396 4060
rect 16062 4029 16074 4032
rect 16016 4023 16074 4029
rect 16390 4020 16396 4032
rect 16448 4020 16454 4072
rect 19245 4063 19303 4069
rect 19245 4029 19257 4063
rect 19291 4060 19303 4063
rect 19904 4060 19932 4091
rect 20622 4088 20628 4100
rect 20680 4088 20686 4140
rect 21836 4137 21864 4168
rect 22738 4156 22744 4168
rect 22796 4156 22802 4208
rect 23106 4196 23112 4208
rect 23019 4168 23112 4196
rect 23106 4156 23112 4168
rect 23164 4196 23170 4208
rect 23164 4168 25084 4196
rect 23164 4156 23170 4168
rect 25056 4140 25084 4168
rect 21821 4131 21879 4137
rect 21821 4097 21833 4131
rect 21867 4097 21879 4131
rect 21821 4091 21879 4097
rect 23750 4088 23756 4140
rect 23808 4128 23814 4140
rect 24210 4128 24216 4140
rect 23808 4100 24216 4128
rect 23808 4088 23814 4100
rect 24210 4088 24216 4100
rect 24268 4088 24274 4140
rect 25038 4128 25044 4140
rect 24999 4100 25044 4128
rect 25038 4088 25044 4100
rect 25096 4088 25102 4140
rect 19291 4032 19932 4060
rect 19291 4029 19303 4032
rect 19245 4023 19303 4029
rect 20346 4020 20352 4072
rect 20404 4060 20410 4072
rect 23937 4063 23995 4069
rect 23937 4060 23949 4063
rect 20404 4032 23949 4060
rect 20404 4020 20410 4032
rect 23937 4029 23949 4032
rect 23983 4060 23995 4063
rect 24857 4063 24915 4069
rect 24857 4060 24869 4063
rect 23983 4032 24869 4060
rect 23983 4029 23995 4032
rect 23937 4023 23995 4029
rect 24857 4029 24869 4032
rect 24903 4029 24915 4063
rect 24857 4023 24915 4029
rect 9953 3995 10011 4001
rect 9953 3961 9965 3995
rect 9999 3992 10011 3995
rect 10134 3992 10140 4004
rect 9999 3964 10140 3992
rect 9999 3961 10011 3964
rect 9953 3955 10011 3961
rect 10134 3952 10140 3964
rect 10192 3952 10198 4004
rect 19150 3992 19156 4004
rect 19063 3964 19156 3992
rect 19150 3952 19156 3964
rect 19208 3992 19214 4004
rect 20165 3995 20223 4001
rect 20165 3992 20177 3995
rect 19208 3964 20177 3992
rect 19208 3952 19214 3964
rect 20165 3961 20177 3964
rect 20211 3961 20223 3995
rect 20714 3992 20720 4004
rect 20675 3964 20720 3992
rect 20165 3955 20223 3961
rect 20714 3952 20720 3964
rect 20772 3992 20778 4004
rect 21637 3995 21695 4001
rect 21637 3992 21649 3995
rect 20772 3964 21649 3992
rect 20772 3952 20778 3964
rect 21637 3961 21649 3964
rect 21683 3992 21695 3995
rect 21818 3992 21824 4004
rect 21683 3964 21824 3992
rect 21683 3961 21695 3964
rect 21637 3955 21695 3961
rect 21818 3952 21824 3964
rect 21876 3952 21882 4004
rect 7834 3924 7840 3936
rect 7795 3896 7840 3924
rect 7834 3884 7840 3896
rect 7892 3884 7898 3936
rect 8757 3927 8815 3933
rect 8757 3893 8769 3927
rect 8803 3924 8815 3927
rect 8938 3924 8944 3936
rect 8803 3896 8944 3924
rect 8803 3893 8815 3896
rect 8757 3887 8815 3893
rect 8938 3884 8944 3896
rect 8996 3884 9002 3936
rect 10042 3884 10048 3936
rect 10100 3924 10106 3936
rect 10321 3927 10379 3933
rect 10321 3924 10333 3927
rect 10100 3896 10333 3924
rect 10100 3884 10106 3896
rect 10321 3893 10333 3896
rect 10367 3893 10379 3927
rect 10686 3924 10692 3936
rect 10647 3896 10692 3924
rect 10321 3887 10379 3893
rect 10686 3884 10692 3896
rect 10744 3884 10750 3936
rect 10778 3884 10784 3936
rect 10836 3924 10842 3936
rect 11422 3924 11428 3936
rect 10836 3896 11428 3924
rect 10836 3884 10842 3896
rect 11422 3884 11428 3896
rect 11480 3884 11486 3936
rect 11698 3924 11704 3936
rect 11659 3896 11704 3924
rect 11698 3884 11704 3896
rect 11756 3884 11762 3936
rect 12066 3924 12072 3936
rect 12027 3896 12072 3924
rect 12066 3884 12072 3896
rect 12124 3884 12130 3936
rect 13262 3924 13268 3936
rect 13223 3896 13268 3924
rect 13262 3884 13268 3896
rect 13320 3884 13326 3936
rect 13538 3884 13544 3936
rect 13596 3924 13602 3936
rect 13725 3927 13783 3933
rect 13725 3924 13737 3927
rect 13596 3896 13737 3924
rect 13596 3884 13602 3896
rect 13725 3893 13737 3896
rect 13771 3893 13783 3927
rect 17126 3924 17132 3936
rect 17087 3896 17132 3924
rect 13725 3887 13783 3893
rect 17126 3884 17132 3896
rect 17184 3884 17190 3936
rect 17402 3924 17408 3936
rect 17363 3896 17408 3924
rect 17402 3884 17408 3896
rect 17460 3884 17466 3936
rect 18782 3924 18788 3936
rect 18743 3896 18788 3924
rect 18782 3884 18788 3896
rect 18840 3884 18846 3936
rect 21269 3927 21327 3933
rect 21269 3893 21281 3927
rect 21315 3924 21327 3927
rect 21450 3924 21456 3936
rect 21315 3896 21456 3924
rect 21315 3893 21327 3896
rect 21269 3887 21327 3893
rect 21450 3884 21456 3896
rect 21508 3884 21514 3936
rect 21542 3884 21548 3936
rect 21600 3924 21606 3936
rect 21729 3927 21787 3933
rect 21729 3924 21741 3927
rect 21600 3896 21741 3924
rect 21600 3884 21606 3896
rect 21729 3893 21741 3896
rect 21775 3893 21787 3927
rect 22278 3924 22284 3936
rect 22239 3896 22284 3924
rect 21729 3887 21787 3893
rect 22278 3884 22284 3896
rect 22336 3884 22342 3936
rect 24210 3924 24216 3936
rect 24171 3896 24216 3924
rect 24210 3884 24216 3896
rect 24268 3924 24274 3936
rect 24765 3927 24823 3933
rect 24765 3924 24777 3927
rect 24268 3896 24777 3924
rect 24268 3884 24274 3896
rect 24765 3893 24777 3896
rect 24811 3893 24823 3927
rect 24765 3887 24823 3893
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 8021 3723 8079 3729
rect 8021 3689 8033 3723
rect 8067 3720 8079 3723
rect 8846 3720 8852 3732
rect 8067 3692 8852 3720
rect 8067 3689 8079 3692
rect 8021 3683 8079 3689
rect 8846 3680 8852 3692
rect 8904 3680 8910 3732
rect 9490 3720 9496 3732
rect 9451 3692 9496 3720
rect 9490 3680 9496 3692
rect 9548 3680 9554 3732
rect 12434 3680 12440 3732
rect 12492 3720 12498 3732
rect 12989 3723 13047 3729
rect 12492 3692 12537 3720
rect 12492 3680 12498 3692
rect 12989 3689 13001 3723
rect 13035 3720 13047 3723
rect 13262 3720 13268 3732
rect 13035 3692 13268 3720
rect 13035 3689 13047 3692
rect 12989 3683 13047 3689
rect 13262 3680 13268 3692
rect 13320 3720 13326 3732
rect 14001 3723 14059 3729
rect 14001 3720 14013 3723
rect 13320 3692 14013 3720
rect 13320 3680 13326 3692
rect 14001 3689 14013 3692
rect 14047 3689 14059 3723
rect 14001 3683 14059 3689
rect 14182 3680 14188 3732
rect 14240 3720 14246 3732
rect 15013 3723 15071 3729
rect 15013 3720 15025 3723
rect 14240 3692 15025 3720
rect 14240 3680 14246 3692
rect 15013 3689 15025 3692
rect 15059 3720 15071 3723
rect 15470 3720 15476 3732
rect 15059 3692 15476 3720
rect 15059 3689 15071 3692
rect 15013 3683 15071 3689
rect 15470 3680 15476 3692
rect 15528 3680 15534 3732
rect 15657 3723 15715 3729
rect 15657 3689 15669 3723
rect 15703 3720 15715 3723
rect 17218 3720 17224 3732
rect 15703 3692 17224 3720
rect 15703 3689 15715 3692
rect 15657 3683 15715 3689
rect 17218 3680 17224 3692
rect 17276 3720 17282 3732
rect 17681 3723 17739 3729
rect 17681 3720 17693 3723
rect 17276 3692 17693 3720
rect 17276 3680 17282 3692
rect 17681 3689 17693 3692
rect 17727 3689 17739 3723
rect 17681 3683 17739 3689
rect 17862 3680 17868 3732
rect 17920 3720 17926 3732
rect 18046 3720 18052 3732
rect 17920 3692 18052 3720
rect 17920 3680 17926 3692
rect 18046 3680 18052 3692
rect 18104 3720 18110 3732
rect 18417 3723 18475 3729
rect 18417 3720 18429 3723
rect 18104 3692 18429 3720
rect 18104 3680 18110 3692
rect 18417 3689 18429 3692
rect 18463 3689 18475 3723
rect 18417 3683 18475 3689
rect 18785 3723 18843 3729
rect 18785 3689 18797 3723
rect 18831 3720 18843 3723
rect 19150 3720 19156 3732
rect 18831 3692 19156 3720
rect 18831 3689 18843 3692
rect 18785 3683 18843 3689
rect 8478 3612 8484 3664
rect 8536 3652 8542 3664
rect 8938 3652 8944 3664
rect 8536 3624 8944 3652
rect 8536 3612 8542 3624
rect 8938 3612 8944 3624
rect 8996 3652 9002 3664
rect 9033 3655 9091 3661
rect 9033 3652 9045 3655
rect 8996 3624 9045 3652
rect 8996 3612 9002 3624
rect 9033 3621 9045 3624
rect 9079 3621 9091 3655
rect 9033 3615 9091 3621
rect 13357 3655 13415 3661
rect 13357 3621 13369 3655
rect 13403 3652 13415 3655
rect 13538 3652 13544 3664
rect 13403 3624 13544 3652
rect 13403 3621 13415 3624
rect 13357 3615 13415 3621
rect 13538 3612 13544 3624
rect 13596 3612 13602 3664
rect 13814 3612 13820 3664
rect 13872 3652 13878 3664
rect 13909 3655 13967 3661
rect 13909 3652 13921 3655
rect 13872 3624 13921 3652
rect 13872 3612 13878 3624
rect 13909 3621 13921 3624
rect 13955 3621 13967 3655
rect 13909 3615 13967 3621
rect 15378 3612 15384 3664
rect 15436 3652 15442 3664
rect 16025 3655 16083 3661
rect 16025 3652 16037 3655
rect 15436 3624 16037 3652
rect 15436 3612 15442 3624
rect 16025 3621 16037 3624
rect 16071 3621 16083 3655
rect 17586 3652 17592 3664
rect 17547 3624 17592 3652
rect 16025 3615 16083 3621
rect 17586 3612 17592 3624
rect 17644 3612 17650 3664
rect 18432 3652 18460 3683
rect 19150 3680 19156 3692
rect 19208 3680 19214 3732
rect 23750 3720 23756 3732
rect 23711 3692 23756 3720
rect 23750 3680 23756 3692
rect 23808 3680 23814 3732
rect 19889 3655 19947 3661
rect 19889 3652 19901 3655
rect 18432 3624 19901 3652
rect 19889 3621 19901 3624
rect 19935 3652 19947 3655
rect 20717 3655 20775 3661
rect 20717 3652 20729 3655
rect 19935 3624 20729 3652
rect 19935 3621 19947 3624
rect 19889 3615 19947 3621
rect 20717 3621 20729 3624
rect 20763 3652 20775 3655
rect 21174 3652 21180 3664
rect 20763 3624 21180 3652
rect 20763 3621 20775 3624
rect 20717 3615 20775 3621
rect 21174 3612 21180 3624
rect 21232 3652 21238 3664
rect 24296 3655 24354 3661
rect 21232 3624 24072 3652
rect 21232 3612 21238 3624
rect 6914 3584 6920 3596
rect 6875 3556 6920 3584
rect 6914 3544 6920 3556
rect 6972 3544 6978 3596
rect 8386 3584 8392 3596
rect 8347 3556 8392 3584
rect 8386 3544 8392 3556
rect 8444 3544 8450 3596
rect 9950 3584 9956 3596
rect 9911 3556 9956 3584
rect 9950 3544 9956 3556
rect 10008 3544 10014 3596
rect 11330 3593 11336 3596
rect 11324 3584 11336 3593
rect 11291 3556 11336 3584
rect 11324 3547 11336 3556
rect 11330 3544 11336 3547
rect 11388 3544 11394 3596
rect 15470 3544 15476 3596
rect 15528 3584 15534 3596
rect 16669 3587 16727 3593
rect 16669 3584 16681 3587
rect 15528 3556 16681 3584
rect 15528 3544 15534 3556
rect 16669 3553 16681 3556
rect 16715 3584 16727 3587
rect 17402 3584 17408 3596
rect 16715 3556 17408 3584
rect 16715 3553 16727 3556
rect 16669 3547 16727 3553
rect 17402 3544 17408 3556
rect 17460 3544 17466 3596
rect 19150 3584 19156 3596
rect 19111 3556 19156 3584
rect 19150 3544 19156 3556
rect 19208 3544 19214 3596
rect 21634 3584 21640 3596
rect 21595 3556 21640 3584
rect 21634 3544 21640 3556
rect 21692 3544 21698 3596
rect 21836 3593 21864 3624
rect 21821 3587 21879 3593
rect 21821 3553 21833 3587
rect 21867 3553 21879 3587
rect 21821 3547 21879 3553
rect 21910 3544 21916 3596
rect 21968 3584 21974 3596
rect 22077 3587 22135 3593
rect 22077 3584 22089 3587
rect 21968 3556 22089 3584
rect 21968 3544 21974 3556
rect 22077 3553 22089 3556
rect 22123 3553 22135 3587
rect 22077 3547 22135 3553
rect 24044 3528 24072 3624
rect 24296 3621 24308 3655
rect 24342 3652 24354 3655
rect 24762 3652 24768 3664
rect 24342 3624 24768 3652
rect 24342 3621 24354 3624
rect 24296 3615 24354 3621
rect 24762 3612 24768 3624
rect 24820 3612 24826 3664
rect 8478 3516 8484 3528
rect 8439 3488 8484 3516
rect 8478 3476 8484 3488
rect 8536 3476 8542 3528
rect 8662 3516 8668 3528
rect 8623 3488 8668 3516
rect 8662 3476 8668 3488
rect 8720 3476 8726 3528
rect 11057 3519 11115 3525
rect 11057 3485 11069 3519
rect 11103 3485 11115 3519
rect 11057 3479 11115 3485
rect 14185 3519 14243 3525
rect 14185 3485 14197 3519
rect 14231 3516 14243 3519
rect 14642 3516 14648 3528
rect 14231 3488 14648 3516
rect 14231 3485 14243 3488
rect 14185 3479 14243 3485
rect 7929 3451 7987 3457
rect 7929 3417 7941 3451
rect 7975 3448 7987 3451
rect 8680 3448 8708 3476
rect 7975 3420 8708 3448
rect 7975 3417 7987 3420
rect 7929 3411 7987 3417
rect 9766 3408 9772 3460
rect 9824 3448 9830 3460
rect 10505 3451 10563 3457
rect 10505 3448 10517 3451
rect 9824 3420 10517 3448
rect 9824 3408 9830 3420
rect 10505 3417 10517 3420
rect 10551 3448 10563 3451
rect 10686 3448 10692 3460
rect 10551 3420 10692 3448
rect 10551 3417 10563 3420
rect 10505 3411 10563 3417
rect 10686 3408 10692 3420
rect 10744 3408 10750 3460
rect 7098 3380 7104 3392
rect 7059 3352 7104 3380
rect 7098 3340 7104 3352
rect 7156 3340 7162 3392
rect 7561 3383 7619 3389
rect 7561 3349 7573 3383
rect 7607 3380 7619 3383
rect 9030 3380 9036 3392
rect 7607 3352 9036 3380
rect 7607 3349 7619 3352
rect 7561 3343 7619 3349
rect 9030 3340 9036 3352
rect 9088 3340 9094 3392
rect 10137 3383 10195 3389
rect 10137 3349 10149 3383
rect 10183 3380 10195 3383
rect 10778 3380 10784 3392
rect 10183 3352 10784 3380
rect 10183 3349 10195 3352
rect 10137 3343 10195 3349
rect 10778 3340 10784 3352
rect 10836 3340 10842 3392
rect 10962 3380 10968 3392
rect 10923 3352 10968 3380
rect 10962 3340 10968 3352
rect 11020 3340 11026 3392
rect 11072 3380 11100 3479
rect 14642 3476 14648 3488
rect 14700 3476 14706 3528
rect 16114 3516 16120 3528
rect 16075 3488 16120 3516
rect 16114 3476 16120 3488
rect 16172 3476 16178 3528
rect 16301 3519 16359 3525
rect 16301 3485 16313 3519
rect 16347 3516 16359 3519
rect 16482 3516 16488 3528
rect 16347 3488 16488 3516
rect 16347 3485 16359 3488
rect 16301 3479 16359 3485
rect 13541 3451 13599 3457
rect 13541 3417 13553 3451
rect 13587 3448 13599 3451
rect 13630 3448 13636 3460
rect 13587 3420 13636 3448
rect 13587 3417 13599 3420
rect 13541 3411 13599 3417
rect 13630 3408 13636 3420
rect 13688 3408 13694 3460
rect 15565 3451 15623 3457
rect 15565 3417 15577 3451
rect 15611 3448 15623 3451
rect 16316 3448 16344 3479
rect 16482 3476 16488 3488
rect 16540 3476 16546 3528
rect 17862 3516 17868 3528
rect 17823 3488 17868 3516
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 19242 3516 19248 3528
rect 19203 3488 19248 3516
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 19334 3476 19340 3528
rect 19392 3516 19398 3528
rect 19429 3519 19487 3525
rect 19429 3516 19441 3519
rect 19392 3488 19441 3516
rect 19392 3476 19398 3488
rect 19429 3485 19441 3488
rect 19475 3516 19487 3519
rect 20622 3516 20628 3528
rect 19475 3488 20628 3516
rect 19475 3485 19487 3488
rect 19429 3479 19487 3485
rect 20622 3476 20628 3488
rect 20680 3476 20686 3528
rect 24026 3516 24032 3528
rect 23987 3488 24032 3516
rect 24026 3476 24032 3488
rect 24084 3476 24090 3528
rect 15611 3420 16344 3448
rect 15611 3417 15623 3420
rect 15565 3411 15623 3417
rect 17034 3408 17040 3460
rect 17092 3448 17098 3460
rect 17221 3451 17279 3457
rect 17221 3448 17233 3451
rect 17092 3420 17233 3448
rect 17092 3408 17098 3420
rect 17221 3417 17233 3420
rect 17267 3417 17279 3451
rect 17221 3411 17279 3417
rect 11422 3380 11428 3392
rect 11072 3352 11428 3380
rect 11422 3340 11428 3352
rect 11480 3340 11486 3392
rect 21361 3383 21419 3389
rect 21361 3349 21373 3383
rect 21407 3380 21419 3383
rect 21450 3380 21456 3392
rect 21407 3352 21456 3380
rect 21407 3349 21419 3352
rect 21361 3343 21419 3349
rect 21450 3340 21456 3352
rect 21508 3340 21514 3392
rect 21634 3340 21640 3392
rect 21692 3380 21698 3392
rect 23201 3383 23259 3389
rect 23201 3380 23213 3383
rect 21692 3352 23213 3380
rect 21692 3340 21698 3352
rect 23201 3349 23213 3352
rect 23247 3349 23259 3383
rect 25406 3380 25412 3392
rect 25367 3352 25412 3380
rect 23201 3343 23259 3349
rect 25406 3340 25412 3352
rect 25464 3340 25470 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 5813 3179 5871 3185
rect 5813 3145 5825 3179
rect 5859 3176 5871 3179
rect 5994 3176 6000 3188
rect 5859 3148 6000 3176
rect 5859 3145 5871 3148
rect 5813 3139 5871 3145
rect 5994 3136 6000 3148
rect 6052 3136 6058 3188
rect 6270 3176 6276 3188
rect 6231 3148 6276 3176
rect 6270 3136 6276 3148
rect 6328 3136 6334 3188
rect 6638 3176 6644 3188
rect 6599 3148 6644 3176
rect 6638 3136 6644 3148
rect 6696 3136 6702 3188
rect 6914 3136 6920 3188
rect 6972 3176 6978 3188
rect 7009 3179 7067 3185
rect 7009 3176 7021 3179
rect 6972 3148 7021 3176
rect 6972 3136 6978 3148
rect 7009 3145 7021 3148
rect 7055 3145 7067 3179
rect 7009 3139 7067 3145
rect 8018 3136 8024 3188
rect 8076 3176 8082 3188
rect 9766 3176 9772 3188
rect 8076 3148 9772 3176
rect 8076 3136 8082 3148
rect 9766 3136 9772 3148
rect 9824 3136 9830 3188
rect 9861 3179 9919 3185
rect 9861 3145 9873 3179
rect 9907 3176 9919 3179
rect 11330 3176 11336 3188
rect 9907 3148 11336 3176
rect 9907 3145 9919 3148
rect 9861 3139 9919 3145
rect 11330 3136 11336 3148
rect 11388 3176 11394 3188
rect 11517 3179 11575 3185
rect 11517 3176 11529 3179
rect 11388 3148 11529 3176
rect 11388 3136 11394 3148
rect 11517 3145 11529 3148
rect 11563 3176 11575 3179
rect 11793 3179 11851 3185
rect 11793 3176 11805 3179
rect 11563 3148 11805 3176
rect 11563 3145 11575 3148
rect 11517 3139 11575 3145
rect 11793 3145 11805 3148
rect 11839 3145 11851 3179
rect 11793 3139 11851 3145
rect 13814 3136 13820 3188
rect 13872 3176 13878 3188
rect 14093 3179 14151 3185
rect 14093 3176 14105 3179
rect 13872 3148 14105 3176
rect 13872 3136 13878 3148
rect 14093 3145 14105 3148
rect 14139 3145 14151 3179
rect 15378 3176 15384 3188
rect 15339 3148 15384 3176
rect 14093 3139 14151 3145
rect 15378 3136 15384 3148
rect 15436 3136 15442 3188
rect 16114 3176 16120 3188
rect 15488 3148 16120 3176
rect 7653 3111 7711 3117
rect 7653 3077 7665 3111
rect 7699 3108 7711 3111
rect 8294 3108 8300 3120
rect 7699 3080 8300 3108
rect 7699 3077 7711 3080
rect 7653 3071 7711 3077
rect 8294 3068 8300 3080
rect 8352 3068 8358 3120
rect 8570 3108 8576 3120
rect 8531 3080 8576 3108
rect 8570 3068 8576 3080
rect 8628 3068 8634 3120
rect 9674 3068 9680 3120
rect 9732 3108 9738 3120
rect 15013 3111 15071 3117
rect 9732 3080 10180 3108
rect 9732 3068 9738 3080
rect 8110 3040 8116 3052
rect 7484 3012 8116 3040
rect 5629 2975 5687 2981
rect 5629 2941 5641 2975
rect 5675 2972 5687 2975
rect 6270 2972 6276 2984
rect 5675 2944 6276 2972
rect 5675 2941 5687 2944
rect 5629 2935 5687 2941
rect 6270 2932 6276 2944
rect 6328 2932 6334 2984
rect 7484 2981 7512 3012
rect 8110 3000 8116 3012
rect 8168 3000 8174 3052
rect 10152 3049 10180 3080
rect 15013 3077 15025 3111
rect 15059 3108 15071 3111
rect 15488 3108 15516 3148
rect 16114 3136 16120 3148
rect 16172 3136 16178 3188
rect 16850 3176 16856 3188
rect 16763 3148 16856 3176
rect 16850 3136 16856 3148
rect 16908 3176 16914 3188
rect 17681 3179 17739 3185
rect 17681 3176 17693 3179
rect 16908 3148 17693 3176
rect 16908 3136 16914 3148
rect 17681 3145 17693 3148
rect 17727 3176 17739 3179
rect 17862 3176 17868 3188
rect 17727 3148 17868 3176
rect 17727 3145 17739 3148
rect 17681 3139 17739 3145
rect 17862 3136 17868 3148
rect 17920 3136 17926 3188
rect 19150 3136 19156 3188
rect 19208 3176 19214 3188
rect 20073 3179 20131 3185
rect 20073 3176 20085 3179
rect 19208 3148 20085 3176
rect 19208 3136 19214 3148
rect 20073 3145 20085 3148
rect 20119 3145 20131 3179
rect 20073 3139 20131 3145
rect 20533 3179 20591 3185
rect 20533 3145 20545 3179
rect 20579 3176 20591 3179
rect 20622 3176 20628 3188
rect 20579 3148 20628 3176
rect 20579 3145 20591 3148
rect 20533 3139 20591 3145
rect 20622 3136 20628 3148
rect 20680 3136 20686 3188
rect 21085 3179 21143 3185
rect 21085 3145 21097 3179
rect 21131 3176 21143 3179
rect 21910 3176 21916 3188
rect 21131 3148 21916 3176
rect 21131 3145 21143 3148
rect 21085 3139 21143 3145
rect 21910 3136 21916 3148
rect 21968 3176 21974 3188
rect 21968 3148 23152 3176
rect 21968 3136 21974 3148
rect 15059 3080 15516 3108
rect 17313 3111 17371 3117
rect 15059 3077 15071 3080
rect 15013 3071 15071 3077
rect 17313 3077 17325 3111
rect 17359 3108 17371 3111
rect 17586 3108 17592 3120
rect 17359 3080 17592 3108
rect 17359 3077 17371 3080
rect 17313 3071 17371 3077
rect 17586 3068 17592 3080
rect 17644 3068 17650 3120
rect 19242 3068 19248 3120
rect 19300 3108 19306 3120
rect 19705 3111 19763 3117
rect 19705 3108 19717 3111
rect 19300 3080 19717 3108
rect 19300 3068 19306 3080
rect 19705 3077 19717 3080
rect 19751 3077 19763 3111
rect 19705 3071 19763 3077
rect 9217 3043 9275 3049
rect 9217 3009 9229 3043
rect 9263 3040 9275 3043
rect 9861 3043 9919 3049
rect 9861 3040 9873 3043
rect 9263 3012 9873 3040
rect 9263 3009 9275 3012
rect 9217 3003 9275 3009
rect 9861 3009 9873 3012
rect 9907 3040 9919 3043
rect 9953 3043 10011 3049
rect 9953 3040 9965 3043
rect 9907 3012 9965 3040
rect 9907 3009 9919 3012
rect 9861 3003 9919 3009
rect 9953 3009 9965 3012
rect 9999 3009 10011 3043
rect 9953 3003 10011 3009
rect 10137 3043 10195 3049
rect 10137 3009 10149 3043
rect 10183 3009 10195 3043
rect 10137 3003 10195 3009
rect 11422 3000 11428 3052
rect 11480 3040 11486 3052
rect 12434 3040 12440 3052
rect 11480 3012 12440 3040
rect 11480 3000 11486 3012
rect 12434 3000 12440 3012
rect 12492 3040 12498 3052
rect 15470 3040 15476 3052
rect 12492 3012 12585 3040
rect 15431 3012 15476 3040
rect 12492 3000 12498 3012
rect 15470 3000 15476 3012
rect 15528 3000 15534 3052
rect 17034 3000 17040 3052
rect 17092 3040 17098 3052
rect 17494 3040 17500 3052
rect 17092 3012 17500 3040
rect 17092 3000 17098 3012
rect 17494 3000 17500 3012
rect 17552 3000 17558 3052
rect 18046 3040 18052 3052
rect 18007 3012 18052 3040
rect 18046 3000 18052 3012
rect 18104 3000 18110 3052
rect 21174 3040 21180 3052
rect 21135 3012 21180 3040
rect 21174 3000 21180 3012
rect 21232 3000 21238 3052
rect 23124 3049 23152 3148
rect 24026 3136 24032 3188
rect 24084 3176 24090 3188
rect 25041 3179 25099 3185
rect 25041 3176 25053 3179
rect 24084 3148 25053 3176
rect 24084 3136 24090 3148
rect 25041 3145 25053 3148
rect 25087 3145 25099 3179
rect 25041 3139 25099 3145
rect 23477 3111 23535 3117
rect 23477 3077 23489 3111
rect 23523 3108 23535 3111
rect 24118 3108 24124 3120
rect 23523 3080 24124 3108
rect 23523 3077 23535 3080
rect 23477 3071 23535 3077
rect 24118 3068 24124 3080
rect 24176 3068 24182 3120
rect 24762 3108 24768 3120
rect 24723 3080 24768 3108
rect 24762 3068 24768 3080
rect 24820 3068 24826 3120
rect 23109 3043 23167 3049
rect 23109 3009 23121 3043
rect 23155 3040 23167 3043
rect 24305 3043 24363 3049
rect 24305 3040 24317 3043
rect 23155 3012 24317 3040
rect 23155 3009 23167 3012
rect 23109 3003 23167 3009
rect 24305 3009 24317 3012
rect 24351 3040 24363 3043
rect 24578 3040 24584 3052
rect 24351 3012 24584 3040
rect 24351 3009 24363 3012
rect 24305 3003 24363 3009
rect 24578 3000 24584 3012
rect 24636 3040 24642 3052
rect 25406 3040 25412 3052
rect 24636 3012 25412 3040
rect 24636 3000 24642 3012
rect 25406 3000 25412 3012
rect 25464 3000 25470 3052
rect 7469 2975 7527 2981
rect 7469 2941 7481 2975
rect 7515 2941 7527 2975
rect 8478 2972 8484 2984
rect 8439 2944 8484 2972
rect 7469 2935 7527 2941
rect 8478 2932 8484 2944
rect 8536 2932 8542 2984
rect 8938 2972 8944 2984
rect 8899 2944 8944 2972
rect 8938 2932 8944 2944
rect 8996 2932 9002 2984
rect 9030 2932 9036 2984
rect 9088 2972 9094 2984
rect 10042 2972 10048 2984
rect 9088 2944 10048 2972
rect 9088 2932 9094 2944
rect 10042 2932 10048 2944
rect 10100 2932 10106 2984
rect 10870 2972 10876 2984
rect 10244 2944 10876 2972
rect 8386 2864 8392 2916
rect 8444 2904 8450 2916
rect 9585 2907 9643 2913
rect 9585 2904 9597 2907
rect 8444 2876 9597 2904
rect 8444 2864 8450 2876
rect 9585 2873 9597 2876
rect 9631 2904 9643 2907
rect 10244 2904 10272 2944
rect 10870 2932 10876 2944
rect 10928 2932 10934 2984
rect 24118 2972 24124 2984
rect 24079 2944 24124 2972
rect 24118 2932 24124 2944
rect 24176 2932 24182 2984
rect 9631 2876 10272 2904
rect 10404 2907 10462 2913
rect 9631 2873 9643 2876
rect 9585 2867 9643 2873
rect 10404 2873 10416 2907
rect 10450 2904 10462 2907
rect 12250 2904 12256 2916
rect 10450 2876 10484 2904
rect 12163 2876 12256 2904
rect 10450 2873 10462 2876
rect 10404 2867 10462 2873
rect 9674 2796 9680 2848
rect 9732 2836 9738 2848
rect 10419 2836 10447 2867
rect 12250 2864 12256 2876
rect 12308 2904 12314 2916
rect 12704 2907 12762 2913
rect 12704 2904 12716 2907
rect 12308 2876 12716 2904
rect 12308 2864 12314 2876
rect 12704 2873 12716 2876
rect 12750 2904 12762 2907
rect 13722 2904 13728 2916
rect 12750 2876 13728 2904
rect 12750 2873 12762 2876
rect 12704 2867 12762 2873
rect 13722 2864 13728 2876
rect 13780 2864 13786 2916
rect 14645 2907 14703 2913
rect 14645 2873 14657 2907
rect 14691 2904 14703 2907
rect 15740 2907 15798 2913
rect 15740 2904 15752 2907
rect 14691 2876 15752 2904
rect 14691 2873 14703 2876
rect 14645 2867 14703 2873
rect 15740 2873 15752 2876
rect 15786 2904 15798 2907
rect 16482 2904 16488 2916
rect 15786 2876 16488 2904
rect 15786 2873 15798 2876
rect 15740 2867 15798 2873
rect 16482 2864 16488 2876
rect 16540 2864 16546 2916
rect 18138 2864 18144 2916
rect 18196 2904 18202 2916
rect 18294 2907 18352 2913
rect 18294 2904 18306 2907
rect 18196 2876 18306 2904
rect 18196 2864 18202 2876
rect 18294 2873 18306 2876
rect 18340 2873 18352 2907
rect 18294 2867 18352 2873
rect 21444 2907 21502 2913
rect 21444 2873 21456 2907
rect 21490 2904 21502 2907
rect 21634 2904 21640 2916
rect 21490 2876 21640 2904
rect 21490 2873 21502 2876
rect 21444 2867 21502 2873
rect 21634 2864 21640 2876
rect 21692 2864 21698 2916
rect 23750 2864 23756 2916
rect 23808 2904 23814 2916
rect 24029 2907 24087 2913
rect 24029 2904 24041 2907
rect 23808 2876 24041 2904
rect 23808 2864 23814 2876
rect 24029 2873 24041 2876
rect 24075 2873 24087 2907
rect 24029 2867 24087 2873
rect 10962 2836 10968 2848
rect 9732 2808 10968 2836
rect 9732 2796 9738 2808
rect 10962 2796 10968 2808
rect 11020 2796 11026 2848
rect 13814 2836 13820 2848
rect 13775 2808 13820 2836
rect 13814 2796 13820 2808
rect 13872 2796 13878 2848
rect 19426 2836 19432 2848
rect 19387 2808 19432 2836
rect 19426 2796 19432 2808
rect 19484 2796 19490 2848
rect 22554 2836 22560 2848
rect 22515 2808 22560 2836
rect 22554 2796 22560 2808
rect 22612 2796 22618 2848
rect 23474 2796 23480 2848
rect 23532 2836 23538 2848
rect 23661 2839 23719 2845
rect 23661 2836 23673 2839
rect 23532 2808 23673 2836
rect 23532 2796 23538 2808
rect 23661 2805 23673 2808
rect 23707 2805 23719 2839
rect 25406 2836 25412 2848
rect 25367 2808 25412 2836
rect 23661 2799 23719 2805
rect 25406 2796 25412 2808
rect 25464 2796 25470 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 5626 2632 5632 2644
rect 5587 2604 5632 2632
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 6362 2632 6368 2644
rect 6323 2604 6368 2632
rect 6362 2592 6368 2604
rect 6420 2592 6426 2644
rect 8110 2632 8116 2644
rect 8071 2604 8116 2632
rect 8110 2592 8116 2604
rect 8168 2592 8174 2644
rect 10962 2592 10968 2644
rect 11020 2632 11026 2644
rect 11517 2635 11575 2641
rect 11517 2632 11529 2635
rect 11020 2604 11529 2632
rect 11020 2592 11026 2604
rect 11517 2601 11529 2604
rect 11563 2601 11575 2635
rect 11882 2632 11888 2644
rect 11843 2604 11888 2632
rect 11517 2595 11575 2601
rect 11882 2592 11888 2604
rect 11940 2592 11946 2644
rect 13814 2592 13820 2644
rect 13872 2632 13878 2644
rect 14001 2635 14059 2641
rect 14001 2632 14013 2635
rect 13872 2604 14013 2632
rect 13872 2592 13878 2604
rect 14001 2601 14013 2604
rect 14047 2601 14059 2635
rect 14734 2632 14740 2644
rect 14695 2604 14740 2632
rect 14001 2595 14059 2601
rect 14734 2592 14740 2604
rect 14792 2592 14798 2644
rect 16482 2592 16488 2644
rect 16540 2632 16546 2644
rect 16853 2635 16911 2641
rect 16853 2632 16865 2635
rect 16540 2604 16865 2632
rect 16540 2592 16546 2604
rect 16853 2601 16865 2604
rect 16899 2601 16911 2635
rect 17218 2632 17224 2644
rect 17179 2604 17224 2632
rect 16853 2595 16911 2601
rect 17218 2592 17224 2604
rect 17276 2592 17282 2644
rect 17402 2592 17408 2644
rect 17460 2632 17466 2644
rect 17589 2635 17647 2641
rect 17589 2632 17601 2635
rect 17460 2604 17601 2632
rect 17460 2592 17466 2604
rect 17589 2601 17601 2604
rect 17635 2601 17647 2635
rect 18138 2632 18144 2644
rect 18099 2604 18144 2632
rect 17589 2595 17647 2601
rect 18138 2592 18144 2604
rect 18196 2632 18202 2644
rect 19334 2632 19340 2644
rect 18196 2604 19340 2632
rect 18196 2592 18202 2604
rect 19334 2592 19340 2604
rect 19392 2632 19398 2644
rect 20257 2635 20315 2641
rect 20257 2632 20269 2635
rect 19392 2604 20269 2632
rect 19392 2592 19398 2604
rect 20257 2601 20269 2604
rect 20303 2601 20315 2635
rect 20257 2595 20315 2601
rect 20993 2635 21051 2641
rect 20993 2601 21005 2635
rect 21039 2632 21051 2635
rect 22189 2635 22247 2641
rect 21039 2604 22140 2632
rect 21039 2601 21051 2604
rect 20993 2595 21051 2601
rect 5721 2499 5779 2505
rect 5721 2465 5733 2499
rect 5767 2496 5779 2499
rect 6380 2496 6408 2592
rect 8021 2567 8079 2573
rect 8021 2533 8033 2567
rect 8067 2564 8079 2567
rect 8481 2567 8539 2573
rect 8481 2564 8493 2567
rect 8067 2536 8493 2564
rect 8067 2533 8079 2536
rect 8021 2527 8079 2533
rect 8481 2533 8493 2536
rect 8527 2564 8539 2567
rect 8662 2564 8668 2576
rect 8527 2536 8668 2564
rect 8527 2533 8539 2536
rect 8481 2527 8539 2533
rect 8662 2524 8668 2536
rect 8720 2524 8726 2576
rect 9582 2564 9588 2576
rect 9543 2536 9588 2564
rect 9582 2524 9588 2536
rect 9640 2524 9646 2576
rect 9950 2524 9956 2576
rect 10008 2564 10014 2576
rect 11422 2564 11428 2576
rect 10008 2536 11428 2564
rect 10008 2524 10014 2536
rect 11422 2524 11428 2536
rect 11480 2524 11486 2576
rect 12434 2524 12440 2576
rect 12492 2564 12498 2576
rect 14752 2564 14780 2592
rect 12492 2536 14780 2564
rect 15289 2567 15347 2573
rect 12492 2524 12498 2536
rect 5767 2468 6408 2496
rect 6733 2499 6791 2505
rect 5767 2465 5779 2468
rect 5721 2459 5779 2465
rect 6733 2465 6745 2499
rect 6779 2496 6791 2499
rect 7006 2496 7012 2508
rect 6779 2468 7012 2496
rect 6779 2465 6791 2468
rect 6733 2459 6791 2465
rect 7006 2456 7012 2468
rect 7064 2456 7070 2508
rect 10045 2499 10103 2505
rect 10045 2465 10057 2499
rect 10091 2496 10103 2499
rect 10404 2499 10462 2505
rect 10404 2496 10416 2499
rect 10091 2468 10416 2496
rect 10091 2465 10103 2468
rect 10045 2459 10103 2465
rect 10404 2465 10416 2468
rect 10450 2496 10462 2499
rect 10962 2496 10968 2508
rect 10450 2468 10968 2496
rect 10450 2465 10462 2468
rect 10404 2459 10462 2465
rect 10962 2456 10968 2468
rect 11020 2456 11026 2508
rect 12636 2505 12664 2536
rect 15289 2533 15301 2567
rect 15335 2564 15347 2567
rect 15740 2567 15798 2573
rect 15740 2564 15752 2567
rect 15335 2536 15752 2564
rect 15335 2533 15347 2536
rect 15289 2527 15347 2533
rect 15740 2533 15752 2536
rect 15786 2564 15798 2567
rect 15930 2564 15936 2576
rect 15786 2536 15936 2564
rect 15786 2533 15798 2536
rect 15740 2527 15798 2533
rect 15930 2524 15936 2536
rect 15988 2524 15994 2576
rect 19150 2573 19156 2576
rect 18785 2567 18843 2573
rect 18785 2533 18797 2567
rect 18831 2564 18843 2567
rect 19144 2564 19156 2573
rect 18831 2536 19156 2564
rect 18831 2533 18843 2536
rect 18785 2527 18843 2533
rect 19144 2527 19156 2536
rect 19150 2524 19156 2527
rect 19208 2524 19214 2576
rect 12894 2505 12900 2508
rect 12621 2499 12679 2505
rect 12621 2465 12633 2499
rect 12667 2465 12679 2499
rect 12888 2496 12900 2505
rect 12621 2459 12679 2465
rect 12728 2468 12900 2496
rect 4706 2428 4712 2440
rect 4667 2400 4712 2428
rect 4706 2388 4712 2400
rect 4764 2388 4770 2440
rect 7653 2431 7711 2437
rect 7653 2397 7665 2431
rect 7699 2428 7711 2431
rect 8570 2428 8576 2440
rect 7699 2400 8576 2428
rect 7699 2397 7711 2400
rect 7653 2391 7711 2397
rect 8570 2388 8576 2400
rect 8628 2388 8634 2440
rect 8757 2431 8815 2437
rect 8757 2397 8769 2431
rect 8803 2428 8815 2431
rect 8803 2400 9260 2428
rect 8803 2397 8815 2400
rect 8757 2391 8815 2397
rect 9232 2304 9260 2400
rect 9950 2388 9956 2440
rect 10008 2428 10014 2440
rect 10137 2431 10195 2437
rect 10137 2428 10149 2431
rect 10008 2400 10149 2428
rect 10008 2388 10014 2400
rect 10137 2397 10149 2400
rect 10183 2397 10195 2431
rect 10137 2391 10195 2397
rect 12437 2431 12495 2437
rect 12437 2397 12449 2431
rect 12483 2428 12495 2431
rect 12728 2428 12756 2468
rect 12888 2459 12900 2468
rect 12894 2456 12900 2459
rect 12952 2456 12958 2508
rect 14369 2499 14427 2505
rect 14369 2465 14381 2499
rect 14415 2496 14427 2499
rect 14642 2496 14648 2508
rect 14415 2468 14648 2496
rect 14415 2465 14427 2468
rect 14369 2459 14427 2465
rect 14642 2456 14648 2468
rect 14700 2456 14706 2508
rect 15470 2496 15476 2508
rect 15431 2468 15476 2496
rect 15470 2456 15476 2468
rect 15528 2456 15534 2508
rect 18877 2499 18935 2505
rect 18877 2465 18889 2499
rect 18923 2496 18935 2499
rect 20625 2499 20683 2505
rect 20625 2496 20637 2499
rect 18923 2468 20637 2496
rect 18923 2465 18935 2468
rect 18877 2459 18935 2465
rect 20625 2465 20637 2468
rect 20671 2496 20683 2499
rect 21174 2496 21180 2508
rect 20671 2468 21180 2496
rect 20671 2465 20683 2468
rect 20625 2459 20683 2465
rect 21174 2456 21180 2468
rect 21232 2456 21238 2508
rect 22112 2496 22140 2604
rect 22189 2601 22201 2635
rect 22235 2632 22247 2635
rect 22925 2635 22983 2641
rect 22925 2632 22937 2635
rect 22235 2604 22937 2632
rect 22235 2601 22247 2604
rect 22189 2595 22247 2601
rect 22925 2601 22937 2604
rect 22971 2632 22983 2635
rect 23382 2632 23388 2644
rect 22971 2604 23388 2632
rect 22971 2601 22983 2604
rect 22925 2595 22983 2601
rect 23382 2592 23388 2604
rect 23440 2592 23446 2644
rect 25590 2632 25596 2644
rect 25551 2604 25596 2632
rect 25590 2592 25596 2604
rect 25648 2592 25654 2644
rect 24397 2567 24455 2573
rect 24397 2533 24409 2567
rect 24443 2564 24455 2567
rect 24762 2564 24768 2576
rect 24443 2536 24768 2564
rect 24443 2533 24455 2536
rect 24397 2527 24455 2533
rect 22281 2499 22339 2505
rect 22281 2496 22293 2499
rect 22112 2468 22293 2496
rect 22281 2465 22293 2468
rect 22327 2496 22339 2499
rect 23477 2499 23535 2505
rect 22327 2468 22784 2496
rect 22327 2465 22339 2468
rect 22281 2459 22339 2465
rect 21634 2428 21640 2440
rect 12483 2400 12756 2428
rect 21595 2400 21640 2428
rect 12483 2397 12495 2400
rect 12437 2391 12495 2397
rect 21634 2388 21640 2400
rect 21692 2428 21698 2440
rect 22373 2431 22431 2437
rect 22373 2428 22385 2431
rect 21692 2400 22385 2428
rect 21692 2388 21698 2400
rect 22373 2397 22385 2400
rect 22419 2397 22431 2431
rect 22373 2391 22431 2397
rect 21818 2360 21824 2372
rect 21779 2332 21824 2360
rect 21818 2320 21824 2332
rect 21876 2320 21882 2372
rect 22756 2360 22784 2468
rect 23477 2465 23489 2499
rect 23523 2496 23535 2499
rect 23566 2496 23572 2508
rect 23523 2468 23572 2496
rect 23523 2465 23535 2468
rect 23477 2459 23535 2465
rect 23566 2456 23572 2468
rect 23624 2496 23630 2508
rect 24412 2496 24440 2527
rect 24762 2524 24768 2536
rect 24820 2524 24826 2576
rect 23624 2468 24440 2496
rect 24489 2499 24547 2505
rect 23624 2456 23630 2468
rect 24489 2465 24501 2499
rect 24535 2496 24547 2499
rect 24670 2496 24676 2508
rect 24535 2468 24676 2496
rect 24535 2465 24547 2468
rect 24489 2459 24547 2465
rect 23658 2388 23664 2440
rect 23716 2428 23722 2440
rect 23845 2431 23903 2437
rect 23845 2428 23857 2431
rect 23716 2400 23857 2428
rect 23716 2388 23722 2400
rect 23845 2397 23857 2400
rect 23891 2428 23903 2431
rect 24504 2428 24532 2459
rect 24670 2456 24676 2468
rect 24728 2456 24734 2508
rect 23891 2400 24532 2428
rect 23891 2397 23903 2400
rect 23845 2391 23903 2397
rect 24578 2388 24584 2440
rect 24636 2428 24642 2440
rect 25041 2431 25099 2437
rect 25041 2428 25053 2431
rect 24636 2400 25053 2428
rect 24636 2388 24642 2400
rect 25041 2397 25053 2400
rect 25087 2397 25099 2431
rect 25041 2391 25099 2397
rect 24029 2363 24087 2369
rect 24029 2360 24041 2363
rect 22756 2332 24041 2360
rect 24029 2329 24041 2332
rect 24075 2329 24087 2363
rect 24029 2323 24087 2329
rect 5905 2295 5963 2301
rect 5905 2261 5917 2295
rect 5951 2292 5963 2295
rect 6822 2292 6828 2304
rect 5951 2264 6828 2292
rect 5951 2261 5963 2264
rect 5905 2255 5963 2261
rect 6822 2252 6828 2264
rect 6880 2252 6886 2304
rect 7190 2292 7196 2304
rect 7151 2264 7196 2292
rect 7190 2252 7196 2264
rect 7248 2252 7254 2304
rect 9214 2292 9220 2304
rect 9175 2264 9220 2292
rect 9214 2252 9220 2264
rect 9272 2252 9278 2304
rect 13262 2252 13268 2304
rect 13320 2292 13326 2304
rect 18506 2292 18512 2304
rect 13320 2264 18512 2292
rect 13320 2252 13326 2264
rect 18506 2252 18512 2264
rect 18564 2252 18570 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 10042 1776 10048 1828
rect 10100 1816 10106 1828
rect 16758 1816 16764 1828
rect 10100 1788 16764 1816
rect 10100 1776 10106 1788
rect 16758 1776 16764 1788
rect 16816 1776 16822 1828
rect 10778 1232 10784 1284
rect 10836 1272 10842 1284
rect 13906 1272 13912 1284
rect 10836 1244 13912 1272
rect 10836 1232 10842 1244
rect 13906 1232 13912 1244
rect 13964 1232 13970 1284
rect 20070 552 20076 604
rect 20128 592 20134 604
rect 20438 592 20444 604
rect 20128 564 20444 592
rect 20128 552 20134 564
rect 20438 552 20444 564
rect 20496 552 20502 604
<< via1 >>
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 24768 24352 24820 24404
rect 25228 24216 25280 24268
rect 24768 24123 24820 24132
rect 24768 24089 24777 24123
rect 24777 24089 24811 24123
rect 24811 24089 24820 24123
rect 24768 24080 24820 24089
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 24676 23808 24728 23860
rect 24400 23715 24452 23724
rect 24400 23681 24409 23715
rect 24409 23681 24443 23715
rect 24443 23681 24452 23715
rect 24400 23672 24452 23681
rect 25228 23511 25280 23520
rect 25228 23477 25237 23511
rect 25237 23477 25271 23511
rect 25271 23477 25280 23511
rect 25228 23468 25280 23477
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 24124 23264 24176 23316
rect 12808 23239 12860 23248
rect 12808 23205 12817 23239
rect 12817 23205 12851 23239
rect 12851 23205 12860 23239
rect 12808 23196 12860 23205
rect 12532 23171 12584 23180
rect 12532 23137 12541 23171
rect 12541 23137 12575 23171
rect 12575 23137 12584 23171
rect 12532 23128 12584 23137
rect 23848 23128 23900 23180
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 24768 22763 24820 22772
rect 24768 22729 24777 22763
rect 24777 22729 24811 22763
rect 24811 22729 24820 22763
rect 24768 22720 24820 22729
rect 25228 22584 25280 22636
rect 26240 22584 26292 22636
rect 24584 22559 24636 22568
rect 24584 22525 24593 22559
rect 24593 22525 24627 22559
rect 24627 22525 24636 22559
rect 24584 22516 24636 22525
rect 11980 22380 12032 22432
rect 12532 22380 12584 22432
rect 23848 22380 23900 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 23848 22151 23900 22160
rect 23848 22117 23857 22151
rect 23857 22117 23891 22151
rect 23891 22117 23900 22151
rect 23848 22108 23900 22117
rect 23480 22040 23532 22092
rect 24860 22083 24912 22092
rect 24860 22049 24869 22083
rect 24869 22049 24903 22083
rect 24903 22049 24912 22083
rect 24860 22040 24912 22049
rect 23388 21972 23440 22024
rect 24216 21972 24268 22024
rect 25044 21947 25096 21956
rect 25044 21913 25053 21947
rect 25053 21913 25087 21947
rect 25087 21913 25096 21947
rect 25044 21904 25096 21913
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 24860 21675 24912 21684
rect 24860 21641 24869 21675
rect 24869 21641 24903 21675
rect 24903 21641 24912 21675
rect 24860 21632 24912 21641
rect 25136 21675 25188 21684
rect 25136 21641 25145 21675
rect 25145 21641 25179 21675
rect 25179 21641 25188 21675
rect 25136 21632 25188 21641
rect 14556 21539 14608 21548
rect 14556 21505 14565 21539
rect 14565 21505 14599 21539
rect 14599 21505 14608 21539
rect 14556 21496 14608 21505
rect 14004 21428 14056 21480
rect 23480 21471 23532 21480
rect 23480 21437 23489 21471
rect 23489 21437 23523 21471
rect 23523 21437 23532 21471
rect 23480 21428 23532 21437
rect 23572 21428 23624 21480
rect 23756 21428 23808 21480
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 25228 21088 25280 21140
rect 23848 20952 23900 21004
rect 24860 20995 24912 21004
rect 24860 20961 24869 20995
rect 24869 20961 24903 20995
rect 24903 20961 24912 20995
rect 24860 20952 24912 20961
rect 23756 20927 23808 20936
rect 23756 20893 23765 20927
rect 23765 20893 23799 20927
rect 23799 20893 23808 20927
rect 23756 20884 23808 20893
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 16856 20587 16908 20596
rect 16856 20553 16865 20587
rect 16865 20553 16899 20587
rect 16899 20553 16908 20587
rect 16856 20544 16908 20553
rect 24676 20544 24728 20596
rect 16580 20340 16632 20392
rect 23940 20340 23992 20392
rect 23848 20247 23900 20256
rect 23848 20213 23857 20247
rect 23857 20213 23891 20247
rect 23891 20213 23900 20247
rect 23848 20204 23900 20213
rect 25504 20247 25556 20256
rect 25504 20213 25513 20247
rect 25513 20213 25547 20247
rect 25547 20213 25556 20247
rect 25504 20204 25556 20213
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 17500 19932 17552 19984
rect 24860 19932 24912 19984
rect 25504 19932 25556 19984
rect 23480 19907 23532 19916
rect 23480 19873 23489 19907
rect 23489 19873 23523 19907
rect 23523 19873 23532 19907
rect 23480 19864 23532 19873
rect 17040 19839 17092 19848
rect 17040 19805 17049 19839
rect 17049 19805 17083 19839
rect 17083 19805 17092 19839
rect 17040 19796 17092 19805
rect 18236 19660 18288 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 17500 19456 17552 19508
rect 17040 19388 17092 19440
rect 17868 19388 17920 19440
rect 23940 19363 23992 19372
rect 23940 19329 23949 19363
rect 23949 19329 23983 19363
rect 23983 19329 23992 19363
rect 23940 19320 23992 19329
rect 15292 19252 15344 19304
rect 16488 19252 16540 19304
rect 23664 19295 23716 19304
rect 23664 19261 23673 19295
rect 23673 19261 23707 19295
rect 23707 19261 23716 19295
rect 23664 19252 23716 19261
rect 24952 19295 25004 19304
rect 24952 19261 24961 19295
rect 24961 19261 24995 19295
rect 24995 19261 25004 19295
rect 24952 19252 25004 19261
rect 26240 19252 26292 19304
rect 26884 19252 26936 19304
rect 23480 19159 23532 19168
rect 23480 19125 23489 19159
rect 23489 19125 23523 19159
rect 23523 19125 23532 19159
rect 23480 19116 23532 19125
rect 24860 19116 24912 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 24676 18912 24728 18964
rect 24584 18819 24636 18828
rect 24584 18785 24593 18819
rect 24593 18785 24627 18819
rect 24627 18785 24636 18819
rect 24584 18776 24636 18785
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 14832 18368 14884 18420
rect 24676 18411 24728 18420
rect 24676 18377 24685 18411
rect 24685 18377 24719 18411
rect 24719 18377 24728 18411
rect 24676 18368 24728 18377
rect 13544 18207 13596 18216
rect 13544 18173 13553 18207
rect 13553 18173 13587 18207
rect 13587 18173 13596 18207
rect 13544 18164 13596 18173
rect 13820 18139 13872 18148
rect 13820 18105 13829 18139
rect 13829 18105 13863 18139
rect 13863 18105 13872 18139
rect 13820 18096 13872 18105
rect 13912 18096 13964 18148
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 24768 17867 24820 17876
rect 24768 17833 24777 17867
rect 24777 17833 24811 17867
rect 24811 17833 24820 17867
rect 24768 17824 24820 17833
rect 11612 17799 11664 17808
rect 11612 17765 11621 17799
rect 11621 17765 11655 17799
rect 11655 17765 11664 17799
rect 11612 17756 11664 17765
rect 11428 17688 11480 17740
rect 25044 17688 25096 17740
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 24676 17280 24728 17332
rect 13728 17144 13780 17196
rect 13176 17119 13228 17128
rect 13176 17085 13185 17119
rect 13185 17085 13219 17119
rect 13219 17085 13228 17119
rect 13176 17076 13228 17085
rect 11520 16940 11572 16992
rect 23940 16940 23992 16992
rect 25044 16940 25096 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 22928 16779 22980 16788
rect 22928 16745 22937 16779
rect 22937 16745 22971 16779
rect 22971 16745 22980 16779
rect 22928 16736 22980 16745
rect 16580 16643 16632 16652
rect 16580 16609 16589 16643
rect 16589 16609 16623 16643
rect 16623 16609 16632 16643
rect 16580 16600 16632 16609
rect 22744 16643 22796 16652
rect 22744 16609 22753 16643
rect 22753 16609 22787 16643
rect 22787 16609 22796 16643
rect 22744 16600 22796 16609
rect 16488 16532 16540 16584
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 25136 16235 25188 16244
rect 25136 16201 25145 16235
rect 25145 16201 25179 16235
rect 25179 16201 25188 16235
rect 25136 16192 25188 16201
rect 23940 16099 23992 16108
rect 23940 16065 23949 16099
rect 23949 16065 23983 16099
rect 23983 16065 23992 16099
rect 23940 16056 23992 16065
rect 23664 16031 23716 16040
rect 23664 15997 23673 16031
rect 23673 15997 23707 16031
rect 23707 15997 23716 16031
rect 23664 15988 23716 15997
rect 24860 15988 24912 16040
rect 16488 15852 16540 15904
rect 22192 15852 22244 15904
rect 22744 15895 22796 15904
rect 22744 15861 22753 15895
rect 22753 15861 22787 15895
rect 22787 15861 22796 15895
rect 22744 15852 22796 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 23388 15691 23440 15700
rect 23388 15657 23397 15691
rect 23397 15657 23431 15691
rect 23431 15657 23440 15691
rect 23388 15648 23440 15657
rect 22192 15623 22244 15632
rect 22192 15589 22201 15623
rect 22201 15589 22235 15623
rect 22235 15589 22244 15623
rect 22192 15580 22244 15589
rect 21916 15555 21968 15564
rect 21916 15521 21925 15555
rect 21925 15521 21959 15555
rect 21959 15521 21968 15555
rect 21916 15512 21968 15521
rect 23204 15555 23256 15564
rect 23204 15521 23213 15555
rect 23213 15521 23247 15555
rect 23247 15521 23256 15555
rect 23204 15512 23256 15521
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 25872 15147 25924 15156
rect 25872 15113 25881 15147
rect 25881 15113 25915 15147
rect 25915 15113 25924 15147
rect 25872 15104 25924 15113
rect 24768 14968 24820 15020
rect 23848 14900 23900 14952
rect 25872 14900 25924 14952
rect 21916 14807 21968 14816
rect 21916 14773 21925 14807
rect 21925 14773 21959 14807
rect 21959 14773 21968 14807
rect 21916 14764 21968 14773
rect 22468 14764 22520 14816
rect 23204 14807 23256 14816
rect 23204 14773 23213 14807
rect 23213 14773 23247 14807
rect 23247 14773 23256 14807
rect 23204 14764 23256 14773
rect 25688 14764 25740 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 24676 14560 24728 14612
rect 22468 14535 22520 14544
rect 22468 14501 22477 14535
rect 22477 14501 22511 14535
rect 22511 14501 22520 14535
rect 22468 14492 22520 14501
rect 22744 14424 22796 14476
rect 24676 14424 24728 14476
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 17868 14016 17920 14068
rect 18328 14016 18380 14068
rect 24676 14059 24728 14068
rect 24676 14025 24685 14059
rect 24685 14025 24719 14059
rect 24719 14025 24728 14059
rect 24676 14016 24728 14025
rect 25596 14059 25648 14068
rect 25596 14025 25605 14059
rect 25605 14025 25639 14059
rect 25639 14025 25648 14059
rect 25596 14016 25648 14025
rect 25136 13991 25188 14000
rect 25136 13957 25145 13991
rect 25145 13957 25179 13991
rect 25179 13957 25188 13991
rect 25136 13948 25188 13957
rect 22744 13812 22796 13864
rect 24032 13812 24084 13864
rect 25596 13812 25648 13864
rect 19248 13719 19300 13728
rect 19248 13685 19257 13719
rect 19257 13685 19291 13719
rect 19291 13685 19300 13719
rect 19248 13676 19300 13685
rect 19524 13676 19576 13728
rect 21640 13676 21692 13728
rect 22100 13719 22152 13728
rect 22100 13685 22109 13719
rect 22109 13685 22143 13719
rect 22143 13685 22152 13719
rect 22100 13676 22152 13685
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 19156 13472 19208 13524
rect 24216 13472 24268 13524
rect 18512 13336 18564 13388
rect 19524 13336 19576 13388
rect 23480 13379 23532 13388
rect 23480 13345 23489 13379
rect 23489 13345 23523 13379
rect 23523 13345 23532 13379
rect 23480 13336 23532 13345
rect 24676 13336 24728 13388
rect 19248 13268 19300 13320
rect 20076 13268 20128 13320
rect 21548 13268 21600 13320
rect 22560 13268 22612 13320
rect 19524 13200 19576 13252
rect 23664 13243 23716 13252
rect 23664 13209 23673 13243
rect 23673 13209 23707 13243
rect 23707 13209 23716 13243
rect 23664 13200 23716 13209
rect 19432 13132 19484 13184
rect 21180 13175 21232 13184
rect 21180 13141 21189 13175
rect 21189 13141 21223 13175
rect 21223 13141 21232 13175
rect 21180 13132 21232 13141
rect 23940 13132 23992 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 18512 12971 18564 12980
rect 18512 12937 18521 12971
rect 18521 12937 18555 12971
rect 18555 12937 18564 12971
rect 18512 12928 18564 12937
rect 19248 12928 19300 12980
rect 21272 12928 21324 12980
rect 23480 12971 23532 12980
rect 23480 12937 23489 12971
rect 23489 12937 23523 12971
rect 23523 12937 23532 12971
rect 23480 12928 23532 12937
rect 19340 12860 19392 12912
rect 22652 12903 22704 12912
rect 19524 12835 19576 12844
rect 19524 12801 19533 12835
rect 19533 12801 19567 12835
rect 19567 12801 19576 12835
rect 19524 12792 19576 12801
rect 21180 12792 21232 12844
rect 22652 12869 22661 12903
rect 22661 12869 22695 12903
rect 22695 12869 22704 12903
rect 22652 12860 22704 12869
rect 23940 12928 23992 12980
rect 24676 12971 24728 12980
rect 24676 12937 24685 12971
rect 24685 12937 24719 12971
rect 24719 12937 24728 12971
rect 24676 12928 24728 12937
rect 24952 12928 25004 12980
rect 19156 12724 19208 12776
rect 19432 12767 19484 12776
rect 19432 12733 19441 12767
rect 19441 12733 19475 12767
rect 19475 12733 19484 12767
rect 19432 12724 19484 12733
rect 18788 12699 18840 12708
rect 18788 12665 18797 12699
rect 18797 12665 18831 12699
rect 18831 12665 18840 12699
rect 18788 12656 18840 12665
rect 21364 12656 21416 12708
rect 16212 12588 16264 12640
rect 20536 12588 20588 12640
rect 21272 12588 21324 12640
rect 21732 12631 21784 12640
rect 21732 12597 21741 12631
rect 21741 12597 21775 12631
rect 21775 12597 21784 12631
rect 21732 12588 21784 12597
rect 24952 12767 25004 12776
rect 24952 12733 24961 12767
rect 24961 12733 24995 12767
rect 24995 12733 25004 12767
rect 24952 12724 25004 12733
rect 23388 12588 23440 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 17132 12427 17184 12436
rect 17132 12393 17141 12427
rect 17141 12393 17175 12427
rect 17175 12393 17184 12427
rect 17132 12384 17184 12393
rect 18328 12384 18380 12436
rect 19064 12427 19116 12436
rect 19064 12393 19073 12427
rect 19073 12393 19107 12427
rect 19107 12393 19116 12427
rect 19064 12384 19116 12393
rect 22744 12384 22796 12436
rect 19248 12316 19300 12368
rect 19340 12316 19392 12368
rect 20076 12316 20128 12368
rect 21180 12359 21232 12368
rect 21180 12325 21214 12359
rect 21214 12325 21232 12359
rect 21180 12316 21232 12325
rect 24952 12359 25004 12368
rect 24952 12325 24961 12359
rect 24961 12325 24995 12359
rect 24995 12325 25004 12359
rect 24952 12316 25004 12325
rect 17408 12248 17460 12300
rect 17592 12291 17644 12300
rect 17592 12257 17601 12291
rect 17601 12257 17635 12291
rect 17635 12257 17644 12291
rect 19432 12291 19484 12300
rect 17592 12248 17644 12257
rect 19432 12257 19441 12291
rect 19441 12257 19475 12291
rect 19475 12257 19484 12291
rect 19432 12248 19484 12257
rect 17684 12223 17736 12232
rect 17684 12189 17693 12223
rect 17693 12189 17727 12223
rect 17727 12189 17736 12223
rect 17684 12180 17736 12189
rect 19616 12223 19668 12232
rect 19616 12189 19625 12223
rect 19625 12189 19659 12223
rect 19659 12189 19668 12223
rect 21732 12248 21784 12300
rect 24676 12291 24728 12300
rect 24676 12257 24685 12291
rect 24685 12257 24719 12291
rect 24719 12257 24728 12291
rect 24676 12248 24728 12257
rect 19616 12180 19668 12189
rect 18604 12087 18656 12096
rect 18604 12053 18613 12087
rect 18613 12053 18647 12087
rect 18647 12053 18656 12087
rect 18604 12044 18656 12053
rect 20168 12044 20220 12096
rect 21272 12044 21324 12096
rect 22284 12087 22336 12096
rect 22284 12053 22293 12087
rect 22293 12053 22327 12087
rect 22327 12053 22336 12087
rect 22284 12044 22336 12053
rect 22928 12087 22980 12096
rect 22928 12053 22937 12087
rect 22937 12053 22971 12087
rect 22971 12053 22980 12087
rect 23664 12223 23716 12232
rect 23664 12189 23673 12223
rect 23673 12189 23707 12223
rect 23707 12189 23716 12223
rect 23664 12180 23716 12189
rect 24216 12087 24268 12096
rect 22928 12044 22980 12053
rect 24216 12053 24225 12087
rect 24225 12053 24259 12087
rect 24259 12053 24268 12087
rect 24216 12044 24268 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 16856 11883 16908 11892
rect 16856 11849 16865 11883
rect 16865 11849 16899 11883
rect 16899 11849 16908 11883
rect 16856 11840 16908 11849
rect 17592 11840 17644 11892
rect 17684 11840 17736 11892
rect 17960 11840 18012 11892
rect 21180 11840 21232 11892
rect 21364 11840 21416 11892
rect 22376 11840 22428 11892
rect 24676 11840 24728 11892
rect 19432 11704 19484 11756
rect 22652 11747 22704 11756
rect 22652 11713 22661 11747
rect 22661 11713 22695 11747
rect 22695 11713 22704 11747
rect 22652 11704 22704 11713
rect 15660 11636 15712 11688
rect 16120 11636 16172 11688
rect 18328 11636 18380 11688
rect 18880 11636 18932 11688
rect 20168 11636 20220 11688
rect 15476 11611 15528 11620
rect 15476 11577 15485 11611
rect 15485 11577 15519 11611
rect 15519 11577 15528 11611
rect 15476 11568 15528 11577
rect 19340 11568 19392 11620
rect 19616 11568 19668 11620
rect 20260 11568 20312 11620
rect 24216 11636 24268 11688
rect 16028 11543 16080 11552
rect 16028 11509 16037 11543
rect 16037 11509 16071 11543
rect 16071 11509 16080 11543
rect 16028 11500 16080 11509
rect 16120 11500 16172 11552
rect 17408 11543 17460 11552
rect 17408 11509 17417 11543
rect 17417 11509 17451 11543
rect 17451 11509 17460 11543
rect 17408 11500 17460 11509
rect 22192 11500 22244 11552
rect 22376 11543 22428 11552
rect 22376 11509 22385 11543
rect 22385 11509 22419 11543
rect 22419 11509 22428 11543
rect 22376 11500 22428 11509
rect 23388 11500 23440 11552
rect 24768 11500 24820 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 15292 11339 15344 11348
rect 15292 11305 15301 11339
rect 15301 11305 15335 11339
rect 15335 11305 15344 11339
rect 15292 11296 15344 11305
rect 20260 11339 20312 11348
rect 20260 11305 20269 11339
rect 20269 11305 20303 11339
rect 20303 11305 20312 11339
rect 20260 11296 20312 11305
rect 20536 11339 20588 11348
rect 20536 11305 20545 11339
rect 20545 11305 20579 11339
rect 20579 11305 20588 11339
rect 20536 11296 20588 11305
rect 21180 11339 21232 11348
rect 21180 11305 21189 11339
rect 21189 11305 21223 11339
rect 21223 11305 21232 11339
rect 21180 11296 21232 11305
rect 22652 11339 22704 11348
rect 22652 11305 22661 11339
rect 22661 11305 22695 11339
rect 22695 11305 22704 11339
rect 22652 11296 22704 11305
rect 23664 11296 23716 11348
rect 24216 11228 24268 11280
rect 15384 11160 15436 11212
rect 17040 11203 17092 11212
rect 17040 11169 17049 11203
rect 17049 11169 17083 11203
rect 17083 11169 17092 11203
rect 17040 11160 17092 11169
rect 18880 11203 18932 11212
rect 18880 11169 18889 11203
rect 18889 11169 18923 11203
rect 18923 11169 18932 11203
rect 18880 11160 18932 11169
rect 19156 11203 19208 11212
rect 19156 11169 19190 11203
rect 19190 11169 19208 11203
rect 19156 11160 19208 11169
rect 21364 11160 21416 11212
rect 22284 11160 22336 11212
rect 23480 11203 23532 11212
rect 23480 11169 23489 11203
rect 23489 11169 23523 11203
rect 23523 11169 23532 11203
rect 23480 11160 23532 11169
rect 23572 11160 23624 11212
rect 24768 11160 24820 11212
rect 13728 11092 13780 11144
rect 15292 11092 15344 11144
rect 15844 11135 15896 11144
rect 15844 11101 15853 11135
rect 15853 11101 15887 11135
rect 15887 11101 15896 11135
rect 15844 11092 15896 11101
rect 20168 11092 20220 11144
rect 14740 11024 14792 11076
rect 22376 11024 22428 11076
rect 16672 10956 16724 11008
rect 17132 10956 17184 11008
rect 18052 10956 18104 11008
rect 24216 10956 24268 11008
rect 24860 10999 24912 11008
rect 24860 10965 24869 10999
rect 24869 10965 24903 10999
rect 24903 10965 24912 10999
rect 24860 10956 24912 10965
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 16212 10752 16264 10804
rect 16672 10752 16724 10804
rect 16856 10795 16908 10804
rect 16856 10761 16865 10795
rect 16865 10761 16899 10795
rect 16899 10761 16908 10795
rect 16856 10752 16908 10761
rect 19156 10752 19208 10804
rect 15292 10684 15344 10736
rect 16396 10684 16448 10736
rect 14924 10659 14976 10668
rect 14924 10625 14933 10659
rect 14933 10625 14967 10659
rect 14967 10625 14976 10659
rect 14924 10616 14976 10625
rect 17408 10659 17460 10668
rect 13084 10591 13136 10600
rect 13084 10557 13093 10591
rect 13093 10557 13127 10591
rect 13127 10557 13136 10591
rect 13084 10548 13136 10557
rect 16212 10548 16264 10600
rect 12624 10480 12676 10532
rect 17408 10625 17417 10659
rect 17417 10625 17451 10659
rect 17451 10625 17460 10659
rect 17408 10616 17460 10625
rect 19340 10684 19392 10736
rect 17592 10548 17644 10600
rect 18880 10548 18932 10600
rect 18696 10480 18748 10532
rect 20536 10616 20588 10668
rect 21364 10752 21416 10804
rect 22100 10752 22152 10804
rect 24768 10795 24820 10804
rect 24768 10761 24777 10795
rect 24777 10761 24811 10795
rect 24811 10761 24820 10795
rect 24768 10752 24820 10761
rect 25412 10795 25464 10804
rect 25412 10761 25421 10795
rect 25421 10761 25455 10795
rect 25455 10761 25464 10795
rect 25412 10752 25464 10761
rect 20904 10684 20956 10736
rect 22192 10616 22244 10668
rect 22560 10616 22612 10668
rect 23572 10684 23624 10736
rect 23480 10616 23532 10668
rect 24860 10616 24912 10668
rect 22100 10548 22152 10600
rect 24124 10591 24176 10600
rect 24124 10557 24133 10591
rect 24133 10557 24167 10591
rect 24167 10557 24176 10591
rect 24124 10548 24176 10557
rect 25228 10591 25280 10600
rect 25228 10557 25237 10591
rect 25237 10557 25271 10591
rect 25271 10557 25280 10591
rect 25228 10548 25280 10557
rect 13820 10455 13872 10464
rect 13820 10421 13829 10455
rect 13829 10421 13863 10455
rect 13863 10421 13872 10455
rect 13820 10412 13872 10421
rect 14280 10455 14332 10464
rect 14280 10421 14289 10455
rect 14289 10421 14323 10455
rect 14323 10421 14332 10455
rect 14280 10412 14332 10421
rect 15384 10455 15436 10464
rect 15384 10421 15393 10455
rect 15393 10421 15427 10455
rect 15427 10421 15436 10455
rect 15384 10412 15436 10421
rect 16120 10412 16172 10464
rect 17132 10412 17184 10464
rect 20260 10455 20312 10464
rect 20260 10421 20269 10455
rect 20269 10421 20303 10455
rect 20303 10421 20312 10455
rect 20260 10412 20312 10421
rect 23940 10412 23992 10464
rect 24124 10412 24176 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 12900 10251 12952 10260
rect 12900 10217 12909 10251
rect 12909 10217 12943 10251
rect 12943 10217 12952 10251
rect 12900 10208 12952 10217
rect 14924 10208 14976 10260
rect 15292 10208 15344 10260
rect 15844 10208 15896 10260
rect 17040 10208 17092 10260
rect 17960 10208 18012 10260
rect 18604 10251 18656 10260
rect 13912 10115 13964 10124
rect 13912 10081 13921 10115
rect 13921 10081 13955 10115
rect 13955 10081 13964 10115
rect 13912 10072 13964 10081
rect 14188 10115 14240 10124
rect 14188 10081 14197 10115
rect 14197 10081 14231 10115
rect 14231 10081 14240 10115
rect 14188 10072 14240 10081
rect 17592 10140 17644 10192
rect 18604 10217 18613 10251
rect 18613 10217 18647 10251
rect 18647 10217 18656 10251
rect 18604 10208 18656 10217
rect 18696 10208 18748 10260
rect 20168 10251 20220 10260
rect 20168 10217 20177 10251
rect 20177 10217 20211 10251
rect 20211 10217 20220 10251
rect 20168 10208 20220 10217
rect 21272 10251 21324 10260
rect 21272 10217 21281 10251
rect 21281 10217 21315 10251
rect 21315 10217 21324 10251
rect 21272 10208 21324 10217
rect 21640 10251 21692 10260
rect 21640 10217 21649 10251
rect 21649 10217 21683 10251
rect 21683 10217 21692 10251
rect 21640 10208 21692 10217
rect 22192 10208 22244 10260
rect 20260 10140 20312 10192
rect 16396 10115 16448 10124
rect 16396 10081 16430 10115
rect 16430 10081 16448 10115
rect 16396 10072 16448 10081
rect 18052 10072 18104 10124
rect 18604 10072 18656 10124
rect 19064 10115 19116 10124
rect 19064 10081 19073 10115
rect 19073 10081 19107 10115
rect 19107 10081 19116 10115
rect 21916 10140 21968 10192
rect 22560 10140 22612 10192
rect 23480 10140 23532 10192
rect 19064 10072 19116 10081
rect 23296 10115 23348 10124
rect 23296 10081 23305 10115
rect 23305 10081 23339 10115
rect 23339 10081 23348 10115
rect 23296 10072 23348 10081
rect 19156 10047 19208 10056
rect 19156 10013 19165 10047
rect 19165 10013 19199 10047
rect 19199 10013 19208 10047
rect 19156 10004 19208 10013
rect 19708 10004 19760 10056
rect 18696 9936 18748 9988
rect 22008 10004 22060 10056
rect 19156 9868 19208 9920
rect 24216 9868 24268 9920
rect 24952 9911 25004 9920
rect 24952 9877 24961 9911
rect 24961 9877 24995 9911
rect 24995 9877 25004 9911
rect 24952 9868 25004 9877
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 13912 9664 13964 9716
rect 16948 9707 17000 9716
rect 16948 9673 16957 9707
rect 16957 9673 16991 9707
rect 16991 9673 17000 9707
rect 16948 9664 17000 9673
rect 17408 9664 17460 9716
rect 19248 9664 19300 9716
rect 19708 9707 19760 9716
rect 19708 9673 19717 9707
rect 19717 9673 19751 9707
rect 19751 9673 19760 9707
rect 19708 9664 19760 9673
rect 14740 9596 14792 9648
rect 13360 9528 13412 9580
rect 13728 9460 13780 9512
rect 18052 9596 18104 9648
rect 19524 9596 19576 9648
rect 20076 9639 20128 9648
rect 20076 9605 20085 9639
rect 20085 9605 20119 9639
rect 20119 9605 20128 9639
rect 20076 9596 20128 9605
rect 23112 9639 23164 9648
rect 23112 9605 23121 9639
rect 23121 9605 23155 9639
rect 23155 9605 23164 9639
rect 23112 9596 23164 9605
rect 17868 9571 17920 9580
rect 17868 9537 17877 9571
rect 17877 9537 17911 9571
rect 17911 9537 17920 9571
rect 17868 9528 17920 9537
rect 14924 9460 14976 9512
rect 17224 9503 17276 9512
rect 17224 9469 17233 9503
rect 17233 9469 17267 9503
rect 17267 9469 17276 9503
rect 17224 9460 17276 9469
rect 17684 9460 17736 9512
rect 19156 9460 19208 9512
rect 20168 9460 20220 9512
rect 20352 9460 20404 9512
rect 21640 9460 21692 9512
rect 23296 9528 23348 9580
rect 24952 9460 25004 9512
rect 14740 9435 14792 9444
rect 14740 9401 14749 9435
rect 14749 9401 14783 9435
rect 14783 9401 14792 9435
rect 14740 9392 14792 9401
rect 17960 9392 18012 9444
rect 24768 9392 24820 9444
rect 12992 9324 13044 9376
rect 16396 9324 16448 9376
rect 16580 9367 16632 9376
rect 16580 9333 16589 9367
rect 16589 9333 16623 9367
rect 16623 9333 16632 9367
rect 16580 9324 16632 9333
rect 17040 9367 17092 9376
rect 17040 9333 17049 9367
rect 17049 9333 17083 9367
rect 17083 9333 17092 9367
rect 17040 9324 17092 9333
rect 21640 9367 21692 9376
rect 21640 9333 21649 9367
rect 21649 9333 21683 9367
rect 21683 9333 21692 9367
rect 21640 9324 21692 9333
rect 21916 9367 21968 9376
rect 21916 9333 21925 9367
rect 21925 9333 21959 9367
rect 21959 9333 21968 9367
rect 21916 9324 21968 9333
rect 22652 9367 22704 9376
rect 22652 9333 22661 9367
rect 22661 9333 22695 9367
rect 22695 9333 22704 9367
rect 22652 9324 22704 9333
rect 23204 9324 23256 9376
rect 23756 9324 23808 9376
rect 25136 9367 25188 9376
rect 25136 9333 25145 9367
rect 25145 9333 25179 9367
rect 25179 9333 25188 9367
rect 25136 9324 25188 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 11980 9163 12032 9172
rect 11980 9129 11989 9163
rect 11989 9129 12023 9163
rect 12023 9129 12032 9163
rect 11980 9120 12032 9129
rect 13360 9163 13412 9172
rect 13360 9129 13369 9163
rect 13369 9129 13403 9163
rect 13403 9129 13412 9163
rect 13360 9120 13412 9129
rect 13544 9163 13596 9172
rect 13544 9129 13553 9163
rect 13553 9129 13587 9163
rect 13587 9129 13596 9163
rect 13544 9120 13596 9129
rect 17960 9120 18012 9172
rect 20260 9163 20312 9172
rect 20260 9129 20269 9163
rect 20269 9129 20303 9163
rect 20303 9129 20312 9163
rect 20260 9120 20312 9129
rect 21180 9163 21232 9172
rect 21180 9129 21189 9163
rect 21189 9129 21223 9163
rect 21223 9129 21232 9163
rect 21180 9120 21232 9129
rect 23388 9120 23440 9172
rect 16948 9095 17000 9104
rect 16948 9061 16982 9095
rect 16982 9061 17000 9095
rect 16948 9052 17000 9061
rect 19432 9052 19484 9104
rect 22468 9052 22520 9104
rect 24676 9052 24728 9104
rect 12348 9027 12400 9036
rect 12348 8993 12357 9027
rect 12357 8993 12391 9027
rect 12391 8993 12400 9027
rect 12348 8984 12400 8993
rect 13452 8984 13504 9036
rect 14556 8984 14608 9036
rect 15476 8984 15528 9036
rect 17684 8984 17736 9036
rect 18972 8984 19024 9036
rect 21272 8984 21324 9036
rect 23296 8984 23348 9036
rect 24216 8984 24268 9036
rect 11244 8916 11296 8968
rect 12256 8848 12308 8900
rect 13176 8848 13228 8900
rect 14924 8848 14976 8900
rect 15752 8891 15804 8900
rect 15752 8857 15761 8891
rect 15761 8857 15795 8891
rect 15795 8857 15804 8891
rect 15752 8848 15804 8857
rect 19248 8848 19300 8900
rect 21456 8916 21508 8968
rect 22008 8916 22060 8968
rect 13544 8780 13596 8832
rect 15292 8780 15344 8832
rect 16028 8780 16080 8832
rect 16672 8780 16724 8832
rect 17868 8780 17920 8832
rect 18604 8823 18656 8832
rect 18604 8789 18613 8823
rect 18613 8789 18647 8823
rect 18647 8789 18656 8823
rect 18604 8780 18656 8789
rect 18880 8823 18932 8832
rect 18880 8789 18889 8823
rect 18889 8789 18923 8823
rect 18923 8789 18932 8823
rect 18880 8780 18932 8789
rect 19340 8780 19392 8832
rect 23572 8780 23624 8832
rect 25136 8848 25188 8900
rect 24768 8823 24820 8832
rect 24768 8789 24777 8823
rect 24777 8789 24811 8823
rect 24811 8789 24820 8823
rect 24768 8780 24820 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 10968 8576 11020 8628
rect 11244 8619 11296 8628
rect 11244 8585 11253 8619
rect 11253 8585 11287 8619
rect 11287 8585 11296 8619
rect 11244 8576 11296 8585
rect 12348 8576 12400 8628
rect 13176 8619 13228 8628
rect 13176 8585 13185 8619
rect 13185 8585 13219 8619
rect 13219 8585 13228 8619
rect 13176 8576 13228 8585
rect 14740 8576 14792 8628
rect 16120 8619 16172 8628
rect 16120 8585 16129 8619
rect 16129 8585 16163 8619
rect 16163 8585 16172 8619
rect 16120 8576 16172 8585
rect 16948 8576 17000 8628
rect 19432 8576 19484 8628
rect 20352 8576 20404 8628
rect 20720 8619 20772 8628
rect 20720 8585 20729 8619
rect 20729 8585 20763 8619
rect 20763 8585 20772 8619
rect 20720 8576 20772 8585
rect 21272 8619 21324 8628
rect 21272 8585 21281 8619
rect 21281 8585 21315 8619
rect 21315 8585 21324 8619
rect 21272 8576 21324 8585
rect 23480 8619 23532 8628
rect 23480 8585 23489 8619
rect 23489 8585 23523 8619
rect 23523 8585 23532 8619
rect 23480 8576 23532 8585
rect 24216 8576 24268 8628
rect 12532 8440 12584 8492
rect 13544 8440 13596 8492
rect 16580 8440 16632 8492
rect 20352 8440 20404 8492
rect 21272 8440 21324 8492
rect 13452 8415 13504 8424
rect 13452 8381 13461 8415
rect 13461 8381 13495 8415
rect 13495 8381 13504 8415
rect 13452 8372 13504 8381
rect 15016 8372 15068 8424
rect 15292 8372 15344 8424
rect 11980 8304 12032 8356
rect 14004 8304 14056 8356
rect 15476 8304 15528 8356
rect 15752 8304 15804 8356
rect 16120 8372 16172 8424
rect 19156 8372 19208 8424
rect 20720 8372 20772 8424
rect 21732 8372 21784 8424
rect 23940 8440 23992 8492
rect 24216 8483 24268 8492
rect 24216 8449 24225 8483
rect 24225 8449 24259 8483
rect 24259 8449 24268 8483
rect 24216 8440 24268 8449
rect 17040 8304 17092 8356
rect 18972 8347 19024 8356
rect 18972 8313 18981 8347
rect 18981 8313 19015 8347
rect 19015 8313 19024 8347
rect 18972 8304 19024 8313
rect 19524 8304 19576 8356
rect 15292 8236 15344 8288
rect 16672 8236 16724 8288
rect 18052 8279 18104 8288
rect 18052 8245 18061 8279
rect 18061 8245 18095 8279
rect 18095 8245 18104 8279
rect 18052 8236 18104 8245
rect 21456 8304 21508 8356
rect 23480 8304 23532 8356
rect 25504 8347 25556 8356
rect 25504 8313 25513 8347
rect 25513 8313 25547 8347
rect 25547 8313 25556 8347
rect 25504 8304 25556 8313
rect 21916 8236 21968 8288
rect 25136 8279 25188 8288
rect 25136 8245 25145 8279
rect 25145 8245 25179 8279
rect 25179 8245 25188 8279
rect 25136 8236 25188 8245
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 10692 8032 10744 8084
rect 10968 8075 11020 8084
rect 10968 8041 10977 8075
rect 10977 8041 11011 8075
rect 11011 8041 11020 8075
rect 10968 8032 11020 8041
rect 14372 8032 14424 8084
rect 16948 8075 17000 8084
rect 12256 7964 12308 8016
rect 15844 8007 15896 8016
rect 15844 7973 15878 8007
rect 15878 7973 15896 8007
rect 15844 7964 15896 7973
rect 16948 8041 16957 8075
rect 16957 8041 16991 8075
rect 16991 8041 17000 8075
rect 16948 8032 17000 8041
rect 17224 8075 17276 8084
rect 17224 8041 17233 8075
rect 17233 8041 17267 8075
rect 17267 8041 17276 8075
rect 17224 8032 17276 8041
rect 17684 8075 17736 8084
rect 17684 8041 17693 8075
rect 17693 8041 17727 8075
rect 17727 8041 17736 8075
rect 17684 8032 17736 8041
rect 18512 8075 18564 8084
rect 18512 8041 18521 8075
rect 18521 8041 18555 8075
rect 18555 8041 18564 8075
rect 18512 8032 18564 8041
rect 19524 8075 19576 8084
rect 19524 8041 19533 8075
rect 19533 8041 19567 8075
rect 19567 8041 19576 8075
rect 19524 8032 19576 8041
rect 21732 8032 21784 8084
rect 22008 8075 22060 8084
rect 22008 8041 22017 8075
rect 22017 8041 22051 8075
rect 22051 8041 22060 8075
rect 22008 8032 22060 8041
rect 22744 8032 22796 8084
rect 25136 8075 25188 8084
rect 25136 8041 25145 8075
rect 25145 8041 25179 8075
rect 25179 8041 25188 8075
rect 25136 8032 25188 8041
rect 20812 7964 20864 8016
rect 21640 7964 21692 8016
rect 22836 7964 22888 8016
rect 24216 7964 24268 8016
rect 11796 7896 11848 7948
rect 14648 7896 14700 7948
rect 15016 7939 15068 7948
rect 15016 7905 15025 7939
rect 15025 7905 15059 7939
rect 15059 7905 15068 7939
rect 15016 7896 15068 7905
rect 17960 7896 18012 7948
rect 20260 7939 20312 7948
rect 20260 7905 20269 7939
rect 20269 7905 20303 7939
rect 20303 7905 20312 7939
rect 20260 7896 20312 7905
rect 11060 7828 11112 7880
rect 11612 7871 11664 7880
rect 11612 7837 11621 7871
rect 11621 7837 11655 7871
rect 11655 7837 11664 7871
rect 11612 7828 11664 7837
rect 12532 7871 12584 7880
rect 11336 7692 11388 7744
rect 12532 7837 12541 7871
rect 12541 7837 12575 7871
rect 12575 7837 12584 7871
rect 12532 7828 12584 7837
rect 15476 7828 15528 7880
rect 18972 7871 19024 7880
rect 18972 7837 18981 7871
rect 18981 7837 19015 7871
rect 19015 7837 19024 7871
rect 18972 7828 19024 7837
rect 19064 7871 19116 7880
rect 19064 7837 19073 7871
rect 19073 7837 19107 7871
rect 19107 7837 19116 7871
rect 19064 7828 19116 7837
rect 20352 7828 20404 7880
rect 23204 7896 23256 7948
rect 23480 7896 23532 7948
rect 24124 7896 24176 7948
rect 25412 7896 25464 7948
rect 21640 7828 21692 7880
rect 23020 7828 23072 7880
rect 24768 7871 24820 7880
rect 24768 7837 24777 7871
rect 24777 7837 24811 7871
rect 24811 7837 24820 7871
rect 24768 7828 24820 7837
rect 19984 7803 20036 7812
rect 19984 7769 19993 7803
rect 19993 7769 20027 7803
rect 20027 7769 20036 7803
rect 19984 7760 20036 7769
rect 21088 7760 21140 7812
rect 14004 7692 14056 7744
rect 14556 7735 14608 7744
rect 14556 7701 14565 7735
rect 14565 7701 14599 7735
rect 14599 7701 14608 7735
rect 14556 7692 14608 7701
rect 17960 7735 18012 7744
rect 17960 7701 17969 7735
rect 17969 7701 18003 7735
rect 18003 7701 18012 7735
rect 17960 7692 18012 7701
rect 19248 7692 19300 7744
rect 20720 7692 20772 7744
rect 22192 7692 22244 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 4160 7488 4212 7540
rect 5448 7488 5500 7540
rect 12256 7531 12308 7540
rect 12256 7497 12265 7531
rect 12265 7497 12299 7531
rect 12299 7497 12308 7531
rect 12256 7488 12308 7497
rect 12992 7531 13044 7540
rect 12992 7497 13001 7531
rect 13001 7497 13035 7531
rect 13035 7497 13044 7531
rect 12992 7488 13044 7497
rect 14004 7531 14056 7540
rect 14004 7497 14013 7531
rect 14013 7497 14047 7531
rect 14047 7497 14056 7531
rect 14004 7488 14056 7497
rect 15844 7488 15896 7540
rect 17408 7531 17460 7540
rect 17408 7497 17417 7531
rect 17417 7497 17451 7531
rect 17451 7497 17460 7531
rect 17408 7488 17460 7497
rect 19064 7488 19116 7540
rect 19524 7488 19576 7540
rect 20628 7531 20680 7540
rect 20628 7497 20637 7531
rect 20637 7497 20671 7531
rect 20671 7497 20680 7531
rect 20628 7488 20680 7497
rect 22836 7488 22888 7540
rect 23020 7531 23072 7540
rect 23020 7497 23029 7531
rect 23029 7497 23063 7531
rect 23063 7497 23072 7531
rect 23020 7488 23072 7497
rect 25412 7531 25464 7540
rect 25412 7497 25421 7531
rect 25421 7497 25455 7531
rect 25455 7497 25464 7531
rect 25412 7488 25464 7497
rect 12808 7395 12860 7404
rect 12808 7361 12817 7395
rect 12817 7361 12851 7395
rect 12851 7361 12860 7395
rect 12808 7352 12860 7361
rect 19432 7420 19484 7472
rect 14372 7284 14424 7336
rect 14832 7327 14884 7336
rect 14832 7293 14866 7327
rect 14866 7293 14884 7327
rect 14832 7284 14884 7293
rect 17408 7284 17460 7336
rect 17592 7284 17644 7336
rect 19156 7284 19208 7336
rect 19984 7284 20036 7336
rect 21180 7395 21232 7404
rect 21180 7361 21189 7395
rect 21189 7361 21223 7395
rect 21223 7361 21232 7395
rect 21180 7352 21232 7361
rect 22376 7395 22428 7404
rect 22376 7361 22385 7395
rect 22385 7361 22419 7395
rect 22419 7361 22428 7395
rect 22376 7352 22428 7361
rect 23204 7352 23256 7404
rect 23572 7352 23624 7404
rect 22192 7327 22244 7336
rect 22192 7293 22201 7327
rect 22201 7293 22235 7327
rect 22235 7293 22244 7327
rect 22192 7284 22244 7293
rect 10784 7216 10836 7268
rect 11336 7148 11388 7200
rect 11612 7148 11664 7200
rect 11796 7191 11848 7200
rect 11796 7157 11805 7191
rect 11805 7157 11839 7191
rect 11839 7157 11848 7191
rect 11796 7148 11848 7157
rect 13452 7191 13504 7200
rect 13452 7157 13461 7191
rect 13461 7157 13495 7191
rect 13495 7157 13504 7191
rect 13452 7148 13504 7157
rect 16580 7191 16632 7200
rect 16580 7157 16589 7191
rect 16589 7157 16623 7191
rect 16623 7157 16632 7191
rect 16580 7148 16632 7157
rect 16672 7148 16724 7200
rect 17684 7148 17736 7200
rect 23664 7216 23716 7268
rect 20352 7148 20404 7200
rect 20996 7191 21048 7200
rect 20996 7157 21005 7191
rect 21005 7157 21039 7191
rect 21039 7157 21048 7191
rect 20996 7148 21048 7157
rect 21732 7191 21784 7200
rect 21732 7157 21741 7191
rect 21741 7157 21775 7191
rect 21775 7157 21784 7191
rect 21732 7148 21784 7157
rect 23480 7191 23532 7200
rect 23480 7157 23489 7191
rect 23489 7157 23523 7191
rect 23523 7157 23532 7191
rect 23480 7148 23532 7157
rect 25044 7191 25096 7200
rect 25044 7157 25053 7191
rect 25053 7157 25087 7191
rect 25087 7157 25096 7191
rect 25044 7148 25096 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 12256 6944 12308 6996
rect 13452 6944 13504 6996
rect 14372 6944 14424 6996
rect 14556 6944 14608 6996
rect 14648 6944 14700 6996
rect 16488 6944 16540 6996
rect 20168 6944 20220 6996
rect 10324 6851 10376 6860
rect 10324 6817 10333 6851
rect 10333 6817 10367 6851
rect 10367 6817 10376 6851
rect 10324 6808 10376 6817
rect 11612 6808 11664 6860
rect 12164 6808 12216 6860
rect 14096 6851 14148 6860
rect 14096 6817 14105 6851
rect 14105 6817 14139 6851
rect 14139 6817 14148 6851
rect 14096 6808 14148 6817
rect 19340 6876 19392 6928
rect 21180 6944 21232 6996
rect 22008 6944 22060 6996
rect 22744 6987 22796 6996
rect 22744 6953 22753 6987
rect 22753 6953 22787 6987
rect 22787 6953 22796 6987
rect 22744 6944 22796 6953
rect 24768 6944 24820 6996
rect 23480 6919 23532 6928
rect 23480 6885 23492 6919
rect 23492 6885 23532 6919
rect 23480 6876 23532 6885
rect 10140 6740 10192 6792
rect 10784 6740 10836 6792
rect 11336 6740 11388 6792
rect 15936 6740 15988 6792
rect 10048 6672 10100 6724
rect 13268 6672 13320 6724
rect 15476 6672 15528 6724
rect 16304 6740 16356 6792
rect 16580 6808 16632 6860
rect 17408 6808 17460 6860
rect 17592 6808 17644 6860
rect 17960 6851 18012 6860
rect 17960 6817 17994 6851
rect 17994 6817 18012 6851
rect 17960 6808 18012 6817
rect 18236 6808 18288 6860
rect 21088 6808 21140 6860
rect 21272 6851 21324 6860
rect 21272 6817 21306 6851
rect 21306 6817 21324 6851
rect 21272 6808 21324 6817
rect 23204 6851 23256 6860
rect 23204 6817 23213 6851
rect 23213 6817 23247 6851
rect 23247 6817 23256 6851
rect 23204 6808 23256 6817
rect 24952 6740 25004 6792
rect 9864 6604 9916 6656
rect 11060 6647 11112 6656
rect 11060 6613 11069 6647
rect 11069 6613 11103 6647
rect 11103 6613 11112 6647
rect 11060 6604 11112 6613
rect 14280 6647 14332 6656
rect 14280 6613 14289 6647
rect 14289 6613 14323 6647
rect 14323 6613 14332 6647
rect 14280 6604 14332 6613
rect 15936 6604 15988 6656
rect 17592 6647 17644 6656
rect 17592 6613 17601 6647
rect 17601 6613 17635 6647
rect 17635 6613 17644 6647
rect 17592 6604 17644 6613
rect 19064 6647 19116 6656
rect 19064 6613 19073 6647
rect 19073 6613 19107 6647
rect 19107 6613 19116 6647
rect 19064 6604 19116 6613
rect 19340 6647 19392 6656
rect 19340 6613 19349 6647
rect 19349 6613 19383 6647
rect 19383 6613 19392 6647
rect 19340 6604 19392 6613
rect 20996 6604 21048 6656
rect 21364 6604 21416 6656
rect 23572 6604 23624 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 10324 6400 10376 6452
rect 10784 6400 10836 6452
rect 12164 6443 12216 6452
rect 12164 6409 12173 6443
rect 12173 6409 12207 6443
rect 12207 6409 12216 6443
rect 12164 6400 12216 6409
rect 13176 6400 13228 6452
rect 14832 6443 14884 6452
rect 14832 6409 14841 6443
rect 14841 6409 14875 6443
rect 14875 6409 14884 6443
rect 14832 6400 14884 6409
rect 16212 6443 16264 6452
rect 16212 6409 16221 6443
rect 16221 6409 16255 6443
rect 16255 6409 16264 6443
rect 16212 6400 16264 6409
rect 16396 6443 16448 6452
rect 16396 6409 16405 6443
rect 16405 6409 16439 6443
rect 16439 6409 16448 6443
rect 16396 6400 16448 6409
rect 17960 6400 18012 6452
rect 18972 6400 19024 6452
rect 19340 6400 19392 6452
rect 19524 6400 19576 6452
rect 21272 6443 21324 6452
rect 16304 6332 16356 6384
rect 9956 6196 10008 6248
rect 17684 6264 17736 6316
rect 19064 6264 19116 6316
rect 21272 6409 21281 6443
rect 21281 6409 21315 6443
rect 21315 6409 21324 6443
rect 21272 6400 21324 6409
rect 21088 6332 21140 6384
rect 23204 6400 23256 6452
rect 23480 6443 23532 6452
rect 23480 6409 23489 6443
rect 23489 6409 23523 6443
rect 23523 6409 23532 6443
rect 23480 6400 23532 6409
rect 25044 6400 25096 6452
rect 10784 6196 10836 6248
rect 13268 6196 13320 6248
rect 13544 6196 13596 6248
rect 16212 6196 16264 6248
rect 17592 6196 17644 6248
rect 18328 6196 18380 6248
rect 19248 6196 19300 6248
rect 23388 6332 23440 6384
rect 23204 6264 23256 6316
rect 25044 6196 25096 6248
rect 10140 6060 10192 6112
rect 11796 6103 11848 6112
rect 11796 6069 11805 6103
rect 11805 6069 11839 6103
rect 11839 6069 11848 6103
rect 11796 6060 11848 6069
rect 13268 6060 13320 6112
rect 19984 6128 20036 6180
rect 13728 6060 13780 6112
rect 15936 6060 15988 6112
rect 16856 6103 16908 6112
rect 16856 6069 16865 6103
rect 16865 6069 16899 6103
rect 16899 6069 16908 6103
rect 16856 6060 16908 6069
rect 22652 6103 22704 6112
rect 22652 6069 22661 6103
rect 22661 6069 22695 6103
rect 22695 6069 22704 6103
rect 22652 6060 22704 6069
rect 25228 6103 25280 6112
rect 25228 6069 25237 6103
rect 25237 6069 25271 6103
rect 25271 6069 25280 6103
rect 25228 6060 25280 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 8576 5899 8628 5908
rect 8576 5865 8585 5899
rect 8585 5865 8619 5899
rect 8619 5865 8628 5899
rect 8576 5856 8628 5865
rect 10140 5856 10192 5908
rect 13544 5856 13596 5908
rect 14096 5899 14148 5908
rect 14096 5865 14105 5899
rect 14105 5865 14139 5899
rect 14139 5865 14148 5899
rect 14096 5856 14148 5865
rect 15568 5856 15620 5908
rect 17408 5899 17460 5908
rect 17408 5865 17417 5899
rect 17417 5865 17451 5899
rect 17451 5865 17460 5899
rect 17408 5856 17460 5865
rect 17960 5856 18012 5908
rect 18328 5899 18380 5908
rect 18328 5865 18337 5899
rect 18337 5865 18371 5899
rect 18371 5865 18380 5899
rect 18328 5856 18380 5865
rect 19984 5856 20036 5908
rect 21088 5856 21140 5908
rect 23204 5856 23256 5908
rect 12440 5788 12492 5840
rect 19248 5788 19300 5840
rect 9772 5720 9824 5772
rect 16212 5763 16264 5772
rect 16212 5729 16221 5763
rect 16221 5729 16255 5763
rect 16255 5729 16264 5763
rect 16212 5720 16264 5729
rect 18236 5720 18288 5772
rect 19524 5720 19576 5772
rect 20904 5763 20956 5772
rect 20904 5729 20913 5763
rect 20913 5729 20947 5763
rect 20947 5729 20956 5763
rect 20904 5720 20956 5729
rect 22008 5720 22060 5772
rect 23480 5788 23532 5840
rect 25228 5788 25280 5840
rect 10232 5652 10284 5704
rect 9680 5584 9732 5636
rect 10784 5652 10836 5704
rect 10968 5652 11020 5704
rect 11796 5652 11848 5704
rect 15752 5652 15804 5704
rect 18144 5652 18196 5704
rect 22744 5695 22796 5704
rect 9956 5516 10008 5568
rect 11336 5516 11388 5568
rect 15568 5516 15620 5568
rect 18604 5584 18656 5636
rect 22744 5661 22753 5695
rect 22753 5661 22787 5695
rect 22787 5661 22796 5695
rect 22744 5652 22796 5661
rect 23480 5652 23532 5704
rect 23388 5584 23440 5636
rect 16856 5516 16908 5568
rect 17868 5516 17920 5568
rect 20352 5516 20404 5568
rect 21088 5559 21140 5568
rect 21088 5525 21097 5559
rect 21097 5525 21131 5559
rect 21131 5525 21140 5559
rect 21088 5516 21140 5525
rect 22100 5559 22152 5568
rect 22100 5525 22109 5559
rect 22109 5525 22143 5559
rect 22143 5525 22152 5559
rect 22100 5516 22152 5525
rect 24860 5516 24912 5568
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 9588 5312 9640 5364
rect 11796 5312 11848 5364
rect 14648 5355 14700 5364
rect 14648 5321 14657 5355
rect 14657 5321 14691 5355
rect 14691 5321 14700 5355
rect 14648 5312 14700 5321
rect 15752 5355 15804 5364
rect 15752 5321 15761 5355
rect 15761 5321 15795 5355
rect 15795 5321 15804 5355
rect 15752 5312 15804 5321
rect 17960 5312 18012 5364
rect 19340 5312 19392 5364
rect 20904 5355 20956 5364
rect 20904 5321 20913 5355
rect 20913 5321 20947 5355
rect 20947 5321 20956 5355
rect 20904 5312 20956 5321
rect 22008 5355 22060 5364
rect 22008 5321 22017 5355
rect 22017 5321 22051 5355
rect 22051 5321 22060 5355
rect 22008 5312 22060 5321
rect 23480 5355 23532 5364
rect 23480 5321 23489 5355
rect 23489 5321 23523 5355
rect 23523 5321 23532 5355
rect 23480 5312 23532 5321
rect 23848 5312 23900 5364
rect 14464 5244 14516 5296
rect 13268 5219 13320 5228
rect 13268 5185 13277 5219
rect 13277 5185 13311 5219
rect 13311 5185 13320 5219
rect 13268 5176 13320 5185
rect 14372 5176 14424 5228
rect 9956 5151 10008 5160
rect 9956 5117 9965 5151
rect 9965 5117 9999 5151
rect 9999 5117 10008 5151
rect 9956 5108 10008 5117
rect 10232 5151 10284 5160
rect 10232 5117 10266 5151
rect 10266 5117 10284 5151
rect 10232 5108 10284 5117
rect 11336 5108 11388 5160
rect 12348 5108 12400 5160
rect 14464 5108 14516 5160
rect 16212 5244 16264 5296
rect 18052 5244 18104 5296
rect 16396 5219 16448 5228
rect 16396 5185 16405 5219
rect 16405 5185 16439 5219
rect 16439 5185 16448 5219
rect 16396 5176 16448 5185
rect 18604 5176 18656 5228
rect 22652 5219 22704 5228
rect 22652 5185 22661 5219
rect 22661 5185 22695 5219
rect 22695 5185 22704 5219
rect 22652 5176 22704 5185
rect 23480 5176 23532 5228
rect 17684 5108 17736 5160
rect 18972 5108 19024 5160
rect 19524 5108 19576 5160
rect 22100 5108 22152 5160
rect 23388 5108 23440 5160
rect 24768 5176 24820 5228
rect 12532 5040 12584 5092
rect 14372 5040 14424 5092
rect 8484 4972 8536 5024
rect 8852 5015 8904 5024
rect 8852 4981 8861 5015
rect 8861 4981 8895 5015
rect 8895 4981 8904 5015
rect 8852 4972 8904 4981
rect 9588 4972 9640 5024
rect 9772 5015 9824 5024
rect 9772 4981 9781 5015
rect 9781 4981 9815 5015
rect 9815 4981 9824 5015
rect 9772 4972 9824 4981
rect 12440 4972 12492 5024
rect 16120 4972 16172 5024
rect 16948 4972 17000 5024
rect 18144 5040 18196 5092
rect 20444 5040 20496 5092
rect 21824 5083 21876 5092
rect 21824 5049 21833 5083
rect 21833 5049 21867 5083
rect 21867 5049 21876 5083
rect 21824 5040 21876 5049
rect 23664 5040 23716 5092
rect 20352 5015 20404 5024
rect 20352 4981 20361 5015
rect 20361 4981 20395 5015
rect 20395 4981 20404 5015
rect 20352 4972 20404 4981
rect 22928 4972 22980 5024
rect 25596 5015 25648 5024
rect 25596 4981 25605 5015
rect 25605 4981 25639 5015
rect 25639 4981 25648 5015
rect 25596 4972 25648 4981
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 8668 4811 8720 4820
rect 8668 4777 8677 4811
rect 8677 4777 8711 4811
rect 8711 4777 8720 4811
rect 8668 4768 8720 4777
rect 10692 4768 10744 4820
rect 10968 4811 11020 4820
rect 10968 4777 10977 4811
rect 10977 4777 11011 4811
rect 11011 4777 11020 4811
rect 10968 4768 11020 4777
rect 11428 4811 11480 4820
rect 11428 4777 11437 4811
rect 11437 4777 11471 4811
rect 11471 4777 11480 4811
rect 11428 4768 11480 4777
rect 12348 4768 12400 4820
rect 13268 4768 13320 4820
rect 14188 4768 14240 4820
rect 14372 4811 14424 4820
rect 14372 4777 14381 4811
rect 14381 4777 14415 4811
rect 14415 4777 14424 4811
rect 14372 4768 14424 4777
rect 15752 4768 15804 4820
rect 16396 4768 16448 4820
rect 18972 4768 19024 4820
rect 21272 4768 21324 4820
rect 22008 4811 22060 4820
rect 22008 4777 22017 4811
rect 22017 4777 22051 4811
rect 22051 4777 22060 4811
rect 22008 4768 22060 4777
rect 25412 4811 25464 4820
rect 25412 4777 25421 4811
rect 25421 4777 25455 4811
rect 25455 4777 25464 4811
rect 25412 4768 25464 4777
rect 9496 4700 9548 4752
rect 11060 4700 11112 4752
rect 18604 4700 18656 4752
rect 22376 4700 22428 4752
rect 22744 4700 22796 4752
rect 23296 4700 23348 4752
rect 23572 4743 23624 4752
rect 23572 4709 23581 4743
rect 23581 4709 23615 4743
rect 23615 4709 23624 4743
rect 23572 4700 23624 4709
rect 23756 4700 23808 4752
rect 24952 4700 25004 4752
rect 8760 4632 8812 4684
rect 10140 4632 10192 4684
rect 11704 4632 11756 4684
rect 12808 4632 12860 4684
rect 13544 4632 13596 4684
rect 16028 4675 16080 4684
rect 16028 4641 16062 4675
rect 16062 4641 16080 4675
rect 16028 4632 16080 4641
rect 18328 4632 18380 4684
rect 19248 4632 19300 4684
rect 20996 4675 21048 4684
rect 20996 4641 21005 4675
rect 21005 4641 21039 4675
rect 21039 4641 21048 4675
rect 20996 4632 21048 4641
rect 22284 4632 22336 4684
rect 7472 4607 7524 4616
rect 7472 4573 7481 4607
rect 7481 4573 7515 4607
rect 7515 4573 7524 4607
rect 7472 4564 7524 4573
rect 10508 4607 10560 4616
rect 10508 4573 10517 4607
rect 10517 4573 10551 4607
rect 10551 4573 10560 4607
rect 10508 4564 10560 4573
rect 12072 4607 12124 4616
rect 8392 4471 8444 4480
rect 8392 4437 8401 4471
rect 8401 4437 8435 4471
rect 8435 4437 8444 4471
rect 8392 4428 8444 4437
rect 9312 4428 9364 4480
rect 11244 4471 11296 4480
rect 11244 4437 11253 4471
rect 11253 4437 11287 4471
rect 11287 4437 11296 4471
rect 12072 4573 12081 4607
rect 12081 4573 12115 4607
rect 12115 4573 12124 4607
rect 12072 4564 12124 4573
rect 15476 4564 15528 4616
rect 17408 4564 17460 4616
rect 17868 4564 17920 4616
rect 22560 4607 22612 4616
rect 22560 4573 22569 4607
rect 22569 4573 22603 4607
rect 22603 4573 22612 4607
rect 22560 4564 22612 4573
rect 22652 4607 22704 4616
rect 22652 4573 22661 4607
rect 22661 4573 22695 4607
rect 22695 4573 22704 4607
rect 22652 4564 22704 4573
rect 23112 4564 23164 4616
rect 25044 4632 25096 4684
rect 25228 4675 25280 4684
rect 25228 4641 25237 4675
rect 25237 4641 25271 4675
rect 25271 4641 25280 4675
rect 25228 4632 25280 4641
rect 22744 4496 22796 4548
rect 23664 4539 23716 4548
rect 23664 4505 23673 4539
rect 23673 4505 23707 4539
rect 23707 4505 23716 4539
rect 23664 4496 23716 4505
rect 12532 4471 12584 4480
rect 11244 4428 11296 4437
rect 12532 4437 12541 4471
rect 12541 4437 12575 4471
rect 12575 4437 12584 4471
rect 12532 4428 12584 4437
rect 19800 4471 19852 4480
rect 19800 4437 19809 4471
rect 19809 4437 19843 4471
rect 19843 4437 19852 4471
rect 19800 4428 19852 4437
rect 21180 4471 21232 4480
rect 21180 4437 21189 4471
rect 21189 4437 21223 4471
rect 21223 4437 21232 4471
rect 21180 4428 21232 4437
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 8760 4224 8812 4276
rect 9680 4224 9732 4276
rect 11336 4224 11388 4276
rect 12808 4267 12860 4276
rect 12808 4233 12817 4267
rect 12817 4233 12851 4267
rect 12851 4233 12860 4267
rect 12808 4224 12860 4233
rect 14372 4267 14424 4276
rect 14372 4233 14381 4267
rect 14381 4233 14415 4267
rect 14415 4233 14424 4267
rect 14372 4224 14424 4233
rect 16028 4224 16080 4276
rect 20996 4267 21048 4276
rect 8300 4131 8352 4140
rect 8300 4097 8309 4131
rect 8309 4097 8343 4131
rect 8343 4097 8352 4131
rect 8300 4088 8352 4097
rect 8392 4088 8444 4140
rect 8852 4020 8904 4072
rect 9312 4131 9364 4140
rect 9312 4097 9321 4131
rect 9321 4097 9355 4131
rect 9355 4097 9364 4131
rect 10968 4131 11020 4140
rect 9312 4088 9364 4097
rect 10968 4097 10977 4131
rect 10977 4097 11011 4131
rect 11011 4097 11020 4131
rect 10968 4088 11020 4097
rect 13084 4131 13136 4140
rect 13084 4097 13093 4131
rect 13093 4097 13127 4131
rect 13127 4097 13136 4131
rect 13084 4088 13136 4097
rect 9404 4020 9456 4072
rect 18328 4199 18380 4208
rect 18328 4165 18337 4199
rect 18337 4165 18371 4199
rect 18371 4165 18380 4199
rect 18328 4156 18380 4165
rect 20996 4233 21005 4267
rect 21005 4233 21039 4267
rect 21039 4233 21048 4267
rect 20996 4224 21048 4233
rect 23756 4224 23808 4276
rect 24032 4224 24084 4276
rect 25228 4224 25280 4276
rect 14556 4088 14608 4140
rect 14740 4088 14792 4140
rect 17868 4131 17920 4140
rect 15476 4020 15528 4072
rect 17868 4097 17877 4131
rect 17877 4097 17911 4131
rect 17911 4097 17920 4131
rect 17868 4088 17920 4097
rect 19800 4156 19852 4208
rect 21272 4156 21324 4208
rect 22744 4199 22796 4208
rect 16396 4020 16448 4072
rect 20628 4088 20680 4140
rect 22744 4165 22753 4199
rect 22753 4165 22787 4199
rect 22787 4165 22796 4199
rect 22744 4156 22796 4165
rect 23112 4199 23164 4208
rect 23112 4165 23121 4199
rect 23121 4165 23155 4199
rect 23155 4165 23164 4199
rect 23112 4156 23164 4165
rect 23756 4088 23808 4140
rect 24216 4088 24268 4140
rect 25044 4131 25096 4140
rect 25044 4097 25053 4131
rect 25053 4097 25087 4131
rect 25087 4097 25096 4131
rect 25044 4088 25096 4097
rect 20352 4020 20404 4072
rect 10140 3952 10192 4004
rect 19156 3995 19208 4004
rect 19156 3961 19165 3995
rect 19165 3961 19199 3995
rect 19199 3961 19208 3995
rect 19156 3952 19208 3961
rect 20720 3995 20772 4004
rect 20720 3961 20729 3995
rect 20729 3961 20763 3995
rect 20763 3961 20772 3995
rect 20720 3952 20772 3961
rect 21824 3952 21876 4004
rect 7840 3927 7892 3936
rect 7840 3893 7849 3927
rect 7849 3893 7883 3927
rect 7883 3893 7892 3927
rect 7840 3884 7892 3893
rect 8944 3884 8996 3936
rect 10048 3884 10100 3936
rect 10692 3927 10744 3936
rect 10692 3893 10701 3927
rect 10701 3893 10735 3927
rect 10735 3893 10744 3927
rect 10692 3884 10744 3893
rect 10784 3927 10836 3936
rect 10784 3893 10793 3927
rect 10793 3893 10827 3927
rect 10827 3893 10836 3927
rect 11428 3927 11480 3936
rect 10784 3884 10836 3893
rect 11428 3893 11437 3927
rect 11437 3893 11471 3927
rect 11471 3893 11480 3927
rect 11428 3884 11480 3893
rect 11704 3927 11756 3936
rect 11704 3893 11713 3927
rect 11713 3893 11747 3927
rect 11747 3893 11756 3927
rect 11704 3884 11756 3893
rect 12072 3927 12124 3936
rect 12072 3893 12081 3927
rect 12081 3893 12115 3927
rect 12115 3893 12124 3927
rect 12072 3884 12124 3893
rect 13268 3927 13320 3936
rect 13268 3893 13277 3927
rect 13277 3893 13311 3927
rect 13311 3893 13320 3927
rect 13268 3884 13320 3893
rect 13544 3884 13596 3936
rect 17132 3927 17184 3936
rect 17132 3893 17141 3927
rect 17141 3893 17175 3927
rect 17175 3893 17184 3927
rect 17132 3884 17184 3893
rect 17408 3927 17460 3936
rect 17408 3893 17417 3927
rect 17417 3893 17451 3927
rect 17451 3893 17460 3927
rect 17408 3884 17460 3893
rect 18788 3927 18840 3936
rect 18788 3893 18797 3927
rect 18797 3893 18831 3927
rect 18831 3893 18840 3927
rect 18788 3884 18840 3893
rect 21456 3884 21508 3936
rect 21548 3884 21600 3936
rect 22284 3927 22336 3936
rect 22284 3893 22293 3927
rect 22293 3893 22327 3927
rect 22327 3893 22336 3927
rect 22284 3884 22336 3893
rect 24216 3927 24268 3936
rect 24216 3893 24225 3927
rect 24225 3893 24259 3927
rect 24259 3893 24268 3927
rect 24216 3884 24268 3893
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 8852 3680 8904 3732
rect 9496 3723 9548 3732
rect 9496 3689 9505 3723
rect 9505 3689 9539 3723
rect 9539 3689 9548 3723
rect 9496 3680 9548 3689
rect 12440 3723 12492 3732
rect 12440 3689 12449 3723
rect 12449 3689 12483 3723
rect 12483 3689 12492 3723
rect 12440 3680 12492 3689
rect 13268 3680 13320 3732
rect 14188 3680 14240 3732
rect 15476 3680 15528 3732
rect 17224 3680 17276 3732
rect 17868 3680 17920 3732
rect 18052 3680 18104 3732
rect 8484 3612 8536 3664
rect 8944 3612 8996 3664
rect 13544 3612 13596 3664
rect 13820 3612 13872 3664
rect 15384 3612 15436 3664
rect 17592 3655 17644 3664
rect 17592 3621 17601 3655
rect 17601 3621 17635 3655
rect 17635 3621 17644 3655
rect 17592 3612 17644 3621
rect 19156 3680 19208 3732
rect 23756 3723 23808 3732
rect 23756 3689 23765 3723
rect 23765 3689 23799 3723
rect 23799 3689 23808 3723
rect 23756 3680 23808 3689
rect 21180 3612 21232 3664
rect 6920 3587 6972 3596
rect 6920 3553 6929 3587
rect 6929 3553 6963 3587
rect 6963 3553 6972 3587
rect 6920 3544 6972 3553
rect 8392 3587 8444 3596
rect 8392 3553 8401 3587
rect 8401 3553 8435 3587
rect 8435 3553 8444 3587
rect 8392 3544 8444 3553
rect 9956 3587 10008 3596
rect 9956 3553 9965 3587
rect 9965 3553 9999 3587
rect 9999 3553 10008 3587
rect 9956 3544 10008 3553
rect 11336 3587 11388 3596
rect 11336 3553 11370 3587
rect 11370 3553 11388 3587
rect 11336 3544 11388 3553
rect 15476 3544 15528 3596
rect 17408 3544 17460 3596
rect 19156 3587 19208 3596
rect 19156 3553 19165 3587
rect 19165 3553 19199 3587
rect 19199 3553 19208 3587
rect 19156 3544 19208 3553
rect 21640 3587 21692 3596
rect 21640 3553 21649 3587
rect 21649 3553 21683 3587
rect 21683 3553 21692 3587
rect 21640 3544 21692 3553
rect 21916 3544 21968 3596
rect 24768 3612 24820 3664
rect 8484 3519 8536 3528
rect 8484 3485 8493 3519
rect 8493 3485 8527 3519
rect 8527 3485 8536 3519
rect 8484 3476 8536 3485
rect 8668 3519 8720 3528
rect 8668 3485 8677 3519
rect 8677 3485 8711 3519
rect 8711 3485 8720 3519
rect 8668 3476 8720 3485
rect 9772 3408 9824 3460
rect 10692 3408 10744 3460
rect 7104 3383 7156 3392
rect 7104 3349 7113 3383
rect 7113 3349 7147 3383
rect 7147 3349 7156 3383
rect 7104 3340 7156 3349
rect 9036 3340 9088 3392
rect 10784 3340 10836 3392
rect 10968 3383 11020 3392
rect 10968 3349 10977 3383
rect 10977 3349 11011 3383
rect 11011 3349 11020 3383
rect 10968 3340 11020 3349
rect 14648 3476 14700 3528
rect 16120 3519 16172 3528
rect 16120 3485 16129 3519
rect 16129 3485 16163 3519
rect 16163 3485 16172 3519
rect 16120 3476 16172 3485
rect 13636 3408 13688 3460
rect 16488 3476 16540 3528
rect 17868 3519 17920 3528
rect 17868 3485 17877 3519
rect 17877 3485 17911 3519
rect 17911 3485 17920 3519
rect 17868 3476 17920 3485
rect 19248 3519 19300 3528
rect 19248 3485 19257 3519
rect 19257 3485 19291 3519
rect 19291 3485 19300 3519
rect 19248 3476 19300 3485
rect 19340 3476 19392 3528
rect 20628 3476 20680 3528
rect 24032 3519 24084 3528
rect 24032 3485 24041 3519
rect 24041 3485 24075 3519
rect 24075 3485 24084 3519
rect 24032 3476 24084 3485
rect 17040 3408 17092 3460
rect 11428 3340 11480 3392
rect 21456 3340 21508 3392
rect 21640 3340 21692 3392
rect 25412 3383 25464 3392
rect 25412 3349 25421 3383
rect 25421 3349 25455 3383
rect 25455 3349 25464 3383
rect 25412 3340 25464 3349
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 6000 3136 6052 3188
rect 6276 3179 6328 3188
rect 6276 3145 6285 3179
rect 6285 3145 6319 3179
rect 6319 3145 6328 3179
rect 6276 3136 6328 3145
rect 6644 3179 6696 3188
rect 6644 3145 6653 3179
rect 6653 3145 6687 3179
rect 6687 3145 6696 3179
rect 6644 3136 6696 3145
rect 6920 3136 6972 3188
rect 8024 3136 8076 3188
rect 9772 3136 9824 3188
rect 11336 3136 11388 3188
rect 13820 3136 13872 3188
rect 15384 3179 15436 3188
rect 15384 3145 15393 3179
rect 15393 3145 15427 3179
rect 15427 3145 15436 3179
rect 15384 3136 15436 3145
rect 8300 3068 8352 3120
rect 8576 3111 8628 3120
rect 8576 3077 8585 3111
rect 8585 3077 8619 3111
rect 8619 3077 8628 3111
rect 8576 3068 8628 3077
rect 9680 3068 9732 3120
rect 8116 3043 8168 3052
rect 6276 2932 6328 2984
rect 8116 3009 8125 3043
rect 8125 3009 8159 3043
rect 8159 3009 8168 3043
rect 8116 3000 8168 3009
rect 16120 3136 16172 3188
rect 16856 3179 16908 3188
rect 16856 3145 16865 3179
rect 16865 3145 16899 3179
rect 16899 3145 16908 3179
rect 16856 3136 16908 3145
rect 17868 3136 17920 3188
rect 19156 3136 19208 3188
rect 20628 3136 20680 3188
rect 21916 3136 21968 3188
rect 17592 3068 17644 3120
rect 19248 3068 19300 3120
rect 11428 3000 11480 3052
rect 12440 3043 12492 3052
rect 12440 3009 12449 3043
rect 12449 3009 12483 3043
rect 12483 3009 12492 3043
rect 15476 3043 15528 3052
rect 12440 3000 12492 3009
rect 15476 3009 15485 3043
rect 15485 3009 15519 3043
rect 15519 3009 15528 3043
rect 15476 3000 15528 3009
rect 17040 3000 17092 3052
rect 17500 3000 17552 3052
rect 18052 3043 18104 3052
rect 18052 3009 18061 3043
rect 18061 3009 18095 3043
rect 18095 3009 18104 3043
rect 18052 3000 18104 3009
rect 21180 3043 21232 3052
rect 21180 3009 21189 3043
rect 21189 3009 21223 3043
rect 21223 3009 21232 3043
rect 21180 3000 21232 3009
rect 24032 3136 24084 3188
rect 24124 3068 24176 3120
rect 24768 3111 24820 3120
rect 24768 3077 24777 3111
rect 24777 3077 24811 3111
rect 24811 3077 24820 3111
rect 24768 3068 24820 3077
rect 24584 3000 24636 3052
rect 25412 3000 25464 3052
rect 8484 2975 8536 2984
rect 8484 2941 8493 2975
rect 8493 2941 8527 2975
rect 8527 2941 8536 2975
rect 8484 2932 8536 2941
rect 8944 2975 8996 2984
rect 8944 2941 8953 2975
rect 8953 2941 8987 2975
rect 8987 2941 8996 2975
rect 8944 2932 8996 2941
rect 9036 2975 9088 2984
rect 9036 2941 9045 2975
rect 9045 2941 9079 2975
rect 9079 2941 9088 2975
rect 9036 2932 9088 2941
rect 10048 2932 10100 2984
rect 8392 2864 8444 2916
rect 10876 2932 10928 2984
rect 24124 2975 24176 2984
rect 24124 2941 24133 2975
rect 24133 2941 24167 2975
rect 24167 2941 24176 2975
rect 24124 2932 24176 2941
rect 12256 2907 12308 2916
rect 9680 2796 9732 2848
rect 12256 2873 12265 2907
rect 12265 2873 12299 2907
rect 12299 2873 12308 2907
rect 12256 2864 12308 2873
rect 13728 2864 13780 2916
rect 16488 2864 16540 2916
rect 18144 2864 18196 2916
rect 21640 2864 21692 2916
rect 23756 2864 23808 2916
rect 10968 2796 11020 2848
rect 13820 2839 13872 2848
rect 13820 2805 13829 2839
rect 13829 2805 13863 2839
rect 13863 2805 13872 2839
rect 13820 2796 13872 2805
rect 19432 2839 19484 2848
rect 19432 2805 19441 2839
rect 19441 2805 19475 2839
rect 19475 2805 19484 2839
rect 19432 2796 19484 2805
rect 22560 2839 22612 2848
rect 22560 2805 22569 2839
rect 22569 2805 22603 2839
rect 22603 2805 22612 2839
rect 22560 2796 22612 2805
rect 23480 2796 23532 2848
rect 25412 2839 25464 2848
rect 25412 2805 25421 2839
rect 25421 2805 25455 2839
rect 25455 2805 25464 2839
rect 25412 2796 25464 2805
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 5632 2635 5684 2644
rect 5632 2601 5641 2635
rect 5641 2601 5675 2635
rect 5675 2601 5684 2635
rect 5632 2592 5684 2601
rect 6368 2635 6420 2644
rect 6368 2601 6377 2635
rect 6377 2601 6411 2635
rect 6411 2601 6420 2635
rect 6368 2592 6420 2601
rect 8116 2635 8168 2644
rect 8116 2601 8125 2635
rect 8125 2601 8159 2635
rect 8159 2601 8168 2635
rect 8116 2592 8168 2601
rect 10968 2592 11020 2644
rect 11888 2635 11940 2644
rect 11888 2601 11897 2635
rect 11897 2601 11931 2635
rect 11931 2601 11940 2635
rect 11888 2592 11940 2601
rect 13820 2592 13872 2644
rect 14740 2635 14792 2644
rect 14740 2601 14749 2635
rect 14749 2601 14783 2635
rect 14783 2601 14792 2635
rect 14740 2592 14792 2601
rect 16488 2592 16540 2644
rect 17224 2635 17276 2644
rect 17224 2601 17233 2635
rect 17233 2601 17267 2635
rect 17267 2601 17276 2635
rect 17224 2592 17276 2601
rect 17408 2592 17460 2644
rect 18144 2635 18196 2644
rect 18144 2601 18153 2635
rect 18153 2601 18187 2635
rect 18187 2601 18196 2635
rect 18144 2592 18196 2601
rect 19340 2592 19392 2644
rect 8668 2524 8720 2576
rect 9588 2567 9640 2576
rect 9588 2533 9597 2567
rect 9597 2533 9631 2567
rect 9631 2533 9640 2567
rect 9588 2524 9640 2533
rect 9956 2524 10008 2576
rect 11428 2524 11480 2576
rect 12440 2524 12492 2576
rect 7012 2499 7064 2508
rect 7012 2465 7021 2499
rect 7021 2465 7055 2499
rect 7055 2465 7064 2499
rect 7012 2456 7064 2465
rect 10968 2456 11020 2508
rect 15936 2524 15988 2576
rect 19156 2567 19208 2576
rect 19156 2533 19190 2567
rect 19190 2533 19208 2567
rect 19156 2524 19208 2533
rect 12900 2499 12952 2508
rect 4712 2431 4764 2440
rect 4712 2397 4721 2431
rect 4721 2397 4755 2431
rect 4755 2397 4764 2431
rect 4712 2388 4764 2397
rect 8576 2431 8628 2440
rect 8576 2397 8585 2431
rect 8585 2397 8619 2431
rect 8619 2397 8628 2431
rect 8576 2388 8628 2397
rect 9956 2388 10008 2440
rect 12900 2465 12934 2499
rect 12934 2465 12952 2499
rect 12900 2456 12952 2465
rect 14648 2456 14700 2508
rect 15476 2499 15528 2508
rect 15476 2465 15485 2499
rect 15485 2465 15519 2499
rect 15519 2465 15528 2499
rect 15476 2456 15528 2465
rect 21180 2456 21232 2508
rect 23388 2592 23440 2644
rect 25596 2635 25648 2644
rect 25596 2601 25605 2635
rect 25605 2601 25639 2635
rect 25639 2601 25648 2635
rect 25596 2592 25648 2601
rect 21640 2431 21692 2440
rect 21640 2397 21649 2431
rect 21649 2397 21683 2431
rect 21683 2397 21692 2431
rect 21640 2388 21692 2397
rect 21824 2363 21876 2372
rect 21824 2329 21833 2363
rect 21833 2329 21867 2363
rect 21867 2329 21876 2363
rect 21824 2320 21876 2329
rect 23572 2456 23624 2508
rect 24768 2524 24820 2576
rect 23664 2388 23716 2440
rect 24676 2456 24728 2508
rect 24584 2431 24636 2440
rect 24584 2397 24593 2431
rect 24593 2397 24627 2431
rect 24627 2397 24636 2431
rect 24584 2388 24636 2397
rect 6828 2252 6880 2304
rect 7196 2295 7248 2304
rect 7196 2261 7205 2295
rect 7205 2261 7239 2295
rect 7239 2261 7248 2295
rect 7196 2252 7248 2261
rect 9220 2295 9272 2304
rect 9220 2261 9229 2295
rect 9229 2261 9263 2295
rect 9263 2261 9272 2295
rect 9220 2252 9272 2261
rect 13268 2252 13320 2304
rect 18512 2252 18564 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 10048 1776 10100 1828
rect 16764 1776 16816 1828
rect 10784 1232 10836 1284
rect 13912 1232 13964 1284
rect 20076 552 20128 604
rect 20444 552 20496 604
<< metal2 >>
rect 3514 27520 3570 28000
rect 10506 27520 10562 28000
rect 17498 27520 17554 28000
rect 23662 27704 23718 27713
rect 23662 27639 23718 27648
rect 3528 24177 3556 27520
rect 10520 25786 10548 27520
rect 10520 25758 10824 25786
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 3514 24168 3570 24177
rect 3514 24103 3570 24112
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 10046 21448 10102 21457
rect 10046 21383 10102 21392
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 4158 12744 4214 12753
rect 4158 12679 4214 12688
rect 4066 8528 4122 8537
rect 4066 8463 4122 8472
rect 1582 7440 1638 7449
rect 1582 7375 1638 7384
rect 294 6216 350 6225
rect 294 6151 350 6160
rect 308 480 336 6151
rect 938 3496 994 3505
rect 938 3431 994 3440
rect 952 480 980 3431
rect 1596 480 1624 7375
rect 2226 6896 2282 6905
rect 2226 6831 2282 6840
rect 2240 480 2268 6831
rect 2870 4992 2926 5001
rect 2870 4927 2926 4936
rect 2884 480 2912 4927
rect 3514 4176 3570 4185
rect 3514 4111 3570 4120
rect 3528 480 3556 4111
rect 4080 3505 4108 8463
rect 4172 7546 4200 12679
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 8942 11112 8998 11121
rect 8942 11047 8998 11056
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 6274 9480 6330 9489
rect 6274 9415 6330 9424
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 6090 7712 6146 7721
rect 5622 7644 5918 7664
rect 6090 7647 6146 7656
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 4158 6352 4214 6361
rect 4158 6287 4214 6296
rect 4066 3496 4122 3505
rect 4066 3431 4122 3440
rect 4172 480 4200 6287
rect 4802 3088 4858 3097
rect 4802 3023 4858 3032
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 4724 1601 4752 2382
rect 4710 1592 4766 1601
rect 4710 1527 4766 1536
rect 4816 480 4844 3023
rect 5460 480 5488 7482
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5998 5672 6054 5681
rect 5998 5607 6054 5616
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 6012 3194 6040 5607
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 5630 2680 5686 2689
rect 5630 2615 5632 2624
rect 5684 2615 5686 2624
rect 5632 2586 5684 2592
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 6104 480 6132 7647
rect 6288 3194 6316 9415
rect 8574 8392 8630 8401
rect 8574 8327 8630 8336
rect 6734 7984 6790 7993
rect 6734 7919 6790 7928
rect 6366 6760 6422 6769
rect 6366 6695 6422 6704
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 6288 2990 6316 3130
rect 6276 2984 6328 2990
rect 6276 2926 6328 2932
rect 6380 2650 6408 6695
rect 6642 3224 6698 3233
rect 6642 3159 6644 3168
rect 6696 3159 6698 3168
rect 6644 3130 6696 3136
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 6748 480 6776 7919
rect 7010 7576 7066 7585
rect 7010 7511 7066 7520
rect 6918 5264 6974 5273
rect 6918 5199 6974 5208
rect 6932 3602 6960 5199
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 6932 3194 6960 3538
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 7024 2514 7052 7511
rect 8114 7304 8170 7313
rect 8114 7239 8170 7248
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7484 4049 7512 4558
rect 7470 4040 7526 4049
rect 7470 3975 7526 3984
rect 7840 3936 7892 3942
rect 7840 3878 7892 3884
rect 7104 3392 7156 3398
rect 7104 3334 7156 3340
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 6828 2304 6880 2310
rect 6828 2246 6880 2252
rect 6840 1737 6868 2246
rect 6826 1728 6882 1737
rect 6826 1663 6882 1672
rect 7116 1329 7144 3334
rect 7196 2304 7248 2310
rect 7196 2246 7248 2252
rect 7102 1320 7158 1329
rect 7102 1255 7158 1264
rect 294 0 350 480
rect 938 0 994 480
rect 1582 0 1638 480
rect 2226 0 2282 480
rect 2870 0 2926 480
rect 3514 0 3570 480
rect 4158 0 4214 480
rect 4802 0 4858 480
rect 5446 0 5502 480
rect 6090 0 6146 480
rect 6734 0 6790 480
rect 7208 241 7236 2246
rect 7378 1456 7434 1465
rect 7378 1391 7434 1400
rect 7392 480 7420 1391
rect 7194 232 7250 241
rect 7194 167 7250 176
rect 7378 0 7434 480
rect 7852 105 7880 3878
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 8036 480 8064 3130
rect 8128 3058 8156 7239
rect 8588 5914 8616 8327
rect 8758 6216 8814 6225
rect 8758 6151 8814 6160
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8666 5808 8722 5817
rect 8666 5743 8722 5752
rect 8484 5024 8536 5030
rect 8484 4966 8536 4972
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 8298 4312 8354 4321
rect 8298 4247 8354 4256
rect 8312 4146 8340 4247
rect 8404 4146 8432 4422
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 8496 3670 8524 4966
rect 8680 4826 8708 5743
rect 8668 4820 8720 4826
rect 8668 4762 8720 4768
rect 8772 4690 8800 6151
rect 8852 5024 8904 5030
rect 8852 4966 8904 4972
rect 8760 4684 8812 4690
rect 8760 4626 8812 4632
rect 8772 4282 8800 4626
rect 8760 4276 8812 4282
rect 8760 4218 8812 4224
rect 8864 4078 8892 4966
rect 8852 4072 8904 4078
rect 8852 4014 8904 4020
rect 8864 3738 8892 4014
rect 8956 3942 8984 11047
rect 10060 6730 10088 21383
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10796 20505 10824 25758
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 12806 23760 12862 23769
rect 12806 23695 12862 23704
rect 12820 23254 12848 23695
rect 12808 23248 12860 23254
rect 12808 23190 12860 23196
rect 12532 23180 12584 23186
rect 12532 23122 12584 23128
rect 12544 22438 12572 23122
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 14554 22672 14610 22681
rect 14554 22607 14610 22616
rect 11980 22432 12032 22438
rect 11980 22374 12032 22380
rect 12532 22432 12584 22438
rect 12532 22374 12584 22380
rect 10782 20496 10838 20505
rect 10782 20431 10838 20440
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 11610 18864 11666 18873
rect 11610 18799 11666 18808
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 11624 17814 11652 18799
rect 11612 17808 11664 17814
rect 11612 17750 11664 17756
rect 11428 17740 11480 17746
rect 11428 17682 11480 17688
rect 11440 17626 11468 17682
rect 11440 17598 11560 17626
rect 11426 17096 11482 17105
rect 11426 17031 11482 17040
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 11256 8634 11284 8910
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 10690 8256 10746 8265
rect 10289 8188 10585 8208
rect 10690 8191 10746 8200
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10704 8090 10732 8191
rect 10782 8120 10838 8129
rect 10692 8084 10744 8090
rect 10980 8090 11008 8570
rect 10782 8055 10838 8064
rect 10968 8084 11020 8090
rect 10692 8026 10744 8032
rect 10796 7834 10824 8055
rect 10968 8026 11020 8032
rect 11150 7984 11206 7993
rect 11150 7919 11206 7928
rect 10520 7806 10824 7834
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 10520 7721 10548 7806
rect 10506 7712 10562 7721
rect 10506 7647 10562 7656
rect 10690 7712 10746 7721
rect 10690 7647 10746 7656
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10048 6724 10100 6730
rect 10048 6666 10100 6672
rect 9864 6656 9916 6662
rect 9916 6604 9996 6610
rect 9864 6598 9996 6604
rect 9876 6582 9996 6598
rect 9968 6254 9996 6582
rect 9956 6248 10008 6254
rect 9956 6190 10008 6196
rect 9772 5772 9824 5778
rect 9772 5714 9824 5720
rect 9680 5636 9732 5642
rect 9680 5578 9732 5584
rect 9692 5386 9720 5578
rect 9600 5370 9720 5386
rect 9588 5364 9720 5370
rect 9640 5358 9720 5364
rect 9588 5306 9640 5312
rect 9784 5030 9812 5714
rect 9968 5574 9996 6190
rect 10152 6118 10180 6734
rect 10336 6458 10364 6802
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 10140 6112 10192 6118
rect 10140 6054 10192 6060
rect 10152 5914 10180 6054
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 9956 5568 10008 5574
rect 9956 5510 10008 5516
rect 9968 5166 9996 5510
rect 10244 5409 10272 5646
rect 10230 5400 10286 5409
rect 10230 5335 10286 5344
rect 10244 5166 10272 5335
rect 9956 5160 10008 5166
rect 9956 5102 10008 5108
rect 10232 5160 10284 5166
rect 10232 5102 10284 5108
rect 9588 5024 9640 5030
rect 9772 5024 9824 5030
rect 9588 4966 9640 4972
rect 9770 4992 9772 5001
rect 9824 4992 9826 5001
rect 9496 4752 9548 4758
rect 9496 4694 9548 4700
rect 9218 4584 9274 4593
rect 9218 4519 9274 4528
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 8852 3732 8904 3738
rect 8852 3674 8904 3680
rect 8484 3664 8536 3670
rect 8944 3664 8996 3670
rect 8484 3606 8536 3612
rect 8666 3632 8722 3641
rect 8392 3596 8444 3602
rect 8944 3606 8996 3612
rect 8666 3567 8722 3576
rect 8392 3538 8444 3544
rect 8300 3120 8352 3126
rect 8300 3062 8352 3068
rect 8116 3052 8168 3058
rect 8116 2994 8168 3000
rect 8116 2644 8168 2650
rect 8116 2586 8168 2592
rect 8128 2553 8156 2586
rect 8114 2544 8170 2553
rect 8114 2479 8170 2488
rect 8312 2009 8340 3062
rect 8404 2922 8432 3538
rect 8680 3534 8708 3567
rect 8484 3528 8536 3534
rect 8668 3528 8720 3534
rect 8484 3470 8536 3476
rect 8574 3496 8630 3505
rect 8496 2990 8524 3470
rect 8668 3470 8720 3476
rect 8574 3431 8630 3440
rect 8588 3126 8616 3431
rect 8576 3120 8628 3126
rect 8576 3062 8628 3068
rect 8956 2990 8984 3606
rect 9036 3392 9088 3398
rect 9036 3334 9088 3340
rect 9048 2990 9076 3334
rect 8484 2984 8536 2990
rect 8482 2952 8484 2961
rect 8944 2984 8996 2990
rect 8536 2952 8538 2961
rect 8392 2916 8444 2922
rect 8944 2926 8996 2932
rect 9036 2984 9088 2990
rect 9036 2926 9088 2932
rect 9232 2938 9260 4519
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 9324 4146 9352 4422
rect 9312 4140 9364 4146
rect 9312 4082 9364 4088
rect 9324 3097 9352 4082
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 9310 3088 9366 3097
rect 9310 3023 9366 3032
rect 9232 2910 9352 2938
rect 8482 2887 8538 2896
rect 8392 2858 8444 2864
rect 8668 2576 8720 2582
rect 8668 2518 8720 2524
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 8588 2145 8616 2382
rect 8574 2136 8630 2145
rect 8574 2071 8630 2080
rect 8298 2000 8354 2009
rect 8298 1935 8354 1944
rect 8680 480 8708 2518
rect 9220 2304 9272 2310
rect 9218 2272 9220 2281
rect 9272 2272 9274 2281
rect 9218 2207 9274 2216
rect 9324 480 9352 2910
rect 9416 2417 9444 4014
rect 9508 3738 9536 4694
rect 9496 3732 9548 3738
rect 9496 3674 9548 3680
rect 9600 3369 9628 4966
rect 9770 4927 9826 4936
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10704 4826 10732 7647
rect 10874 7576 10930 7585
rect 10874 7511 10930 7520
rect 10888 7313 10916 7511
rect 10874 7304 10930 7313
rect 10784 7268 10836 7274
rect 10874 7239 10930 7248
rect 10784 7210 10836 7216
rect 10796 6798 10824 7210
rect 10784 6792 10836 6798
rect 10784 6734 10836 6740
rect 10796 6458 10824 6734
rect 11072 6662 11100 7822
rect 11164 7585 11192 7919
rect 11336 7744 11388 7750
rect 11336 7686 11388 7692
rect 11150 7576 11206 7585
rect 11150 7511 11206 7520
rect 11348 7206 11376 7686
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11348 6798 11376 7142
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 10784 6452 10836 6458
rect 10784 6394 10836 6400
rect 10796 6254 10824 6394
rect 10784 6248 10836 6254
rect 10784 6190 10836 6196
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 10968 5704 11020 5710
rect 10968 5646 11020 5652
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 10506 4720 10562 4729
rect 10140 4684 10192 4690
rect 10506 4655 10562 4664
rect 10140 4626 10192 4632
rect 9680 4276 9732 4282
rect 9680 4218 9732 4224
rect 9586 3360 9642 3369
rect 9586 3295 9642 3304
rect 9692 3233 9720 4218
rect 10152 4010 10180 4626
rect 10520 4622 10548 4655
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10140 4004 10192 4010
rect 10140 3946 10192 3952
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 9772 3460 9824 3466
rect 9772 3402 9824 3408
rect 9678 3224 9734 3233
rect 9784 3194 9812 3402
rect 9968 3233 9996 3538
rect 9954 3224 10010 3233
rect 9678 3159 9734 3168
rect 9772 3188 9824 3194
rect 9692 3126 9720 3159
rect 9954 3159 10010 3168
rect 9772 3130 9824 3136
rect 9680 3120 9732 3126
rect 9680 3062 9732 3068
rect 10060 2990 10088 3878
rect 10048 2984 10100 2990
rect 10048 2926 10100 2932
rect 9680 2848 9732 2854
rect 10152 2836 10180 3946
rect 10796 3942 10824 5646
rect 10874 4856 10930 4865
rect 10980 4826 11008 5646
rect 10874 4791 10930 4800
rect 10968 4820 11020 4826
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 10784 3936 10836 3942
rect 10784 3878 10836 3884
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10704 3466 10732 3878
rect 10692 3460 10744 3466
rect 10692 3402 10744 3408
rect 10784 3392 10836 3398
rect 10784 3334 10836 3340
rect 10690 2952 10746 2961
rect 10690 2887 10746 2896
rect 9680 2790 9732 2796
rect 10060 2808 10180 2836
rect 9588 2576 9640 2582
rect 9692 2564 9720 2790
rect 9954 2680 10010 2689
rect 9954 2615 10010 2624
rect 9968 2582 9996 2615
rect 9640 2536 9720 2564
rect 9956 2576 10008 2582
rect 9588 2518 9640 2524
rect 9956 2518 10008 2524
rect 9968 2446 9996 2518
rect 9956 2440 10008 2446
rect 9402 2408 9458 2417
rect 9956 2382 10008 2388
rect 9402 2343 9458 2352
rect 10060 2292 10088 2808
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 9876 2264 10088 2292
rect 9876 1465 9904 2264
rect 10048 1828 10100 1834
rect 10048 1770 10100 1776
rect 9862 1456 9918 1465
rect 9862 1391 9918 1400
rect 10060 480 10088 1770
rect 10704 480 10732 2887
rect 10796 1290 10824 3334
rect 10888 2990 10916 4791
rect 10968 4762 11020 4768
rect 11072 4758 11100 6598
rect 11348 5574 11376 6734
rect 11336 5568 11388 5574
rect 11336 5510 11388 5516
rect 11348 5166 11376 5510
rect 11336 5160 11388 5166
rect 11336 5102 11388 5108
rect 11060 4752 11112 4758
rect 11060 4694 11112 4700
rect 11072 4457 11100 4694
rect 11244 4480 11296 4486
rect 11058 4448 11114 4457
rect 11244 4422 11296 4428
rect 11058 4383 11114 4392
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 10980 3398 11008 4082
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 11058 3360 11114 3369
rect 10876 2984 10928 2990
rect 10876 2926 10928 2932
rect 10980 2854 11008 3334
rect 11058 3295 11114 3304
rect 11072 3097 11100 3295
rect 11058 3088 11114 3097
rect 11058 3023 11114 3032
rect 10968 2848 11020 2854
rect 10968 2790 11020 2796
rect 11150 2816 11206 2825
rect 10980 2650 11008 2790
rect 11150 2751 11206 2760
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 11164 2530 11192 2751
rect 11256 2553 11284 4422
rect 11348 4282 11376 5102
rect 11440 4826 11468 17031
rect 11532 16998 11560 17598
rect 11520 16992 11572 16998
rect 11520 16934 11572 16940
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11336 4276 11388 4282
rect 11336 4218 11388 4224
rect 11428 3936 11480 3942
rect 11426 3904 11428 3913
rect 11480 3904 11482 3913
rect 11426 3839 11482 3848
rect 11336 3596 11388 3602
rect 11336 3538 11388 3544
rect 11348 3194 11376 3538
rect 11532 3505 11560 16934
rect 11992 9178 12020 22374
rect 14568 21554 14596 22607
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 16854 21584 16910 21593
rect 14556 21548 14608 21554
rect 16854 21519 16910 21528
rect 14556 21490 14608 21496
rect 14004 21480 14056 21486
rect 14004 21422 14056 21428
rect 13544 18216 13596 18222
rect 13544 18158 13596 18164
rect 13818 18184 13874 18193
rect 13176 17128 13228 17134
rect 13174 17096 13176 17105
rect 13228 17096 13230 17105
rect 13174 17031 13230 17040
rect 12438 14512 12494 14521
rect 12438 14447 12494 14456
rect 12452 11121 12480 14447
rect 12898 11520 12954 11529
rect 12898 11455 12954 11464
rect 12438 11112 12494 11121
rect 12438 11047 12494 11056
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 11980 9172 12032 9178
rect 11980 9114 12032 9120
rect 12070 9072 12126 9081
rect 12070 9007 12126 9016
rect 12348 9036 12400 9042
rect 11980 8356 12032 8362
rect 11980 8298 12032 8304
rect 11796 7948 11848 7954
rect 11796 7890 11848 7896
rect 11612 7880 11664 7886
rect 11612 7822 11664 7828
rect 11624 7206 11652 7822
rect 11808 7206 11836 7890
rect 11612 7200 11664 7206
rect 11612 7142 11664 7148
rect 11796 7200 11848 7206
rect 11796 7142 11848 7148
rect 11624 6866 11652 7142
rect 11808 6905 11836 7142
rect 11992 6905 12020 8298
rect 11794 6896 11850 6905
rect 11612 6860 11664 6866
rect 11794 6831 11850 6840
rect 11978 6896 12034 6905
rect 11978 6831 12034 6840
rect 11612 6802 11664 6808
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11808 5710 11836 6054
rect 12084 5930 12112 9007
rect 12348 8978 12400 8984
rect 12256 8900 12308 8906
rect 12256 8842 12308 8848
rect 12268 8022 12296 8842
rect 12360 8634 12388 8978
rect 12348 8628 12400 8634
rect 12348 8570 12400 8576
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12256 8016 12308 8022
rect 12256 7958 12308 7964
rect 12268 7546 12296 7958
rect 12544 7886 12572 8434
rect 12532 7880 12584 7886
rect 12532 7822 12584 7828
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12268 7002 12296 7482
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 12164 6860 12216 6866
rect 12164 6802 12216 6808
rect 12176 6458 12204 6802
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 11992 5902 12112 5930
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11808 5370 11836 5646
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11704 4684 11756 4690
rect 11704 4626 11756 4632
rect 11716 3942 11744 4626
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 11518 3496 11574 3505
rect 11518 3431 11574 3440
rect 11428 3392 11480 3398
rect 11428 3334 11480 3340
rect 11336 3188 11388 3194
rect 11336 3130 11388 3136
rect 11440 3058 11468 3334
rect 11428 3052 11480 3058
rect 11428 2994 11480 3000
rect 11440 2582 11468 2994
rect 11428 2576 11480 2582
rect 10980 2514 11192 2530
rect 10968 2508 11192 2514
rect 11020 2502 11192 2508
rect 11242 2544 11298 2553
rect 11428 2518 11480 2524
rect 11242 2479 11298 2488
rect 10968 2450 11020 2456
rect 11334 1864 11390 1873
rect 11334 1799 11390 1808
rect 10784 1284 10836 1290
rect 10784 1226 10836 1232
rect 11348 480 11376 1799
rect 11716 1465 11744 3878
rect 11886 3224 11942 3233
rect 11886 3159 11942 3168
rect 11900 2650 11928 3159
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 11702 1456 11758 1465
rect 11702 1391 11758 1400
rect 11992 480 12020 5902
rect 12440 5840 12492 5846
rect 12440 5782 12492 5788
rect 12348 5160 12400 5166
rect 12348 5102 12400 5108
rect 12360 4826 12388 5102
rect 12452 5030 12480 5782
rect 12532 5092 12584 5098
rect 12532 5034 12584 5040
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 12452 4729 12480 4966
rect 12438 4720 12494 4729
rect 12438 4655 12494 4664
rect 12072 4616 12124 4622
rect 12072 4558 12124 4564
rect 12084 3942 12112 4558
rect 12072 3936 12124 3942
rect 12072 3878 12124 3884
rect 12084 2825 12112 3878
rect 12452 3738 12480 4655
rect 12544 4486 12572 5034
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12544 3618 12572 4422
rect 12452 3590 12572 3618
rect 12452 3058 12480 3590
rect 12636 3233 12664 10474
rect 12912 10266 12940 11455
rect 13084 10600 13136 10606
rect 13082 10568 13084 10577
rect 13136 10568 13138 10577
rect 13082 10503 13138 10512
rect 12900 10260 12952 10266
rect 12900 10202 12952 10208
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 13004 7546 13032 9318
rect 13372 9178 13400 9522
rect 13556 9178 13584 18158
rect 13818 18119 13820 18128
rect 13872 18119 13874 18128
rect 13912 18148 13964 18154
rect 13820 18090 13872 18096
rect 13912 18090 13964 18096
rect 13924 18034 13952 18090
rect 13740 18006 13952 18034
rect 13740 17202 13768 18006
rect 13728 17196 13780 17202
rect 13728 17138 13780 17144
rect 14016 16674 14044 21422
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 16868 20602 16896 21519
rect 16856 20596 16908 20602
rect 16856 20538 16908 20544
rect 17130 20496 17186 20505
rect 17130 20431 17186 20440
rect 16580 20392 16632 20398
rect 16500 20340 16580 20346
rect 16500 20334 16632 20340
rect 16500 20318 16620 20334
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14830 19408 14886 19417
rect 14830 19343 14886 19352
rect 14844 18426 14872 19343
rect 16500 19310 16528 20318
rect 17040 19848 17092 19854
rect 17040 19790 17092 19796
rect 17052 19446 17080 19790
rect 17040 19440 17092 19446
rect 17040 19382 17092 19388
rect 15292 19304 15344 19310
rect 15292 19246 15344 19252
rect 16488 19304 16540 19310
rect 17144 19258 17172 20431
rect 17512 19990 17540 27520
rect 23478 27160 23534 27169
rect 23478 27095 23534 27104
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 23492 22250 23520 27095
rect 23400 22222 23520 22250
rect 23400 22030 23428 22222
rect 23480 22092 23532 22098
rect 23480 22034 23532 22040
rect 23388 22024 23440 22030
rect 23388 21966 23440 21972
rect 23492 21486 23520 22034
rect 23480 21480 23532 21486
rect 23478 21448 23480 21457
rect 23572 21480 23624 21486
rect 23532 21448 23534 21457
rect 23572 21422 23624 21428
rect 23478 21383 23534 21392
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 17500 19984 17552 19990
rect 17500 19926 17552 19932
rect 18694 19952 18750 19961
rect 17512 19514 17540 19926
rect 18694 19887 18750 19896
rect 23480 19916 23532 19922
rect 18236 19712 18288 19718
rect 18236 19654 18288 19660
rect 17500 19508 17552 19514
rect 17500 19450 17552 19456
rect 17868 19440 17920 19446
rect 17868 19382 17920 19388
rect 16488 19246 16540 19252
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14832 18420 14884 18426
rect 14832 18362 14884 18368
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 13648 16646 14044 16674
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 13544 9172 13596 9178
rect 13544 9114 13596 9120
rect 13452 9036 13504 9042
rect 13452 8978 13504 8984
rect 13176 8900 13228 8906
rect 13176 8842 13228 8848
rect 13188 8634 13216 8842
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 12992 7540 13044 7546
rect 12992 7482 13044 7488
rect 12806 7440 12862 7449
rect 12806 7375 12808 7384
rect 12860 7375 12862 7384
rect 12808 7346 12860 7352
rect 13188 6458 13216 8570
rect 13464 8430 13492 8978
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 13556 8498 13584 8774
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 13452 8424 13504 8430
rect 13450 8392 13452 8401
rect 13504 8392 13506 8401
rect 13450 8327 13506 8336
rect 13452 7200 13504 7206
rect 13452 7142 13504 7148
rect 13464 7041 13492 7142
rect 13450 7032 13506 7041
rect 13450 6967 13452 6976
rect 13504 6967 13506 6976
rect 13452 6938 13504 6944
rect 13464 6907 13492 6938
rect 13268 6724 13320 6730
rect 13268 6666 13320 6672
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 13280 6254 13308 6666
rect 13268 6248 13320 6254
rect 13268 6190 13320 6196
rect 13544 6248 13596 6254
rect 13544 6190 13596 6196
rect 13280 6118 13308 6190
rect 13268 6112 13320 6118
rect 13268 6054 13320 6060
rect 13280 5234 13308 6054
rect 13556 5914 13584 6190
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 13268 5228 13320 5234
rect 13268 5170 13320 5176
rect 12714 5128 12770 5137
rect 12714 5063 12770 5072
rect 12622 3224 12678 3233
rect 12622 3159 12678 3168
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 12256 2916 12308 2922
rect 12256 2858 12308 2864
rect 12070 2816 12126 2825
rect 12070 2751 12126 2760
rect 12268 2281 12296 2858
rect 12452 2582 12480 2994
rect 12440 2576 12492 2582
rect 12440 2518 12492 2524
rect 12254 2272 12310 2281
rect 12254 2207 12310 2216
rect 12728 626 12756 5063
rect 13280 4826 13308 5170
rect 13542 4992 13598 5001
rect 13542 4927 13598 4936
rect 13268 4820 13320 4826
rect 13268 4762 13320 4768
rect 13556 4690 13584 4927
rect 12808 4684 12860 4690
rect 12808 4626 12860 4632
rect 13544 4684 13596 4690
rect 13544 4626 13596 4632
rect 12820 4282 12848 4626
rect 12808 4276 12860 4282
rect 12808 4218 12860 4224
rect 13082 4176 13138 4185
rect 13082 4111 13084 4120
rect 13136 4111 13138 4120
rect 13084 4082 13136 4088
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 13280 3738 13308 3878
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 13556 3670 13584 3878
rect 13544 3664 13596 3670
rect 13544 3606 13596 3612
rect 13556 3505 13584 3606
rect 13542 3496 13598 3505
rect 13464 3454 13542 3482
rect 12898 2544 12954 2553
rect 12898 2479 12900 2488
rect 12952 2479 12954 2488
rect 12900 2450 12952 2456
rect 13268 2304 13320 2310
rect 13268 2246 13320 2252
rect 12636 598 12756 626
rect 12636 480 12664 598
rect 13280 480 13308 2246
rect 13464 2145 13492 3454
rect 13648 3466 13676 16646
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15304 11354 15332 19246
rect 17052 19230 17172 19258
rect 16578 16688 16634 16697
rect 16578 16623 16580 16632
rect 16632 16623 16634 16632
rect 16580 16594 16632 16600
rect 16488 16584 16540 16590
rect 16488 16526 16540 16532
rect 15566 16144 15622 16153
rect 15566 16079 15622 16088
rect 15476 11620 15528 11626
rect 15476 11562 15528 11568
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15384 11212 15436 11218
rect 15384 11154 15436 11160
rect 13728 11144 13780 11150
rect 15292 11144 15344 11150
rect 13728 11086 13780 11092
rect 14462 11112 14518 11121
rect 13740 9518 13768 11086
rect 15292 11086 15344 11092
rect 14462 11047 14518 11056
rect 14740 11076 14792 11082
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 14280 10464 14332 10470
rect 14280 10406 14332 10412
rect 13728 9512 13780 9518
rect 13728 9454 13780 9460
rect 13832 7041 13860 10406
rect 14186 10160 14242 10169
rect 13912 10124 13964 10130
rect 14186 10095 14188 10104
rect 13912 10066 13964 10072
rect 14240 10095 14242 10104
rect 14188 10066 14240 10072
rect 13924 9722 13952 10066
rect 14094 10024 14150 10033
rect 14094 9959 14150 9968
rect 13912 9716 13964 9722
rect 13912 9658 13964 9664
rect 14004 8356 14056 8362
rect 14004 8298 14056 8304
rect 14016 7750 14044 8298
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 14016 7546 14044 7686
rect 14004 7540 14056 7546
rect 14004 7482 14056 7488
rect 13818 7032 13874 7041
rect 13818 6967 13874 6976
rect 14108 6866 14136 9959
rect 14292 7585 14320 10406
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14278 7576 14334 7585
rect 14278 7511 14334 7520
rect 14384 7342 14412 8026
rect 14372 7336 14424 7342
rect 14372 7278 14424 7284
rect 14384 7002 14412 7278
rect 14372 6996 14424 7002
rect 14372 6938 14424 6944
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 13740 3754 13768 6054
rect 14108 5914 14136 6802
rect 14280 6656 14332 6662
rect 14476 6610 14504 11047
rect 14740 11018 14792 11024
rect 14752 9654 14780 11018
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15304 10742 15332 11086
rect 15292 10736 15344 10742
rect 15292 10678 15344 10684
rect 14924 10668 14976 10674
rect 14924 10610 14976 10616
rect 14936 10266 14964 10610
rect 15304 10266 15332 10678
rect 15396 10470 15424 11154
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 14924 10260 14976 10266
rect 14844 10220 14924 10248
rect 14740 9648 14792 9654
rect 14740 9590 14792 9596
rect 14740 9444 14792 9450
rect 14740 9386 14792 9392
rect 14556 9036 14608 9042
rect 14556 8978 14608 8984
rect 14568 7750 14596 8978
rect 14752 8634 14780 9386
rect 14740 8628 14792 8634
rect 14740 8570 14792 8576
rect 14648 7948 14700 7954
rect 14648 7890 14700 7896
rect 14556 7744 14608 7750
rect 14554 7712 14556 7721
rect 14608 7712 14610 7721
rect 14554 7647 14610 7656
rect 14660 7002 14688 7890
rect 14738 7440 14794 7449
rect 14738 7375 14794 7384
rect 14556 6996 14608 7002
rect 14556 6938 14608 6944
rect 14648 6996 14700 7002
rect 14648 6938 14700 6944
rect 14280 6598 14332 6604
rect 14096 5908 14148 5914
rect 14096 5850 14148 5856
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 13740 3726 13860 3754
rect 14200 3738 14228 4762
rect 14292 4049 14320 6598
rect 14384 6582 14504 6610
rect 14384 5234 14412 6582
rect 14462 6488 14518 6497
rect 14462 6423 14518 6432
rect 14476 5302 14504 6423
rect 14464 5296 14516 5302
rect 14464 5238 14516 5244
rect 14372 5228 14424 5234
rect 14372 5170 14424 5176
rect 14464 5160 14516 5166
rect 14464 5102 14516 5108
rect 14372 5092 14424 5098
rect 14372 5034 14424 5040
rect 14384 4826 14412 5034
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 14384 4282 14412 4762
rect 14372 4276 14424 4282
rect 14372 4218 14424 4224
rect 14278 4040 14334 4049
rect 14278 3975 14334 3984
rect 13832 3670 13860 3726
rect 14188 3732 14240 3738
rect 14188 3674 14240 3680
rect 13820 3664 13872 3670
rect 13820 3606 13872 3612
rect 13542 3431 13598 3440
rect 13636 3460 13688 3466
rect 13636 3402 13688 3408
rect 13832 3194 13860 3606
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 13728 2916 13780 2922
rect 13728 2858 13780 2864
rect 13740 2666 13768 2858
rect 13820 2848 13872 2854
rect 13818 2816 13820 2825
rect 13872 2816 13874 2825
rect 14476 2802 14504 5102
rect 14568 4146 14596 6938
rect 14752 6361 14780 7375
rect 14844 7342 14872 10220
rect 14924 10202 14976 10208
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14924 9512 14976 9518
rect 14924 9454 14976 9460
rect 14936 8906 14964 9454
rect 14924 8900 14976 8906
rect 14924 8842 14976 8848
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15304 8430 15332 8774
rect 15016 8424 15068 8430
rect 15016 8366 15068 8372
rect 15292 8424 15344 8430
rect 15292 8366 15344 8372
rect 15028 7954 15056 8366
rect 15292 8288 15344 8294
rect 15396 8265 15424 10406
rect 15488 10033 15516 11562
rect 15474 10024 15530 10033
rect 15474 9959 15530 9968
rect 15476 9036 15528 9042
rect 15476 8978 15528 8984
rect 15488 8362 15516 8978
rect 15476 8356 15528 8362
rect 15476 8298 15528 8304
rect 15292 8230 15344 8236
rect 15382 8256 15438 8265
rect 15016 7948 15068 7954
rect 15016 7890 15068 7896
rect 15304 7868 15332 8230
rect 15382 8191 15438 8200
rect 15476 7880 15528 7886
rect 15304 7840 15476 7868
rect 15476 7822 15528 7828
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14832 7336 14884 7342
rect 14832 7278 14884 7284
rect 14844 6458 14872 7278
rect 15488 6730 15516 7822
rect 15476 6724 15528 6730
rect 15476 6666 15528 6672
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14832 6452 14884 6458
rect 14832 6394 14884 6400
rect 14738 6352 14794 6361
rect 14738 6287 14794 6296
rect 15580 5914 15608 16079
rect 15934 16008 15990 16017
rect 15934 15943 15990 15952
rect 15660 11688 15712 11694
rect 15660 11630 15712 11636
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 15568 5568 15620 5574
rect 15568 5510 15620 5516
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14646 5400 14702 5409
rect 14956 5392 15252 5412
rect 14646 5335 14648 5344
rect 14700 5335 14702 5344
rect 14648 5306 14700 5312
rect 14556 4140 14608 4146
rect 14556 4082 14608 4088
rect 14660 3534 14688 5306
rect 15580 5001 15608 5510
rect 15566 4992 15622 5001
rect 15566 4927 15622 4936
rect 14738 4720 14794 4729
rect 15672 4706 15700 11630
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15856 10266 15884 11086
rect 15844 10260 15896 10266
rect 15844 10202 15896 10208
rect 15750 8936 15806 8945
rect 15750 8871 15752 8880
rect 15804 8871 15806 8880
rect 15752 8842 15804 8848
rect 15752 8356 15804 8362
rect 15752 8298 15804 8304
rect 15764 6633 15792 8298
rect 15856 8022 15884 10202
rect 15844 8016 15896 8022
rect 15844 7958 15896 7964
rect 15856 7546 15884 7958
rect 15844 7540 15896 7546
rect 15844 7482 15896 7488
rect 15948 6798 15976 15943
rect 16500 15910 16528 16526
rect 16488 15904 16540 15910
rect 16488 15846 16540 15852
rect 16118 13288 16174 13297
rect 16118 13223 16174 13232
rect 16132 11694 16160 13223
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 16120 11688 16172 11694
rect 16120 11630 16172 11636
rect 16028 11552 16080 11558
rect 16028 11494 16080 11500
rect 16120 11552 16172 11558
rect 16120 11494 16172 11500
rect 16040 11257 16068 11494
rect 16026 11248 16082 11257
rect 16026 11183 16082 11192
rect 16132 10470 16160 11494
rect 16224 10810 16252 12582
rect 16394 12336 16450 12345
rect 16394 12271 16450 12280
rect 16212 10804 16264 10810
rect 16212 10746 16264 10752
rect 16224 10606 16252 10746
rect 16408 10742 16436 12271
rect 16396 10736 16448 10742
rect 16396 10678 16448 10684
rect 16212 10600 16264 10606
rect 16212 10542 16264 10548
rect 16120 10464 16172 10470
rect 16120 10406 16172 10412
rect 16028 8832 16080 8838
rect 16028 8774 16080 8780
rect 16040 8537 16068 8774
rect 16132 8634 16160 10406
rect 16396 10124 16448 10130
rect 16396 10066 16448 10072
rect 16408 9382 16436 10066
rect 16500 9761 16528 15846
rect 16856 11892 16908 11898
rect 16856 11834 16908 11840
rect 16672 11008 16724 11014
rect 16672 10950 16724 10956
rect 16684 10810 16712 10950
rect 16868 10810 16896 11834
rect 17052 11218 17080 19230
rect 17130 17640 17186 17649
rect 17130 17575 17186 17584
rect 17144 12442 17172 17575
rect 17880 14074 17908 19382
rect 17868 14068 17920 14074
rect 17868 14010 17920 14016
rect 17866 13832 17922 13841
rect 17866 13767 17922 13776
rect 17774 12880 17830 12889
rect 17774 12815 17830 12824
rect 17132 12436 17184 12442
rect 17132 12378 17184 12384
rect 17408 12300 17460 12306
rect 17408 12242 17460 12248
rect 17592 12300 17644 12306
rect 17592 12242 17644 12248
rect 17420 11558 17448 12242
rect 17604 11898 17632 12242
rect 17684 12232 17736 12238
rect 17684 12174 17736 12180
rect 17696 11898 17724 12174
rect 17592 11892 17644 11898
rect 17592 11834 17644 11840
rect 17684 11892 17736 11898
rect 17684 11834 17736 11840
rect 17408 11552 17460 11558
rect 17406 11520 17408 11529
rect 17460 11520 17462 11529
rect 17406 11455 17462 11464
rect 17040 11212 17092 11218
rect 17040 11154 17092 11160
rect 16672 10804 16724 10810
rect 16672 10746 16724 10752
rect 16856 10804 16908 10810
rect 16856 10746 16908 10752
rect 16486 9752 16542 9761
rect 16486 9687 16542 9696
rect 16396 9376 16448 9382
rect 16396 9318 16448 9324
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 16026 8528 16082 8537
rect 16082 8486 16160 8514
rect 16592 8498 16620 9318
rect 16684 8838 16712 10746
rect 17052 10266 17080 11154
rect 17132 11008 17184 11014
rect 17132 10950 17184 10956
rect 17144 10470 17172 10950
rect 17408 10668 17460 10674
rect 17408 10610 17460 10616
rect 17132 10464 17184 10470
rect 17132 10406 17184 10412
rect 17040 10260 17092 10266
rect 17040 10202 17092 10208
rect 16948 9716 17000 9722
rect 16948 9658 17000 9664
rect 16854 9616 16910 9625
rect 16854 9551 16910 9560
rect 16672 8832 16724 8838
rect 16672 8774 16724 8780
rect 16026 8463 16082 8472
rect 16132 8430 16160 8486
rect 16580 8492 16632 8498
rect 16580 8434 16632 8440
rect 16120 8424 16172 8430
rect 16120 8366 16172 8372
rect 16486 8392 16542 8401
rect 16486 8327 16542 8336
rect 16302 7848 16358 7857
rect 16302 7783 16358 7792
rect 16210 6896 16266 6905
rect 16210 6831 16266 6840
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 15936 6656 15988 6662
rect 15750 6624 15806 6633
rect 15936 6598 15988 6604
rect 15750 6559 15806 6568
rect 15948 6118 15976 6598
rect 16224 6458 16252 6831
rect 16316 6798 16344 7783
rect 16394 7712 16450 7721
rect 16394 7647 16450 7656
rect 16304 6792 16356 6798
rect 16304 6734 16356 6740
rect 16212 6452 16264 6458
rect 16212 6394 16264 6400
rect 16224 6254 16252 6394
rect 16316 6390 16344 6734
rect 16408 6458 16436 7647
rect 16500 7002 16528 8327
rect 16684 8294 16712 8774
rect 16672 8288 16724 8294
rect 16672 8230 16724 8236
rect 16762 8120 16818 8129
rect 16762 8055 16818 8064
rect 16580 7200 16632 7206
rect 16580 7142 16632 7148
rect 16672 7200 16724 7206
rect 16672 7142 16724 7148
rect 16488 6996 16540 7002
rect 16488 6938 16540 6944
rect 16592 6866 16620 7142
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16396 6452 16448 6458
rect 16396 6394 16448 6400
rect 16304 6384 16356 6390
rect 16304 6326 16356 6332
rect 16212 6248 16264 6254
rect 16212 6190 16264 6196
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 15752 5704 15804 5710
rect 15752 5646 15804 5652
rect 15764 5370 15792 5646
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 15764 4826 15792 5306
rect 15752 4820 15804 4826
rect 15752 4762 15804 4768
rect 15672 4678 15884 4706
rect 14738 4655 14794 4664
rect 14752 4457 14780 4655
rect 15476 4616 15528 4622
rect 15382 4584 15438 4593
rect 15476 4558 15528 4564
rect 15382 4519 15438 4528
rect 14738 4448 14794 4457
rect 14738 4383 14794 4392
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14740 4140 14792 4146
rect 14740 4082 14792 4088
rect 14648 3528 14700 3534
rect 14648 3470 14700 3476
rect 13818 2751 13874 2760
rect 14384 2774 14504 2802
rect 14384 2666 14412 2774
rect 13740 2650 13860 2666
rect 13740 2644 13872 2650
rect 13740 2638 13820 2644
rect 14384 2638 14596 2666
rect 13820 2586 13872 2592
rect 13450 2136 13506 2145
rect 13450 2071 13506 2080
rect 13912 1284 13964 1290
rect 13912 1226 13964 1232
rect 13924 480 13952 1226
rect 14568 480 14596 2638
rect 14660 2514 14688 3470
rect 14752 2650 14780 4082
rect 15290 4040 15346 4049
rect 15290 3975 15346 3984
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14740 2644 14792 2650
rect 14740 2586 14792 2592
rect 14648 2508 14700 2514
rect 14648 2450 14700 2456
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 15304 1170 15332 3975
rect 15396 3670 15424 4519
rect 15488 4078 15516 4558
rect 15476 4072 15528 4078
rect 15476 4014 15528 4020
rect 15488 3738 15516 4014
rect 15476 3732 15528 3738
rect 15476 3674 15528 3680
rect 15384 3664 15436 3670
rect 15384 3606 15436 3612
rect 15396 3194 15424 3606
rect 15488 3602 15516 3674
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15488 3058 15516 3538
rect 15476 3052 15528 3058
rect 15476 2994 15528 3000
rect 15488 2514 15516 2994
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 15212 1142 15332 1170
rect 15212 480 15240 1142
rect 15856 480 15884 4678
rect 15948 2825 15976 6054
rect 16212 5772 16264 5778
rect 16212 5714 16264 5720
rect 16224 5302 16252 5714
rect 16212 5296 16264 5302
rect 16212 5238 16264 5244
rect 16396 5228 16448 5234
rect 16396 5170 16448 5176
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 16028 4684 16080 4690
rect 16028 4626 16080 4632
rect 16040 4282 16068 4626
rect 16028 4276 16080 4282
rect 16028 4218 16080 4224
rect 16132 3534 16160 4966
rect 16408 4826 16436 5170
rect 16396 4820 16448 4826
rect 16396 4762 16448 4768
rect 16408 4078 16436 4762
rect 16684 4298 16712 7142
rect 16500 4270 16712 4298
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16500 3924 16528 4270
rect 16408 3896 16528 3924
rect 16120 3528 16172 3534
rect 16118 3496 16120 3505
rect 16172 3496 16174 3505
rect 16118 3431 16174 3440
rect 16132 3194 16160 3431
rect 16120 3188 16172 3194
rect 16120 3130 16172 3136
rect 15934 2816 15990 2825
rect 15934 2751 15990 2760
rect 15948 2582 15976 2751
rect 15936 2576 15988 2582
rect 15936 2518 15988 2524
rect 16408 1034 16436 3896
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 16500 2922 16528 3470
rect 16488 2916 16540 2922
rect 16488 2858 16540 2864
rect 16500 2650 16528 2858
rect 16488 2644 16540 2650
rect 16488 2586 16540 2592
rect 16776 1834 16804 8055
rect 16868 6202 16896 9551
rect 16960 9110 16988 9658
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 16948 9104 17000 9110
rect 16948 9046 17000 9052
rect 16960 8634 16988 9046
rect 16948 8628 17000 8634
rect 16948 8570 17000 8576
rect 16960 8090 16988 8570
rect 17052 8362 17080 9318
rect 17040 8356 17092 8362
rect 17040 8298 17092 8304
rect 17144 8265 17172 10406
rect 17420 9722 17448 10610
rect 17592 10600 17644 10606
rect 17592 10542 17644 10548
rect 17604 10198 17632 10542
rect 17592 10192 17644 10198
rect 17592 10134 17644 10140
rect 17408 9716 17460 9722
rect 17408 9658 17460 9664
rect 17224 9512 17276 9518
rect 17224 9454 17276 9460
rect 17684 9512 17736 9518
rect 17684 9454 17736 9460
rect 17130 8256 17186 8265
rect 17130 8191 17186 8200
rect 17236 8090 17264 9454
rect 17696 9042 17724 9454
rect 17684 9036 17736 9042
rect 17684 8978 17736 8984
rect 17498 8528 17554 8537
rect 17498 8463 17554 8472
rect 16948 8084 17000 8090
rect 16948 8026 17000 8032
rect 17224 8084 17276 8090
rect 17224 8026 17276 8032
rect 17406 7984 17462 7993
rect 17406 7919 17462 7928
rect 17222 7576 17278 7585
rect 17420 7546 17448 7919
rect 17222 7511 17278 7520
rect 17408 7540 17460 7546
rect 17236 7177 17264 7511
rect 17408 7482 17460 7488
rect 17420 7342 17448 7482
rect 17408 7336 17460 7342
rect 17408 7278 17460 7284
rect 17222 7168 17278 7177
rect 17406 7168 17462 7177
rect 17222 7103 17278 7112
rect 17328 7126 17406 7154
rect 17038 7032 17094 7041
rect 17328 7018 17356 7126
rect 17406 7103 17462 7112
rect 17094 6990 17356 7018
rect 17038 6967 17094 6976
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 17222 6352 17278 6361
rect 17222 6287 17278 6296
rect 16868 6174 17080 6202
rect 16856 6112 16908 6118
rect 16856 6054 16908 6060
rect 16868 5574 16896 6054
rect 16856 5568 16908 5574
rect 16856 5510 16908 5516
rect 16948 5024 17000 5030
rect 16948 4966 17000 4972
rect 16960 4729 16988 4966
rect 16946 4720 17002 4729
rect 16946 4655 17002 4664
rect 17052 3466 17080 6174
rect 17236 5817 17264 6287
rect 17420 5914 17448 6802
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 17222 5808 17278 5817
rect 17222 5743 17278 5752
rect 17130 4992 17186 5001
rect 17130 4927 17186 4936
rect 17144 3942 17172 4927
rect 17420 4622 17448 5850
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 17132 3936 17184 3942
rect 17132 3878 17184 3884
rect 17408 3936 17460 3942
rect 17408 3878 17460 3884
rect 17224 3732 17276 3738
rect 17224 3674 17276 3680
rect 17040 3460 17092 3466
rect 17040 3402 17092 3408
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 16868 2553 16896 3130
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 16854 2544 16910 2553
rect 16854 2479 16910 2488
rect 16764 1828 16816 1834
rect 16764 1770 16816 1776
rect 16408 1006 16528 1034
rect 16500 480 16528 1006
rect 17052 626 17080 2994
rect 17236 2650 17264 3674
rect 17420 3602 17448 3878
rect 17408 3596 17460 3602
rect 17408 3538 17460 3544
rect 17420 2650 17448 3538
rect 17512 3058 17540 8463
rect 17696 8090 17724 8978
rect 17684 8084 17736 8090
rect 17684 8026 17736 8032
rect 17592 7336 17644 7342
rect 17592 7278 17644 7284
rect 17604 6866 17632 7278
rect 17684 7200 17736 7206
rect 17684 7142 17736 7148
rect 17592 6860 17644 6866
rect 17592 6802 17644 6808
rect 17592 6656 17644 6662
rect 17592 6598 17644 6604
rect 17604 6254 17632 6598
rect 17696 6322 17724 7142
rect 17684 6316 17736 6322
rect 17684 6258 17736 6264
rect 17592 6248 17644 6254
rect 17592 6190 17644 6196
rect 17684 5160 17736 5166
rect 17682 5128 17684 5137
rect 17736 5128 17738 5137
rect 17682 5063 17738 5072
rect 17590 3768 17646 3777
rect 17590 3703 17646 3712
rect 17604 3670 17632 3703
rect 17592 3664 17644 3670
rect 17592 3606 17644 3612
rect 17604 3126 17632 3606
rect 17592 3120 17644 3126
rect 17592 3062 17644 3068
rect 17500 3052 17552 3058
rect 17500 2994 17552 3000
rect 17224 2644 17276 2650
rect 17224 2586 17276 2592
rect 17408 2644 17460 2650
rect 17408 2586 17460 2592
rect 17052 598 17172 626
rect 17144 480 17172 598
rect 17788 480 17816 12815
rect 17880 11121 17908 13767
rect 17960 11892 18012 11898
rect 17960 11834 18012 11840
rect 17866 11112 17922 11121
rect 17866 11047 17922 11056
rect 17972 10266 18000 11834
rect 18052 11008 18104 11014
rect 18052 10950 18104 10956
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 17866 9616 17922 9625
rect 17866 9551 17868 9560
rect 17920 9551 17922 9560
rect 17868 9522 17920 9528
rect 17972 9450 18000 10202
rect 18064 10130 18092 10950
rect 18052 10124 18104 10130
rect 18052 10066 18104 10072
rect 18064 9654 18092 10066
rect 18052 9648 18104 9654
rect 18052 9590 18104 9596
rect 17960 9444 18012 9450
rect 17960 9386 18012 9392
rect 17972 9178 18000 9386
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 17868 8832 17920 8838
rect 17920 8780 18184 8786
rect 17868 8774 18184 8780
rect 17880 8758 18184 8774
rect 18052 8288 18104 8294
rect 18052 8230 18104 8236
rect 17960 7948 18012 7954
rect 17960 7890 18012 7896
rect 17972 7750 18000 7890
rect 17960 7744 18012 7750
rect 17958 7712 17960 7721
rect 18012 7712 18014 7721
rect 17958 7647 18014 7656
rect 17960 6860 18012 6866
rect 17960 6802 18012 6808
rect 17972 6458 18000 6802
rect 17960 6452 18012 6458
rect 17960 6394 18012 6400
rect 17972 5914 18000 6394
rect 17960 5908 18012 5914
rect 17960 5850 18012 5856
rect 17868 5568 17920 5574
rect 17920 5528 18000 5556
rect 17868 5510 17920 5516
rect 17972 5370 18000 5528
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 18064 5302 18092 8230
rect 18156 6746 18184 8758
rect 18248 6866 18276 19654
rect 18328 14068 18380 14074
rect 18328 14010 18380 14016
rect 18340 12442 18368 14010
rect 18512 13388 18564 13394
rect 18512 13330 18564 13336
rect 18524 12986 18552 13330
rect 18512 12980 18564 12986
rect 18512 12922 18564 12928
rect 18708 12594 18736 19887
rect 23480 19858 23532 19864
rect 23492 19174 23520 19858
rect 23480 19168 23532 19174
rect 23480 19110 23532 19116
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 22926 17912 22982 17921
rect 22926 17847 22982 17856
rect 19154 17776 19210 17785
rect 19154 17711 19210 17720
rect 19168 13530 19196 17711
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 22940 16794 22968 17847
rect 23492 17785 23520 19110
rect 23478 17776 23534 17785
rect 23478 17711 23534 17720
rect 23478 16824 23534 16833
rect 22928 16788 22980 16794
rect 23478 16759 23534 16768
rect 22928 16730 22980 16736
rect 22744 16652 22796 16658
rect 22744 16594 22796 16600
rect 22756 15910 22784 16594
rect 23492 16130 23520 16759
rect 23584 16153 23612 21422
rect 23676 19394 23704 27639
rect 24490 27520 24546 28000
rect 24504 27418 24532 27520
rect 24504 27390 24808 27418
rect 24674 25392 24730 25401
rect 24674 25327 24730 25336
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24122 24848 24178 24857
rect 24122 24783 24178 24792
rect 24136 23322 24164 24783
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24688 23866 24716 25327
rect 24780 24410 24808 27390
rect 24950 26616 25006 26625
rect 24950 26551 25006 26560
rect 24768 24404 24820 24410
rect 24768 24346 24820 24352
rect 24766 24168 24822 24177
rect 24766 24103 24768 24112
rect 24820 24103 24822 24112
rect 24768 24074 24820 24080
rect 24766 23896 24822 23905
rect 24676 23860 24728 23866
rect 24766 23831 24822 23840
rect 24676 23802 24728 23808
rect 24398 23760 24454 23769
rect 24398 23695 24400 23704
rect 24452 23695 24454 23704
rect 24400 23666 24452 23672
rect 24124 23316 24176 23322
rect 24124 23258 24176 23264
rect 23848 23180 23900 23186
rect 23848 23122 23900 23128
rect 23860 22438 23888 23122
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24780 22778 24808 23831
rect 24768 22772 24820 22778
rect 24768 22714 24820 22720
rect 24582 22672 24638 22681
rect 24582 22607 24638 22616
rect 24596 22574 24624 22607
rect 24584 22568 24636 22574
rect 24584 22510 24636 22516
rect 23848 22432 23900 22438
rect 23848 22374 23900 22380
rect 23860 22166 23888 22374
rect 23848 22160 23900 22166
rect 23848 22102 23900 22108
rect 24860 22092 24912 22098
rect 24860 22034 24912 22040
rect 24216 22024 24268 22030
rect 24216 21966 24268 21972
rect 24674 21992 24730 22001
rect 23756 21480 23808 21486
rect 23756 21422 23808 21428
rect 23768 20942 23796 21422
rect 23848 21004 23900 21010
rect 23848 20946 23900 20952
rect 23756 20936 23808 20942
rect 23756 20878 23808 20884
rect 23860 20262 23888 20946
rect 23940 20392 23992 20398
rect 23940 20334 23992 20340
rect 23848 20256 23900 20262
rect 23848 20198 23900 20204
rect 23860 19961 23888 20198
rect 23846 19952 23902 19961
rect 23846 19887 23902 19896
rect 23676 19366 23796 19394
rect 23952 19378 23980 20334
rect 23664 19304 23716 19310
rect 23664 19246 23716 19252
rect 23676 17649 23704 19246
rect 23662 17640 23718 17649
rect 23662 17575 23718 17584
rect 23400 16102 23520 16130
rect 23570 16144 23626 16153
rect 22192 15904 22244 15910
rect 22192 15846 22244 15852
rect 22744 15904 22796 15910
rect 22744 15846 22796 15852
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 22204 15638 22232 15846
rect 23400 15706 23428 16102
rect 23570 16079 23626 16088
rect 23664 16040 23716 16046
rect 23662 16008 23664 16017
rect 23716 16008 23718 16017
rect 23662 15943 23718 15952
rect 23388 15700 23440 15706
rect 23388 15642 23440 15648
rect 22192 15632 22244 15638
rect 22192 15574 22244 15580
rect 21916 15564 21968 15570
rect 21916 15506 21968 15512
rect 23204 15564 23256 15570
rect 23204 15506 23256 15512
rect 21928 14822 21956 15506
rect 23216 14822 23244 15506
rect 21916 14816 21968 14822
rect 21916 14758 21968 14764
rect 22468 14816 22520 14822
rect 22468 14758 22520 14764
rect 23204 14816 23256 14822
rect 23204 14758 23256 14764
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 21928 14521 21956 14758
rect 22480 14550 22508 14758
rect 22468 14544 22520 14550
rect 21914 14512 21970 14521
rect 22468 14486 22520 14492
rect 21914 14447 21970 14456
rect 22744 14476 22796 14482
rect 22744 14418 22796 14424
rect 22756 13870 22784 14418
rect 23018 14376 23074 14385
rect 23018 14311 23074 14320
rect 22744 13864 22796 13870
rect 22744 13806 22796 13812
rect 19248 13728 19300 13734
rect 19248 13670 19300 13676
rect 19524 13728 19576 13734
rect 19524 13670 19576 13676
rect 21640 13728 21692 13734
rect 21640 13670 21692 13676
rect 22100 13728 22152 13734
rect 22100 13670 22152 13676
rect 19156 13524 19208 13530
rect 19156 13466 19208 13472
rect 19260 13326 19288 13670
rect 19536 13394 19564 13670
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19524 13388 19576 13394
rect 19524 13330 19576 13336
rect 19248 13320 19300 13326
rect 19248 13262 19300 13268
rect 20076 13320 20128 13326
rect 20076 13262 20128 13268
rect 21548 13320 21600 13326
rect 21548 13262 21600 13268
rect 19260 12986 19288 13262
rect 19524 13252 19576 13258
rect 19524 13194 19576 13200
rect 19432 13184 19484 13190
rect 19432 13126 19484 13132
rect 19248 12980 19300 12986
rect 19248 12922 19300 12928
rect 19340 12912 19392 12918
rect 19340 12854 19392 12860
rect 19156 12776 19208 12782
rect 18786 12744 18842 12753
rect 19156 12718 19208 12724
rect 18786 12679 18788 12688
rect 18840 12679 18842 12688
rect 18788 12650 18840 12656
rect 19062 12608 19118 12617
rect 18708 12566 18828 12594
rect 18328 12436 18380 12442
rect 18328 12378 18380 12384
rect 18340 11694 18368 12378
rect 18604 12096 18656 12102
rect 18604 12038 18656 12044
rect 18328 11688 18380 11694
rect 18328 11630 18380 11636
rect 18510 10976 18566 10985
rect 18510 10911 18566 10920
rect 18524 8090 18552 10911
rect 18616 10266 18644 12038
rect 18696 10532 18748 10538
rect 18696 10474 18748 10480
rect 18708 10266 18736 10474
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 18604 10124 18656 10130
rect 18604 10066 18656 10072
rect 18616 8838 18644 10066
rect 18708 9994 18736 10202
rect 18696 9988 18748 9994
rect 18696 9930 18748 9936
rect 18604 8832 18656 8838
rect 18604 8774 18656 8780
rect 18512 8084 18564 8090
rect 18512 8026 18564 8032
rect 18326 7712 18382 7721
rect 18326 7647 18382 7656
rect 18340 7177 18368 7647
rect 18326 7168 18382 7177
rect 18326 7103 18382 7112
rect 18236 6860 18288 6866
rect 18236 6802 18288 6808
rect 18156 6718 18276 6746
rect 18248 5778 18276 6718
rect 18616 6644 18644 8774
rect 18524 6616 18644 6644
rect 18328 6248 18380 6254
rect 18328 6190 18380 6196
rect 18340 5914 18368 6190
rect 18328 5908 18380 5914
rect 18328 5850 18380 5856
rect 18236 5772 18288 5778
rect 18236 5714 18288 5720
rect 18144 5704 18196 5710
rect 18144 5646 18196 5652
rect 18052 5296 18104 5302
rect 18052 5238 18104 5244
rect 18156 5137 18184 5646
rect 18142 5128 18198 5137
rect 18142 5063 18144 5072
rect 18196 5063 18198 5072
rect 18144 5034 18196 5040
rect 18156 5003 18184 5034
rect 18418 4720 18474 4729
rect 18328 4684 18380 4690
rect 18418 4655 18474 4664
rect 18328 4626 18380 4632
rect 17868 4616 17920 4622
rect 17868 4558 17920 4564
rect 17880 4146 17908 4558
rect 18340 4214 18368 4626
rect 18328 4208 18380 4214
rect 18328 4150 18380 4156
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 17880 3738 17908 4082
rect 17868 3732 17920 3738
rect 17868 3674 17920 3680
rect 18052 3732 18104 3738
rect 18052 3674 18104 3680
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 17880 3194 17908 3470
rect 17868 3188 17920 3194
rect 17868 3130 17920 3136
rect 18064 3058 18092 3674
rect 18052 3052 18104 3058
rect 18052 2994 18104 3000
rect 18144 2916 18196 2922
rect 18144 2858 18196 2864
rect 18156 2650 18184 2858
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 18432 480 18460 4655
rect 18524 2310 18552 6616
rect 18604 5636 18656 5642
rect 18604 5578 18656 5584
rect 18616 5234 18644 5578
rect 18604 5228 18656 5234
rect 18604 5170 18656 5176
rect 18616 4758 18644 5170
rect 18604 4752 18656 4758
rect 18604 4694 18656 4700
rect 18800 3942 18828 12566
rect 19062 12543 19118 12552
rect 19076 12442 19104 12543
rect 19064 12436 19116 12442
rect 19064 12378 19116 12384
rect 18880 11688 18932 11694
rect 18880 11630 18932 11636
rect 18892 11218 18920 11630
rect 19168 11370 19196 12718
rect 19352 12617 19380 12854
rect 19444 12782 19472 13126
rect 19536 12850 19564 13194
rect 19524 12844 19576 12850
rect 19524 12786 19576 12792
rect 19432 12776 19484 12782
rect 19432 12718 19484 12724
rect 19338 12608 19394 12617
rect 19338 12543 19394 12552
rect 19248 12368 19300 12374
rect 19340 12368 19392 12374
rect 19300 12328 19340 12356
rect 19248 12310 19300 12316
rect 19340 12310 19392 12316
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 19444 11762 19472 12242
rect 19432 11756 19484 11762
rect 19432 11698 19484 11704
rect 19340 11620 19392 11626
rect 19340 11562 19392 11568
rect 19076 11342 19196 11370
rect 18880 11212 18932 11218
rect 18880 11154 18932 11160
rect 18892 10606 18920 11154
rect 18880 10600 18932 10606
rect 18880 10542 18932 10548
rect 19076 10130 19104 11342
rect 19156 11212 19208 11218
rect 19156 11154 19208 11160
rect 19168 10810 19196 11154
rect 19156 10804 19208 10810
rect 19156 10746 19208 10752
rect 19064 10124 19116 10130
rect 19064 10066 19116 10072
rect 19076 9625 19104 10066
rect 19168 10062 19196 10746
rect 19352 10742 19380 11562
rect 19340 10736 19392 10742
rect 19340 10678 19392 10684
rect 19156 10056 19208 10062
rect 19156 9998 19208 10004
rect 19156 9920 19208 9926
rect 19156 9862 19208 9868
rect 19062 9616 19118 9625
rect 19062 9551 19118 9560
rect 19168 9518 19196 9862
rect 19248 9716 19300 9722
rect 19248 9658 19300 9664
rect 19156 9512 19208 9518
rect 19156 9454 19208 9460
rect 19260 9160 19288 9658
rect 19536 9654 19564 12786
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 20088 12374 20116 13262
rect 21180 13184 21232 13190
rect 21180 13126 21232 13132
rect 21192 12850 21220 13126
rect 21270 13016 21326 13025
rect 21270 12951 21272 12960
rect 21324 12951 21326 12960
rect 21272 12922 21324 12928
rect 21180 12844 21232 12850
rect 21180 12786 21232 12792
rect 20536 12640 20588 12646
rect 20536 12582 20588 12588
rect 20076 12368 20128 12374
rect 20076 12310 20128 12316
rect 19616 12232 19668 12238
rect 19616 12174 19668 12180
rect 19628 11626 19656 12174
rect 19616 11620 19668 11626
rect 19616 11562 19668 11568
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19708 10056 19760 10062
rect 19708 9998 19760 10004
rect 19720 9722 19748 9998
rect 19708 9716 19760 9722
rect 19708 9658 19760 9664
rect 20088 9654 20116 12310
rect 20168 12096 20220 12102
rect 20168 12038 20220 12044
rect 20180 11694 20208 12038
rect 20168 11688 20220 11694
rect 20168 11630 20220 11636
rect 20180 11150 20208 11630
rect 20260 11620 20312 11626
rect 20260 11562 20312 11568
rect 20272 11354 20300 11562
rect 20548 11354 20576 12582
rect 21192 12374 21220 12786
rect 21284 12646 21312 12922
rect 21364 12708 21416 12714
rect 21364 12650 21416 12656
rect 21272 12640 21324 12646
rect 21272 12582 21324 12588
rect 21180 12368 21232 12374
rect 21180 12310 21232 12316
rect 21192 11898 21220 12310
rect 21272 12096 21324 12102
rect 21272 12038 21324 12044
rect 21180 11892 21232 11898
rect 21180 11834 21232 11840
rect 21192 11354 21220 11834
rect 20260 11348 20312 11354
rect 20260 11290 20312 11296
rect 20536 11348 20588 11354
rect 20536 11290 20588 11296
rect 21180 11348 21232 11354
rect 21180 11290 21232 11296
rect 20168 11144 20220 11150
rect 20168 11086 20220 11092
rect 20180 10266 20208 11086
rect 20548 10674 20576 11290
rect 20902 11248 20958 11257
rect 20902 11183 20958 11192
rect 21178 11248 21234 11257
rect 21178 11183 21234 11192
rect 20916 10742 20944 11183
rect 20904 10736 20956 10742
rect 20904 10678 20956 10684
rect 20536 10668 20588 10674
rect 20536 10610 20588 10616
rect 20258 10568 20314 10577
rect 20258 10503 20314 10512
rect 20272 10470 20300 10503
rect 20260 10464 20312 10470
rect 20260 10406 20312 10412
rect 20168 10260 20220 10266
rect 20168 10202 20220 10208
rect 20180 9761 20208 10202
rect 20260 10192 20312 10198
rect 20260 10134 20312 10140
rect 20166 9752 20222 9761
rect 20166 9687 20222 9696
rect 19524 9648 19576 9654
rect 19524 9590 19576 9596
rect 20076 9648 20128 9654
rect 20076 9590 20128 9596
rect 19260 9132 19380 9160
rect 18972 9036 19024 9042
rect 18972 8978 19024 8984
rect 18880 8832 18932 8838
rect 18880 8774 18932 8780
rect 18892 8401 18920 8774
rect 18878 8392 18934 8401
rect 18984 8362 19012 8978
rect 19248 8900 19300 8906
rect 19248 8842 19300 8848
rect 19156 8424 19208 8430
rect 19156 8366 19208 8372
rect 18878 8327 18934 8336
rect 18972 8356 19024 8362
rect 18972 8298 19024 8304
rect 18984 7970 19012 8298
rect 18892 7942 19012 7970
rect 18892 5386 18920 7942
rect 18972 7880 19024 7886
rect 18972 7822 19024 7828
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 18984 6458 19012 7822
rect 19076 7546 19104 7822
rect 19064 7540 19116 7546
rect 19064 7482 19116 7488
rect 19168 7342 19196 8366
rect 19260 7750 19288 8842
rect 19352 8838 19380 9132
rect 19432 9104 19484 9110
rect 19432 9046 19484 9052
rect 19340 8832 19392 8838
rect 19340 8774 19392 8780
rect 19444 8634 19472 9046
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 19536 8362 19564 9590
rect 20180 9518 20208 9687
rect 20168 9512 20220 9518
rect 20168 9454 20220 9460
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 20272 9178 20300 10134
rect 20718 9616 20774 9625
rect 20718 9551 20774 9560
rect 20352 9512 20404 9518
rect 20352 9454 20404 9460
rect 20260 9172 20312 9178
rect 20260 9114 20312 9120
rect 19524 8356 19576 8362
rect 19524 8298 19576 8304
rect 19430 8120 19486 8129
rect 19536 8090 19564 8298
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19430 8055 19486 8064
rect 19524 8084 19576 8090
rect 19248 7744 19300 7750
rect 19248 7686 19300 7692
rect 19156 7336 19208 7342
rect 19260 7324 19288 7686
rect 19444 7478 19472 8055
rect 19524 8026 19576 8032
rect 20272 7954 20300 9114
rect 20364 8634 20392 9454
rect 20732 8634 20760 9551
rect 21192 9178 21220 11183
rect 21284 10266 21312 12038
rect 21376 11898 21404 12650
rect 21364 11892 21416 11898
rect 21364 11834 21416 11840
rect 21364 11212 21416 11218
rect 21364 11154 21416 11160
rect 21376 10810 21404 11154
rect 21364 10804 21416 10810
rect 21364 10746 21416 10752
rect 21272 10260 21324 10266
rect 21272 10202 21324 10208
rect 21180 9172 21232 9178
rect 21180 9114 21232 9120
rect 21272 9036 21324 9042
rect 21272 8978 21324 8984
rect 21284 8634 21312 8978
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 20720 8628 20772 8634
rect 20720 8570 20772 8576
rect 21272 8628 21324 8634
rect 21272 8570 21324 8576
rect 20352 8492 20404 8498
rect 20352 8434 20404 8440
rect 20260 7948 20312 7954
rect 20260 7890 20312 7896
rect 19984 7812 20036 7818
rect 19984 7754 20036 7760
rect 19524 7540 19576 7546
rect 19524 7482 19576 7488
rect 19432 7472 19484 7478
rect 19432 7414 19484 7420
rect 19260 7296 19380 7324
rect 19156 7278 19208 7284
rect 19352 6934 19380 7296
rect 19340 6928 19392 6934
rect 19392 6888 19472 6916
rect 19340 6870 19392 6876
rect 19064 6656 19116 6662
rect 19064 6598 19116 6604
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 18972 6452 19024 6458
rect 18972 6394 19024 6400
rect 19076 6322 19104 6598
rect 19352 6458 19380 6598
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19064 6316 19116 6322
rect 19064 6258 19116 6264
rect 19248 6248 19300 6254
rect 19248 6190 19300 6196
rect 19260 6066 19288 6190
rect 19260 6038 19380 6066
rect 19260 5846 19288 6038
rect 19248 5840 19300 5846
rect 19248 5782 19300 5788
rect 18970 5400 19026 5409
rect 18892 5358 18970 5386
rect 19352 5370 19380 6038
rect 18970 5335 19026 5344
rect 19340 5364 19392 5370
rect 18984 5166 19012 5335
rect 19340 5306 19392 5312
rect 18972 5160 19024 5166
rect 18972 5102 19024 5108
rect 18984 4826 19012 5102
rect 18972 4820 19024 4826
rect 18972 4762 19024 4768
rect 19248 4684 19300 4690
rect 19300 4644 19380 4672
rect 19248 4626 19300 4632
rect 19062 4312 19118 4321
rect 19062 4247 19118 4256
rect 18788 3936 18840 3942
rect 18788 3878 18840 3884
rect 18512 2304 18564 2310
rect 18512 2246 18564 2252
rect 19076 1034 19104 4247
rect 19156 4004 19208 4010
rect 19156 3946 19208 3952
rect 19168 3738 19196 3946
rect 19156 3732 19208 3738
rect 19156 3674 19208 3680
rect 19156 3596 19208 3602
rect 19156 3538 19208 3544
rect 19168 3233 19196 3538
rect 19352 3534 19380 4644
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 19154 3224 19210 3233
rect 19154 3159 19156 3168
rect 19208 3159 19210 3168
rect 19156 3130 19208 3136
rect 19168 3099 19196 3130
rect 19260 3126 19288 3470
rect 19248 3120 19300 3126
rect 19246 3088 19248 3097
rect 19300 3088 19302 3097
rect 19246 3023 19302 3032
rect 19260 2997 19288 3023
rect 19154 2952 19210 2961
rect 19444 2938 19472 6888
rect 19536 6458 19564 7482
rect 19996 7342 20024 7754
rect 20272 7562 20300 7890
rect 20364 7886 20392 8434
rect 20732 8430 20760 8570
rect 21272 8492 21324 8498
rect 21272 8434 21324 8440
rect 20720 8424 20772 8430
rect 20720 8366 20772 8372
rect 20812 8016 20864 8022
rect 20812 7958 20864 7964
rect 20902 7984 20958 7993
rect 20352 7880 20404 7886
rect 20352 7822 20404 7828
rect 20626 7848 20682 7857
rect 20180 7534 20300 7562
rect 19984 7336 20036 7342
rect 19984 7278 20036 7284
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 20180 7002 20208 7534
rect 20258 7440 20314 7449
rect 20258 7375 20314 7384
rect 20272 7041 20300 7375
rect 20364 7206 20392 7822
rect 20626 7783 20682 7792
rect 20640 7546 20668 7783
rect 20720 7744 20772 7750
rect 20720 7686 20772 7692
rect 20628 7540 20680 7546
rect 20628 7482 20680 7488
rect 20352 7200 20404 7206
rect 20352 7142 20404 7148
rect 20258 7032 20314 7041
rect 20168 6996 20220 7002
rect 20258 6967 20314 6976
rect 20168 6938 20220 6944
rect 19524 6452 19576 6458
rect 19524 6394 19576 6400
rect 19984 6180 20036 6186
rect 19984 6122 20036 6128
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19996 5914 20024 6122
rect 19984 5908 20036 5914
rect 19984 5850 20036 5856
rect 19982 5808 20038 5817
rect 19524 5772 19576 5778
rect 19982 5743 20038 5752
rect 19524 5714 19576 5720
rect 19536 5166 19564 5714
rect 19524 5160 19576 5166
rect 19524 5102 19576 5108
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19800 4480 19852 4486
rect 19800 4422 19852 4428
rect 19812 4214 19840 4422
rect 19800 4208 19852 4214
rect 19800 4150 19852 4156
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19154 2887 19210 2896
rect 19352 2910 19472 2938
rect 19168 2582 19196 2887
rect 19352 2650 19380 2910
rect 19432 2848 19484 2854
rect 19430 2816 19432 2825
rect 19484 2816 19486 2825
rect 19430 2751 19486 2760
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19340 2644 19392 2650
rect 19340 2586 19392 2592
rect 19156 2576 19208 2582
rect 19156 2518 19208 2524
rect 19076 1006 19196 1034
rect 19168 480 19196 1006
rect 19996 762 20024 5743
rect 20074 5672 20130 5681
rect 20074 5607 20130 5616
rect 19812 734 20024 762
rect 19812 480 19840 734
rect 20088 610 20116 5607
rect 20364 5574 20392 7142
rect 20352 5568 20404 5574
rect 20352 5510 20404 5516
rect 20364 5030 20392 5510
rect 20444 5092 20496 5098
rect 20444 5034 20496 5040
rect 20352 5024 20404 5030
rect 20352 4966 20404 4972
rect 20364 4078 20392 4966
rect 20352 4072 20404 4078
rect 20352 4014 20404 4020
rect 20456 3913 20484 5034
rect 20732 4162 20760 7686
rect 20640 4146 20760 4162
rect 20628 4140 20760 4146
rect 20680 4134 20760 4140
rect 20628 4082 20680 4088
rect 20718 4040 20774 4049
rect 20718 3975 20720 3984
rect 20772 3975 20774 3984
rect 20720 3946 20772 3952
rect 20442 3904 20498 3913
rect 20824 3890 20852 7958
rect 20902 7919 20958 7928
rect 20916 5778 20944 7919
rect 21088 7812 21140 7818
rect 21088 7754 21140 7760
rect 20996 7200 21048 7206
rect 20996 7142 21048 7148
rect 21008 6662 21036 7142
rect 21100 6866 21128 7754
rect 21180 7404 21232 7410
rect 21180 7346 21232 7352
rect 21192 7002 21220 7346
rect 21180 6996 21232 7002
rect 21180 6938 21232 6944
rect 21284 6866 21312 8434
rect 21468 8362 21496 8910
rect 21560 8673 21588 13262
rect 21652 10266 21680 13670
rect 21732 12640 21784 12646
rect 21732 12582 21784 12588
rect 21744 12306 21772 12582
rect 21732 12300 21784 12306
rect 21732 12242 21784 12248
rect 22112 10810 22140 13670
rect 22560 13320 22612 13326
rect 22560 13262 22612 13268
rect 22284 12096 22336 12102
rect 22284 12038 22336 12044
rect 22192 11552 22244 11558
rect 22192 11494 22244 11500
rect 22100 10804 22152 10810
rect 22100 10746 22152 10752
rect 22112 10606 22140 10746
rect 22204 10674 22232 11494
rect 22296 11218 22324 12038
rect 22376 11892 22428 11898
rect 22376 11834 22428 11840
rect 22388 11558 22416 11834
rect 22376 11552 22428 11558
rect 22376 11494 22428 11500
rect 22284 11212 22336 11218
rect 22284 11154 22336 11160
rect 22388 11082 22416 11494
rect 22572 11234 22600 13262
rect 22652 12912 22704 12918
rect 22650 12880 22652 12889
rect 22704 12880 22706 12889
rect 22650 12815 22706 12824
rect 22756 12442 22784 13806
rect 22744 12436 22796 12442
rect 22744 12378 22796 12384
rect 22928 12096 22980 12102
rect 22928 12038 22980 12044
rect 22652 11756 22704 11762
rect 22652 11698 22704 11704
rect 22664 11354 22692 11698
rect 22652 11348 22704 11354
rect 22652 11290 22704 11296
rect 22940 11257 22968 12038
rect 22926 11248 22982 11257
rect 22572 11206 22876 11234
rect 22376 11076 22428 11082
rect 22376 11018 22428 11024
rect 22192 10668 22244 10674
rect 22192 10610 22244 10616
rect 22560 10668 22612 10674
rect 22560 10610 22612 10616
rect 22100 10600 22152 10606
rect 22100 10542 22152 10548
rect 22204 10266 22232 10610
rect 21640 10260 21692 10266
rect 21640 10202 21692 10208
rect 22192 10260 22244 10266
rect 22192 10202 22244 10208
rect 21652 9518 21680 10202
rect 22572 10198 22600 10610
rect 21916 10192 21968 10198
rect 21916 10134 21968 10140
rect 22560 10192 22612 10198
rect 22560 10134 22612 10140
rect 21640 9512 21692 9518
rect 21640 9454 21692 9460
rect 21928 9382 21956 10134
rect 22008 10056 22060 10062
rect 22008 9998 22060 10004
rect 21640 9376 21692 9382
rect 21640 9318 21692 9324
rect 21916 9376 21968 9382
rect 21916 9318 21968 9324
rect 21546 8664 21602 8673
rect 21546 8599 21602 8608
rect 21456 8356 21508 8362
rect 21456 8298 21508 8304
rect 21088 6860 21140 6866
rect 21088 6802 21140 6808
rect 21272 6860 21324 6866
rect 21272 6802 21324 6808
rect 20996 6656 21048 6662
rect 20996 6598 21048 6604
rect 21100 6390 21128 6802
rect 21284 6458 21312 6802
rect 21364 6656 21416 6662
rect 21364 6598 21416 6604
rect 21272 6452 21324 6458
rect 21272 6394 21324 6400
rect 21088 6384 21140 6390
rect 21088 6326 21140 6332
rect 21100 5914 21128 6326
rect 21088 5908 21140 5914
rect 21088 5850 21140 5856
rect 20904 5772 20956 5778
rect 20904 5714 20956 5720
rect 20916 5370 20944 5714
rect 21088 5568 21140 5574
rect 21088 5510 21140 5516
rect 20904 5364 20956 5370
rect 20904 5306 20956 5312
rect 20996 4684 21048 4690
rect 20996 4626 21048 4632
rect 21008 4282 21036 4626
rect 20996 4276 21048 4282
rect 20996 4218 21048 4224
rect 20442 3839 20498 3848
rect 20640 3862 20852 3890
rect 20456 3369 20484 3839
rect 20640 3534 20668 3862
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 20442 3360 20498 3369
rect 20442 3295 20498 3304
rect 20640 3194 20668 3470
rect 20628 3188 20680 3194
rect 20628 3130 20680 3136
rect 20076 604 20128 610
rect 20076 546 20128 552
rect 20444 604 20496 610
rect 20444 546 20496 552
rect 20456 480 20484 546
rect 21100 480 21128 5510
rect 21284 4826 21312 6394
rect 21272 4820 21324 4826
rect 21272 4762 21324 4768
rect 21180 4480 21232 4486
rect 21180 4422 21232 4428
rect 21192 4321 21220 4422
rect 21178 4312 21234 4321
rect 21178 4247 21234 4256
rect 21284 4214 21312 4762
rect 21272 4208 21324 4214
rect 21272 4150 21324 4156
rect 21180 3664 21232 3670
rect 21180 3606 21232 3612
rect 21192 3058 21220 3606
rect 21180 3052 21232 3058
rect 21180 2994 21232 3000
rect 21192 2514 21220 2994
rect 21376 2689 21404 6598
rect 21468 3942 21496 8298
rect 21652 8022 21680 9318
rect 21928 9081 21956 9318
rect 21914 9072 21970 9081
rect 21914 9007 21970 9016
rect 22020 8974 22048 9998
rect 22652 9376 22704 9382
rect 22652 9318 22704 9324
rect 22468 9104 22520 9110
rect 22468 9046 22520 9052
rect 22008 8968 22060 8974
rect 22008 8910 22060 8916
rect 21732 8424 21784 8430
rect 21730 8392 21732 8401
rect 21784 8392 21786 8401
rect 21730 8327 21786 8336
rect 21916 8288 21968 8294
rect 21916 8230 21968 8236
rect 21732 8084 21784 8090
rect 21732 8026 21784 8032
rect 21640 8016 21692 8022
rect 21640 7958 21692 7964
rect 21652 7886 21680 7958
rect 21640 7880 21692 7886
rect 21640 7822 21692 7828
rect 21744 7206 21772 8026
rect 21928 7857 21956 8230
rect 22020 8090 22048 8910
rect 22008 8084 22060 8090
rect 22008 8026 22060 8032
rect 21914 7848 21970 7857
rect 21914 7783 21970 7792
rect 21732 7200 21784 7206
rect 21732 7142 21784 7148
rect 21744 5409 21772 7142
rect 22020 7002 22048 8026
rect 22192 7744 22244 7750
rect 22192 7686 22244 7692
rect 22204 7342 22232 7686
rect 22376 7404 22428 7410
rect 22376 7346 22428 7352
rect 22192 7336 22244 7342
rect 22388 7313 22416 7346
rect 22192 7278 22244 7284
rect 22374 7304 22430 7313
rect 22374 7239 22430 7248
rect 22008 6996 22060 7002
rect 22008 6938 22060 6944
rect 22008 5772 22060 5778
rect 22008 5714 22060 5720
rect 21730 5400 21786 5409
rect 22020 5370 22048 5714
rect 22480 5658 22508 9046
rect 22664 8537 22692 9318
rect 22650 8528 22706 8537
rect 22650 8463 22706 8472
rect 22848 8344 22876 11206
rect 22926 11183 22982 11192
rect 23032 9353 23060 14311
rect 23570 13968 23626 13977
rect 23570 13903 23626 13912
rect 23478 13424 23534 13433
rect 23478 13359 23480 13368
rect 23532 13359 23534 13368
rect 23480 13330 23532 13336
rect 23492 12986 23520 13330
rect 23480 12980 23532 12986
rect 23480 12922 23532 12928
rect 23388 12640 23440 12646
rect 23440 12600 23520 12628
rect 23388 12582 23440 12588
rect 23110 12200 23166 12209
rect 23110 12135 23166 12144
rect 23124 9654 23152 12135
rect 23492 11801 23520 12600
rect 23478 11792 23534 11801
rect 23478 11727 23534 11736
rect 23584 11642 23612 13903
rect 23662 13288 23718 13297
rect 23662 13223 23664 13232
rect 23716 13223 23718 13232
rect 23664 13194 23716 13200
rect 23664 12232 23716 12238
rect 23664 12174 23716 12180
rect 23400 11614 23612 11642
rect 23400 11558 23428 11614
rect 23388 11552 23440 11558
rect 23388 11494 23440 11500
rect 23676 11354 23704 12174
rect 23664 11348 23716 11354
rect 23664 11290 23716 11296
rect 23480 11212 23532 11218
rect 23480 11154 23532 11160
rect 23572 11212 23624 11218
rect 23572 11154 23624 11160
rect 23492 10826 23520 11154
rect 23308 10798 23520 10826
rect 23308 10130 23336 10798
rect 23584 10742 23612 11154
rect 23572 10736 23624 10742
rect 23572 10678 23624 10684
rect 23480 10668 23532 10674
rect 23480 10610 23532 10616
rect 23492 10198 23520 10610
rect 23480 10192 23532 10198
rect 23400 10152 23480 10180
rect 23296 10124 23348 10130
rect 23296 10066 23348 10072
rect 23308 9761 23336 10066
rect 23294 9752 23350 9761
rect 23294 9687 23350 9696
rect 23112 9648 23164 9654
rect 23112 9590 23164 9596
rect 23308 9586 23336 9687
rect 23296 9580 23348 9586
rect 23296 9522 23348 9528
rect 23204 9376 23256 9382
rect 23018 9344 23074 9353
rect 23204 9318 23256 9324
rect 23018 9279 23074 9288
rect 22756 8316 22876 8344
rect 22756 8242 22784 8316
rect 22756 8214 22876 8242
rect 22744 8084 22796 8090
rect 22744 8026 22796 8032
rect 22756 7002 22784 8026
rect 22848 8022 22876 8214
rect 22836 8016 22888 8022
rect 22836 7958 22888 7964
rect 22848 7546 22876 7958
rect 23032 7886 23060 9279
rect 23216 7954 23244 9318
rect 23308 9042 23336 9522
rect 23400 9178 23428 10152
rect 23480 10134 23532 10140
rect 23478 10024 23534 10033
rect 23478 9959 23534 9968
rect 23388 9172 23440 9178
rect 23388 9114 23440 9120
rect 23296 9036 23348 9042
rect 23296 8978 23348 8984
rect 23492 8786 23520 9959
rect 23400 8758 23520 8786
rect 23572 8832 23624 8838
rect 23572 8774 23624 8780
rect 23204 7948 23256 7954
rect 23204 7890 23256 7896
rect 23020 7880 23072 7886
rect 23020 7822 23072 7828
rect 23032 7546 23060 7822
rect 22836 7540 22888 7546
rect 22836 7482 22888 7488
rect 23020 7540 23072 7546
rect 23020 7482 23072 7488
rect 23204 7404 23256 7410
rect 23204 7346 23256 7352
rect 22744 6996 22796 7002
rect 22744 6938 22796 6944
rect 23216 6866 23244 7346
rect 23204 6860 23256 6866
rect 23204 6802 23256 6808
rect 23216 6458 23244 6802
rect 23204 6452 23256 6458
rect 23204 6394 23256 6400
rect 23216 6322 23244 6394
rect 23400 6390 23428 8758
rect 23478 8664 23534 8673
rect 23478 8599 23480 8608
rect 23532 8599 23534 8608
rect 23480 8570 23532 8576
rect 23492 8362 23520 8570
rect 23480 8356 23532 8362
rect 23480 8298 23532 8304
rect 23480 7948 23532 7954
rect 23480 7890 23532 7896
rect 23492 7206 23520 7890
rect 23584 7410 23612 8774
rect 23572 7404 23624 7410
rect 23572 7346 23624 7352
rect 23676 7274 23704 11290
rect 23768 9382 23796 19366
rect 23940 19372 23992 19378
rect 23940 19314 23992 19320
rect 23940 16992 23992 16998
rect 23940 16934 23992 16940
rect 23952 16114 23980 16934
rect 23940 16108 23992 16114
rect 23940 16050 23992 16056
rect 24122 15056 24178 15065
rect 24122 14991 24178 15000
rect 23848 14952 23900 14958
rect 23848 14894 23900 14900
rect 23860 12594 23888 14894
rect 24032 13864 24084 13870
rect 24032 13806 24084 13812
rect 23940 13184 23992 13190
rect 23940 13126 23992 13132
rect 23952 12986 23980 13126
rect 23940 12980 23992 12986
rect 23940 12922 23992 12928
rect 23860 12566 23949 12594
rect 23921 12356 23949 12566
rect 23860 12328 23949 12356
rect 23756 9376 23808 9382
rect 23756 9318 23808 9324
rect 23754 8936 23810 8945
rect 23754 8871 23810 8880
rect 23664 7268 23716 7274
rect 23664 7210 23716 7216
rect 23480 7200 23532 7206
rect 23480 7142 23532 7148
rect 23492 7041 23520 7142
rect 23478 7032 23534 7041
rect 23478 6967 23534 6976
rect 23480 6928 23532 6934
rect 23480 6870 23532 6876
rect 23492 6458 23520 6870
rect 23676 6746 23704 7210
rect 23584 6718 23704 6746
rect 23584 6662 23612 6718
rect 23572 6656 23624 6662
rect 23572 6598 23624 6604
rect 23480 6452 23532 6458
rect 23480 6394 23532 6400
rect 23388 6384 23440 6390
rect 23388 6326 23440 6332
rect 23204 6316 23256 6322
rect 23204 6258 23256 6264
rect 22652 6112 22704 6118
rect 22652 6054 22704 6060
rect 22664 5817 22692 6054
rect 23216 5914 23244 6258
rect 23204 5908 23256 5914
rect 23204 5850 23256 5856
rect 23480 5840 23532 5846
rect 22650 5808 22706 5817
rect 23480 5782 23532 5788
rect 22650 5743 22706 5752
rect 23492 5710 23520 5782
rect 22388 5630 22508 5658
rect 22744 5704 22796 5710
rect 22744 5646 22796 5652
rect 23480 5704 23532 5710
rect 23480 5646 23532 5652
rect 22100 5568 22152 5574
rect 22100 5510 22152 5516
rect 21730 5335 21786 5344
rect 22008 5364 22060 5370
rect 21744 4865 21772 5335
rect 22008 5306 22060 5312
rect 21822 5128 21878 5137
rect 21822 5063 21824 5072
rect 21876 5063 21878 5072
rect 21824 5034 21876 5040
rect 21730 4856 21786 4865
rect 22020 4826 22048 5306
rect 22112 5166 22140 5510
rect 22100 5160 22152 5166
rect 22100 5102 22152 5108
rect 21730 4791 21786 4800
rect 22008 4820 22060 4826
rect 22008 4762 22060 4768
rect 22388 4758 22416 5630
rect 22652 5228 22704 5234
rect 22652 5170 22704 5176
rect 22466 4992 22522 5001
rect 22466 4927 22522 4936
rect 22376 4752 22428 4758
rect 22376 4694 22428 4700
rect 22284 4684 22336 4690
rect 22284 4626 22336 4632
rect 21824 4004 21876 4010
rect 21824 3946 21876 3952
rect 21456 3936 21508 3942
rect 21456 3878 21508 3884
rect 21548 3936 21600 3942
rect 21548 3878 21600 3884
rect 21560 3754 21588 3878
rect 21468 3726 21588 3754
rect 21468 3505 21496 3726
rect 21638 3632 21694 3641
rect 21638 3567 21640 3576
rect 21692 3567 21694 3576
rect 21640 3538 21692 3544
rect 21454 3496 21510 3505
rect 21454 3431 21510 3440
rect 21468 3398 21496 3431
rect 21652 3398 21680 3538
rect 21456 3392 21508 3398
rect 21456 3334 21508 3340
rect 21640 3392 21692 3398
rect 21640 3334 21692 3340
rect 21468 3233 21496 3334
rect 21454 3224 21510 3233
rect 21454 3159 21510 3168
rect 21652 2922 21680 3334
rect 21640 2916 21692 2922
rect 21640 2858 21692 2864
rect 21362 2680 21418 2689
rect 21362 2615 21418 2624
rect 21180 2508 21232 2514
rect 21180 2450 21232 2456
rect 21652 2446 21680 2858
rect 21836 2825 21864 3946
rect 22296 3942 22324 4626
rect 22480 4185 22508 4927
rect 22558 4856 22614 4865
rect 22558 4791 22614 4800
rect 22572 4622 22600 4791
rect 22664 4622 22692 5170
rect 22756 4758 22784 5646
rect 23388 5636 23440 5642
rect 23388 5578 23440 5584
rect 23400 5250 23428 5578
rect 23492 5370 23520 5646
rect 23480 5364 23532 5370
rect 23532 5324 23612 5352
rect 23480 5306 23532 5312
rect 23400 5234 23520 5250
rect 23400 5228 23532 5234
rect 23400 5222 23480 5228
rect 23480 5170 23532 5176
rect 23388 5160 23440 5166
rect 23388 5102 23440 5108
rect 22928 5024 22980 5030
rect 22928 4966 22980 4972
rect 22744 4752 22796 4758
rect 22744 4694 22796 4700
rect 22560 4616 22612 4622
rect 22560 4558 22612 4564
rect 22652 4616 22704 4622
rect 22652 4558 22704 4564
rect 22744 4548 22796 4554
rect 22744 4490 22796 4496
rect 22756 4214 22784 4490
rect 22744 4208 22796 4214
rect 22466 4176 22522 4185
rect 22466 4111 22522 4120
rect 22742 4176 22744 4185
rect 22796 4176 22798 4185
rect 22742 4111 22798 4120
rect 22284 3936 22336 3942
rect 22284 3878 22336 3884
rect 21916 3596 21968 3602
rect 21916 3538 21968 3544
rect 21928 3194 21956 3538
rect 21916 3188 21968 3194
rect 21916 3130 21968 3136
rect 21822 2816 21878 2825
rect 21822 2751 21878 2760
rect 21640 2440 21692 2446
rect 21640 2382 21692 2388
rect 21822 2408 21878 2417
rect 21822 2343 21824 2352
rect 21876 2343 21878 2352
rect 21824 2314 21876 2320
rect 22296 1873 22324 3878
rect 22558 2952 22614 2961
rect 22558 2887 22614 2896
rect 22572 2854 22600 2887
rect 22560 2848 22612 2854
rect 22560 2790 22612 2796
rect 22940 2009 22968 4966
rect 23296 4752 23348 4758
rect 23296 4694 23348 4700
rect 23112 4616 23164 4622
rect 23112 4558 23164 4564
rect 23124 4214 23152 4558
rect 23308 4321 23336 4694
rect 23294 4312 23350 4321
rect 23294 4247 23350 4256
rect 23112 4208 23164 4214
rect 23112 4150 23164 4156
rect 23400 3890 23428 5102
rect 23584 4758 23612 5324
rect 23768 5250 23796 8871
rect 23860 5370 23888 12328
rect 24044 11234 24072 13806
rect 24136 13025 24164 14991
rect 24228 13530 24256 21966
rect 24674 21927 24730 21936
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24688 20602 24716 21927
rect 24872 21690 24900 22034
rect 24860 21684 24912 21690
rect 24860 21626 24912 21632
rect 24860 21004 24912 21010
rect 24860 20946 24912 20952
rect 24766 20904 24822 20913
rect 24766 20839 24822 20848
rect 24676 20596 24728 20602
rect 24676 20538 24728 20544
rect 24674 20360 24730 20369
rect 24674 20295 24730 20304
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24688 18970 24716 20295
rect 24780 19258 24808 20839
rect 24872 19990 24900 20946
rect 24860 19984 24912 19990
rect 24860 19926 24912 19932
rect 24964 19394 24992 26551
rect 25410 26072 25466 26081
rect 25410 26007 25466 26016
rect 25228 24268 25280 24274
rect 25228 24210 25280 24216
rect 25042 23760 25098 23769
rect 25042 23695 25098 23704
rect 25056 21962 25084 23695
rect 25240 23526 25268 24210
rect 25228 23520 25280 23526
rect 25228 23462 25280 23468
rect 25134 23216 25190 23225
rect 25134 23151 25190 23160
rect 25044 21956 25096 21962
rect 25044 21898 25096 21904
rect 25148 21690 25176 23151
rect 25240 22642 25268 23462
rect 25228 22636 25280 22642
rect 25228 22578 25280 22584
rect 25226 22536 25282 22545
rect 25226 22471 25282 22480
rect 25136 21684 25188 21690
rect 25136 21626 25188 21632
rect 25240 21146 25268 22471
rect 25228 21140 25280 21146
rect 25228 21082 25280 21088
rect 24964 19366 25084 19394
rect 24952 19304 25004 19310
rect 24780 19230 24900 19258
rect 24952 19246 25004 19252
rect 24872 19174 24900 19230
rect 24860 19168 24912 19174
rect 24766 19136 24822 19145
rect 24860 19110 24912 19116
rect 24766 19071 24822 19080
rect 24676 18964 24728 18970
rect 24676 18906 24728 18912
rect 24582 18864 24638 18873
rect 24582 18799 24584 18808
rect 24636 18799 24638 18808
rect 24584 18770 24636 18776
rect 24596 18714 24624 18770
rect 24596 18686 24716 18714
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24688 18426 24716 18686
rect 24676 18420 24728 18426
rect 24676 18362 24728 18368
rect 24674 18320 24730 18329
rect 24674 18255 24730 18264
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24688 17338 24716 18255
rect 24780 17882 24808 19071
rect 24964 18193 24992 19246
rect 24950 18184 25006 18193
rect 24950 18119 25006 18128
rect 25056 17898 25084 19366
rect 24768 17876 24820 17882
rect 24768 17818 24820 17824
rect 24964 17870 25084 17898
rect 24676 17332 24728 17338
rect 24676 17274 24728 17280
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24674 16280 24730 16289
rect 24674 16215 24730 16224
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24688 14618 24716 16215
rect 24860 16040 24912 16046
rect 24780 15988 24860 15994
rect 24780 15982 24912 15988
rect 24780 15966 24900 15982
rect 24780 15026 24808 15966
rect 24768 15020 24820 15026
rect 24768 14962 24820 14968
rect 24676 14612 24728 14618
rect 24676 14554 24728 14560
rect 24676 14476 24728 14482
rect 24676 14418 24728 14424
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24688 14074 24716 14418
rect 24676 14068 24728 14074
rect 24676 14010 24728 14016
rect 24216 13524 24268 13530
rect 24216 13466 24268 13472
rect 24676 13388 24728 13394
rect 24676 13330 24728 13336
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24122 13016 24178 13025
rect 24289 13008 24585 13028
rect 24688 12986 24716 13330
rect 24964 12986 24992 17870
rect 25044 17740 25096 17746
rect 25044 17682 25096 17688
rect 25056 16998 25084 17682
rect 25134 17504 25190 17513
rect 25134 17439 25190 17448
rect 25044 16992 25096 16998
rect 25044 16934 25096 16940
rect 25056 16697 25084 16934
rect 25042 16688 25098 16697
rect 25042 16623 25098 16632
rect 25148 16250 25176 17439
rect 25136 16244 25188 16250
rect 25136 16186 25188 16192
rect 25136 14000 25188 14006
rect 25136 13942 25188 13948
rect 25148 13841 25176 13942
rect 25134 13832 25190 13841
rect 25134 13767 25190 13776
rect 24122 12951 24178 12960
rect 24676 12980 24728 12986
rect 24676 12922 24728 12928
rect 24952 12980 25004 12986
rect 24952 12922 25004 12928
rect 24122 12880 24178 12889
rect 24122 12815 24178 12824
rect 23952 11206 24072 11234
rect 23952 10985 23980 11206
rect 24030 11112 24086 11121
rect 24030 11047 24086 11056
rect 23938 10976 23994 10985
rect 23938 10911 23994 10920
rect 23940 10464 23992 10470
rect 23940 10406 23992 10412
rect 23952 8498 23980 10406
rect 23940 8492 23992 8498
rect 23940 8434 23992 8440
rect 23938 6352 23994 6361
rect 23938 6287 23994 6296
rect 23848 5364 23900 5370
rect 23848 5306 23900 5312
rect 23768 5222 23888 5250
rect 23664 5092 23716 5098
rect 23664 5034 23716 5040
rect 23572 4752 23624 4758
rect 23572 4694 23624 4700
rect 23676 4554 23704 5034
rect 23756 4752 23808 4758
rect 23756 4694 23808 4700
rect 23664 4548 23716 4554
rect 23664 4490 23716 4496
rect 23768 4282 23796 4694
rect 23756 4276 23808 4282
rect 23756 4218 23808 4224
rect 23756 4140 23808 4146
rect 23756 4082 23808 4088
rect 23400 3862 23520 3890
rect 23492 3505 23520 3862
rect 23768 3777 23796 4082
rect 23754 3768 23810 3777
rect 23754 3703 23756 3712
rect 23808 3703 23810 3712
rect 23756 3674 23808 3680
rect 23478 3496 23534 3505
rect 23478 3431 23534 3440
rect 23662 3224 23718 3233
rect 23662 3159 23718 3168
rect 23480 2848 23532 2854
rect 23400 2796 23480 2802
rect 23400 2790 23532 2796
rect 23570 2816 23626 2825
rect 23400 2774 23520 2790
rect 23400 2650 23428 2774
rect 23570 2751 23626 2760
rect 23388 2644 23440 2650
rect 23388 2586 23440 2592
rect 23584 2514 23612 2751
rect 23572 2508 23624 2514
rect 23572 2450 23624 2456
rect 23676 2446 23704 3159
rect 23768 2922 23796 3674
rect 23756 2916 23808 2922
rect 23756 2858 23808 2864
rect 23664 2440 23716 2446
rect 23664 2382 23716 2388
rect 22374 2000 22430 2009
rect 22374 1935 22430 1944
rect 22926 2000 22982 2009
rect 22926 1935 22982 1944
rect 22282 1864 22338 1873
rect 22282 1799 22338 1808
rect 21652 598 21772 626
rect 7838 96 7894 105
rect 7838 31 7894 40
rect 8022 0 8078 480
rect 8666 0 8722 480
rect 9310 0 9366 480
rect 10046 0 10102 480
rect 10690 0 10746 480
rect 11334 0 11390 480
rect 11978 0 12034 480
rect 12622 0 12678 480
rect 13266 0 13322 480
rect 13910 0 13966 480
rect 14554 0 14610 480
rect 15198 0 15254 480
rect 15842 0 15898 480
rect 16486 0 16542 480
rect 17130 0 17186 480
rect 17774 0 17830 480
rect 18418 0 18474 480
rect 19154 0 19210 480
rect 19798 0 19854 480
rect 20442 0 20498 480
rect 21086 0 21142 480
rect 21652 241 21680 598
rect 21744 480 21772 598
rect 22388 480 22416 1935
rect 23018 1728 23074 1737
rect 23018 1663 23074 1672
rect 23032 480 23060 1663
rect 23860 898 23888 5222
rect 23952 1306 23980 6287
rect 24044 5681 24072 11047
rect 24136 10606 24164 12815
rect 24952 12776 25004 12782
rect 24952 12718 25004 12724
rect 24964 12374 24992 12718
rect 24952 12368 25004 12374
rect 24674 12336 24730 12345
rect 24952 12310 25004 12316
rect 24674 12271 24676 12280
rect 24728 12271 24730 12280
rect 24676 12242 24728 12248
rect 24216 12096 24268 12102
rect 24216 12038 24268 12044
rect 24228 11694 24256 12038
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24688 11898 24716 12242
rect 24676 11892 24728 11898
rect 24676 11834 24728 11840
rect 24216 11688 24268 11694
rect 24216 11630 24268 11636
rect 24228 11286 24256 11630
rect 24768 11552 24820 11558
rect 24768 11494 24820 11500
rect 24216 11280 24268 11286
rect 24216 11222 24268 11228
rect 24780 11218 24808 11494
rect 24768 11212 24820 11218
rect 24768 11154 24820 11160
rect 24216 11008 24268 11014
rect 24216 10950 24268 10956
rect 24124 10600 24176 10606
rect 24124 10542 24176 10548
rect 24124 10464 24176 10470
rect 24228 10418 24256 10950
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24780 10810 24808 11154
rect 24860 11008 24912 11014
rect 24860 10950 24912 10956
rect 24768 10804 24820 10810
rect 24768 10746 24820 10752
rect 24872 10674 24900 10950
rect 25424 10810 25452 26007
rect 26240 22636 26292 22642
rect 26240 22578 26292 22584
rect 25504 20256 25556 20262
rect 25504 20198 25556 20204
rect 25516 19990 25544 20198
rect 25504 19984 25556 19990
rect 25504 19926 25556 19932
rect 26252 19310 26280 22578
rect 26240 19304 26292 19310
rect 26240 19246 26292 19252
rect 26884 19304 26936 19310
rect 26884 19246 26936 19252
rect 25870 15736 25926 15745
rect 25870 15671 25926 15680
rect 25884 15162 25912 15671
rect 25872 15156 25924 15162
rect 25872 15098 25924 15104
rect 25884 14958 25912 15098
rect 25872 14952 25924 14958
rect 25872 14894 25924 14900
rect 25688 14816 25740 14822
rect 25688 14758 25740 14764
rect 25594 14648 25650 14657
rect 25594 14583 25650 14592
rect 25608 14074 25636 14583
rect 25596 14068 25648 14074
rect 25596 14010 25648 14016
rect 25608 13870 25636 14010
rect 25596 13864 25648 13870
rect 25596 13806 25648 13812
rect 25412 10804 25464 10810
rect 25412 10746 25464 10752
rect 24860 10668 24912 10674
rect 24860 10610 24912 10616
rect 25228 10600 25280 10606
rect 24674 10568 24730 10577
rect 25228 10542 25280 10548
rect 24674 10503 24730 10512
rect 24176 10412 24256 10418
rect 24124 10406 24256 10412
rect 24136 10390 24256 10406
rect 24136 7954 24164 10390
rect 24216 9920 24268 9926
rect 24216 9862 24268 9868
rect 24228 9042 24256 9862
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24688 9110 24716 10503
rect 25240 10169 25268 10542
rect 25226 10160 25282 10169
rect 25226 10095 25282 10104
rect 24952 9920 25004 9926
rect 24952 9862 25004 9868
rect 24964 9518 24992 9862
rect 24952 9512 25004 9518
rect 24952 9454 25004 9460
rect 24768 9444 24820 9450
rect 24768 9386 24820 9392
rect 24676 9104 24728 9110
rect 24676 9046 24728 9052
rect 24216 9036 24268 9042
rect 24216 8978 24268 8984
rect 24228 8634 24256 8978
rect 24674 8936 24730 8945
rect 24674 8871 24730 8880
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24216 8628 24268 8634
rect 24216 8570 24268 8576
rect 24228 8498 24256 8570
rect 24216 8492 24268 8498
rect 24216 8434 24268 8440
rect 24228 8022 24256 8434
rect 24306 8392 24362 8401
rect 24306 8327 24362 8336
rect 24216 8016 24268 8022
rect 24216 7958 24268 7964
rect 24124 7948 24176 7954
rect 24124 7890 24176 7896
rect 24122 7848 24178 7857
rect 24122 7783 24178 7792
rect 24030 5672 24086 5681
rect 24030 5607 24086 5616
rect 24030 4312 24086 4321
rect 24030 4247 24032 4256
rect 24084 4247 24086 4256
rect 24032 4218 24084 4224
rect 24032 3528 24084 3534
rect 24032 3470 24084 3476
rect 24044 3194 24072 3470
rect 24032 3188 24084 3194
rect 24032 3130 24084 3136
rect 24136 3126 24164 7783
rect 24320 7732 24348 8327
rect 24688 7993 24716 8871
rect 24780 8838 24808 9386
rect 25136 9376 25188 9382
rect 25134 9344 25136 9353
rect 25188 9344 25190 9353
rect 25134 9279 25190 9288
rect 25136 8900 25188 8906
rect 25136 8842 25188 8848
rect 24768 8832 24820 8838
rect 24768 8774 24820 8780
rect 24674 7984 24730 7993
rect 24674 7919 24730 7928
rect 24780 7886 24808 8774
rect 25148 8294 25176 8842
rect 25504 8356 25556 8362
rect 25504 8298 25556 8304
rect 25136 8288 25188 8294
rect 25136 8230 25188 8236
rect 25410 8256 25466 8265
rect 25148 8090 25176 8230
rect 25410 8191 25466 8200
rect 25136 8084 25188 8090
rect 25136 8026 25188 8032
rect 25424 7954 25452 8191
rect 25516 8129 25544 8298
rect 25502 8120 25558 8129
rect 25502 8055 25558 8064
rect 25412 7948 25464 7954
rect 25412 7890 25464 7896
rect 24768 7880 24820 7886
rect 24768 7822 24820 7828
rect 24228 7704 24348 7732
rect 24228 4146 24256 7704
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24780 7002 24808 7822
rect 25424 7546 25452 7890
rect 25412 7540 25464 7546
rect 25412 7482 25464 7488
rect 25044 7200 25096 7206
rect 25044 7142 25096 7148
rect 24768 6996 24820 7002
rect 24768 6938 24820 6944
rect 24952 6792 25004 6798
rect 24952 6734 25004 6740
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24860 5568 24912 5574
rect 24860 5510 24912 5516
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24674 5400 24730 5409
rect 24674 5335 24730 5344
rect 24688 5001 24716 5335
rect 24872 5250 24900 5510
rect 24780 5234 24900 5250
rect 24768 5228 24900 5234
rect 24820 5222 24900 5228
rect 24768 5170 24820 5176
rect 24674 4992 24730 5001
rect 24674 4927 24730 4936
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24216 4140 24268 4146
rect 24216 4082 24268 4088
rect 24216 3936 24268 3942
rect 24214 3904 24216 3913
rect 24268 3904 24270 3913
rect 24214 3839 24270 3848
rect 24124 3120 24176 3126
rect 24124 3062 24176 3068
rect 24136 2990 24164 3062
rect 24124 2984 24176 2990
rect 24124 2926 24176 2932
rect 24136 2553 24164 2926
rect 24122 2544 24178 2553
rect 24122 2479 24178 2488
rect 24228 1850 24256 3839
rect 24780 3670 24808 5170
rect 24964 4758 24992 6734
rect 25056 6458 25084 7142
rect 25044 6452 25096 6458
rect 25044 6394 25096 6400
rect 25056 6254 25084 6394
rect 25044 6248 25096 6254
rect 25044 6190 25096 6196
rect 24952 4752 25004 4758
rect 24952 4694 25004 4700
rect 25056 4690 25084 6190
rect 25228 6112 25280 6118
rect 25228 6054 25280 6060
rect 25240 5846 25268 6054
rect 25228 5840 25280 5846
rect 25228 5782 25280 5788
rect 25226 5672 25282 5681
rect 25226 5607 25282 5616
rect 25240 4690 25268 5607
rect 25596 5024 25648 5030
rect 25596 4966 25648 4972
rect 25412 4820 25464 4826
rect 25412 4762 25464 4768
rect 25424 4729 25452 4762
rect 25410 4720 25466 4729
rect 25044 4684 25096 4690
rect 25044 4626 25096 4632
rect 25228 4684 25280 4690
rect 25410 4655 25466 4664
rect 25228 4626 25280 4632
rect 25056 4146 25084 4626
rect 25240 4282 25268 4626
rect 25608 4593 25636 4966
rect 25594 4584 25650 4593
rect 25594 4519 25650 4528
rect 25228 4276 25280 4282
rect 25228 4218 25280 4224
rect 25044 4140 25096 4146
rect 25044 4082 25096 4088
rect 25700 4049 25728 14758
rect 25686 4040 25742 4049
rect 25686 3975 25742 3984
rect 26238 4040 26294 4049
rect 26238 3975 26294 3984
rect 24768 3664 24820 3670
rect 24768 3606 24820 3612
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24780 3126 24808 3606
rect 25412 3392 25464 3398
rect 25412 3334 25464 3340
rect 24768 3120 24820 3126
rect 24768 3062 24820 3068
rect 25424 3058 25452 3334
rect 24584 3052 24636 3058
rect 24584 2994 24636 3000
rect 25412 3052 25464 3058
rect 25412 2994 25464 3000
rect 24596 2446 24624 2994
rect 25412 2848 25464 2854
rect 25410 2816 25412 2825
rect 25464 2816 25466 2825
rect 25410 2751 25466 2760
rect 25594 2680 25650 2689
rect 25594 2615 25596 2624
rect 25648 2615 25650 2624
rect 25596 2586 25648 2592
rect 24768 2576 24820 2582
rect 24768 2518 24820 2524
rect 24676 2508 24728 2514
rect 24676 2450 24728 2456
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24228 1822 24440 1850
rect 23952 1278 24348 1306
rect 23676 870 23888 898
rect 23676 480 23704 870
rect 24320 480 24348 1278
rect 24412 921 24440 1822
rect 24398 912 24454 921
rect 24398 847 24454 856
rect 21638 232 21694 241
rect 21638 167 21694 176
rect 21730 0 21786 480
rect 22374 0 22430 480
rect 23018 0 23074 480
rect 23662 0 23718 480
rect 24306 0 24362 480
rect 24688 377 24716 2450
rect 24780 1465 24808 2518
rect 24766 1456 24822 1465
rect 24766 1391 24822 1400
rect 25594 1320 25650 1329
rect 25594 1255 25650 1264
rect 24872 598 24992 626
rect 24674 368 24730 377
rect 24674 303 24730 312
rect 24872 105 24900 598
rect 24964 480 24992 598
rect 25608 480 25636 1255
rect 26252 480 26280 3975
rect 26896 480 26924 19246
rect 27526 2816 27582 2825
rect 27526 2751 27582 2760
rect 27540 480 27568 2751
rect 24858 96 24914 105
rect 24858 31 24914 40
rect 24950 0 25006 480
rect 25594 0 25650 480
rect 26238 0 26294 480
rect 26882 0 26938 480
rect 27526 0 27582 480
<< via2 >>
rect 23662 27648 23718 27704
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 3514 24112 3570 24168
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 10046 21392 10102 21448
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 4158 12688 4214 12744
rect 4066 8472 4122 8528
rect 1582 7384 1638 7440
rect 294 6160 350 6216
rect 938 3440 994 3496
rect 2226 6840 2282 6896
rect 2870 4936 2926 4992
rect 3514 4120 3570 4176
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 8942 11056 8998 11112
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 6274 9424 6330 9480
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 6090 7656 6146 7712
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 4158 6296 4214 6352
rect 4066 3440 4122 3496
rect 4802 3032 4858 3088
rect 4710 1536 4766 1592
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5998 5616 6054 5672
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5630 2644 5686 2680
rect 5630 2624 5632 2644
rect 5632 2624 5684 2644
rect 5684 2624 5686 2644
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 8574 8336 8630 8392
rect 6734 7928 6790 7984
rect 6366 6704 6422 6760
rect 6642 3188 6698 3224
rect 6642 3168 6644 3188
rect 6644 3168 6696 3188
rect 6696 3168 6698 3188
rect 7010 7520 7066 7576
rect 6918 5208 6974 5264
rect 8114 7248 8170 7304
rect 7470 3984 7526 4040
rect 6826 1672 6882 1728
rect 7102 1264 7158 1320
rect 7378 1400 7434 1456
rect 7194 176 7250 232
rect 8758 6160 8814 6216
rect 8666 5752 8722 5808
rect 8298 4256 8354 4312
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 12806 23704 12862 23760
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14554 22616 14610 22672
rect 10782 20440 10838 20496
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 11610 18808 11666 18864
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 11426 17040 11482 17096
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10690 8200 10746 8256
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10782 8064 10838 8120
rect 11150 7928 11206 7984
rect 10506 7656 10562 7712
rect 10690 7656 10746 7712
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10230 5344 10286 5400
rect 9770 4972 9772 4992
rect 9772 4972 9824 4992
rect 9824 4972 9826 4992
rect 9218 4528 9274 4584
rect 8666 3576 8722 3632
rect 8114 2488 8170 2544
rect 8574 3440 8630 3496
rect 8482 2932 8484 2952
rect 8484 2932 8536 2952
rect 8536 2932 8538 2952
rect 8482 2896 8538 2932
rect 9310 3032 9366 3088
rect 8574 2080 8630 2136
rect 8298 1944 8354 2000
rect 9218 2252 9220 2272
rect 9220 2252 9272 2272
rect 9272 2252 9274 2272
rect 9218 2216 9274 2252
rect 9770 4936 9826 4972
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10874 7520 10930 7576
rect 10874 7248 10930 7304
rect 11150 7520 11206 7576
rect 10506 4664 10562 4720
rect 9586 3304 9642 3360
rect 9678 3168 9734 3224
rect 9954 3168 10010 3224
rect 10874 4800 10930 4856
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10690 2896 10746 2952
rect 9954 2624 10010 2680
rect 9402 2352 9458 2408
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 9862 1400 9918 1456
rect 11058 4392 11114 4448
rect 11058 3304 11114 3360
rect 11058 3032 11114 3088
rect 11150 2760 11206 2816
rect 11426 3884 11428 3904
rect 11428 3884 11480 3904
rect 11480 3884 11482 3904
rect 11426 3848 11482 3884
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 16854 21528 16910 21584
rect 13174 17076 13176 17096
rect 13176 17076 13228 17096
rect 13228 17076 13230 17096
rect 13174 17040 13230 17076
rect 12438 14456 12494 14512
rect 12898 11464 12954 11520
rect 12438 11056 12494 11112
rect 12070 9016 12126 9072
rect 11794 6840 11850 6896
rect 11978 6840 12034 6896
rect 11518 3440 11574 3496
rect 11242 2488 11298 2544
rect 11334 1808 11390 1864
rect 11886 3168 11942 3224
rect 11702 1400 11758 1456
rect 12438 4664 12494 4720
rect 13082 10548 13084 10568
rect 13084 10548 13136 10568
rect 13136 10548 13138 10568
rect 13082 10512 13138 10548
rect 13818 18148 13874 18184
rect 13818 18128 13820 18148
rect 13820 18128 13872 18148
rect 13872 18128 13874 18148
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 17130 20440 17186 20496
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14830 19352 14886 19408
rect 23478 27104 23534 27160
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 23478 21428 23480 21448
rect 23480 21428 23532 21448
rect 23532 21428 23534 21448
rect 23478 21392 23534 21428
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 18694 19896 18750 19952
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 12806 7404 12862 7440
rect 12806 7384 12808 7404
rect 12808 7384 12860 7404
rect 12860 7384 12862 7404
rect 13450 8372 13452 8392
rect 13452 8372 13504 8392
rect 13504 8372 13506 8392
rect 13450 8336 13506 8372
rect 13450 6996 13506 7032
rect 13450 6976 13452 6996
rect 13452 6976 13504 6996
rect 13504 6976 13506 6996
rect 12714 5072 12770 5128
rect 12622 3168 12678 3224
rect 12070 2760 12126 2816
rect 12254 2216 12310 2272
rect 13542 4936 13598 4992
rect 13082 4140 13138 4176
rect 13082 4120 13084 4140
rect 13084 4120 13136 4140
rect 13136 4120 13138 4140
rect 12898 2508 12954 2544
rect 12898 2488 12900 2508
rect 12900 2488 12952 2508
rect 12952 2488 12954 2508
rect 13542 3440 13598 3496
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 16578 16652 16634 16688
rect 16578 16632 16580 16652
rect 16580 16632 16632 16652
rect 16632 16632 16634 16652
rect 15566 16088 15622 16144
rect 14462 11056 14518 11112
rect 14186 10124 14242 10160
rect 14186 10104 14188 10124
rect 14188 10104 14240 10124
rect 14240 10104 14242 10124
rect 14094 9968 14150 10024
rect 13818 6976 13874 7032
rect 14278 7520 14334 7576
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14554 7692 14556 7712
rect 14556 7692 14608 7712
rect 14608 7692 14610 7712
rect 14554 7656 14610 7692
rect 14738 7384 14794 7440
rect 14462 6432 14518 6488
rect 14278 3984 14334 4040
rect 13818 2796 13820 2816
rect 13820 2796 13872 2816
rect 13872 2796 13874 2816
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 15474 9968 15530 10024
rect 15382 8200 15438 8256
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14738 6296 14794 6352
rect 15934 15952 15990 16008
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14646 5364 14702 5400
rect 14646 5344 14648 5364
rect 14648 5344 14700 5364
rect 14700 5344 14702 5364
rect 15566 4936 15622 4992
rect 14738 4664 14794 4720
rect 15750 8900 15806 8936
rect 15750 8880 15752 8900
rect 15752 8880 15804 8900
rect 15804 8880 15806 8900
rect 16118 13232 16174 13288
rect 16026 11192 16082 11248
rect 16394 12280 16450 12336
rect 17130 17584 17186 17640
rect 17866 13776 17922 13832
rect 17774 12824 17830 12880
rect 17406 11500 17408 11520
rect 17408 11500 17460 11520
rect 17460 11500 17462 11520
rect 17406 11464 17462 11500
rect 16486 9696 16542 9752
rect 16026 8472 16082 8528
rect 16854 9560 16910 9616
rect 16486 8336 16542 8392
rect 16302 7792 16358 7848
rect 16210 6840 16266 6896
rect 15750 6568 15806 6624
rect 16394 7656 16450 7712
rect 16762 8064 16818 8120
rect 15382 4528 15438 4584
rect 14738 4392 14794 4448
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 13818 2760 13874 2796
rect 13450 2080 13506 2136
rect 15290 3984 15346 4040
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 16118 3476 16120 3496
rect 16120 3476 16172 3496
rect 16172 3476 16174 3496
rect 16118 3440 16174 3476
rect 15934 2760 15990 2816
rect 17130 8200 17186 8256
rect 17498 8472 17554 8528
rect 17406 7928 17462 7984
rect 17222 7520 17278 7576
rect 17222 7112 17278 7168
rect 17038 6976 17094 7032
rect 17406 7112 17462 7168
rect 17222 6296 17278 6352
rect 16946 4664 17002 4720
rect 17222 5752 17278 5808
rect 17130 4936 17186 4992
rect 16854 2488 16910 2544
rect 17682 5108 17684 5128
rect 17684 5108 17736 5128
rect 17736 5108 17738 5128
rect 17682 5072 17738 5108
rect 17590 3712 17646 3768
rect 17866 11056 17922 11112
rect 17866 9580 17922 9616
rect 17866 9560 17868 9580
rect 17868 9560 17920 9580
rect 17920 9560 17922 9580
rect 17958 7692 17960 7712
rect 17960 7692 18012 7712
rect 18012 7692 18014 7712
rect 17958 7656 18014 7692
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 22926 17856 22982 17912
rect 19154 17720 19210 17776
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 23478 17720 23534 17776
rect 23478 16768 23534 16824
rect 24674 25336 24730 25392
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24122 24792 24178 24848
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24950 26560 25006 26616
rect 24766 24132 24822 24168
rect 24766 24112 24768 24132
rect 24768 24112 24820 24132
rect 24820 24112 24822 24132
rect 24766 23840 24822 23896
rect 24398 23724 24454 23760
rect 24398 23704 24400 23724
rect 24400 23704 24452 23724
rect 24452 23704 24454 23724
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24582 22616 24638 22672
rect 23846 19896 23902 19952
rect 23662 17584 23718 17640
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 23570 16088 23626 16144
rect 23662 15988 23664 16008
rect 23664 15988 23716 16008
rect 23716 15988 23718 16008
rect 23662 15952 23718 15988
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 21914 14456 21970 14512
rect 23018 14320 23074 14376
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 18786 12708 18842 12744
rect 18786 12688 18788 12708
rect 18788 12688 18840 12708
rect 18840 12688 18842 12708
rect 18510 10920 18566 10976
rect 18326 7656 18382 7712
rect 18326 7112 18382 7168
rect 18142 5092 18198 5128
rect 18142 5072 18144 5092
rect 18144 5072 18196 5092
rect 18196 5072 18198 5092
rect 18418 4664 18474 4720
rect 19062 12552 19118 12608
rect 19338 12552 19394 12608
rect 19062 9560 19118 9616
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 21270 12980 21326 13016
rect 21270 12960 21272 12980
rect 21272 12960 21324 12980
rect 21324 12960 21326 12980
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 20902 11192 20958 11248
rect 21178 11192 21234 11248
rect 20258 10512 20314 10568
rect 20166 9696 20222 9752
rect 18878 8336 18934 8392
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 20718 9560 20774 9616
rect 19430 8064 19486 8120
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 18970 5344 19026 5400
rect 19062 4256 19118 4312
rect 19154 3188 19210 3224
rect 19154 3168 19156 3188
rect 19156 3168 19208 3188
rect 19208 3168 19210 3188
rect 19246 3068 19248 3088
rect 19248 3068 19300 3088
rect 19300 3068 19302 3088
rect 19246 3032 19302 3068
rect 19154 2896 19210 2952
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 20258 7384 20314 7440
rect 20626 7792 20682 7848
rect 20258 6976 20314 7032
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19982 5752 20038 5808
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19430 2796 19432 2816
rect 19432 2796 19484 2816
rect 19484 2796 19486 2816
rect 19430 2760 19486 2796
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 20074 5616 20130 5672
rect 20718 4004 20774 4040
rect 20718 3984 20720 4004
rect 20720 3984 20772 4004
rect 20772 3984 20774 4004
rect 20442 3848 20498 3904
rect 20902 7928 20958 7984
rect 22650 12860 22652 12880
rect 22652 12860 22704 12880
rect 22704 12860 22706 12880
rect 22650 12824 22706 12860
rect 21546 8608 21602 8664
rect 20442 3304 20498 3360
rect 21178 4256 21234 4312
rect 21914 9016 21970 9072
rect 21730 8372 21732 8392
rect 21732 8372 21784 8392
rect 21784 8372 21786 8392
rect 21730 8336 21786 8372
rect 21914 7792 21970 7848
rect 22374 7248 22430 7304
rect 21730 5344 21786 5400
rect 22650 8472 22706 8528
rect 22926 11192 22982 11248
rect 23570 13912 23626 13968
rect 23478 13388 23534 13424
rect 23478 13368 23480 13388
rect 23480 13368 23532 13388
rect 23532 13368 23534 13388
rect 23110 12144 23166 12200
rect 23478 11736 23534 11792
rect 23662 13252 23718 13288
rect 23662 13232 23664 13252
rect 23664 13232 23716 13252
rect 23716 13232 23718 13252
rect 23294 9696 23350 9752
rect 23018 9288 23074 9344
rect 23478 9968 23534 10024
rect 23478 8628 23534 8664
rect 23478 8608 23480 8628
rect 23480 8608 23532 8628
rect 23532 8608 23534 8628
rect 24122 15000 24178 15056
rect 23754 8880 23810 8936
rect 23478 6976 23534 7032
rect 22650 5752 22706 5808
rect 21822 5092 21878 5128
rect 21822 5072 21824 5092
rect 21824 5072 21876 5092
rect 21876 5072 21878 5092
rect 21730 4800 21786 4856
rect 22466 4936 22522 4992
rect 21638 3596 21694 3632
rect 21638 3576 21640 3596
rect 21640 3576 21692 3596
rect 21692 3576 21694 3596
rect 21454 3440 21510 3496
rect 21454 3168 21510 3224
rect 21362 2624 21418 2680
rect 22558 4800 22614 4856
rect 22466 4120 22522 4176
rect 22742 4156 22744 4176
rect 22744 4156 22796 4176
rect 22796 4156 22798 4176
rect 22742 4120 22798 4156
rect 21822 2760 21878 2816
rect 21822 2372 21878 2408
rect 21822 2352 21824 2372
rect 21824 2352 21876 2372
rect 21876 2352 21878 2372
rect 22558 2896 22614 2952
rect 23294 4256 23350 4312
rect 24674 21936 24730 21992
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24766 20848 24822 20904
rect 24674 20304 24730 20360
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 25410 26016 25466 26072
rect 25042 23704 25098 23760
rect 25134 23160 25190 23216
rect 25226 22480 25282 22536
rect 24766 19080 24822 19136
rect 24582 18828 24638 18864
rect 24582 18808 24584 18828
rect 24584 18808 24636 18828
rect 24636 18808 24638 18828
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24674 18264 24730 18320
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24950 18128 25006 18184
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24674 16224 24730 16280
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24122 12960 24178 13016
rect 25134 17448 25190 17504
rect 25042 16632 25098 16688
rect 25134 13776 25190 13832
rect 24122 12824 24178 12880
rect 24030 11056 24086 11112
rect 23938 10920 23994 10976
rect 23938 6296 23994 6352
rect 23754 3732 23810 3768
rect 23754 3712 23756 3732
rect 23756 3712 23808 3732
rect 23808 3712 23810 3732
rect 23478 3440 23534 3496
rect 23662 3168 23718 3224
rect 23570 2760 23626 2816
rect 22374 1944 22430 2000
rect 22926 1944 22982 2000
rect 22282 1808 22338 1864
rect 7838 40 7894 96
rect 23018 1672 23074 1728
rect 24674 12300 24730 12336
rect 24674 12280 24676 12300
rect 24676 12280 24728 12300
rect 24728 12280 24730 12300
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 25870 15680 25926 15736
rect 25594 14592 25650 14648
rect 24674 10512 24730 10568
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 25226 10104 25282 10160
rect 24674 8880 24730 8936
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24306 8336 24362 8392
rect 24122 7792 24178 7848
rect 24030 5616 24086 5672
rect 24030 4276 24086 4312
rect 24030 4256 24032 4276
rect 24032 4256 24084 4276
rect 24084 4256 24086 4276
rect 25134 9324 25136 9344
rect 25136 9324 25188 9344
rect 25188 9324 25190 9344
rect 25134 9288 25190 9324
rect 24674 7928 24730 7984
rect 25410 8200 25466 8256
rect 25502 8064 25558 8120
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24674 5344 24730 5400
rect 24674 4936 24730 4992
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24214 3884 24216 3904
rect 24216 3884 24268 3904
rect 24268 3884 24270 3904
rect 24214 3848 24270 3884
rect 24122 2488 24178 2544
rect 25226 5616 25282 5672
rect 25410 4664 25466 4720
rect 25594 4528 25650 4584
rect 25686 3984 25742 4040
rect 26238 3984 26294 4040
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 25410 2796 25412 2816
rect 25412 2796 25464 2816
rect 25464 2796 25466 2816
rect 25410 2760 25466 2796
rect 25594 2644 25650 2680
rect 25594 2624 25596 2644
rect 25596 2624 25648 2644
rect 25648 2624 25650 2644
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 24398 856 24454 912
rect 21638 176 21694 232
rect 24766 1400 24822 1456
rect 25594 1264 25650 1320
rect 24674 312 24730 368
rect 27526 2760 27582 2816
rect 24858 40 24914 96
<< metal3 >>
rect 23657 27706 23723 27709
rect 27520 27706 28000 27736
rect 23657 27704 28000 27706
rect 23657 27648 23662 27704
rect 23718 27648 28000 27704
rect 23657 27646 28000 27648
rect 23657 27643 23723 27646
rect 27520 27616 28000 27646
rect 23473 27162 23539 27165
rect 27520 27162 28000 27192
rect 23473 27160 28000 27162
rect 23473 27104 23478 27160
rect 23534 27104 28000 27160
rect 23473 27102 28000 27104
rect 23473 27099 23539 27102
rect 27520 27072 28000 27102
rect 24945 26618 25011 26621
rect 27520 26618 28000 26648
rect 24945 26616 28000 26618
rect 24945 26560 24950 26616
rect 25006 26560 28000 26616
rect 24945 26558 28000 26560
rect 24945 26555 25011 26558
rect 27520 26528 28000 26558
rect 25405 26074 25471 26077
rect 27520 26074 28000 26104
rect 25405 26072 28000 26074
rect 25405 26016 25410 26072
rect 25466 26016 28000 26072
rect 25405 26014 28000 26016
rect 25405 26011 25471 26014
rect 27520 25984 28000 26014
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 24669 25394 24735 25397
rect 27520 25394 28000 25424
rect 24669 25392 28000 25394
rect 24669 25336 24674 25392
rect 24730 25336 28000 25392
rect 24669 25334 28000 25336
rect 24669 25331 24735 25334
rect 27520 25304 28000 25334
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 24117 24850 24183 24853
rect 27520 24850 28000 24880
rect 24117 24848 28000 24850
rect 24117 24792 24122 24848
rect 24178 24792 28000 24848
rect 24117 24790 28000 24792
rect 24117 24787 24183 24790
rect 27520 24760 28000 24790
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 27520 24306 28000 24336
rect 24902 24246 28000 24306
rect 3509 24170 3575 24173
rect 24761 24170 24827 24173
rect 3509 24168 24827 24170
rect 3509 24112 3514 24168
rect 3570 24112 24766 24168
rect 24822 24112 24827 24168
rect 3509 24110 24827 24112
rect 3509 24107 3575 24110
rect 24761 24107 24827 24110
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 24761 23898 24827 23901
rect 24902 23898 24962 24246
rect 27520 24216 28000 24246
rect 24761 23896 24962 23898
rect 24761 23840 24766 23896
rect 24822 23840 24962 23896
rect 24761 23838 24962 23840
rect 24761 23835 24827 23838
rect 12801 23762 12867 23765
rect 24393 23762 24459 23765
rect 12801 23760 24459 23762
rect 12801 23704 12806 23760
rect 12862 23704 24398 23760
rect 24454 23704 24459 23760
rect 12801 23702 24459 23704
rect 12801 23699 12867 23702
rect 24393 23699 24459 23702
rect 25037 23762 25103 23765
rect 27520 23762 28000 23792
rect 25037 23760 28000 23762
rect 25037 23704 25042 23760
rect 25098 23704 28000 23760
rect 25037 23702 28000 23704
rect 25037 23699 25103 23702
rect 27520 23672 28000 23702
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 25129 23218 25195 23221
rect 27520 23218 28000 23248
rect 25129 23216 28000 23218
rect 25129 23160 25134 23216
rect 25190 23160 28000 23216
rect 25129 23158 28000 23160
rect 25129 23155 25195 23158
rect 27520 23128 28000 23158
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 14549 22674 14615 22677
rect 24577 22674 24643 22677
rect 14549 22672 24643 22674
rect 14549 22616 14554 22672
rect 14610 22616 24582 22672
rect 24638 22616 24643 22672
rect 14549 22614 24643 22616
rect 14549 22611 14615 22614
rect 24577 22611 24643 22614
rect 25221 22538 25287 22541
rect 27520 22538 28000 22568
rect 25221 22536 28000 22538
rect 25221 22480 25226 22536
rect 25282 22480 28000 22536
rect 25221 22478 28000 22480
rect 25221 22475 25287 22478
rect 27520 22448 28000 22478
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 24669 21994 24735 21997
rect 27520 21994 28000 22024
rect 24669 21992 28000 21994
rect 24669 21936 24674 21992
rect 24730 21936 28000 21992
rect 24669 21934 28000 21936
rect 24669 21931 24735 21934
rect 27520 21904 28000 21934
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 16849 21586 16915 21589
rect 16849 21584 24962 21586
rect 16849 21528 16854 21584
rect 16910 21528 24962 21584
rect 16849 21526 24962 21528
rect 16849 21523 16915 21526
rect 10041 21450 10107 21453
rect 23473 21450 23539 21453
rect 10041 21448 23539 21450
rect 10041 21392 10046 21448
rect 10102 21392 23478 21448
rect 23534 21392 23539 21448
rect 10041 21390 23539 21392
rect 24902 21450 24962 21526
rect 27520 21450 28000 21480
rect 24902 21390 28000 21450
rect 10041 21387 10107 21390
rect 23473 21387 23539 21390
rect 27520 21360 28000 21390
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 24761 20906 24827 20909
rect 27520 20906 28000 20936
rect 24761 20904 28000 20906
rect 24761 20848 24766 20904
rect 24822 20848 28000 20904
rect 24761 20846 28000 20848
rect 24761 20843 24827 20846
rect 27520 20816 28000 20846
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 10777 20498 10843 20501
rect 17125 20498 17191 20501
rect 10777 20496 17191 20498
rect 10777 20440 10782 20496
rect 10838 20440 17130 20496
rect 17186 20440 17191 20496
rect 10777 20438 17191 20440
rect 10777 20435 10843 20438
rect 17125 20435 17191 20438
rect 24669 20362 24735 20365
rect 27520 20362 28000 20392
rect 24669 20360 28000 20362
rect 24669 20304 24674 20360
rect 24730 20304 28000 20360
rect 24669 20302 28000 20304
rect 24669 20299 24735 20302
rect 27520 20272 28000 20302
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 18689 19954 18755 19957
rect 23841 19954 23907 19957
rect 18689 19952 23907 19954
rect 18689 19896 18694 19952
rect 18750 19896 23846 19952
rect 23902 19896 23907 19952
rect 18689 19894 23907 19896
rect 18689 19891 18755 19894
rect 23841 19891 23907 19894
rect 27520 19682 28000 19712
rect 24902 19622 28000 19682
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 14825 19410 14891 19413
rect 24902 19410 24962 19622
rect 27520 19592 28000 19622
rect 14825 19408 24962 19410
rect 14825 19352 14830 19408
rect 14886 19352 24962 19408
rect 14825 19350 24962 19352
rect 14825 19347 14891 19350
rect 24761 19138 24827 19141
rect 27520 19138 28000 19168
rect 24761 19136 28000 19138
rect 24761 19080 24766 19136
rect 24822 19080 28000 19136
rect 24761 19078 28000 19080
rect 24761 19075 24827 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 27520 19048 28000 19078
rect 19610 19007 19930 19008
rect 11605 18866 11671 18869
rect 24577 18866 24643 18869
rect 11605 18864 24643 18866
rect 11605 18808 11610 18864
rect 11666 18808 24582 18864
rect 24638 18808 24643 18864
rect 11605 18806 24643 18808
rect 11605 18803 11671 18806
rect 24577 18803 24643 18806
rect 27520 18594 28000 18624
rect 24672 18534 28000 18594
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 24672 18325 24732 18534
rect 27520 18504 28000 18534
rect 24669 18320 24735 18325
rect 24669 18264 24674 18320
rect 24730 18264 24735 18320
rect 24669 18259 24735 18264
rect 13813 18186 13879 18189
rect 24945 18186 25011 18189
rect 13813 18184 25011 18186
rect 13813 18128 13818 18184
rect 13874 18128 24950 18184
rect 25006 18128 25011 18184
rect 13813 18126 25011 18128
rect 13813 18123 13879 18126
rect 24945 18123 25011 18126
rect 27520 18050 28000 18080
rect 23430 17990 28000 18050
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 22921 17914 22987 17917
rect 23430 17914 23490 17990
rect 27520 17960 28000 17990
rect 22921 17912 23490 17914
rect 22921 17856 22926 17912
rect 22982 17856 23490 17912
rect 22921 17854 23490 17856
rect 22921 17851 22987 17854
rect 19149 17778 19215 17781
rect 23473 17778 23539 17781
rect 19149 17776 23539 17778
rect 19149 17720 19154 17776
rect 19210 17720 23478 17776
rect 23534 17720 23539 17776
rect 19149 17718 23539 17720
rect 19149 17715 19215 17718
rect 23473 17715 23539 17718
rect 17125 17642 17191 17645
rect 23657 17642 23723 17645
rect 17125 17640 23723 17642
rect 17125 17584 17130 17640
rect 17186 17584 23662 17640
rect 23718 17584 23723 17640
rect 17125 17582 23723 17584
rect 17125 17579 17191 17582
rect 23657 17579 23723 17582
rect 25129 17506 25195 17509
rect 27520 17506 28000 17536
rect 25129 17504 28000 17506
rect 25129 17448 25134 17504
rect 25190 17448 28000 17504
rect 25129 17446 28000 17448
rect 25129 17443 25195 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 27520 17416 28000 17446
rect 24277 17375 24597 17376
rect 11421 17098 11487 17101
rect 13169 17098 13235 17101
rect 11421 17096 13235 17098
rect 11421 17040 11426 17096
rect 11482 17040 13174 17096
rect 13230 17040 13235 17096
rect 11421 17038 13235 17040
rect 11421 17035 11487 17038
rect 13169 17035 13235 17038
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 23473 16826 23539 16829
rect 27520 16826 28000 16856
rect 23473 16824 28000 16826
rect 23473 16768 23478 16824
rect 23534 16768 28000 16824
rect 23473 16766 28000 16768
rect 23473 16763 23539 16766
rect 27520 16736 28000 16766
rect 16573 16690 16639 16693
rect 25037 16690 25103 16693
rect 16573 16688 25103 16690
rect 16573 16632 16578 16688
rect 16634 16632 25042 16688
rect 25098 16632 25103 16688
rect 16573 16630 25103 16632
rect 16573 16627 16639 16630
rect 25037 16627 25103 16630
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 24669 16282 24735 16285
rect 27520 16282 28000 16312
rect 24669 16280 28000 16282
rect 24669 16224 24674 16280
rect 24730 16224 28000 16280
rect 24669 16222 28000 16224
rect 24669 16219 24735 16222
rect 27520 16192 28000 16222
rect 15561 16146 15627 16149
rect 23565 16146 23631 16149
rect 15561 16144 23631 16146
rect 15561 16088 15566 16144
rect 15622 16088 23570 16144
rect 23626 16088 23631 16144
rect 15561 16086 23631 16088
rect 15561 16083 15627 16086
rect 23565 16083 23631 16086
rect 15929 16010 15995 16013
rect 23657 16010 23723 16013
rect 15929 16008 23723 16010
rect 15929 15952 15934 16008
rect 15990 15952 23662 16008
rect 23718 15952 23723 16008
rect 15929 15950 23723 15952
rect 15929 15947 15995 15950
rect 23657 15947 23723 15950
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 25865 15738 25931 15741
rect 27520 15738 28000 15768
rect 25865 15736 28000 15738
rect 25865 15680 25870 15736
rect 25926 15680 28000 15736
rect 25865 15678 28000 15680
rect 25865 15675 25931 15678
rect 27520 15648 28000 15678
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 27520 15194 28000 15224
rect 24672 15134 28000 15194
rect 24117 15058 24183 15061
rect 24672 15058 24732 15134
rect 27520 15104 28000 15134
rect 24117 15056 24732 15058
rect 24117 15000 24122 15056
rect 24178 15000 24732 15056
rect 24117 14998 24732 15000
rect 24117 14995 24183 14998
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 25589 14650 25655 14653
rect 27520 14650 28000 14680
rect 25589 14648 28000 14650
rect 25589 14592 25594 14648
rect 25650 14592 28000 14648
rect 25589 14590 28000 14592
rect 25589 14587 25655 14590
rect 27520 14560 28000 14590
rect 12433 14514 12499 14517
rect 21909 14514 21975 14517
rect 12433 14512 21975 14514
rect 12433 14456 12438 14512
rect 12494 14456 21914 14512
rect 21970 14456 21975 14512
rect 12433 14454 21975 14456
rect 12433 14451 12499 14454
rect 21909 14451 21975 14454
rect 23013 14378 23079 14381
rect 3374 14376 23079 14378
rect 3374 14320 23018 14376
rect 23074 14320 23079 14376
rect 3374 14318 23079 14320
rect 0 14106 480 14136
rect 3374 14106 3434 14318
rect 23013 14315 23079 14318
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 0 14046 3434 14106
rect 0 14016 480 14046
rect 23565 13970 23631 13973
rect 27520 13970 28000 14000
rect 23565 13968 28000 13970
rect 23565 13912 23570 13968
rect 23626 13912 28000 13968
rect 23565 13910 28000 13912
rect 23565 13907 23631 13910
rect 27520 13880 28000 13910
rect 17861 13834 17927 13837
rect 25129 13834 25195 13837
rect 17861 13832 25195 13834
rect 17861 13776 17866 13832
rect 17922 13776 25134 13832
rect 25190 13776 25195 13832
rect 17861 13774 25195 13776
rect 17861 13771 17927 13774
rect 25129 13771 25195 13774
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 23473 13426 23539 13429
rect 27520 13426 28000 13456
rect 23473 13424 28000 13426
rect 23473 13368 23478 13424
rect 23534 13368 28000 13424
rect 23473 13366 28000 13368
rect 23473 13363 23539 13366
rect 27520 13336 28000 13366
rect 16113 13290 16179 13293
rect 23657 13290 23723 13293
rect 16113 13288 23723 13290
rect 16113 13232 16118 13288
rect 16174 13232 23662 13288
rect 23718 13232 23723 13288
rect 16113 13230 23723 13232
rect 16113 13227 16179 13230
rect 23657 13227 23723 13230
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 21265 13018 21331 13021
rect 24117 13018 24183 13021
rect 21265 13016 24183 13018
rect 21265 12960 21270 13016
rect 21326 12960 24122 13016
rect 24178 12960 24183 13016
rect 21265 12958 24183 12960
rect 21265 12955 21331 12958
rect 24117 12955 24183 12958
rect 17769 12882 17835 12885
rect 22645 12882 22711 12885
rect 17769 12880 22711 12882
rect 17769 12824 17774 12880
rect 17830 12824 22650 12880
rect 22706 12824 22711 12880
rect 17769 12822 22711 12824
rect 17769 12819 17835 12822
rect 22645 12819 22711 12822
rect 24117 12882 24183 12885
rect 27520 12882 28000 12912
rect 24117 12880 28000 12882
rect 24117 12824 24122 12880
rect 24178 12824 28000 12880
rect 24117 12822 28000 12824
rect 24117 12819 24183 12822
rect 27520 12792 28000 12822
rect 4153 12746 4219 12749
rect 18781 12746 18847 12749
rect 4153 12744 18847 12746
rect 4153 12688 4158 12744
rect 4214 12688 18786 12744
rect 18842 12688 18847 12744
rect 4153 12686 18847 12688
rect 4153 12683 4219 12686
rect 18781 12683 18847 12686
rect 19057 12610 19123 12613
rect 19333 12610 19399 12613
rect 19057 12608 19399 12610
rect 19057 12552 19062 12608
rect 19118 12552 19338 12608
rect 19394 12552 19399 12608
rect 19057 12550 19399 12552
rect 19057 12547 19123 12550
rect 19333 12547 19399 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 16389 12338 16455 12341
rect 24669 12338 24735 12341
rect 27520 12338 28000 12368
rect 16389 12336 24735 12338
rect 16389 12280 16394 12336
rect 16450 12280 24674 12336
rect 24730 12280 24735 12336
rect 16389 12278 24735 12280
rect 16389 12275 16455 12278
rect 24669 12275 24735 12278
rect 24902 12278 28000 12338
rect 23105 12202 23171 12205
rect 24902 12202 24962 12278
rect 27520 12248 28000 12278
rect 23105 12200 24962 12202
rect 23105 12144 23110 12200
rect 23166 12144 24962 12200
rect 23105 12142 24962 12144
rect 23105 12139 23171 12142
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 23473 11794 23539 11797
rect 27520 11794 28000 11824
rect 23473 11792 28000 11794
rect 23473 11736 23478 11792
rect 23534 11736 28000 11792
rect 23473 11734 28000 11736
rect 23473 11731 23539 11734
rect 27520 11704 28000 11734
rect 12893 11522 12959 11525
rect 17401 11522 17467 11525
rect 12893 11520 17467 11522
rect 12893 11464 12898 11520
rect 12954 11464 17406 11520
rect 17462 11464 17467 11520
rect 12893 11462 17467 11464
rect 12893 11459 12959 11462
rect 17401 11459 17467 11462
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 16021 11250 16087 11253
rect 20897 11250 20963 11253
rect 16021 11248 20963 11250
rect 16021 11192 16026 11248
rect 16082 11192 20902 11248
rect 20958 11192 20963 11248
rect 16021 11190 20963 11192
rect 16021 11187 16087 11190
rect 20897 11187 20963 11190
rect 21173 11250 21239 11253
rect 22921 11250 22987 11253
rect 21173 11248 22987 11250
rect 21173 11192 21178 11248
rect 21234 11192 22926 11248
rect 22982 11192 22987 11248
rect 21173 11190 22987 11192
rect 21173 11187 21239 11190
rect 22921 11187 22987 11190
rect 8937 11114 9003 11117
rect 12433 11114 12499 11117
rect 8937 11112 12499 11114
rect 8937 11056 8942 11112
rect 8998 11056 12438 11112
rect 12494 11056 12499 11112
rect 8937 11054 12499 11056
rect 8937 11051 9003 11054
rect 12433 11051 12499 11054
rect 14457 11114 14523 11117
rect 17861 11114 17927 11117
rect 14457 11112 17927 11114
rect 14457 11056 14462 11112
rect 14518 11056 17866 11112
rect 17922 11056 17927 11112
rect 14457 11054 17927 11056
rect 14457 11051 14523 11054
rect 17861 11051 17927 11054
rect 24025 11114 24091 11117
rect 27520 11114 28000 11144
rect 24025 11112 28000 11114
rect 24025 11056 24030 11112
rect 24086 11056 28000 11112
rect 24025 11054 28000 11056
rect 24025 11051 24091 11054
rect 27520 11024 28000 11054
rect 18505 10978 18571 10981
rect 23933 10978 23999 10981
rect 18505 10976 23999 10978
rect 18505 10920 18510 10976
rect 18566 10920 23938 10976
rect 23994 10920 23999 10976
rect 18505 10918 23999 10920
rect 18505 10915 18571 10918
rect 23933 10915 23999 10918
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 13077 10570 13143 10573
rect 20253 10570 20319 10573
rect 13077 10568 20319 10570
rect 13077 10512 13082 10568
rect 13138 10512 20258 10568
rect 20314 10512 20319 10568
rect 13077 10510 20319 10512
rect 13077 10507 13143 10510
rect 20253 10507 20319 10510
rect 24669 10570 24735 10573
rect 27520 10570 28000 10600
rect 24669 10568 28000 10570
rect 24669 10512 24674 10568
rect 24730 10512 28000 10568
rect 24669 10510 28000 10512
rect 24669 10507 24735 10510
rect 27520 10480 28000 10510
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 14181 10162 14247 10165
rect 25221 10162 25287 10165
rect 14181 10160 25287 10162
rect 14181 10104 14186 10160
rect 14242 10104 25226 10160
rect 25282 10104 25287 10160
rect 14181 10102 25287 10104
rect 14181 10099 14247 10102
rect 25221 10099 25287 10102
rect 14089 10026 14155 10029
rect 15469 10026 15535 10029
rect 14089 10024 15535 10026
rect 14089 9968 14094 10024
rect 14150 9968 15474 10024
rect 15530 9968 15535 10024
rect 14089 9966 15535 9968
rect 14089 9963 14155 9966
rect 15469 9963 15535 9966
rect 23473 10026 23539 10029
rect 27520 10026 28000 10056
rect 23473 10024 28000 10026
rect 23473 9968 23478 10024
rect 23534 9968 28000 10024
rect 23473 9966 28000 9968
rect 23473 9963 23539 9966
rect 27520 9936 28000 9966
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 16481 9754 16547 9757
rect 16300 9752 16547 9754
rect 16300 9696 16486 9752
rect 16542 9696 16547 9752
rect 16300 9694 16547 9696
rect 16300 9618 16360 9694
rect 16481 9691 16547 9694
rect 20161 9754 20227 9757
rect 23289 9754 23355 9757
rect 20161 9752 23355 9754
rect 20161 9696 20166 9752
rect 20222 9696 23294 9752
rect 23350 9696 23355 9752
rect 20161 9694 23355 9696
rect 20161 9691 20227 9694
rect 23289 9691 23355 9694
rect 16849 9618 16915 9621
rect 16300 9616 16915 9618
rect 16300 9560 16854 9616
rect 16910 9560 16915 9616
rect 16300 9558 16915 9560
rect 16849 9555 16915 9558
rect 17861 9618 17927 9621
rect 19057 9618 19123 9621
rect 20713 9618 20779 9621
rect 17861 9616 20779 9618
rect 17861 9560 17866 9616
rect 17922 9560 19062 9616
rect 19118 9560 20718 9616
rect 20774 9560 20779 9616
rect 17861 9558 20779 9560
rect 17861 9555 17927 9558
rect 19057 9555 19123 9558
rect 20713 9555 20779 9558
rect 6269 9482 6335 9485
rect 27520 9482 28000 9512
rect 6269 9480 28000 9482
rect 6269 9424 6274 9480
rect 6330 9424 28000 9480
rect 6269 9422 28000 9424
rect 6269 9419 6335 9422
rect 27520 9392 28000 9422
rect 23013 9346 23079 9349
rect 25129 9346 25195 9349
rect 23013 9344 25195 9346
rect 23013 9288 23018 9344
rect 23074 9288 25134 9344
rect 25190 9288 25195 9344
rect 23013 9286 25195 9288
rect 23013 9283 23079 9286
rect 25129 9283 25195 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 12065 9074 12131 9077
rect 21909 9074 21975 9077
rect 12065 9072 21975 9074
rect 12065 9016 12070 9072
rect 12126 9016 21914 9072
rect 21970 9016 21975 9072
rect 12065 9014 21975 9016
rect 12065 9011 12131 9014
rect 21909 9011 21975 9014
rect 15745 8938 15811 8941
rect 23749 8938 23815 8941
rect 15745 8936 23815 8938
rect 15745 8880 15750 8936
rect 15806 8880 23754 8936
rect 23810 8880 23815 8936
rect 15745 8878 23815 8880
rect 15745 8875 15811 8878
rect 23749 8875 23815 8878
rect 24669 8938 24735 8941
rect 27520 8938 28000 8968
rect 24669 8936 28000 8938
rect 24669 8880 24674 8936
rect 24730 8880 28000 8936
rect 24669 8878 28000 8880
rect 24669 8875 24735 8878
rect 27520 8848 28000 8878
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 21541 8666 21607 8669
rect 23473 8666 23539 8669
rect 21541 8664 23539 8666
rect 21541 8608 21546 8664
rect 21602 8608 23478 8664
rect 23534 8608 23539 8664
rect 21541 8606 23539 8608
rect 21541 8603 21607 8606
rect 23473 8603 23539 8606
rect 4061 8530 4127 8533
rect 16021 8530 16087 8533
rect 4061 8528 16087 8530
rect 4061 8472 4066 8528
rect 4122 8472 16026 8528
rect 16082 8472 16087 8528
rect 4061 8470 16087 8472
rect 4061 8467 4127 8470
rect 16021 8467 16087 8470
rect 17493 8530 17559 8533
rect 22645 8530 22711 8533
rect 17493 8528 22711 8530
rect 17493 8472 17498 8528
rect 17554 8472 22650 8528
rect 22706 8472 22711 8528
rect 17493 8470 22711 8472
rect 17493 8467 17559 8470
rect 22645 8467 22711 8470
rect 8569 8394 8635 8397
rect 13445 8394 13511 8397
rect 8569 8392 13511 8394
rect 8569 8336 8574 8392
rect 8630 8336 13450 8392
rect 13506 8336 13511 8392
rect 8569 8334 13511 8336
rect 8569 8331 8635 8334
rect 13445 8331 13511 8334
rect 16481 8394 16547 8397
rect 18873 8394 18939 8397
rect 16481 8392 18939 8394
rect 16481 8336 16486 8392
rect 16542 8336 18878 8392
rect 18934 8336 18939 8392
rect 16481 8334 18939 8336
rect 16481 8331 16547 8334
rect 18873 8331 18939 8334
rect 21725 8394 21791 8397
rect 24301 8394 24367 8397
rect 21725 8392 24367 8394
rect 21725 8336 21730 8392
rect 21786 8336 24306 8392
rect 24362 8336 24367 8392
rect 21725 8334 24367 8336
rect 21725 8331 21791 8334
rect 24301 8331 24367 8334
rect 10685 8258 10751 8261
rect 15377 8258 15443 8261
rect 17125 8258 17191 8261
rect 10685 8256 15443 8258
rect 10685 8200 10690 8256
rect 10746 8200 15382 8256
rect 15438 8200 15443 8256
rect 10685 8198 15443 8200
rect 10685 8195 10751 8198
rect 15377 8195 15443 8198
rect 15886 8256 17191 8258
rect 15886 8200 17130 8256
rect 17186 8200 17191 8256
rect 15886 8198 17191 8200
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 10777 8122 10843 8125
rect 15886 8122 15946 8198
rect 17125 8195 17191 8198
rect 25405 8258 25471 8261
rect 27520 8258 28000 8288
rect 25405 8256 28000 8258
rect 25405 8200 25410 8256
rect 25466 8200 28000 8256
rect 25405 8198 28000 8200
rect 25405 8195 25471 8198
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 27520 8168 28000 8198
rect 19610 8127 19930 8128
rect 10777 8120 15946 8122
rect 10777 8064 10782 8120
rect 10838 8064 15946 8120
rect 10777 8062 15946 8064
rect 16757 8122 16823 8125
rect 19425 8122 19491 8125
rect 25497 8122 25563 8125
rect 16757 8120 19491 8122
rect 16757 8064 16762 8120
rect 16818 8064 19430 8120
rect 19486 8064 19491 8120
rect 16757 8062 19491 8064
rect 10777 8059 10843 8062
rect 16757 8059 16823 8062
rect 19425 8059 19491 8062
rect 20118 8120 25563 8122
rect 20118 8064 25502 8120
rect 25558 8064 25563 8120
rect 20118 8062 25563 8064
rect 6729 7986 6795 7989
rect 11145 7986 11211 7989
rect 6729 7984 11211 7986
rect 6729 7928 6734 7984
rect 6790 7928 11150 7984
rect 11206 7928 11211 7984
rect 6729 7926 11211 7928
rect 6729 7923 6795 7926
rect 11145 7923 11211 7926
rect 17401 7986 17467 7989
rect 20118 7986 20178 8062
rect 25497 8059 25563 8062
rect 17401 7984 20178 7986
rect 17401 7928 17406 7984
rect 17462 7928 20178 7984
rect 17401 7926 20178 7928
rect 20897 7986 20963 7989
rect 24669 7986 24735 7989
rect 20897 7984 24735 7986
rect 20897 7928 20902 7984
rect 20958 7928 24674 7984
rect 24730 7928 24735 7984
rect 20897 7926 24735 7928
rect 17401 7923 17467 7926
rect 20897 7923 20963 7926
rect 24669 7923 24735 7926
rect 16297 7850 16363 7853
rect 20621 7850 20687 7853
rect 21909 7850 21975 7853
rect 24117 7850 24183 7853
rect 16297 7848 20687 7850
rect 16297 7792 16302 7848
rect 16358 7792 20626 7848
rect 20682 7792 20687 7848
rect 16297 7790 20687 7792
rect 16297 7787 16363 7790
rect 20621 7787 20687 7790
rect 20854 7848 24183 7850
rect 20854 7792 21914 7848
rect 21970 7792 24122 7848
rect 24178 7792 24183 7848
rect 20854 7790 24183 7792
rect 6085 7714 6151 7717
rect 10501 7714 10567 7717
rect 6085 7712 10567 7714
rect 6085 7656 6090 7712
rect 6146 7656 10506 7712
rect 10562 7656 10567 7712
rect 6085 7654 10567 7656
rect 6085 7651 6151 7654
rect 10501 7651 10567 7654
rect 10685 7714 10751 7717
rect 14549 7714 14615 7717
rect 10685 7712 14615 7714
rect 10685 7656 10690 7712
rect 10746 7656 14554 7712
rect 14610 7656 14615 7712
rect 10685 7654 14615 7656
rect 10685 7651 10751 7654
rect 14549 7651 14615 7654
rect 16389 7714 16455 7717
rect 17953 7714 18019 7717
rect 16389 7712 18019 7714
rect 16389 7656 16394 7712
rect 16450 7656 17958 7712
rect 18014 7656 18019 7712
rect 16389 7654 18019 7656
rect 16389 7651 16455 7654
rect 17953 7651 18019 7654
rect 18321 7714 18387 7717
rect 20854 7714 20914 7790
rect 21909 7787 21975 7790
rect 24117 7787 24183 7790
rect 27520 7714 28000 7744
rect 18321 7712 20914 7714
rect 18321 7656 18326 7712
rect 18382 7656 20914 7712
rect 18321 7654 20914 7656
rect 21958 7654 23536 7714
rect 18321 7651 18387 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 7005 7578 7071 7581
rect 10869 7578 10935 7581
rect 7005 7576 10935 7578
rect 7005 7520 7010 7576
rect 7066 7520 10874 7576
rect 10930 7520 10935 7576
rect 7005 7518 10935 7520
rect 7005 7515 7071 7518
rect 10869 7515 10935 7518
rect 11145 7578 11211 7581
rect 14273 7578 14339 7581
rect 11145 7576 14339 7578
rect 11145 7520 11150 7576
rect 11206 7520 14278 7576
rect 14334 7520 14339 7576
rect 11145 7518 14339 7520
rect 11145 7515 11211 7518
rect 14273 7515 14339 7518
rect 17217 7578 17283 7581
rect 21958 7578 22018 7654
rect 17217 7576 22018 7578
rect 17217 7520 17222 7576
rect 17278 7520 22018 7576
rect 17217 7518 22018 7520
rect 17217 7515 17283 7518
rect 1577 7442 1643 7445
rect 12801 7442 12867 7445
rect 1577 7440 12867 7442
rect 1577 7384 1582 7440
rect 1638 7384 12806 7440
rect 12862 7384 12867 7440
rect 1577 7382 12867 7384
rect 1577 7379 1643 7382
rect 12801 7379 12867 7382
rect 14733 7442 14799 7445
rect 20253 7442 20319 7445
rect 14733 7440 20319 7442
rect 14733 7384 14738 7440
rect 14794 7384 20258 7440
rect 20314 7384 20319 7440
rect 14733 7382 20319 7384
rect 23476 7442 23536 7654
rect 24672 7654 28000 7714
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 24672 7442 24732 7654
rect 27520 7624 28000 7654
rect 23476 7382 24732 7442
rect 14733 7379 14799 7382
rect 20253 7379 20319 7382
rect 8109 7306 8175 7309
rect 10869 7306 10935 7309
rect 22369 7306 22435 7309
rect 8109 7304 10794 7306
rect 8109 7248 8114 7304
rect 8170 7248 10794 7304
rect 8109 7246 10794 7248
rect 8109 7243 8175 7246
rect 10734 7170 10794 7246
rect 10869 7304 22435 7306
rect 10869 7248 10874 7304
rect 10930 7248 22374 7304
rect 22430 7248 22435 7304
rect 10869 7246 22435 7248
rect 10869 7243 10935 7246
rect 22369 7243 22435 7246
rect 17217 7170 17283 7173
rect 10734 7168 17283 7170
rect 10734 7112 17222 7168
rect 17278 7112 17283 7168
rect 10734 7110 17283 7112
rect 17217 7107 17283 7110
rect 17401 7170 17467 7173
rect 18321 7170 18387 7173
rect 27520 7170 28000 7200
rect 17401 7168 18387 7170
rect 17401 7112 17406 7168
rect 17462 7112 18326 7168
rect 18382 7112 18387 7168
rect 17401 7110 18387 7112
rect 17401 7107 17467 7110
rect 18321 7107 18387 7110
rect 20118 7110 28000 7170
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 13445 7034 13511 7037
rect 13813 7034 13879 7037
rect 17033 7034 17099 7037
rect 13445 7032 17099 7034
rect 13445 6976 13450 7032
rect 13506 6976 13818 7032
rect 13874 6976 17038 7032
rect 17094 6976 17099 7032
rect 13445 6974 17099 6976
rect 13445 6971 13511 6974
rect 13813 6971 13879 6974
rect 17033 6971 17099 6974
rect 17174 6974 19442 7034
rect 2221 6898 2287 6901
rect 11789 6898 11855 6901
rect 2221 6896 11855 6898
rect 2221 6840 2226 6896
rect 2282 6840 11794 6896
rect 11850 6840 11855 6896
rect 2221 6838 11855 6840
rect 2221 6835 2287 6838
rect 11789 6835 11855 6838
rect 11973 6898 12039 6901
rect 16205 6898 16271 6901
rect 11973 6896 16271 6898
rect 11973 6840 11978 6896
rect 12034 6840 16210 6896
rect 16266 6840 16271 6896
rect 11973 6838 16271 6840
rect 11973 6835 12039 6838
rect 16205 6835 16271 6838
rect 6361 6762 6427 6765
rect 17174 6762 17234 6974
rect 19382 6898 19442 6974
rect 20118 6898 20178 7110
rect 27520 7080 28000 7110
rect 20253 7034 20319 7037
rect 23473 7034 23539 7037
rect 20253 7032 23539 7034
rect 20253 6976 20258 7032
rect 20314 6976 23478 7032
rect 23534 6976 23539 7032
rect 20253 6974 23539 6976
rect 20253 6971 20319 6974
rect 23473 6971 23539 6974
rect 19382 6838 20178 6898
rect 6361 6760 17234 6762
rect 6361 6704 6366 6760
rect 6422 6704 17234 6760
rect 6361 6702 17234 6704
rect 22142 6702 24732 6762
rect 6361 6699 6427 6702
rect 22142 6660 22202 6702
rect 15745 6626 15811 6629
rect 21958 6626 22202 6660
rect 15745 6624 22202 6626
rect 15745 6568 15750 6624
rect 15806 6600 22202 6624
rect 24672 6626 24732 6702
rect 27520 6626 28000 6656
rect 15806 6568 22018 6600
rect 15745 6566 22018 6568
rect 24672 6566 28000 6626
rect 15745 6563 15811 6566
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 27520 6536 28000 6566
rect 24277 6495 24597 6496
rect 14457 6490 14523 6493
rect 6134 6488 14523 6490
rect 6134 6432 14462 6488
rect 14518 6432 14523 6488
rect 6134 6430 14523 6432
rect 4153 6354 4219 6357
rect 6134 6354 6194 6430
rect 14457 6427 14523 6430
rect 14733 6354 14799 6357
rect 4153 6352 6194 6354
rect 4153 6296 4158 6352
rect 4214 6296 6194 6352
rect 4153 6294 6194 6296
rect 7606 6352 14799 6354
rect 7606 6296 14738 6352
rect 14794 6296 14799 6352
rect 7606 6294 14799 6296
rect 4153 6291 4219 6294
rect 289 6218 355 6221
rect 7606 6218 7666 6294
rect 14733 6291 14799 6294
rect 17217 6354 17283 6357
rect 23933 6354 23999 6357
rect 17217 6352 23999 6354
rect 17217 6296 17222 6352
rect 17278 6296 23938 6352
rect 23994 6296 23999 6352
rect 17217 6294 23999 6296
rect 17217 6291 17283 6294
rect 23933 6291 23999 6294
rect 289 6216 7666 6218
rect 289 6160 294 6216
rect 350 6160 7666 6216
rect 289 6158 7666 6160
rect 8753 6218 8819 6221
rect 8753 6216 22018 6218
rect 8753 6160 8758 6216
rect 8814 6160 22018 6216
rect 8753 6158 22018 6160
rect 289 6155 355 6158
rect 8753 6155 8819 6158
rect 21958 6116 22018 6158
rect 21958 6082 22202 6116
rect 27520 6082 28000 6112
rect 21958 6056 28000 6082
rect 22142 6022 28000 6056
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 27520 5992 28000 6022
rect 19610 5951 19930 5952
rect 8661 5810 8727 5813
rect 17217 5810 17283 5813
rect 8661 5808 17283 5810
rect 8661 5752 8666 5808
rect 8722 5752 17222 5808
rect 17278 5752 17283 5808
rect 8661 5750 17283 5752
rect 8661 5747 8727 5750
rect 17217 5747 17283 5750
rect 19977 5810 20043 5813
rect 22645 5810 22711 5813
rect 19977 5808 22711 5810
rect 19977 5752 19982 5808
rect 20038 5752 22650 5808
rect 22706 5752 22711 5808
rect 19977 5750 22711 5752
rect 19977 5747 20043 5750
rect 22645 5747 22711 5750
rect 5993 5674 6059 5677
rect 20069 5674 20135 5677
rect 5993 5672 15946 5674
rect 5993 5616 5998 5672
rect 6054 5616 15946 5672
rect 5993 5614 15946 5616
rect 5993 5611 6059 5614
rect 15886 5538 15946 5614
rect 17174 5672 20135 5674
rect 17174 5616 20074 5672
rect 20130 5616 20135 5672
rect 17174 5614 20135 5616
rect 17174 5538 17234 5614
rect 20069 5611 20135 5614
rect 24025 5674 24091 5677
rect 25221 5674 25287 5677
rect 24025 5672 25287 5674
rect 24025 5616 24030 5672
rect 24086 5616 25226 5672
rect 25282 5616 25287 5672
rect 24025 5614 25287 5616
rect 24025 5611 24091 5614
rect 25221 5611 25287 5614
rect 15886 5478 17234 5538
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 10225 5402 10291 5405
rect 14641 5402 14707 5405
rect 10225 5400 14707 5402
rect 10225 5344 10230 5400
rect 10286 5344 14646 5400
rect 14702 5344 14707 5400
rect 10225 5342 14707 5344
rect 10225 5339 10291 5342
rect 14641 5339 14707 5342
rect 18965 5402 19031 5405
rect 21725 5402 21791 5405
rect 18965 5400 21791 5402
rect 18965 5344 18970 5400
rect 19026 5344 21730 5400
rect 21786 5344 21791 5400
rect 18965 5342 21791 5344
rect 18965 5339 19031 5342
rect 21725 5339 21791 5342
rect 24669 5402 24735 5405
rect 27520 5402 28000 5432
rect 24669 5400 28000 5402
rect 24669 5344 24674 5400
rect 24730 5344 28000 5400
rect 24669 5342 28000 5344
rect 24669 5339 24735 5342
rect 27520 5312 28000 5342
rect 6913 5266 6979 5269
rect 6913 5264 24916 5266
rect 6913 5208 6918 5264
rect 6974 5208 24916 5264
rect 6913 5206 24916 5208
rect 6913 5203 6979 5206
rect 12709 5130 12775 5133
rect 17677 5130 17743 5133
rect 12709 5128 17743 5130
rect 12709 5072 12714 5128
rect 12770 5072 17682 5128
rect 17738 5072 17743 5128
rect 12709 5070 17743 5072
rect 12709 5067 12775 5070
rect 17677 5067 17743 5070
rect 18137 5130 18203 5133
rect 21817 5130 21883 5133
rect 18137 5128 21883 5130
rect 18137 5072 18142 5128
rect 18198 5072 21822 5128
rect 21878 5072 21883 5128
rect 18137 5070 21883 5072
rect 18137 5067 18203 5070
rect 21817 5067 21883 5070
rect 2865 4994 2931 4997
rect 9765 4994 9831 4997
rect 2865 4992 9831 4994
rect 2865 4936 2870 4992
rect 2926 4936 9770 4992
rect 9826 4936 9831 4992
rect 2865 4934 9831 4936
rect 2865 4931 2931 4934
rect 9765 4931 9831 4934
rect 13537 4994 13603 4997
rect 15561 4994 15627 4997
rect 17125 4994 17191 4997
rect 13537 4992 17191 4994
rect 13537 4936 13542 4992
rect 13598 4936 15566 4992
rect 15622 4936 17130 4992
rect 17186 4936 17191 4992
rect 13537 4934 17191 4936
rect 13537 4931 13603 4934
rect 15561 4931 15627 4934
rect 17125 4931 17191 4934
rect 22461 4994 22527 4997
rect 24669 4994 24735 4997
rect 22461 4992 24735 4994
rect 22461 4936 22466 4992
rect 22522 4936 24674 4992
rect 24730 4936 24735 4992
rect 22461 4934 24735 4936
rect 22461 4931 22527 4934
rect 24669 4931 24735 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 10869 4858 10935 4861
rect 21725 4858 21791 4861
rect 22553 4858 22619 4861
rect 10869 4856 17234 4858
rect 10869 4800 10874 4856
rect 10930 4800 17234 4856
rect 10869 4798 17234 4800
rect 10869 4795 10935 4798
rect 10501 4722 10567 4725
rect 12433 4722 12499 4725
rect 10501 4720 12499 4722
rect 10501 4664 10506 4720
rect 10562 4664 12438 4720
rect 12494 4664 12499 4720
rect 10501 4662 12499 4664
rect 10501 4659 10567 4662
rect 12433 4659 12499 4662
rect 14733 4722 14799 4725
rect 16941 4722 17007 4725
rect 14733 4720 17007 4722
rect 14733 4664 14738 4720
rect 14794 4664 16946 4720
rect 17002 4664 17007 4720
rect 14733 4662 17007 4664
rect 14733 4659 14799 4662
rect 16941 4659 17007 4662
rect 9213 4586 9279 4589
rect 15377 4586 15443 4589
rect 9213 4584 15443 4586
rect 9213 4528 9218 4584
rect 9274 4528 15382 4584
rect 15438 4528 15443 4584
rect 9213 4526 15443 4528
rect 17174 4586 17234 4798
rect 21725 4856 22619 4858
rect 21725 4800 21730 4856
rect 21786 4800 22558 4856
rect 22614 4800 22619 4856
rect 21725 4798 22619 4800
rect 24856 4858 24916 5206
rect 27520 4858 28000 4888
rect 24856 4798 28000 4858
rect 21725 4795 21791 4798
rect 22553 4795 22619 4798
rect 27520 4768 28000 4798
rect 18413 4722 18479 4725
rect 25405 4722 25471 4725
rect 18413 4720 25471 4722
rect 18413 4664 18418 4720
rect 18474 4664 25410 4720
rect 25466 4664 25471 4720
rect 18413 4662 25471 4664
rect 18413 4659 18479 4662
rect 25405 4659 25471 4662
rect 25589 4586 25655 4589
rect 17174 4584 25655 4586
rect 17174 4528 25594 4584
rect 25650 4528 25655 4584
rect 17174 4526 25655 4528
rect 9213 4523 9279 4526
rect 15377 4523 15443 4526
rect 25589 4523 25655 4526
rect 11053 4450 11119 4453
rect 14733 4450 14799 4453
rect 11053 4448 14799 4450
rect 11053 4392 11058 4448
rect 11114 4392 14738 4448
rect 14794 4392 14799 4448
rect 11053 4390 14799 4392
rect 11053 4387 11119 4390
rect 14733 4387 14799 4390
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 8293 4314 8359 4317
rect 19057 4314 19123 4317
rect 21173 4314 21239 4317
rect 8293 4312 14842 4314
rect 8293 4256 8298 4312
rect 8354 4256 14842 4312
rect 8293 4254 14842 4256
rect 8293 4251 8359 4254
rect 3509 4178 3575 4181
rect 13077 4178 13143 4181
rect 3509 4176 13143 4178
rect 3509 4120 3514 4176
rect 3570 4120 13082 4176
rect 13138 4120 13143 4176
rect 3509 4118 13143 4120
rect 14782 4178 14842 4254
rect 19057 4312 21239 4314
rect 19057 4256 19062 4312
rect 19118 4256 21178 4312
rect 21234 4256 21239 4312
rect 19057 4254 21239 4256
rect 19057 4251 19123 4254
rect 21173 4251 21239 4254
rect 23289 4314 23355 4317
rect 24025 4314 24091 4317
rect 27520 4314 28000 4344
rect 23289 4312 24091 4314
rect 23289 4256 23294 4312
rect 23350 4256 24030 4312
rect 24086 4256 24091 4312
rect 23289 4254 24091 4256
rect 23289 4251 23355 4254
rect 24025 4251 24091 4254
rect 24718 4254 28000 4314
rect 22461 4178 22527 4181
rect 14782 4176 22527 4178
rect 14782 4120 22466 4176
rect 22522 4120 22527 4176
rect 14782 4118 22527 4120
rect 3509 4115 3575 4118
rect 13077 4115 13143 4118
rect 22461 4115 22527 4118
rect 22737 4178 22803 4181
rect 24718 4178 24778 4254
rect 27520 4224 28000 4254
rect 22737 4176 24778 4178
rect 22737 4120 22742 4176
rect 22798 4120 24778 4176
rect 22737 4118 24778 4120
rect 22737 4115 22803 4118
rect 7465 4042 7531 4045
rect 14273 4042 14339 4045
rect 15285 4042 15351 4045
rect 20713 4042 20779 4045
rect 7465 4040 10794 4042
rect 7465 3984 7470 4040
rect 7526 3984 10794 4040
rect 7465 3982 10794 3984
rect 7465 3979 7531 3982
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 10734 3770 10794 3982
rect 14273 4040 15351 4042
rect 14273 3984 14278 4040
rect 14334 3984 15290 4040
rect 15346 3984 15351 4040
rect 14273 3982 15351 3984
rect 14273 3979 14339 3982
rect 15285 3979 15351 3982
rect 19198 4040 20779 4042
rect 19198 3984 20718 4040
rect 20774 3984 20779 4040
rect 19198 3982 20779 3984
rect 11421 3906 11487 3909
rect 19198 3906 19258 3982
rect 20713 3979 20779 3982
rect 25681 4042 25747 4045
rect 26233 4042 26299 4045
rect 25681 4040 26299 4042
rect 25681 3984 25686 4040
rect 25742 3984 26238 4040
rect 26294 3984 26299 4040
rect 25681 3982 26299 3984
rect 25681 3979 25747 3982
rect 26233 3979 26299 3982
rect 11421 3904 19258 3906
rect 11421 3848 11426 3904
rect 11482 3848 19258 3904
rect 11421 3846 19258 3848
rect 20437 3906 20503 3909
rect 24209 3906 24275 3909
rect 20437 3904 24275 3906
rect 20437 3848 20442 3904
rect 20498 3848 24214 3904
rect 24270 3848 24275 3904
rect 20437 3846 24275 3848
rect 11421 3843 11487 3846
rect 20437 3843 20503 3846
rect 24209 3843 24275 3846
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 17585 3770 17651 3773
rect 10734 3768 17651 3770
rect 10734 3712 17590 3768
rect 17646 3712 17651 3768
rect 10734 3710 17651 3712
rect 17585 3707 17651 3710
rect 23749 3770 23815 3773
rect 27520 3770 28000 3800
rect 23749 3768 28000 3770
rect 23749 3712 23754 3768
rect 23810 3712 28000 3768
rect 23749 3710 28000 3712
rect 23749 3707 23815 3710
rect 27520 3680 28000 3710
rect 8661 3634 8727 3637
rect 21633 3634 21699 3637
rect 8661 3632 21699 3634
rect 8661 3576 8666 3632
rect 8722 3576 21638 3632
rect 21694 3576 21699 3632
rect 8661 3574 21699 3576
rect 8661 3571 8727 3574
rect 21633 3571 21699 3574
rect 933 3498 999 3501
rect 4061 3498 4127 3501
rect 933 3496 4127 3498
rect 933 3440 938 3496
rect 994 3440 4066 3496
rect 4122 3440 4127 3496
rect 933 3438 4127 3440
rect 933 3435 999 3438
rect 4061 3435 4127 3438
rect 8569 3498 8635 3501
rect 11513 3498 11579 3501
rect 8569 3496 11579 3498
rect 8569 3440 8574 3496
rect 8630 3440 11518 3496
rect 11574 3440 11579 3496
rect 8569 3438 11579 3440
rect 8569 3435 8635 3438
rect 11513 3435 11579 3438
rect 13537 3498 13603 3501
rect 16113 3498 16179 3501
rect 21449 3498 21515 3501
rect 13537 3496 15394 3498
rect 13537 3440 13542 3496
rect 13598 3440 15394 3496
rect 13537 3438 15394 3440
rect 13537 3435 13603 3438
rect 9581 3362 9647 3365
rect 11053 3362 11119 3365
rect 9581 3360 11119 3362
rect 9581 3304 9586 3360
rect 9642 3304 11058 3360
rect 11114 3304 11119 3360
rect 9581 3302 11119 3304
rect 15334 3362 15394 3438
rect 16113 3496 21515 3498
rect 16113 3440 16118 3496
rect 16174 3440 21454 3496
rect 21510 3440 21515 3496
rect 16113 3438 21515 3440
rect 16113 3435 16179 3438
rect 21449 3435 21515 3438
rect 23473 3498 23539 3501
rect 23473 3496 24778 3498
rect 23473 3440 23478 3496
rect 23534 3440 24778 3496
rect 23473 3438 24778 3440
rect 23473 3435 23539 3438
rect 20437 3362 20503 3365
rect 15334 3360 20503 3362
rect 15334 3304 20442 3360
rect 20498 3304 20503 3360
rect 15334 3302 20503 3304
rect 9581 3299 9647 3302
rect 11053 3299 11119 3302
rect 20437 3299 20503 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 6637 3226 6703 3229
rect 9673 3226 9739 3229
rect 6637 3224 9739 3226
rect 6637 3168 6642 3224
rect 6698 3168 9678 3224
rect 9734 3168 9739 3224
rect 6637 3166 9739 3168
rect 6637 3163 6703 3166
rect 9673 3163 9739 3166
rect 9949 3226 10015 3229
rect 11881 3226 11947 3229
rect 12617 3226 12683 3229
rect 19149 3226 19215 3229
rect 9949 3224 12683 3226
rect 9949 3168 9954 3224
rect 10010 3168 11886 3224
rect 11942 3168 12622 3224
rect 12678 3168 12683 3224
rect 9949 3166 12683 3168
rect 9949 3163 10015 3166
rect 11881 3163 11947 3166
rect 12617 3163 12683 3166
rect 17174 3224 19215 3226
rect 17174 3168 19154 3224
rect 19210 3168 19215 3224
rect 17174 3166 19215 3168
rect 4797 3090 4863 3093
rect 6126 3090 6132 3092
rect 4797 3088 6132 3090
rect 4797 3032 4802 3088
rect 4858 3032 6132 3088
rect 4797 3030 6132 3032
rect 4797 3027 4863 3030
rect 6126 3028 6132 3030
rect 6196 3028 6202 3092
rect 9305 3090 9371 3093
rect 11053 3090 11119 3093
rect 17174 3090 17234 3166
rect 19149 3163 19215 3166
rect 21449 3226 21515 3229
rect 23657 3226 23723 3229
rect 21449 3224 23723 3226
rect 21449 3168 21454 3224
rect 21510 3168 23662 3224
rect 23718 3168 23723 3224
rect 21449 3166 23723 3168
rect 24718 3226 24778 3438
rect 27520 3226 28000 3256
rect 24718 3166 28000 3226
rect 21449 3163 21515 3166
rect 23657 3163 23723 3166
rect 27520 3136 28000 3166
rect 9305 3088 10978 3090
rect 9305 3032 9310 3088
rect 9366 3032 10978 3088
rect 9305 3030 10978 3032
rect 9305 3027 9371 3030
rect 8477 2954 8543 2957
rect 10685 2954 10751 2957
rect 8477 2952 10751 2954
rect 8477 2896 8482 2952
rect 8538 2896 10690 2952
rect 10746 2896 10751 2952
rect 8477 2894 10751 2896
rect 10918 2954 10978 3030
rect 11053 3088 17234 3090
rect 11053 3032 11058 3088
rect 11114 3032 17234 3088
rect 11053 3030 17234 3032
rect 11053 3027 11119 3030
rect 17350 3028 17356 3092
rect 17420 3090 17426 3092
rect 19241 3090 19307 3093
rect 17420 3088 19307 3090
rect 17420 3032 19246 3088
rect 19302 3032 19307 3088
rect 17420 3030 19307 3032
rect 17420 3028 17426 3030
rect 19241 3027 19307 3030
rect 19149 2954 19215 2957
rect 22553 2954 22619 2957
rect 10918 2952 22619 2954
rect 10918 2896 19154 2952
rect 19210 2896 22558 2952
rect 22614 2896 22619 2952
rect 10918 2894 22619 2896
rect 8477 2891 8543 2894
rect 10685 2891 10751 2894
rect 19149 2891 19215 2894
rect 22553 2891 22619 2894
rect 11145 2818 11211 2821
rect 12065 2818 12131 2821
rect 13813 2818 13879 2821
rect 11145 2816 13879 2818
rect 11145 2760 11150 2816
rect 11206 2760 12070 2816
rect 12126 2760 13818 2816
rect 13874 2760 13879 2816
rect 11145 2758 13879 2760
rect 11145 2755 11211 2758
rect 12065 2755 12131 2758
rect 13813 2755 13879 2758
rect 15929 2818 15995 2821
rect 19425 2818 19491 2821
rect 15929 2816 19491 2818
rect 15929 2760 15934 2816
rect 15990 2760 19430 2816
rect 19486 2760 19491 2816
rect 15929 2758 19491 2760
rect 15929 2755 15995 2758
rect 19425 2755 19491 2758
rect 21817 2818 21883 2821
rect 23565 2818 23631 2821
rect 21817 2816 23631 2818
rect 21817 2760 21822 2816
rect 21878 2760 23570 2816
rect 23626 2760 23631 2816
rect 21817 2758 23631 2760
rect 21817 2755 21883 2758
rect 23565 2755 23631 2758
rect 25405 2818 25471 2821
rect 27521 2818 27587 2821
rect 25405 2816 27587 2818
rect 25405 2760 25410 2816
rect 25466 2760 27526 2816
rect 27582 2760 27587 2816
rect 25405 2758 27587 2760
rect 25405 2755 25471 2758
rect 27521 2755 27587 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 5625 2682 5691 2685
rect 9949 2682 10015 2685
rect 5625 2680 10015 2682
rect 5625 2624 5630 2680
rect 5686 2624 9954 2680
rect 10010 2624 10015 2680
rect 5625 2622 10015 2624
rect 5625 2619 5691 2622
rect 9949 2619 10015 2622
rect 21357 2682 21423 2685
rect 25589 2682 25655 2685
rect 21357 2680 25655 2682
rect 21357 2624 21362 2680
rect 21418 2624 25594 2680
rect 25650 2624 25655 2680
rect 21357 2622 25655 2624
rect 21357 2619 21423 2622
rect 25589 2619 25655 2622
rect 8109 2546 8175 2549
rect 11237 2546 11303 2549
rect 8109 2544 11303 2546
rect 8109 2488 8114 2544
rect 8170 2488 11242 2544
rect 11298 2488 11303 2544
rect 8109 2486 11303 2488
rect 8109 2483 8175 2486
rect 11237 2483 11303 2486
rect 12893 2546 12959 2549
rect 16849 2546 16915 2549
rect 12893 2544 16915 2546
rect 12893 2488 12898 2544
rect 12954 2488 16854 2544
rect 16910 2488 16915 2544
rect 12893 2486 16915 2488
rect 12893 2483 12959 2486
rect 16849 2483 16915 2486
rect 24117 2546 24183 2549
rect 27520 2546 28000 2576
rect 24117 2544 28000 2546
rect 24117 2488 24122 2544
rect 24178 2488 28000 2544
rect 24117 2486 28000 2488
rect 24117 2483 24183 2486
rect 27520 2456 28000 2486
rect 9397 2410 9463 2413
rect 21817 2410 21883 2413
rect 9397 2408 21883 2410
rect 9397 2352 9402 2408
rect 9458 2352 21822 2408
rect 21878 2352 21883 2408
rect 9397 2350 21883 2352
rect 9397 2347 9463 2350
rect 21817 2347 21883 2350
rect 9213 2274 9279 2277
rect 12249 2274 12315 2277
rect 9213 2272 12315 2274
rect 9213 2216 9218 2272
rect 9274 2216 12254 2272
rect 12310 2216 12315 2272
rect 9213 2214 12315 2216
rect 9213 2211 9279 2214
rect 12249 2211 12315 2214
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 8569 2138 8635 2141
rect 13445 2138 13511 2141
rect 8569 2136 13511 2138
rect 8569 2080 8574 2136
rect 8630 2080 13450 2136
rect 13506 2080 13511 2136
rect 8569 2078 13511 2080
rect 8569 2075 8635 2078
rect 13445 2075 13511 2078
rect 8293 2002 8359 2005
rect 22369 2002 22435 2005
rect 8293 2000 22435 2002
rect 8293 1944 8298 2000
rect 8354 1944 22374 2000
rect 22430 1944 22435 2000
rect 8293 1942 22435 1944
rect 8293 1939 8359 1942
rect 22369 1939 22435 1942
rect 22921 2002 22987 2005
rect 27520 2002 28000 2032
rect 22921 2000 28000 2002
rect 22921 1944 22926 2000
rect 22982 1944 28000 2000
rect 22921 1942 28000 1944
rect 22921 1939 22987 1942
rect 27520 1912 28000 1942
rect 11329 1866 11395 1869
rect 22277 1866 22343 1869
rect 11329 1864 22343 1866
rect 11329 1808 11334 1864
rect 11390 1808 22282 1864
rect 22338 1808 22343 1864
rect 11329 1806 22343 1808
rect 11329 1803 11395 1806
rect 22277 1803 22343 1806
rect 6821 1730 6887 1733
rect 23013 1730 23079 1733
rect 6821 1728 23079 1730
rect 6821 1672 6826 1728
rect 6882 1672 23018 1728
rect 23074 1672 23079 1728
rect 6821 1670 23079 1672
rect 6821 1667 6887 1670
rect 23013 1667 23079 1670
rect 4705 1594 4771 1597
rect 4705 1592 10058 1594
rect 4705 1536 4710 1592
rect 4766 1536 10058 1592
rect 4705 1534 10058 1536
rect 4705 1531 4771 1534
rect 7373 1458 7439 1461
rect 9857 1458 9923 1461
rect 7373 1456 9923 1458
rect 7373 1400 7378 1456
rect 7434 1400 9862 1456
rect 9918 1400 9923 1456
rect 7373 1398 9923 1400
rect 9998 1458 10058 1534
rect 11697 1458 11763 1461
rect 9998 1456 11763 1458
rect 9998 1400 11702 1456
rect 11758 1400 11763 1456
rect 9998 1398 11763 1400
rect 7373 1395 7439 1398
rect 9857 1395 9923 1398
rect 11697 1395 11763 1398
rect 24761 1458 24827 1461
rect 27520 1458 28000 1488
rect 24761 1456 28000 1458
rect 24761 1400 24766 1456
rect 24822 1400 28000 1456
rect 24761 1398 28000 1400
rect 24761 1395 24827 1398
rect 27520 1368 28000 1398
rect 7097 1322 7163 1325
rect 25589 1322 25655 1325
rect 7097 1320 25655 1322
rect 7097 1264 7102 1320
rect 7158 1264 25594 1320
rect 25650 1264 25655 1320
rect 7097 1262 25655 1264
rect 7097 1259 7163 1262
rect 25589 1259 25655 1262
rect 24393 914 24459 917
rect 27520 914 28000 944
rect 24393 912 28000 914
rect 24393 856 24398 912
rect 24454 856 28000 912
rect 24393 854 28000 856
rect 24393 851 24459 854
rect 27520 824 28000 854
rect 24669 370 24735 373
rect 27520 370 28000 400
rect 24669 368 28000 370
rect 24669 312 24674 368
rect 24730 312 28000 368
rect 24669 310 28000 312
rect 24669 307 24735 310
rect 27520 280 28000 310
rect 7189 234 7255 237
rect 21633 234 21699 237
rect 7189 232 21699 234
rect 7189 176 7194 232
rect 7250 176 21638 232
rect 21694 176 21699 232
rect 7189 174 21699 176
rect 7189 171 7255 174
rect 21633 171 21699 174
rect 7833 98 7899 101
rect 24853 98 24919 101
rect 7833 96 24919 98
rect 7833 40 7838 96
rect 7894 40 24858 96
rect 24914 40 24919 96
rect 7833 38 24919 40
rect 7833 35 7899 38
rect 24853 35 24919 38
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 6132 3028 6196 3092
rect 17356 3028 17420 3092
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
<< via4 >>
rect 6046 3092 6282 3178
rect 6046 3028 6132 3092
rect 6132 3028 6196 3092
rect 6196 3028 6282 3092
rect 6046 2942 6282 3028
rect 17270 3092 17506 3178
rect 17270 3028 17356 3092
rect 17356 3028 17420 3092
rect 17420 3028 17506 3092
rect 17270 2942 17506 3028
<< metal5 >>
rect 6004 3178 17548 3220
rect 6004 2942 6046 3178
rect 6282 2942 17270 3178
rect 17506 2942 17548 3178
rect 6004 2900 17548 2942
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1604681595
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1604681595
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _41_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4692 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4600 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1604681595
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_39 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4692 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_47 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5428 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42
timestamp 1604681595
transform 1 0 4968 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0__CLK tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5520 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_53
timestamp 1604681595
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1604681595
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__80__A
timestamp 1604681595
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _80_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5612 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1604681595
transform 1 0 5704 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_62
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1604681595
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58
timestamp 1604681595
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1604681595
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_66
timestamp 1604681595
transform 1 0 7176 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72
timestamp 1604681595
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68
timestamp 1604681595
transform 1 0 7360 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7544 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1604681595
transform 1 0 6992 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1604681595
transform 1 0 6992 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1604681595
transform 1 0 7452 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_77
timestamp 1604681595
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_73
timestamp 1604681595
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8372 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1604681595
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8556 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8096 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_90
timestamp 1604681595
transform 1 0 9384 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89
timestamp 1604681595
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1604681595
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 9568 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_94
timestamp 1604681595
transform 1 0 9752 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9936 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 9936 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 10120 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10120 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_1_114
timestamp 1604681595
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_114
timestamp 1604681595
transform 1 0 11592 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_118
timestamp 1604681595
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__90__A
timestamp 1604681595
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14076 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14260 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1604681595
transform 1 0 14076 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_145
timestamp 1604681595
transform 1 0 14444 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_139
timestamp 1604681595
transform 1 0 13892 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_143
timestamp 1604681595
transform 1 0 14260 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_152
timestamp 1604681595
transform 1 0 15088 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_148
timestamp 1604681595
transform 1 0 14720 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_149
timestamp 1604681595
transform 1 0 14812 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14904 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 15272 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15456 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_1_177
timestamp 1604681595
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_172
timestamp 1604681595
transform 1 0 16928 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_177
timestamp 1604681595
transform 1 0 17388 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_172
timestamp 1604681595
transform 1 0 16928 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17204 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1604681595
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_181
timestamp 1604681595
transform 1 0 17756 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 17572 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18860 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 19688 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 20056 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 18676 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_200
timestamp 1604681595
transform 1 0 19504 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_204
timestamp 1604681595
transform 1 0 19872 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_208
timestamp 1604681595
transform 1 0 20240 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_212
timestamp 1604681595
transform 1 0 20608 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_218
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_213
timestamp 1604681595
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_209
timestamp 1604681595
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 20976 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 20424 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_222
timestamp 1604681595
transform 1 0 21528 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21620 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21804 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 21160 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_1_234
timestamp 1604681595
transform 1 0 22632 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_238
timestamp 1604681595
transform 1 0 23000 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_234
timestamp 1604681595
transform 1 0 22632 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 22816 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_240
timestamp 1604681595
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_244
timestamp 1604681595
transform 1 0 23552 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_258
timestamp 1604681595
transform 1 0 24840 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_254
timestamp 1604681595
transform 1 0 24472 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_258
timestamp 1604681595
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 24656 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_266
timestamp 1604681595
transform 1 0 25576 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_262
timestamp 1604681595
transform 1 0 25208 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 25024 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1604681595
transform 1 0 25208 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1604681595
transform 1 0 25576 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_269
timestamp 1604681595
transform 1 0 25852 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_274
timestamp 1604681595
transform 1 0 26312 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1604681595
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1604681595
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_56
timestamp 1604681595
transform 1 0 6256 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_62
timestamp 1604681595
transform 1 0 6808 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1604681595
transform 1 0 6900 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8004 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 7820 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_67
timestamp 1604681595
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_71
timestamp 1604681595
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_88
timestamp 1604681595
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_84
timestamp 1604681595
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _90_
timestamp 1604681595
transform 1 0 9936 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_100
timestamp 1604681595
transform 1 0 10304 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_104
timestamp 1604681595
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11040 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10856 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_124
timestamp 1604681595
transform 1 0 12512 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13524 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13248 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12880 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_130
timestamp 1604681595
transform 1 0 13064 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_134
timestamp 1604681595
transform 1 0 13432 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_144
timestamp 1604681595
transform 1 0 14352 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15640 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 15456 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_150
timestamp 1604681595
transform 1 0 14904 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_154
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1604681595
transform 1 0 17204 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 16652 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_167
timestamp 1604681595
transform 1 0 16468 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_171
timestamp 1604681595
transform 1 0 16836 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_184
timestamp 1604681595
transform 1 0 18032 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18768 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 18400 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 19780 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_190
timestamp 1604681595
transform 1 0 18584 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_201
timestamp 1604681595
transform 1 0 19596 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_205
timestamp 1604681595
transform 1 0 19964 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 21804 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21252 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 21620 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_211
timestamp 1604681595
transform 1 0 20516 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_221
timestamp 1604681595
transform 1 0 21436 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 24012 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 23644 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_241
timestamp 1604681595
transform 1 0 23276 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_247
timestamp 1604681595
transform 1 0 23828 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_265
timestamp 1604681595
transform 1 0 25484 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_273
timestamp 1604681595
transform 1 0 26220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_276
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1604681595
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1604681595
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1604681595
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1604681595
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_62
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1604681595
transform 1 0 7636 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8740 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1604681595
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1604681595
transform 1 0 8556 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_70
timestamp 1604681595
transform 1 0 7544 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_75
timestamp 1604681595
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_79
timestamp 1604681595
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10304 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_92
timestamp 1604681595
transform 1 0 9568 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_97
timestamp 1604681595
transform 1 0 10028 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11316 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11684 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12052 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_109
timestamp 1604681595
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1604681595
transform 1 0 11500 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_117
timestamp 1604681595
transform 1 0 11868 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_121
timestamp 1604681595
transform 1 0 12236 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_123
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13248 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13064 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 12696 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14260 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_128
timestamp 1604681595
transform 1 0 12880 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_141
timestamp 1604681595
transform 1 0 14076 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_145
timestamp 1604681595
transform 1 0 14444 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15732 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 15180 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14628 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_149
timestamp 1604681595
transform 1 0 14812 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_155
timestamp 1604681595
transform 1 0 15364 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 18216 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_175
timestamp 1604681595
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_179
timestamp 1604681595
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_184
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18768 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 18584 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19780 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20148 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_188
timestamp 1604681595
transform 1 0 18400 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_201
timestamp 1604681595
transform 1 0 19596 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_205
timestamp 1604681595
transform 1 0 19964 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21252 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__82__A
timestamp 1604681595
transform 1 0 20976 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_209
timestamp 1604681595
transform 1 0 20332 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_214
timestamp 1604681595
transform 1 0 20792 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_218
timestamp 1604681595
transform 1 0 21160 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_228
timestamp 1604681595
transform 1 0 22080 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_232
timestamp 1604681595
transform 1 0 22448 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 22264 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 22632 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_236
timestamp 1604681595
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_240
timestamp 1604681595
transform 1 0 23184 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 23000 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_245
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_249
timestamp 1604681595
transform 1 0 24012 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23828 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24380 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__83__A
timestamp 1604681595
transform 1 0 25392 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 24196 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_262
timestamp 1604681595
transform 1 0 25208 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_266
timestamp 1604681595
transform 1 0 25576 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_274
timestamp 1604681595
transform 1 0 26312 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1604681595
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1604681595
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1604681595
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _40_
timestamp 1604681595
transform 1 0 7452 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1604681595
transform 1 0 8464 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 8280 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_68
timestamp 1604681595
transform 1 0 7360 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_72
timestamp 1604681595
transform 1 0 7728 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9844 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_84
timestamp 1604681595
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_88
timestamp 1604681595
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_93
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_104
timestamp 1604681595
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11408 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10856 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11224 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_108
timestamp 1604681595
transform 1 0 11040 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_121
timestamp 1604681595
transform 1 0 12236 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_125
timestamp 1604681595
transform 1 0 12604 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12972 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 12788 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_145
timestamp 1604681595
transform 1 0 14444 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15732 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 15548 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_154
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 18216 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 17848 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_175
timestamp 1604681595
transform 1 0 17204 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_181
timestamp 1604681595
transform 1 0 17756 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_184
timestamp 1604681595
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18400 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 20056 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_204
timestamp 1604681595
transform 1 0 19872 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_208
timestamp 1604681595
transform 1 0 20240 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1604681595
transform 1 0 20976 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 22080 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21528 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21896 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_215
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_220
timestamp 1604681595
transform 1 0 21344 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_224
timestamp 1604681595
transform 1 0 21712 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 23644 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 23460 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23092 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_237
timestamp 1604681595
transform 1 0 22908 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_241
timestamp 1604681595
transform 1 0 23276 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1604681595
transform 1 0 25208 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24656 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 25024 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_254
timestamp 1604681595
transform 1 0 24472 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_258
timestamp 1604681595
transform 1 0 24840 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_266
timestamp 1604681595
transform 1 0 25576 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_274
timestamp 1604681595
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_276
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1604681595
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1604681595
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1604681595
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1604681595
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _42_
timestamp 1604681595
transform 1 0 7912 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 8740 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_77
timestamp 1604681595
transform 1 0 8188 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1604681595
transform 1 0 8924 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9936 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9752 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_88
timestamp 1604681595
transform 1 0 9200 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_92
timestamp 1604681595
transform 1 0 9568 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 12604 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_112
timestamp 1604681595
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_116
timestamp 1604681595
transform 1 0 11776 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 13248 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 13064 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_127
timestamp 1604681595
transform 1 0 12788 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15732 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 15548 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15180 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_148
timestamp 1604681595
transform 1 0 14720 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_152
timestamp 1604681595
transform 1 0 15088 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_155
timestamp 1604681595
transform 1 0 15364 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_176
timestamp 1604681595
transform 1 0 17296 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_172
timestamp 1604681595
transform 1 0 16928 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_168
timestamp 1604681595
transform 1 0 16560 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16744 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_184
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_179
timestamp 1604681595
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18308 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19872 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19688 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 19320 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_196
timestamp 1604681595
transform 1 0 19136 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_200
timestamp 1604681595
transform 1 0 19504 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 21988 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__79__A
timestamp 1604681595
transform 1 0 20884 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 21804 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 21436 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_213
timestamp 1604681595
transform 1 0 20700 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_217
timestamp 1604681595
transform 1 0 21068 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_223
timestamp 1604681595
transform 1 0 21620 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 24012 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 23828 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_236
timestamp 1604681595
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_240
timestamp 1604681595
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_245
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1604681595
transform 1 0 25576 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 25024 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 25392 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_258
timestamp 1604681595
transform 1 0 24840 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_262
timestamp 1604681595
transform 1 0 25208 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_269
timestamp 1604681595
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1604681595
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1604681595
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1604681595
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1604681595
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1604681595
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1604681595
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1604681595
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1604681595
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1604681595
transform 1 0 8556 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1604681595
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_80
timestamp 1604681595
transform 1 0 8464 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_74
timestamp 1604681595
transform 1 0 7912 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_82
timestamp 1604681595
transform 1 0 8648 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_90
timestamp 1604681595
transform 1 0 9384 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_84
timestamp 1604681595
transform 1 0 8832 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8924 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9568 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1604681595
transform 1 0 9108 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_94
timestamp 1604681595
transform 1 0 9752 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_98
timestamp 1604681595
transform 1 0 10120 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 9936 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10212 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10120 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_114
timestamp 1604681595
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_112
timestamp 1604681595
transform 1 0 11408 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_108
timestamp 1604681595
transform 1 0 11040 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11500 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_118
timestamp 1604681595
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_115
timestamp 1604681595
transform 1 0 11684 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12236 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13432 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__88__A
timestamp 1604681595
transform 1 0 14076 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 12880 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_137
timestamp 1604681595
transform 1 0 13708 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_143
timestamp 1604681595
transform 1 0 14260 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_126
timestamp 1604681595
transform 1 0 12696 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_130
timestamp 1604681595
transform 1 0 13064 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_154
timestamp 1604681595
transform 1 0 15272 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_150
timestamp 1604681595
transform 1 0 14904 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_154
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1604681595
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 15088 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_162
timestamp 1604681595
transform 1 0 16008 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_158
timestamp 1604681595
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15640 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15824 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 16376 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_7_175
timestamp 1604681595
transform 1 0 17204 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_173
timestamp 1604681595
transform 1 0 17020 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_169
timestamp 1604681595
transform 1 0 16652 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 16836 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 17664 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17756 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 17388 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_179
timestamp 1604681595
transform 1 0 17572 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_179
timestamp 1604681595
transform 1 0 17572 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 18124 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_183
timestamp 1604681595
transform 1 0 17940 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_182
timestamp 1604681595
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_184
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18216 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18308 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 19872 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19872 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 19688 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 20240 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_196
timestamp 1604681595
transform 1 0 19136 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_206
timestamp 1604681595
transform 1 0 20056 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_195
timestamp 1604681595
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_199
timestamp 1604681595
transform 1 0 19412 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_210
timestamp 1604681595
transform 1 0 20424 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_224
timestamp 1604681595
transform 1 0 21712 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_220
timestamp 1604681595
transform 1 0 21344 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_219
timestamp 1604681595
transform 1 0 21252 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 21896 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 21528 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_228
timestamp 1604681595
transform 1 0 22080 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_229
timestamp 1604681595
transform 1 0 22172 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 21988 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_236
timestamp 1604681595
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_239
timestamp 1604681595
transform 1 0 23092 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__81__A
timestamp 1604681595
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 22264 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1604681595
transform 1 0 22448 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_245
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_240
timestamp 1604681595
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_243
timestamp 1604681595
transform 1 0 23460 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 23644 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 23276 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 23828 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 23828 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 25484 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 25484 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_263
timestamp 1604681595
transform 1 0 25300 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_267
timestamp 1604681595
transform 1 0 25668 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_263
timestamp 1604681595
transform 1 0 25300 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_267
timestamp 1604681595
transform 1 0 25668 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_275
timestamp 1604681595
transform 1 0 26404 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604681595
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1604681595
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1604681595
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1604681595
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1604681595
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_80
timestamp 1604681595
transform 1 0 8464 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9936 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_88
timestamp 1604681595
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_93
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 11500 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10948 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11316 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_105
timestamp 1604681595
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_109
timestamp 1604681595
transform 1 0 11132 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _88_
timestamp 1604681595
transform 1 0 14076 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13156 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 13892 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_129
timestamp 1604681595
transform 1 0 12972 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1604681595
transform 1 0 13340 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_145
timestamp 1604681595
transform 1 0 14444 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16100 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 15916 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 15548 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1604681595
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_154
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_159
timestamp 1604681595
transform 1 0 15732 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 17664 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17480 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_172
timestamp 1604681595
transform 1 0 16928 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 20240 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 19320 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 19872 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_196
timestamp 1604681595
transform 1 0 19136 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_200
timestamp 1604681595
transform 1 0 19504 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_206
timestamp 1604681595
transform 1 0 20056 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 20976 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_210
timestamp 1604681595
transform 1 0 20424 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_215
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 23184 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 23000 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 22632 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_232
timestamp 1604681595
transform 1 0 22448 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_236
timestamp 1604681595
transform 1 0 22816 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1604681595
transform 1 0 25392 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24840 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_256
timestamp 1604681595
transform 1 0 24656 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_260
timestamp 1604681595
transform 1 0 25024 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_267
timestamp 1604681595
transform 1 0 25668 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1604681595
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1604681595
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1604681595
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1604681595
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1604681595
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1604681595
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10120 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 9568 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_86
timestamp 1604681595
transform 1 0 9016 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_94
timestamp 1604681595
transform 1 0 9752 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_114
timestamp 1604681595
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_118
timestamp 1604681595
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_123
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12972 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12788 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 14352 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13984 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_138
timestamp 1604681595
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_142
timestamp 1604681595
transform 1 0 14168 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 14536 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_162
timestamp 1604681595
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1604681595
transform 1 0 16376 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _86_
timestamp 1604681595
transform 1 0 16744 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 18216 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__86__A
timestamp 1604681595
transform 1 0 17296 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 16560 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_174
timestamp 1604681595
transform 1 0 17112 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_178
timestamp 1604681595
transform 1 0 17480 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_184
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 18400 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20056 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_204
timestamp 1604681595
transform 1 0 19872 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_208
timestamp 1604681595
transform 1 0 20240 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 22172 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 20608 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 20424 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21620 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21988 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_221
timestamp 1604681595
transform 1 0 21436 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1604681595
transform 1 0 21804 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 22908 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_235
timestamp 1604681595
transform 1 0 22724 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_239
timestamp 1604681595
transform 1 0 23092 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 25300 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_261
timestamp 1604681595
transform 1 0 25116 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_265
timestamp 1604681595
transform 1 0 25484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1604681595
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1604681595
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1604681595
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1604681595
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1604681595
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_80
timestamp 1604681595
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1604681595
transform 1 0 9936 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_99
timestamp 1604681595
transform 1 0 10212 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12512 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10948 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11960 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 12328 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_116
timestamp 1604681595
transform 1 0 11776 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_120
timestamp 1604681595
transform 1 0 12144 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 14168 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_140
timestamp 1604681595
transform 1 0 13984 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_144
timestamp 1604681595
transform 1 0 14352 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15548 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 14812 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14536 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_148
timestamp 1604681595
transform 1 0 14720 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_152
timestamp 1604681595
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_154
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18308 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 17940 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 17204 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 17572 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_173
timestamp 1604681595
transform 1 0 17020 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_177
timestamp 1604681595
transform 1 0 17388 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_181
timestamp 1604681595
transform 1 0 17756 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_185
timestamp 1604681595
transform 1 0 18124 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18492 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 20056 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 19504 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 19872 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_198
timestamp 1604681595
transform 1 0 19320 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_202
timestamp 1604681595
transform 1 0 19688 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21896 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_209
timestamp 1604681595
transform 1 0 20332 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_224
timestamp 1604681595
transform 1 0 21712 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_228
timestamp 1604681595
transform 1 0 22080 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24104 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 22540 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23644 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 22264 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_232
timestamp 1604681595
transform 1 0 22448 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_242
timestamp 1604681595
transform 1 0 23368 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_247
timestamp 1604681595
transform 1 0 23828 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 25116 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_259
timestamp 1604681595
transform 1 0 24932 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_263
timestamp 1604681595
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1604681595
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1604681595
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1604681595
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1604681595
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_74
timestamp 1604681595
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_86
timestamp 1604681595
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_98
timestamp 1604681595
transform 1 0 10120 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1604681595
transform 1 0 11316 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_106
timestamp 1604681595
transform 1 0 10856 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_114
timestamp 1604681595
transform 1 0 11592 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1604681595
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 13616 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13064 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_126
timestamp 1604681595
transform 1 0 12696 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_132
timestamp 1604681595
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16100 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 15824 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1604681595
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_152
timestamp 1604681595
transform 1 0 15088 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_156
timestamp 1604681595
transform 1 0 15456 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_159
timestamp 1604681595
transform 1 0 15732 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 17480 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_172
timestamp 1604681595
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_176
timestamp 1604681595
transform 1 0 17296 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_180
timestamp 1604681595
transform 1 0 17664 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_187
timestamp 1604681595
transform 1 0 18308 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 19044 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 18492 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_191
timestamp 1604681595
transform 1 0 18676 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 21252 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 21068 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 20700 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_211
timestamp 1604681595
transform 1 0 20516 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_215
timestamp 1604681595
transform 1 0 20884 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_228
timestamp 1604681595
transform 1 0 22080 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 22264 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 22632 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_232
timestamp 1604681595
transform 1 0 22448 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_236
timestamp 1604681595
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_240
timestamp 1604681595
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 24656 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25944 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 25024 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_254
timestamp 1604681595
transform 1 0 24472 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_258
timestamp 1604681595
transform 1 0 24840 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_268
timestamp 1604681595
transform 1 0 25760 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_272
timestamp 1604681595
transform 1 0 26128 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_276
timestamp 1604681595
transform 1 0 26496 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1604681595
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1604681595
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1604681595
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1604681595
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1604681595
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_80
timestamp 1604681595
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11960 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_12_105
timestamp 1604681595
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_117
timestamp 1604681595
transform 1 0 11868 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13524 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13248 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_127
timestamp 1604681595
transform 1 0 12788 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_131
timestamp 1604681595
transform 1 0 13156 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_134
timestamp 1604681595
transform 1 0 13432 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_144
timestamp 1604681595
transform 1 0 14352 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1604681595
transform 1 0 15548 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 14536 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_148
timestamp 1604681595
transform 1 0 14720 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_154
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_161
timestamp 1604681595
transform 1 0 15916 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_165
timestamp 1604681595
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 16652 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 16468 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_185
timestamp 1604681595
transform 1 0 18124 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18860 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18584 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 19872 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_189
timestamp 1604681595
transform 1 0 18492 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_192
timestamp 1604681595
transform 1 0 18768 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_202
timestamp 1604681595
transform 1 0 19688 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_206
timestamp 1604681595
transform 1 0 20056 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21160 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 22172 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_210
timestamp 1604681595
transform 1 0 20424 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_227
timestamp 1604681595
transform 1 0 21988 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 23368 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 23184 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 22816 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_231
timestamp 1604681595
transform 1 0 22356 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_235
timestamp 1604681595
transform 1 0 22724 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_238
timestamp 1604681595
transform 1 0 23000 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_258
timestamp 1604681595
transform 1 0 24840 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_270
timestamp 1604681595
transform 1 0 25944 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_274
timestamp 1604681595
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_276
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1604681595
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1604681595
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1604681595
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1604681595
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1604681595
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1604681595
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1604681595
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1604681595
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_74
timestamp 1604681595
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1604681595
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_80
timestamp 1604681595
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_86
timestamp 1604681595
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_98
timestamp 1604681595
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_110
timestamp 1604681595
transform 1 0 11224 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_123
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_105
timestamp 1604681595
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_117
timestamp 1604681595
transform 1 0 11868 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_125
timestamp 1604681595
transform 1 0 12604 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_131
timestamp 1604681595
transform 1 0 13156 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_128
timestamp 1604681595
transform 1 0 12880 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12696 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13064 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13248 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1604681595
transform 1 0 12880 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_141
timestamp 1604681595
transform 1 0 14076 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 13708 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13892 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_145
timestamp 1604681595
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_145
timestamp 1604681595
transform 1 0 14444 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_154
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_149
timestamp 1604681595
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 14628 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15456 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_158
timestamp 1604681595
transform 1 0 15640 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_165
timestamp 1604681595
transform 1 0 16284 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15916 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 16100 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 14812 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_13_176
timestamp 1604681595
transform 1 0 17296 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1604681595
transform 1 0 16652 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 16468 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16836 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1604681595
transform 1 0 17020 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_183
timestamp 1604681595
transform 1 0 17940 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_179
timestamp 1604681595
transform 1 0 17572 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_180
timestamp 1604681595
transform 1 0 17664 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 18124 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 17756 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1604681595
transform 1 0 18308 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18584 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_203
timestamp 1604681595
transform 1 0 19780 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_199
timestamp 1604681595
transform 1 0 19412 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_204
timestamp 1604681595
transform 1 0 19872 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_200
timestamp 1604681595
transform 1 0 19504 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 19964 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19688 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 19596 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 20056 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 20148 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 20240 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_210
timestamp 1604681595
transform 1 0 20424 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 21068 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_228
timestamp 1604681595
transform 1 0 22080 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_228
timestamp 1604681595
transform 1 0 22080 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_224
timestamp 1604681595
transform 1 0 21712 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 21896 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 21252 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_236
timestamp 1604681595
transform 1 0 22816 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_232
timestamp 1604681595
transform 1 0 22448 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_236
timestamp 1604681595
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 23000 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 22632 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 22264 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 22264 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__85__A
timestamp 1604681595
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _85_
timestamp 1604681595
transform 1 0 22448 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_240
timestamp 1604681595
transform 1 0 23184 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_245
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_240
timestamp 1604681595
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 23276 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 23736 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 25392 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 24932 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_262
timestamp 1604681595
transform 1 0 25208 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_266
timestamp 1604681595
transform 1 0 25576 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_257
timestamp 1604681595
transform 1 0 24748 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_261
timestamp 1604681595
transform 1 0 25116 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_274
timestamp 1604681595
transform 1 0 26312 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_273
timestamp 1604681595
transform 1 0 26220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_276
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1604681595
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1604681595
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1604681595
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1604681595
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1604681595
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_74
timestamp 1604681595
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_86
timestamp 1604681595
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_98
timestamp 1604681595
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_110
timestamp 1604681595
transform 1 0 11224 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_123
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13064 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14352 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14168 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 12880 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_127
timestamp 1604681595
transform 1 0 12788 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_136
timestamp 1604681595
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_140
timestamp 1604681595
transform 1 0 13984 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16008 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 15364 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_153
timestamp 1604681595
transform 1 0 15180 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_157
timestamp 1604681595
transform 1 0 15548 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16836 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_180
timestamp 1604681595
transform 1 0 17664 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20240 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20056 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19688 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_200
timestamp 1604681595
transform 1 0 19504 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_204
timestamp 1604681595
transform 1 0 19872 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21988 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21804 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 21252 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_217
timestamp 1604681595
transform 1 0 21068 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_221
timestamp 1604681595
transform 1 0 21436 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_236
timestamp 1604681595
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_240
timestamp 1604681595
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1604681595
transform 1 0 25208 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 24656 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 25024 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1604681595
transform 1 0 25760 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_254
timestamp 1604681595
transform 1 0 24472 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_258
timestamp 1604681595
transform 1 0 24840 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_266
timestamp 1604681595
transform 1 0 25576 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_270
timestamp 1604681595
transform 1 0 25944 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_276
timestamp 1604681595
transform 1 0 26496 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1604681595
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1604681595
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1604681595
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1604681595
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1604681595
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_80
timestamp 1604681595
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_105
timestamp 1604681595
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_117
timestamp 1604681595
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1604681595
transform 1 0 14168 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_129
timestamp 1604681595
transform 1 0 12972 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_141
timestamp 1604681595
transform 1 0 14076 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_145
timestamp 1604681595
transform 1 0 14444 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14812 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1604681595
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_163
timestamp 1604681595
transform 1 0 16100 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 17020 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16836 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 16468 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_169
timestamp 1604681595
transform 1 0 16652 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18860 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 21252 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 21068 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20516 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_209
timestamp 1604681595
transform 1 0 20332 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_213
timestamp 1604681595
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 23460 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 23092 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_235
timestamp 1604681595
transform 1 0 22724 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_241
timestamp 1604681595
transform 1 0 23276 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_259
timestamp 1604681595
transform 1 0 24932 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_271
timestamp 1604681595
transform 1 0 26036 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1604681595
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1604681595
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1604681595
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1604681595
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1604681595
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_74
timestamp 1604681595
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_86
timestamp 1604681595
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_98
timestamp 1604681595
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_110
timestamp 1604681595
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_135
timestamp 1604681595
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15180 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16284 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_147
timestamp 1604681595
transform 1 0 14628 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_159
timestamp 1604681595
transform 1 0 15732 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_163
timestamp 1604681595
transform 1 0 16100 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_167
timestamp 1604681595
transform 1 0 16468 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16744 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1604681595
transform 1 0 16928 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_175
timestamp 1604681595
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_179
timestamp 1604681595
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_184
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 18308 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1604681595
transform 1 0 18492 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 19504 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_192
timestamp 1604681595
transform 1 0 18768 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_197
timestamp 1604681595
transform 1 0 19228 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21988 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21804 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21436 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_216
timestamp 1604681595
transform 1 0 20976 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_220
timestamp 1604681595
transform 1 0 21344 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_223
timestamp 1604681595
transform 1 0 21620 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_236
timestamp 1604681595
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_240
timestamp 1604681595
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25300 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_261
timestamp 1604681595
transform 1 0 25116 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_265
timestamp 1604681595
transform 1 0 25484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1604681595
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1604681595
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1604681595
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1604681595
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1604681595
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_80
timestamp 1604681595
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1604681595
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_117
timestamp 1604681595
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_129
timestamp 1604681595
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1604681595
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_154
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_166
timestamp 1604681595
transform 1 0 16376 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1604681595
transform 1 0 17112 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 18124 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_183
timestamp 1604681595
transform 1 0 17940 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_187
timestamp 1604681595
transform 1 0 18308 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19044 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 18860 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18492 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_191
timestamp 1604681595
transform 1 0 18676 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_204
timestamp 1604681595
transform 1 0 19872 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_208
timestamp 1604681595
transform 1 0 20240 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 20424 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1604681595
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 23092 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 22908 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 22540 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 24104 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_231
timestamp 1604681595
transform 1 0 22356 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_235
timestamp 1604681595
transform 1 0 22724 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_248
timestamp 1604681595
transform 1 0 23920 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24656 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_252
timestamp 1604681595
transform 1 0 24288 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_262
timestamp 1604681595
transform 1 0 25208 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_274
timestamp 1604681595
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_276
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1604681595
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1604681595
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1604681595
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1604681595
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1604681595
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1604681595
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1604681595
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1604681595
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1604681595
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1604681595
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_86
timestamp 1604681595
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_98
timestamp 1604681595
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_110
timestamp 1604681595
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1604681595
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1604681595
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1604681595
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_129
timestamp 1604681595
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1604681595
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_147
timestamp 1604681595
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_159
timestamp 1604681595
transform 1 0 15732 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_166
timestamp 1604681595
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1604681595
transform 1 0 16744 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_167
timestamp 1604681595
transform 1 0 16468 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_173
timestamp 1604681595
transform 1 0 17020 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1604681595
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_184
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1604681595
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_196
timestamp 1604681595
transform 1 0 19136 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_192
timestamp 1604681595
transform 1 0 18768 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_190
timestamp 1604681595
transform 1 0 18584 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18584 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 18400 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 18952 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18768 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18952 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_20_206
timestamp 1604681595
transform 1 0 20056 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_203
timestamp 1604681595
transform 1 0 19780 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20148 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_209
timestamp 1604681595
transform 1 0 20332 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21068 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20516 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20700 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_20_224
timestamp 1604681595
transform 1 0 21712 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_219
timestamp 1604681595
transform 1 0 21252 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_226
timestamp 1604681595
transform 1 0 21896 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1604681595
transform 1 0 21528 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 21712 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1604681595
transform 1 0 21436 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_235
timestamp 1604681595
transform 1 0 22724 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_236
timestamp 1604681595
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__84__A
timestamp 1604681595
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _84_
timestamp 1604681595
transform 1 0 22448 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1604681595
transform 1 0 22448 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_240
timestamp 1604681595
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__87__A
timestamp 1604681595
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _87_
timestamp 1604681595
transform 1 0 23460 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_247
timestamp 1604681595
transform 1 0 23828 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24012 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_251
timestamp 1604681595
transform 1 0 24196 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_257
timestamp 1604681595
transform 1 0 24748 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_251
timestamp 1604681595
transform 1 0 24196 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1604681595
transform 1 0 24564 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1604681595
transform 1 0 24932 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1604681595
transform 1 0 24564 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_267
timestamp 1604681595
transform 1 0 25668 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_263
timestamp 1604681595
transform 1 0 25300 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1604681595
transform 1 0 25484 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_259
timestamp 1604681595
transform 1 0 24932 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_275
timestamp 1604681595
transform 1 0 26404 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_271
timestamp 1604681595
transform 1 0 26036 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_276
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1604681595
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1604681595
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1604681595
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1604681595
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_74
timestamp 1604681595
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_86
timestamp 1604681595
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_98
timestamp 1604681595
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_110
timestamp 1604681595
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1604681595
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_147
timestamp 1604681595
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_159
timestamp 1604681595
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_171
timestamp 1604681595
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1604681595
transform 1 0 19596 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19228 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_192
timestamp 1604681595
transform 1 0 18768 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_195
timestamp 1604681595
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_199
timestamp 1604681595
transform 1 0 19412 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_204
timestamp 1604681595
transform 1 0 19872 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1604681595
transform 1 0 22080 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1604681595
transform 1 0 21068 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_216
timestamp 1604681595
transform 1 0 20976 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_220
timestamp 1604681595
transform 1 0 21344 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 22540 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_231
timestamp 1604681595
transform 1 0 22356 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_235
timestamp 1604681595
transform 1 0 22724 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_241
timestamp 1604681595
transform 1 0 23276 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _89_
timestamp 1604681595
transform 1 0 24932 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__89__A
timestamp 1604681595
transform 1 0 25484 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1604681595
transform 1 0 24564 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_251
timestamp 1604681595
transform 1 0 24196 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_257
timestamp 1604681595
transform 1 0 24748 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_263
timestamp 1604681595
transform 1 0 25300 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_267
timestamp 1604681595
transform 1 0 25668 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_275
timestamp 1604681595
transform 1 0 26404 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1604681595
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1604681595
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1604681595
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1604681595
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1604681595
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_80
timestamp 1604681595
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_93
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_105
timestamp 1604681595
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_117
timestamp 1604681595
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_129
timestamp 1604681595
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1604681595
transform 1 0 14076 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1604681595
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1604681595
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1604681595
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_202
timestamp 1604681595
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 22172 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_227
timestamp 1604681595
transform 1 0 21988 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_235
timestamp 1604681595
transform 1 0 22724 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_247
timestamp 1604681595
transform 1 0 23828 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604681595
transform 1 0 24564 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_259
timestamp 1604681595
transform 1 0 24932 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_271
timestamp 1604681595
transform 1 0 26036 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_276
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1604681595
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1604681595
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1604681595
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1604681595
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1604681595
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1604681595
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_98
timestamp 1604681595
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_110
timestamp 1604681595
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1604681595
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1604681595
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_159
timestamp 1604681595
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_171
timestamp 1604681595
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1604681595
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1604681595
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 21896 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_220
timestamp 1604681595
transform 1 0 21344 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_228
timestamp 1604681595
transform 1 0 22080 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23920 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1604681595
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_242
timestamp 1604681595
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_245
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604681595
transform 1 0 25208 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1604681595
transform 1 0 25760 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24656 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_254
timestamp 1604681595
transform 1 0 24472 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_258
timestamp 1604681595
transform 1 0 24840 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_266
timestamp 1604681595
transform 1 0 25576 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_270
timestamp 1604681595
transform 1 0 25944 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_276
timestamp 1604681595
transform 1 0 26496 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1604681595
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1604681595
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1604681595
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1604681595
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1604681595
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_80
timestamp 1604681595
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1604681595
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_117
timestamp 1604681595
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_129
timestamp 1604681595
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1604681595
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1604681595
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1604681595
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1604681595
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_202
timestamp 1604681595
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 21896 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_223
timestamp 1604681595
transform 1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604681595
transform 1 0 23184 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_232
timestamp 1604681595
transform 1 0 22448 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_244
timestamp 1604681595
transform 1 0 23552 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_256
timestamp 1604681595
transform 1 0 24656 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_268
timestamp 1604681595
transform 1 0 25760 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_274
timestamp 1604681595
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_276
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1604681595
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1604681595
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1604681595
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1604681595
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1604681595
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1604681595
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1604681595
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1604681595
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1604681595
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16284 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_147
timestamp 1604681595
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_159
timestamp 1604681595
transform 1 0 15732 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_167
timestamp 1604681595
transform 1 0 16468 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_179
timestamp 1604681595
transform 1 0 17572 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1604681595
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1604681595
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_220
timestamp 1604681595
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1604681595
transform 1 0 22724 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_232
timestamp 1604681595
transform 1 0 22448 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_237
timestamp 1604681595
transform 1 0 22908 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_243
timestamp 1604681595
transform 1 0 23460 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604681595
transform 1 0 24932 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1604681595
transform 1 0 25484 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24380 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_251
timestamp 1604681595
transform 1 0 24196 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_255
timestamp 1604681595
transform 1 0 24564 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_263
timestamp 1604681595
transform 1 0 25300 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_267
timestamp 1604681595
transform 1 0 25668 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_275
timestamp 1604681595
transform 1 0 26404 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1604681595
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1604681595
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1604681595
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1604681595
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1604681595
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1604681595
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1604681595
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1604681595
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1604681595
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1604681595
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_86
timestamp 1604681595
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_98
timestamp 1604681595
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 11316 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1604681595
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1604681595
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_110
timestamp 1604681595
transform 1 0 11224 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_113
timestamp 1604681595
transform 1 0 11500 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_121
timestamp 1604681595
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_123
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13156 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13892 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1604681595
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1604681595
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_137
timestamp 1604681595
transform 1 0 13708 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_141
timestamp 1604681595
transform 1 0 14076 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16284 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_154
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_162
timestamp 1604681595
transform 1 0 16008 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_153
timestamp 1604681595
transform 1 0 15180 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_165
timestamp 1604681595
transform 1 0 16284 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_171
timestamp 1604681595
transform 1 0 16836 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_183
timestamp 1604681595
transform 1 0 17940 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_177
timestamp 1604681595
transform 1 0 17388 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_195
timestamp 1604681595
transform 1 0 19044 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_207
timestamp 1604681595
transform 1 0 20148 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1604681595
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1604681595
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_213
timestamp 1604681595
transform 1 0 20700 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_215
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_227
timestamp 1604681595
transform 1 0 21988 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_220
timestamp 1604681595
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1604681595
transform 1 0 22724 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_239
timestamp 1604681595
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_232
timestamp 1604681595
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_245
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604681595
transform 1 0 24564 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1604681595
transform 1 0 25116 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1604681595
transform 1 0 24380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_251
timestamp 1604681595
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_263
timestamp 1604681595
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_259
timestamp 1604681595
transform 1 0 24932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_263
timestamp 1604681595
transform 1 0 25300 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_275
timestamp 1604681595
transform 1 0 26404 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1604681595
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1604681595
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1604681595
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1604681595
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1604681595
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1604681595
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11316 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_105
timestamp 1604681595
transform 1 0 10764 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_117
timestamp 1604681595
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_129
timestamp 1604681595
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1604681595
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1604681595
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1604681595
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1604681595
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1604681595
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_215
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_227
timestamp 1604681595
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_239
timestamp 1604681595
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604681595
transform 1 0 24564 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_251
timestamp 1604681595
transform 1 0 24196 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_259
timestamp 1604681595
transform 1 0 24932 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_271
timestamp 1604681595
transform 1 0 26036 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1604681595
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1604681595
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1604681595
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1604681595
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1604681595
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1604681595
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_86
timestamp 1604681595
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_98
timestamp 1604681595
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_110
timestamp 1604681595
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13524 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14260 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_141
timestamp 1604681595
transform 1 0 14076 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_145
timestamp 1604681595
transform 1 0 14444 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604681595
transform 1 0 14812 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1604681595
transform 1 0 15364 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_153
timestamp 1604681595
transform 1 0 15180 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_157
timestamp 1604681595
transform 1 0 15548 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_169
timestamp 1604681595
transform 1 0 16652 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_181
timestamp 1604681595
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1604681595
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1604681595
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_220
timestamp 1604681595
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_232
timestamp 1604681595
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_245
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1604681595
transform 1 0 24564 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_253
timestamp 1604681595
transform 1 0 24380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_257
timestamp 1604681595
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_269
timestamp 1604681595
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1604681595
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1604681595
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1604681595
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1604681595
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1604681595
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1604681595
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1604681595
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_117
timestamp 1604681595
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_129
timestamp 1604681595
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1604681595
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1604681595
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_178
timestamp 1604681595
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_190
timestamp 1604681595
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_202
timestamp 1604681595
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_227
timestamp 1604681595
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_239
timestamp 1604681595
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1604681595
transform 1 0 24564 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_251
timestamp 1604681595
transform 1 0 24196 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_259
timestamp 1604681595
transform 1 0 24932 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_271
timestamp 1604681595
transform 1 0 26036 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_276
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1604681595
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1604681595
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1604681595
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1604681595
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1604681595
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1604681595
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1604681595
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1604681595
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1604681595
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15640 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16376 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_147
timestamp 1604681595
transform 1 0 14628 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_155
timestamp 1604681595
transform 1 0 15364 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_164
timestamp 1604681595
transform 1 0 16192 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 17020 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_168
timestamp 1604681595
transform 1 0 16560 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_172
timestamp 1604681595
transform 1 0 16928 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_175
timestamp 1604681595
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_179
timestamp 1604681595
transform 1 0 17572 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1604681595
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1604681595
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_220
timestamp 1604681595
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_232
timestamp 1604681595
transform 1 0 22448 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_240
timestamp 1604681595
transform 1 0 23184 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1604681595
transform 1 0 24932 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1604681595
transform 1 0 25484 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24380 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_251
timestamp 1604681595
transform 1 0 24196 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_255
timestamp 1604681595
transform 1 0 24564 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_263
timestamp 1604681595
transform 1 0 25300 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_267
timestamp 1604681595
transform 1 0 25668 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_275
timestamp 1604681595
transform 1 0 26404 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1604681595
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1604681595
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1604681595
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1604681595
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1604681595
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_80
timestamp 1604681595
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1604681595
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_117
timestamp 1604681595
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_129
timestamp 1604681595
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1604681595
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_154
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_166
timestamp 1604681595
transform 1 0 16376 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 17020 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_32_172
timestamp 1604681595
transform 1 0 16928 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_189
timestamp 1604681595
transform 1 0 18492 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_201
timestamp 1604681595
transform 1 0 19596 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_213
timestamp 1604681595
transform 1 0 20700 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_215
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_227
timestamp 1604681595
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23460 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_239
timestamp 1604681595
transform 1 0 23092 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_249
timestamp 1604681595
transform 1 0 24012 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_261
timestamp 1604681595
transform 1 0 25116 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_273
timestamp 1604681595
transform 1 0 26220 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_276
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1604681595
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1604681595
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1604681595
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1604681595
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1604681595
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_51
timestamp 1604681595
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1604681595
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1604681595
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1604681595
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_74
timestamp 1604681595
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1604681595
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_80
timestamp 1604681595
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_86
timestamp 1604681595
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_98
timestamp 1604681595
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_110
timestamp 1604681595
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_123
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1604681595
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_117
timestamp 1604681595
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_135
timestamp 1604681595
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_129
timestamp 1604681595
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1604681595
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_147
timestamp 1604681595
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_159
timestamp 1604681595
transform 1 0 15732 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_166
timestamp 1604681595
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1604681595
transform 1 0 16652 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1604681595
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_167
timestamp 1604681595
transform 1 0 16468 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_173
timestamp 1604681595
transform 1 0 17020 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_177
timestamp 1604681595
transform 1 0 17388 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_178
timestamp 1604681595
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1604681595
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1604681595
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_190
timestamp 1604681595
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_202
timestamp 1604681595
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_220
timestamp 1604681595
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_227
timestamp 1604681595
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23552 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23828 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_232
timestamp 1604681595
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_245
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_249
timestamp 1604681595
transform 1 0 24012 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_239
timestamp 1604681595
transform 1 0 23092 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_243
timestamp 1604681595
transform 1 0 23460 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_250
timestamp 1604681595
transform 1 0 24104 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1604681595
transform 1 0 24840 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1604681595
transform 1 0 24564 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1604681595
transform 1 0 25116 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1604681595
transform 1 0 25484 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_259
timestamp 1604681595
transform 1 0 24932 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_263
timestamp 1604681595
transform 1 0 25300 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_267
timestamp 1604681595
transform 1 0 25668 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_262
timestamp 1604681595
transform 1 0 25208 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_275
timestamp 1604681595
transform 1 0 26404 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_274
timestamp 1604681595
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604681595
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1604681595
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1604681595
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_51
timestamp 1604681595
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_59
timestamp 1604681595
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_62
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_74
timestamp 1604681595
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_86
timestamp 1604681595
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_98
timestamp 1604681595
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_110
timestamp 1604681595
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_123
timestamp 1604681595
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 14260 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_135
timestamp 1604681595
transform 1 0 13524 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14996 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_149
timestamp 1604681595
transform 1 0 14812 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_153
timestamp 1604681595
transform 1 0 15180 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_165
timestamp 1604681595
transform 1 0 16284 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_177
timestamp 1604681595
transform 1 0 17388 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1604681595
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1604681595
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_208
timestamp 1604681595
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_220
timestamp 1604681595
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23644 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23368 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_232
timestamp 1604681595
transform 1 0 22448 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_240
timestamp 1604681595
transform 1 0 23184 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1604681595
transform 1 0 24932 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1604681595
transform 1 0 25484 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1604681595
transform 1 0 24748 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24380 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_251
timestamp 1604681595
transform 1 0 24196 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_255
timestamp 1604681595
transform 1 0 24564 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_263
timestamp 1604681595
transform 1 0 25300 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_267
timestamp 1604681595
transform 1 0 25668 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_275
timestamp 1604681595
transform 1 0 26404 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1604681595
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1604681595
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1604681595
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1604681595
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_44
timestamp 1604681595
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_56
timestamp 1604681595
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_68
timestamp 1604681595
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_80
timestamp 1604681595
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_93
timestamp 1604681595
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_105
timestamp 1604681595
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_117
timestamp 1604681595
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_129
timestamp 1604681595
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1604681595
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_154
timestamp 1604681595
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_166
timestamp 1604681595
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_178
timestamp 1604681595
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_190
timestamp 1604681595
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_202
timestamp 1604681595
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_215
timestamp 1604681595
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_227
timestamp 1604681595
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23552 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_239
timestamp 1604681595
transform 1 0 23092 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_243
timestamp 1604681595
transform 1 0 23460 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_250
timestamp 1604681595
transform 1 0 24104 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1604681595
transform 1 0 24840 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_262
timestamp 1604681595
transform 1 0 25208 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_274
timestamp 1604681595
transform 1 0 26312 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_276
timestamp 1604681595
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1604681595
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1604681595
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1604681595
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1604681595
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_51
timestamp 1604681595
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_59
timestamp 1604681595
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_62
timestamp 1604681595
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_74
timestamp 1604681595
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_86
timestamp 1604681595
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_98
timestamp 1604681595
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 12604 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_110
timestamp 1604681595
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_123
timestamp 1604681595
transform 1 0 12420 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_127
timestamp 1604681595
transform 1 0 12788 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_139
timestamp 1604681595
transform 1 0 13892 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_151
timestamp 1604681595
transform 1 0 14996 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_163
timestamp 1604681595
transform 1 0 16100 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_175
timestamp 1604681595
transform 1 0 17204 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_184
timestamp 1604681595
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_196
timestamp 1604681595
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_208
timestamp 1604681595
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_220
timestamp 1604681595
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_232
timestamp 1604681595
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_245
timestamp 1604681595
transform 1 0 23644 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1604681595
transform 1 0 24564 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1604681595
transform 1 0 25116 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1604681595
transform 1 0 24380 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_259
timestamp 1604681595
transform 1 0 24932 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_263
timestamp 1604681595
transform 1 0 25300 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_275
timestamp 1604681595
transform 1 0 26404 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1604681595
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1604681595
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1604681595
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1604681595
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_44
timestamp 1604681595
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_56
timestamp 1604681595
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_68
timestamp 1604681595
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_80
timestamp 1604681595
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_93
timestamp 1604681595
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12512 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_105
timestamp 1604681595
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_117
timestamp 1604681595
transform 1 0 11868 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_123
timestamp 1604681595
transform 1 0 12420 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_130
timestamp 1604681595
transform 1 0 13064 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_142
timestamp 1604681595
transform 1 0 14168 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_150
timestamp 1604681595
transform 1 0 14904 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_154
timestamp 1604681595
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_166
timestamp 1604681595
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_178
timestamp 1604681595
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_190
timestamp 1604681595
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_202
timestamp 1604681595
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_215
timestamp 1604681595
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_227
timestamp 1604681595
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_239
timestamp 1604681595
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1604681595
transform 1 0 24564 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_251
timestamp 1604681595
transform 1 0 24196 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_259
timestamp 1604681595
transform 1 0 24932 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604681595
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_271
timestamp 1604681595
transform 1 0 26036 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_276
timestamp 1604681595
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1604681595
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1604681595
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1604681595
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1604681595
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604681595
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1604681595
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1604681595
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1604681595
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_32
timestamp 1604681595
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604681595
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_51
timestamp 1604681595
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_59
timestamp 1604681595
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_62
timestamp 1604681595
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_44
timestamp 1604681595
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_56
timestamp 1604681595
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_74
timestamp 1604681595
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_68
timestamp 1604681595
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_80
timestamp 1604681595
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604681595
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_86
timestamp 1604681595
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_98
timestamp 1604681595
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_93
timestamp 1604681595
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604681595
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_110
timestamp 1604681595
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_123
timestamp 1604681595
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_105
timestamp 1604681595
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_117
timestamp 1604681595
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_135
timestamp 1604681595
transform 1 0 13524 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_129
timestamp 1604681595
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1604681595
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604681595
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_147
timestamp 1604681595
transform 1 0 14628 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_159
timestamp 1604681595
transform 1 0 15732 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_154
timestamp 1604681595
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_166
timestamp 1604681595
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604681595
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_171
timestamp 1604681595
transform 1 0 16836 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_184
timestamp 1604681595
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_178
timestamp 1604681595
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_196
timestamp 1604681595
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_208
timestamp 1604681595
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_190
timestamp 1604681595
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_202
timestamp 1604681595
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604681595
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_220
timestamp 1604681595
transform 1 0 21344 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_215
timestamp 1604681595
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_227
timestamp 1604681595
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1604681595
transform 1 0 23276 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604681595
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_232
timestamp 1604681595
transform 1 0 22448 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_245
timestamp 1604681595
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_239
timestamp 1604681595
transform 1 0 23092 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_245
timestamp 1604681595
transform 1 0 23644 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1604681595
transform 1 0 24564 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1604681595
transform 1 0 24564 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1604681595
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1604681595
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_259
timestamp 1604681595
transform 1 0 24932 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_263
timestamp 1604681595
transform 1 0 25300 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1604681595
transform 1 0 24380 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_259
timestamp 1604681595
transform 1 0 24932 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604681595
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_275
timestamp 1604681595
transform 1 0 26404 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_271
timestamp 1604681595
transform 1 0 26036 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_276
timestamp 1604681595
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1604681595
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1604681595
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1604681595
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1604681595
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604681595
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_51
timestamp 1604681595
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_59
timestamp 1604681595
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_62
timestamp 1604681595
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_74
timestamp 1604681595
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_86
timestamp 1604681595
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_98
timestamp 1604681595
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604681595
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_110
timestamp 1604681595
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_123
timestamp 1604681595
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_135
timestamp 1604681595
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_147
timestamp 1604681595
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_159
timestamp 1604681595
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604681595
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_171
timestamp 1604681595
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1604681595
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_196
timestamp 1604681595
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_208
timestamp 1604681595
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_220
timestamp 1604681595
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604681595
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_232
timestamp 1604681595
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_245
timestamp 1604681595
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_257
timestamp 1604681595
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_269
timestamp 1604681595
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1604681595
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1604681595
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604681595
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1604681595
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1604681595
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604681595
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_44
timestamp 1604681595
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_56
timestamp 1604681595
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_63
timestamp 1604681595
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_75
timestamp 1604681595
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604681595
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_87
timestamp 1604681595
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_94
timestamp 1604681595
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604681595
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_106
timestamp 1604681595
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_118
timestamp 1604681595
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_125
timestamp 1604681595
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_137
timestamp 1604681595
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604681595
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_149
timestamp 1604681595
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_156
timestamp 1604681595
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604681595
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_168
timestamp 1604681595
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_180
timestamp 1604681595
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_187
timestamp 1604681595
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_199
timestamp 1604681595
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604681595
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_211
timestamp 1604681595
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_218
timestamp 1604681595
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604681595
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_230
timestamp 1604681595
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_242
timestamp 1604681595
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_249
timestamp 1604681595
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_261
timestamp 1604681595
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_273
timestamp 1604681595
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 26882 0 26938 480 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 3514 27520 3570 28000 6 SC_IN_TOP
port 1 nsew default input
rlabel metal2 s 27526 0 27582 480 6 SC_OUT_BOT
port 2 nsew default tristate
rlabel metal2 s 24490 27520 24546 28000 6 SC_OUT_TOP
port 3 nsew default tristate
rlabel metal2 s 294 0 350 480 6 bottom_left_grid_pin_1_
port 4 nsew default input
rlabel metal2 s 17498 27520 17554 28000 6 ccff_head
port 5 nsew default input
rlabel metal3 s 0 14016 480 14136 6 ccff_tail
port 6 nsew default tristate
rlabel metal3 s 27520 4768 28000 4888 6 chanx_right_in[0]
port 7 nsew default input
rlabel metal3 s 27520 10480 28000 10600 6 chanx_right_in[10]
port 8 nsew default input
rlabel metal3 s 27520 11024 28000 11144 6 chanx_right_in[11]
port 9 nsew default input
rlabel metal3 s 27520 11704 28000 11824 6 chanx_right_in[12]
port 10 nsew default input
rlabel metal3 s 27520 12248 28000 12368 6 chanx_right_in[13]
port 11 nsew default input
rlabel metal3 s 27520 12792 28000 12912 6 chanx_right_in[14]
port 12 nsew default input
rlabel metal3 s 27520 13336 28000 13456 6 chanx_right_in[15]
port 13 nsew default input
rlabel metal3 s 27520 13880 28000 14000 6 chanx_right_in[16]
port 14 nsew default input
rlabel metal3 s 27520 14560 28000 14680 6 chanx_right_in[17]
port 15 nsew default input
rlabel metal3 s 27520 15104 28000 15224 6 chanx_right_in[18]
port 16 nsew default input
rlabel metal3 s 27520 15648 28000 15768 6 chanx_right_in[19]
port 17 nsew default input
rlabel metal3 s 27520 5312 28000 5432 6 chanx_right_in[1]
port 18 nsew default input
rlabel metal3 s 27520 5992 28000 6112 6 chanx_right_in[2]
port 19 nsew default input
rlabel metal3 s 27520 6536 28000 6656 6 chanx_right_in[3]
port 20 nsew default input
rlabel metal3 s 27520 7080 28000 7200 6 chanx_right_in[4]
port 21 nsew default input
rlabel metal3 s 27520 7624 28000 7744 6 chanx_right_in[5]
port 22 nsew default input
rlabel metal3 s 27520 8168 28000 8288 6 chanx_right_in[6]
port 23 nsew default input
rlabel metal3 s 27520 8848 28000 8968 6 chanx_right_in[7]
port 24 nsew default input
rlabel metal3 s 27520 9392 28000 9512 6 chanx_right_in[8]
port 25 nsew default input
rlabel metal3 s 27520 9936 28000 10056 6 chanx_right_in[9]
port 26 nsew default input
rlabel metal3 s 27520 16192 28000 16312 6 chanx_right_out[0]
port 27 nsew default tristate
rlabel metal3 s 27520 21904 28000 22024 6 chanx_right_out[10]
port 28 nsew default tristate
rlabel metal3 s 27520 22448 28000 22568 6 chanx_right_out[11]
port 29 nsew default tristate
rlabel metal3 s 27520 23128 28000 23248 6 chanx_right_out[12]
port 30 nsew default tristate
rlabel metal3 s 27520 23672 28000 23792 6 chanx_right_out[13]
port 31 nsew default tristate
rlabel metal3 s 27520 24216 28000 24336 6 chanx_right_out[14]
port 32 nsew default tristate
rlabel metal3 s 27520 24760 28000 24880 6 chanx_right_out[15]
port 33 nsew default tristate
rlabel metal3 s 27520 25304 28000 25424 6 chanx_right_out[16]
port 34 nsew default tristate
rlabel metal3 s 27520 25984 28000 26104 6 chanx_right_out[17]
port 35 nsew default tristate
rlabel metal3 s 27520 26528 28000 26648 6 chanx_right_out[18]
port 36 nsew default tristate
rlabel metal3 s 27520 27072 28000 27192 6 chanx_right_out[19]
port 37 nsew default tristate
rlabel metal3 s 27520 16736 28000 16856 6 chanx_right_out[1]
port 38 nsew default tristate
rlabel metal3 s 27520 17416 28000 17536 6 chanx_right_out[2]
port 39 nsew default tristate
rlabel metal3 s 27520 17960 28000 18080 6 chanx_right_out[3]
port 40 nsew default tristate
rlabel metal3 s 27520 18504 28000 18624 6 chanx_right_out[4]
port 41 nsew default tristate
rlabel metal3 s 27520 19048 28000 19168 6 chanx_right_out[5]
port 42 nsew default tristate
rlabel metal3 s 27520 19592 28000 19712 6 chanx_right_out[6]
port 43 nsew default tristate
rlabel metal3 s 27520 20272 28000 20392 6 chanx_right_out[7]
port 44 nsew default tristate
rlabel metal3 s 27520 20816 28000 20936 6 chanx_right_out[8]
port 45 nsew default tristate
rlabel metal3 s 27520 21360 28000 21480 6 chanx_right_out[9]
port 46 nsew default tristate
rlabel metal2 s 938 0 994 480 6 chany_bottom_in[0]
port 47 nsew default input
rlabel metal2 s 7378 0 7434 480 6 chany_bottom_in[10]
port 48 nsew default input
rlabel metal2 s 8022 0 8078 480 6 chany_bottom_in[11]
port 49 nsew default input
rlabel metal2 s 8666 0 8722 480 6 chany_bottom_in[12]
port 50 nsew default input
rlabel metal2 s 9310 0 9366 480 6 chany_bottom_in[13]
port 51 nsew default input
rlabel metal2 s 10046 0 10102 480 6 chany_bottom_in[14]
port 52 nsew default input
rlabel metal2 s 10690 0 10746 480 6 chany_bottom_in[15]
port 53 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_in[16]
port 54 nsew default input
rlabel metal2 s 11978 0 12034 480 6 chany_bottom_in[17]
port 55 nsew default input
rlabel metal2 s 12622 0 12678 480 6 chany_bottom_in[18]
port 56 nsew default input
rlabel metal2 s 13266 0 13322 480 6 chany_bottom_in[19]
port 57 nsew default input
rlabel metal2 s 1582 0 1638 480 6 chany_bottom_in[1]
port 58 nsew default input
rlabel metal2 s 2226 0 2282 480 6 chany_bottom_in[2]
port 59 nsew default input
rlabel metal2 s 2870 0 2926 480 6 chany_bottom_in[3]
port 60 nsew default input
rlabel metal2 s 3514 0 3570 480 6 chany_bottom_in[4]
port 61 nsew default input
rlabel metal2 s 4158 0 4214 480 6 chany_bottom_in[5]
port 62 nsew default input
rlabel metal2 s 4802 0 4858 480 6 chany_bottom_in[6]
port 63 nsew default input
rlabel metal2 s 5446 0 5502 480 6 chany_bottom_in[7]
port 64 nsew default input
rlabel metal2 s 6090 0 6146 480 6 chany_bottom_in[8]
port 65 nsew default input
rlabel metal2 s 6734 0 6790 480 6 chany_bottom_in[9]
port 66 nsew default input
rlabel metal2 s 13910 0 13966 480 6 chany_bottom_out[0]
port 67 nsew default tristate
rlabel metal2 s 20442 0 20498 480 6 chany_bottom_out[10]
port 68 nsew default tristate
rlabel metal2 s 21086 0 21142 480 6 chany_bottom_out[11]
port 69 nsew default tristate
rlabel metal2 s 21730 0 21786 480 6 chany_bottom_out[12]
port 70 nsew default tristate
rlabel metal2 s 22374 0 22430 480 6 chany_bottom_out[13]
port 71 nsew default tristate
rlabel metal2 s 23018 0 23074 480 6 chany_bottom_out[14]
port 72 nsew default tristate
rlabel metal2 s 23662 0 23718 480 6 chany_bottom_out[15]
port 73 nsew default tristate
rlabel metal2 s 24306 0 24362 480 6 chany_bottom_out[16]
port 74 nsew default tristate
rlabel metal2 s 24950 0 25006 480 6 chany_bottom_out[17]
port 75 nsew default tristate
rlabel metal2 s 25594 0 25650 480 6 chany_bottom_out[18]
port 76 nsew default tristate
rlabel metal2 s 26238 0 26294 480 6 chany_bottom_out[19]
port 77 nsew default tristate
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_out[1]
port 78 nsew default tristate
rlabel metal2 s 15198 0 15254 480 6 chany_bottom_out[2]
port 79 nsew default tristate
rlabel metal2 s 15842 0 15898 480 6 chany_bottom_out[3]
port 80 nsew default tristate
rlabel metal2 s 16486 0 16542 480 6 chany_bottom_out[4]
port 81 nsew default tristate
rlabel metal2 s 17130 0 17186 480 6 chany_bottom_out[5]
port 82 nsew default tristate
rlabel metal2 s 17774 0 17830 480 6 chany_bottom_out[6]
port 83 nsew default tristate
rlabel metal2 s 18418 0 18474 480 6 chany_bottom_out[7]
port 84 nsew default tristate
rlabel metal2 s 19154 0 19210 480 6 chany_bottom_out[8]
port 85 nsew default tristate
rlabel metal2 s 19798 0 19854 480 6 chany_bottom_out[9]
port 86 nsew default tristate
rlabel metal2 s 10506 27520 10562 28000 6 prog_clk
port 87 nsew default input
rlabel metal3 s 27520 280 28000 400 6 right_bottom_grid_pin_34_
port 88 nsew default input
rlabel metal3 s 27520 824 28000 944 6 right_bottom_grid_pin_35_
port 89 nsew default input
rlabel metal3 s 27520 1368 28000 1488 6 right_bottom_grid_pin_36_
port 90 nsew default input
rlabel metal3 s 27520 1912 28000 2032 6 right_bottom_grid_pin_37_
port 91 nsew default input
rlabel metal3 s 27520 2456 28000 2576 6 right_bottom_grid_pin_38_
port 92 nsew default input
rlabel metal3 s 27520 3136 28000 3256 6 right_bottom_grid_pin_39_
port 93 nsew default input
rlabel metal3 s 27520 3680 28000 3800 6 right_bottom_grid_pin_40_
port 94 nsew default input
rlabel metal3 s 27520 4224 28000 4344 6 right_bottom_grid_pin_41_
port 95 nsew default input
rlabel metal3 s 27520 27616 28000 27736 6 right_top_grid_pin_1_
port 96 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 VPWR
port 97 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 VGND
port 98 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
