VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tie_array
  CLASS BLOCK ;
  FOREIGN tie_array ;
  ORIGIN 0.000 0.000 ;
  SIZE 52.300 BY 57.360 ;
  PIN x[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 0.020 0.000 0.300 2.400 ;
    END
  END x[0]
  PIN x[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 7.380 0.000 7.660 2.400 ;
    END
  END x[1]
  PIN x[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 14.740 0.000 15.020 2.400 ;
    END
  END x[2]
  PIN x[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 22.100 0.000 22.380 2.400 ;
    END
  END x[3]
  PIN x[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 29.920 0.000 30.200 2.400 ;
    END
  END x[4]
  PIN x[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 37.280 0.000 37.560 2.400 ;
    END
  END x[5]
  PIN x[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 44.640 0.000 44.920 2.400 ;
    END
  END x[6]
  PIN x[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 52.000 0.000 52.280 2.400 ;
    END
  END x[7]
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.130 10.640 10.730 57.360 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 17.290 10.640 18.890 57.360 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.770 10.795 50.530 57.205 ;
      LAYER met1 ;
        RECT 0.000 10.640 52.300 57.360 ;
      LAYER met2 ;
        RECT 0.030 2.680 52.270 57.360 ;
        RECT 0.580 2.400 7.100 2.680 ;
        RECT 7.940 2.400 14.460 2.680 ;
        RECT 15.300 2.400 21.820 2.680 ;
        RECT 22.660 2.400 29.640 2.680 ;
        RECT 30.480 2.400 37.000 2.680 ;
        RECT 37.840 2.400 44.360 2.680 ;
        RECT 45.200 2.400 51.720 2.680 ;
      LAYER met3 ;
        RECT 9.130 10.715 43.370 57.285 ;
      LAYER met4 ;
        RECT 25.450 10.640 43.370 57.360 ;
  END
END tie_array
END LIBRARY

