* NGSPICE file created from sb_0__1_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor4_4 abstract view
.subckt scs8hd_nor4_4 A B C D Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

.subckt sb_0__1_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] bottom_left_grid_pin_11_ bottom_left_grid_pin_13_ bottom_left_grid_pin_15_
+ bottom_left_grid_pin_1_ bottom_left_grid_pin_3_ bottom_left_grid_pin_5_ bottom_left_grid_pin_7_
+ bottom_left_grid_pin_9_ bottom_right_grid_pin_11_ chanx_right_in[0] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_out[0] chanx_right_out[1] chanx_right_out[2]
+ chanx_right_out[3] chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7]
+ chanx_right_out[8] chany_bottom_in[0] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_out[0] chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3]
+ chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7]
+ chany_bottom_out[8] chany_top_in[0] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_out[0] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4]
+ chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8] data_in enable
+ right_bottom_grid_pin_12_ right_top_grid_pin_10_ top_left_grid_pin_11_ top_left_grid_pin_13_
+ top_left_grid_pin_15_ top_left_grid_pin_1_ top_left_grid_pin_3_ top_left_grid_pin_5_
+ top_left_grid_pin_7_ top_left_grid_pin_9_ top_right_grid_pin_11_ vpwr vgnd
Xmem_right_track_12.LATCH_1_.latch data_in _067_/A _133_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_188 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[4] mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_115 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__113__B _113_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_3_ mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_192 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_258 vpwr vgnd scs8hd_fill_2
XFILLER_27_236 vpwr vgnd scs8hd_fill_2
XFILLER_12_32 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB _102_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _067_/A mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_12_98 vpwr vgnd scs8hd_fill_2
XFILLER_37_62 vgnd vpwr scs8hd_decap_12
XFILLER_33_239 vgnd vpwr scs8hd_decap_4
XANTENNA__108__B _105_/B vgnd vpwr scs8hd_diode_2
XANTENNA__124__A _094_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _146_/HI _062_/Y mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _140_/HI mem_bottom_track_17.LATCH_2_.latch/Q
+ mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_062_ _062_/A _062_/Y vgnd vpwr scs8hd_inv_8
X_131_ _135_/A address[6] _132_/C _135_/D _131_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_2_165 vpwr vgnd scs8hd_fill_2
XFILLER_2_110 vpwr vgnd scs8hd_fill_2
XANTENNA__110__C _110_/C vgnd vpwr scs8hd_diode_2
XFILLER_9_44 vpwr vgnd scs8hd_fill_2
XANTENNA__119__A _076_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _165_/A vgnd vpwr scs8hd_inv_1
Xmem_bottom_track_17.LATCH_2_.latch data_in mem_bottom_track_17.LATCH_2_.latch/Q _122_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_11_253 vpwr vgnd scs8hd_fill_2
XFILLER_11_264 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB _082_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_235 vgnd vpwr scs8hd_decap_3
X_114_ _080_/B _113_/B _114_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_22_7 vgnd vpwr scs8hd_decap_12
XANTENNA__121__B _119_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_6_.scs8hd_inv_1 bottom_left_grid_pin_7_ mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_top_track_0.LATCH_4_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_4_238 vgnd vpwr scs8hd_decap_6
XFILLER_20_32 vgnd vpwr scs8hd_decap_12
XFILLER_28_172 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[6] mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_23 vgnd vpwr scs8hd_decap_8
XANTENNA__116__B _113_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_56 vgnd vpwr scs8hd_decap_3
XANTENNA__132__A _135_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_172 vpwr vgnd scs8hd_fill_2
XFILLER_13_3 vgnd vpwr scs8hd_decap_12
Xmem_right_track_8.LATCH_1_.latch data_in _069_/A _135_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_175 vpwr vgnd scs8hd_fill_2
XFILLER_17_109 vgnd vpwr scs8hd_decap_3
XFILLER_40_178 vgnd vpwr scs8hd_decap_12
XFILLER_25_197 vgnd vpwr scs8hd_decap_4
XFILLER_31_86 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ _064_/A mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_0_263 vgnd vpwr scs8hd_decap_12
XFILLER_31_123 vgnd vpwr scs8hd_decap_3
XANTENNA__127__A _135_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_175 vgnd vpwr scs8hd_decap_3
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _066_/Y vgnd
+ vpwr scs8hd_diode_2
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _140_/HI vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _143_/HI _068_/Y mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_9_149 vpwr vgnd scs8hd_fill_2
XFILLER_13_178 vgnd vpwr scs8hd_decap_3
Xmux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_57 vpwr vgnd scs8hd_fill_2
XFILLER_36_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_3_.scs8hd_inv_1 chanx_right_in[1] mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _147_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
XFILLER_12_77 vpwr vgnd scs8hd_fill_2
XFILLER_37_74 vgnd vpwr scs8hd_decap_12
XFILLER_18_215 vgnd vpwr scs8hd_decap_3
XFILLER_18_248 vgnd vpwr scs8hd_decap_4
XFILLER_5_141 vgnd vpwr scs8hd_fill_1
XFILLER_5_163 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__124__B _119_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_32_251 vgnd vpwr scs8hd_decap_12
X_130_ _135_/A address[6] _138_/C address[0] _130_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_23_87 vpwr vgnd scs8hd_fill_2
X_061_ _061_/A _061_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_199 vpwr vgnd scs8hd_fill_2
XFILLER_2_144 vpwr vgnd scs8hd_fill_2
XFILLER_0_58 vpwr vgnd scs8hd_fill_2
XANTENNA__119__B _119_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_2_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_78 vgnd vpwr scs8hd_decap_3
XANTENNA__135__A _135_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A top_left_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
XFILLER_20_254 vgnd vpwr scs8hd_decap_12
XFILLER_20_243 vpwr vgnd scs8hd_fill_2
XFILLER_18_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_214 vgnd vpwr scs8hd_decap_6
XFILLER_11_276 vgnd vpwr scs8hd_fill_1
X_113_ _078_/B _113_/B _113_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_258 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _068_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ _072_/A mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_29_118 vpwr vgnd scs8hd_fill_2
XFILLER_37_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A bottom_right_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_206 vgnd vpwr scs8hd_decap_4
XFILLER_20_44 vgnd vpwr scs8hd_decap_3
XFILLER_20_88 vpwr vgnd scs8hd_fill_2
XFILLER_29_75 vgnd vpwr scs8hd_decap_12
XFILLER_6_46 vgnd vpwr scs8hd_fill_1
XANTENNA__132__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_19_184 vgnd vpwr scs8hd_decap_4
XFILLER_19_151 vgnd vpwr scs8hd_decap_4
XFILLER_34_198 vgnd vpwr scs8hd_decap_3
XFILLER_34_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A bottom_left_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_154 vpwr vgnd scs8hd_fill_2
XFILLER_15_33 vgnd vpwr scs8hd_fill_1
XFILLER_15_88 vpwr vgnd scs8hd_fill_2
XFILLER_31_98 vgnd vpwr scs8hd_decap_12
XFILLER_0_242 vgnd vpwr scs8hd_decap_6
XFILLER_0_231 vgnd vpwr scs8hd_decap_4
XFILLER_0_275 vpwr vgnd scs8hd_fill_2
XFILLER_31_157 vpwr vgnd scs8hd_fill_2
XFILLER_31_135 vpwr vgnd scs8hd_fill_2
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__B address[6] vgnd vpwr scs8hd_diode_2
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_143 vgnd vpwr scs8hd_decap_8
XFILLER_16_187 vpwr vgnd scs8hd_fill_2
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__053__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _059_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_9 vpwr vgnd scs8hd_fill_2
XFILLER_26_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_102 vpwr vgnd scs8hd_fill_2
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _066_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.INVTX1_2_.scs8hd_inv_1_A right_bottom_grid_pin_12_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A bottom_left_grid_pin_3_ vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _161_/A vgnd vpwr scs8hd_inv_1
XFILLER_36_227 vgnd vpwr scs8hd_decap_12
XANTENNA__138__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_8_172 vgnd vpwr scs8hd_decap_4
XFILLER_12_190 vgnd vpwr scs8hd_decap_4
XFILLER_27_205 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_127 vgnd vpwr scs8hd_decap_4
XFILLER_10_149 vpwr vgnd scs8hd_fill_2
XFILLER_12_56 vpwr vgnd scs8hd_fill_2
XFILLER_12_89 vgnd vpwr scs8hd_fill_1
XFILLER_37_86 vgnd vpwr scs8hd_decap_12
XFILLER_26_260 vgnd vpwr scs8hd_decap_12
XFILLER_18_227 vpwr vgnd scs8hd_fill_2
XFILLER_5_153 vgnd vpwr scs8hd_decap_4
XFILLER_5_175 vgnd vpwr scs8hd_decap_3
XFILLER_5_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_263 vgnd vpwr scs8hd_decap_12
XFILLER_24_219 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB _137_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_219 vpwr vgnd scs8hd_fill_2
XFILLER_23_66 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_3 vgnd vpwr scs8hd_decap_12
X_060_ _060_/A _060_/Y vgnd vpwr scs8hd_inv_8
XFILLER_0_15 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_37 vpwr vgnd scs8hd_fill_2
XFILLER_14_230 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
XANTENNA__135__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
XFILLER_20_266 vgnd vpwr scs8hd_decap_8
XANTENNA__061__A _061_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_44 vgnd vpwr scs8hd_decap_8
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_112_ _076_/A _113_/B _112_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _061_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__056__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_29_10 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_track_1.LATCH_5_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _059_/A mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_4_218 vpwr vgnd scs8hd_fill_2
XFILLER_20_67 vgnd vpwr scs8hd_decap_6
XFILLER_29_87 vgnd vpwr scs8hd_decap_4
XFILLER_3_262 vgnd vpwr scs8hd_decap_12
XFILLER_3_240 vgnd vpwr scs8hd_decap_4
XANTENNA__132__C _132_/C vgnd vpwr scs8hd_diode_2
XFILLER_34_166 vgnd vpwr scs8hd_decap_12
XFILLER_31_11 vgnd vpwr scs8hd_decap_12
XFILLER_31_147 vgnd vpwr scs8hd_fill_1
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__C _075_/C vgnd vpwr scs8hd_diode_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_125 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_22_169 vpwr vgnd scs8hd_fill_2
Xmem_right_track_4.LATCH_1_.latch data_in _061_/A _127_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB _126_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_44 vgnd vpwr scs8hd_decap_12
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_114 vpwr vgnd scs8hd_fill_2
XFILLER_13_136 vgnd vpwr scs8hd_decap_4
Xmux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _063_/Y mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_3_15 vgnd vpwr scs8hd_decap_12
XFILLER_36_239 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.INVTX1_4_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__138__B _138_/B vgnd vpwr scs8hd_diode_2
XANTENNA__154__A _154_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_14.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__064__A _064_/A vgnd vpwr scs8hd_diode_2
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XFILLER_37_98 vgnd vpwr scs8hd_decap_8
XFILLER_26_272 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_132 vgnd vpwr scs8hd_decap_3
Xmem_top_track_0.LATCH_0_.latch data_in mem_top_track_0.LATCH_0_.latch/Q _086_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_track_17.LATCH_3_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_231 vpwr vgnd scs8hd_fill_2
XFILLER_23_220 vpwr vgnd scs8hd_fill_2
XANTENNA__059__A _059_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_0_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__135__C _096_/C vgnd vpwr scs8hd_diode_2
Xmux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _065_/A mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _145_/HI _060_/Y mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_67 vgnd vpwr scs8hd_decap_4
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
X_111_ address[5] _138_/B _132_/C _113_/B vgnd vpwr scs8hd_or3_4
XANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_38_109 vgnd vpwr scs8hd_decap_12
XANTENNA__162__A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_6_260 vgnd vpwr scs8hd_decap_12
XFILLER_37_120 vpwr vgnd scs8hd_fill_2
XANTENNA__072__A _072_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_14.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_99 vpwr vgnd scs8hd_fill_2
XFILLER_28_131 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _148_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__132__D address[0] vgnd vpwr scs8hd_diode_2
XFILLER_3_274 vgnd vpwr scs8hd_decap_3
XFILLER_20_7 vgnd vpwr scs8hd_decap_12
XANTENNA__157__A _157_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_178 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _144_/HI _071_/Y mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_track_1.LATCH_2_.latch data_in mem_bottom_track_1.LATCH_2_.latch/Q _107_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_25_123 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_8.LATCH_3_.latch_SLEEPB _091_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__067__A _067_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_57 vpwr vgnd scs8hd_fill_2
XFILLER_31_23 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_222 vgnd vpwr scs8hd_fill_1
XFILLER_0_200 vgnd vpwr scs8hd_fill_1
XFILLER_16_167 vpwr vgnd scs8hd_fill_2
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__D _135_/D vgnd vpwr scs8hd_diode_2
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_259 vpwr vgnd scs8hd_fill_2
XFILLER_39_248 vpwr vgnd scs8hd_fill_2
XFILLER_39_237 vgnd vpwr scs8hd_decap_6
XFILLER_11_3 vgnd vpwr scs8hd_decap_12
XFILLER_22_104 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_181 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_56 vgnd vpwr scs8hd_decap_12
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_9_119 vgnd vpwr scs8hd_decap_3
XFILLER_13_159 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_27 vgnd vpwr scs8hd_decap_12
XANTENNA__138__C _138_/C vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ _062_/A mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__170__A _170_/A vgnd vpwr scs8hd_diode_2
XANTENNA__080__A _080_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_37_11 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_16.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_207 vgnd vpwr scs8hd_decap_6
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
Xmux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _142_/HI _066_/Y mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XANTENNA__165__A _165_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_243 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__075__A address[5] vgnd vpwr scs8hd_diode_2
Xmux_right_track_12.INVTX1_0_.scs8hd_inv_1 chany_top_in[6] mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_169 vpwr vgnd scs8hd_fill_2
XFILLER_2_114 vpwr vgnd scs8hd_fill_2
XFILLER_9_15 vgnd vpwr scs8hd_decap_12
XFILLER_9_48 vgnd vpwr scs8hd_decap_3
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
XANTENNA__135__D _135_/D vgnd vpwr scs8hd_diode_2
XFILLER_20_202 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ _070_/Y mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_9.INVTX1_3_.scs8hd_inv_1 chanx_right_in[3] mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
X_110_ _110_/A _110_/B _110_/C _132_/C vgnd vpwr scs8hd_or3_4
XFILLER_11_213 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _065_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XFILLER_6_272 vgnd vpwr scs8hd_decap_3
Xmux_top_track_16.INVTX1_4_.scs8hd_inv_1 chanx_right_in[3] mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_82 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_176 vgnd vpwr scs8hd_decap_4
XFILLER_28_154 vgnd vpwr scs8hd_decap_6
XFILLER_3_253 vpwr vgnd scs8hd_fill_2
XFILLER_19_176 vpwr vgnd scs8hd_fill_2
XANTENNA__173__A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_25_113 vpwr vgnd scs8hd_fill_2
XFILLER_40_105 vgnd vpwr scs8hd_decap_12
XFILLER_31_35 vgnd vpwr scs8hd_decap_12
XFILLER_25_179 vpwr vgnd scs8hd_fill_2
XANTENNA__083__A address[1] vgnd vpwr scs8hd_diode_2
Xmux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ _068_/A mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_15_36 vpwr vgnd scs8hd_fill_2
XFILLER_0_212 vgnd vpwr scs8hd_decap_3
Xmux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__168__A chany_top_in[0] vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_1_ mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__078__A _080_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_68 vgnd vpwr scs8hd_decap_12
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XFILLER_21_160 vgnd vpwr scs8hd_decap_4
XFILLER_3_39 vgnd vpwr scs8hd_decap_3
XANTENNA__138__D address[0] vgnd vpwr scs8hd_diode_2
XFILLER_16_90 vpwr vgnd scs8hd_fill_2
XFILLER_8_131 vgnd vpwr scs8hd_decap_3
XFILLER_8_164 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A top_right_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_219 vpwr vgnd scs8hd_fill_2
XFILLER_10_108 vpwr vgnd scs8hd_fill_2
XFILLER_12_15 vgnd vpwr scs8hd_decap_12
XANTENNA__080__B _080_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_9 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_23 vgnd vpwr scs8hd_decap_12
XFILLER_26_230 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[4] mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_top_track_8.LATCH_1_.latch data_in mem_top_track_8.LATCH_1_.latch/Q _093_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_101 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _067_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_32_211 vgnd vpwr scs8hd_decap_3
Xmux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_241 vgnd vpwr scs8hd_decap_3
XFILLER_17_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_93 vgnd vpwr scs8hd_fill_1
XANTENNA__075__B address[6] vgnd vpwr scs8hd_diode_2
XANTENNA__091__A _080_/B vgnd vpwr scs8hd_diode_2
XFILLER_2_148 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_1.LATCH_3_.latch_SLEEPB _106_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _062_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__176__A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_247 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_1.INVTX1_6_.scs8hd_inv_1 bottom_left_grid_pin_5_ mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XFILLER_11_236 vpwr vgnd scs8hd_fill_2
XANTENNA__086__A _080_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_169_ _169_/A chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
Xmux_right_track_10.INVTX1_0_.scs8hd_inv_1 chany_top_in[5] mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB _097_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_39 vgnd vpwr scs8hd_decap_4
XFILLER_3_232 vpwr vgnd scs8hd_fill_2
XFILLER_3_210 vpwr vgnd scs8hd_fill_2
XFILLER_19_100 vpwr vgnd scs8hd_fill_2
XFILLER_19_111 vpwr vgnd scs8hd_fill_2
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
Xmem_bottom_track_9.LATCH_3_.latch data_in mem_bottom_track_9.LATCH_3_.latch/Q _114_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_40_117 vgnd vpwr scs8hd_decap_12
XFILLER_25_158 vpwr vgnd scs8hd_fill_2
XFILLER_15_15 vgnd vpwr scs8hd_decap_12
XFILLER_31_47 vgnd vpwr scs8hd_decap_12
XANTENNA__083__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_103 vgnd vpwr scs8hd_decap_4
XFILLER_31_139 vgnd vpwr scs8hd_decap_8
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_91 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _060_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_39_228 vpwr vgnd scs8hd_fill_2
XPHY_0 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_38_250 vgnd vpwr scs8hd_decap_12
XANTENNA__078__B _078_/B vgnd vpwr scs8hd_diode_2
XANTENNA__094__A _094_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_106 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _064_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_110 vpwr vgnd scs8hd_fill_2
XFILLER_8_154 vgnd vpwr scs8hd_fill_1
XFILLER_8_198 vpwr vgnd scs8hd_fill_2
XFILLER_35_220 vgnd vpwr scs8hd_decap_12
XFILLER_12_27 vgnd vpwr scs8hd_decap_4
Xmux_right_track_12.tap_buf4_0_.scs8hd_inv_1 mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ _154_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_track_17.LATCH_4_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_35 vgnd vpwr scs8hd_decap_12
Xmem_top_track_16.LATCH_3_.latch data_in mem_top_track_16.LATCH_3_.latch/Q _099_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__089__A _076_/A vgnd vpwr scs8hd_diode_2
XFILLER_41_245 vgnd vpwr scs8hd_decap_12
XFILLER_17_220 vpwr vgnd scs8hd_fill_2
XFILLER_17_275 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ _061_/Y mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_23_245 vgnd vpwr scs8hd_decap_12
XFILLER_23_59 vpwr vgnd scs8hd_fill_2
XFILLER_23_15 vgnd vpwr scs8hd_decap_12
XANTENNA__075__C _075_/C vgnd vpwr scs8hd_diode_2
XANTENNA__091__B _091_/B vgnd vpwr scs8hd_diode_2
XFILLER_2_127 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_0_19 vgnd vpwr scs8hd_fill_1
XFILLER_14_201 vpwr vgnd scs8hd_fill_2
XFILLER_9_39 vpwr vgnd scs8hd_fill_2
Xmux_right_track_6.INVTX1_1_.scs8hd_inv_1 chany_top_in[8] mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_6 vpwr vgnd scs8hd_fill_2
XFILLER_1_193 vpwr vgnd scs8hd_fill_2
XFILLER_20_226 vpwr vgnd scs8hd_fill_2
XANTENNA__086__B _094_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _062_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_230 vgnd vpwr scs8hd_decap_4
X_168_ chany_top_in[0] chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
X_099_ _080_/B _099_/B _099_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_27_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_123 vgnd vpwr scs8hd_decap_12
XFILLER_1_40 vpwr vgnd scs8hd_fill_2
XFILLER_1_62 vgnd vpwr scs8hd_decap_4
XFILLER_1_95 vpwr vgnd scs8hd_fill_2
XFILLER_29_58 vgnd vpwr scs8hd_decap_3
XFILLER_29_14 vgnd vpwr scs8hd_decap_12
XFILLER_28_145 vgnd vpwr scs8hd_decap_8
XFILLER_28_112 vpwr vgnd scs8hd_fill_2
XFILLER_28_189 vgnd vpwr scs8hd_decap_12
XANTENNA__097__A _076_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_123 vpwr vgnd scs8hd_fill_2
XFILLER_19_134 vpwr vgnd scs8hd_fill_2
XFILLER_40_129 vgnd vpwr scs8hd_decap_12
XFILLER_25_137 vpwr vgnd scs8hd_fill_2
XFILLER_15_27 vgnd vpwr scs8hd_decap_6
XFILLER_31_59 vpwr vgnd scs8hd_fill_2
XANTENNA__083__C _135_/D vgnd vpwr scs8hd_diode_2
XFILLER_0_203 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_17.LATCH_3_.latch data_in mem_bottom_track_17.LATCH_3_.latch/Q _121_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_31_118 vpwr vgnd scs8hd_fill_2
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_30_140 vpwr vgnd scs8hd_fill_2
XFILLER_38_262 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.tap_buf4_0_.scs8hd_inv_1 mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ _157_/A vgnd vpwr scs8hd_inv_1
XFILLER_26_15 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.INVTX1_1_.scs8hd_inv_1 chany_top_in[6] mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_140 vpwr vgnd scs8hd_fill_2
XANTENNA__094__B _091_/B vgnd vpwr scs8hd_diode_2
XFILLER_13_118 vpwr vgnd scs8hd_fill_2
XFILLER_21_184 vgnd vpwr scs8hd_decap_4
Xmux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _067_/Y mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_32_80 vgnd vpwr scs8hd_decap_12
XFILLER_12_140 vpwr vgnd scs8hd_fill_2
XFILLER_12_173 vpwr vgnd scs8hd_fill_2
XFILLER_35_232 vgnd vpwr scs8hd_decap_12
XANTENNA__089__B _091_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_47 vgnd vpwr scs8hd_decap_12
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_26_243 vgnd vpwr scs8hd_decap_8
XFILLER_41_257 vgnd vpwr scs8hd_decap_12
XFILLER_5_114 vpwr vgnd scs8hd_fill_2
XFILLER_17_254 vpwr vgnd scs8hd_fill_2
XFILLER_4_180 vgnd vpwr scs8hd_decap_3
XFILLER_4_84 vpwr vgnd scs8hd_fill_2
XFILLER_23_257 vgnd vpwr scs8hd_decap_12
XFILLER_23_235 vgnd vpwr scs8hd_decap_8
XFILLER_23_224 vpwr vgnd scs8hd_fill_2
XFILLER_23_27 vgnd vpwr scs8hd_decap_12
Xmux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ _060_/A mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_2_.latch/Q mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB _132_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_213 vgnd vpwr scs8hd_fill_1
Xmux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_track_0.LATCH_5_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_9.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XFILLER_11_249 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_80 vgnd vpwr scs8hd_decap_12
X_098_ _078_/B _099_/B _098_/Y vgnd vpwr scs8hd_nor2_4
X_167_ chany_top_in[1] chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_37_135 vgnd vpwr scs8hd_decap_12
Xmux_right_track_4.INVTX1_1_.scs8hd_inv_1 chany_top_in[7] mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_26 vgnd vpwr scs8hd_decap_12
XFILLER_28_135 vgnd vpwr scs8hd_fill_1
XANTENNA__097__B _099_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_190 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ _064_/Y mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB _094_/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_50 vgnd vpwr scs8hd_fill_1
XFILLER_34_105 vgnd vpwr scs8hd_decap_12
XFILLER_19_157 vpwr vgnd scs8hd_fill_2
XFILLER_19_70 vpwr vgnd scs8hd_fill_2
XFILLER_33_193 vpwr vgnd scs8hd_fill_2
XFILLER_33_171 vgnd vpwr scs8hd_decap_12
XFILLER_0_259 vpwr vgnd scs8hd_fill_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_116 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _150_/HI mem_top_track_16.LATCH_2_.latch/Q
+ mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_208 vgnd vpwr scs8hd_decap_12
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_15_160 vpwr vgnd scs8hd_fill_2
XFILLER_15_171 vpwr vgnd scs8hd_fill_2
XFILLER_15_193 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_152 vgnd vpwr scs8hd_fill_1
XFILLER_7_40 vpwr vgnd scs8hd_fill_2
XFILLER_7_62 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_274 vgnd vpwr scs8hd_fill_1
XFILLER_26_27 vgnd vpwr scs8hd_decap_4
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_8.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _068_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_16_71 vgnd vpwr scs8hd_decap_8
XFILLER_16_82 vgnd vpwr scs8hd_decap_8
XFILLER_16_93 vgnd vpwr scs8hd_decap_3
XFILLER_8_145 vgnd vpwr scs8hd_decap_6
XFILLER_8_178 vgnd vpwr scs8hd_decap_3
XFILLER_12_130 vgnd vpwr scs8hd_fill_1
XFILLER_12_152 vgnd vpwr scs8hd_fill_1
Xmux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ _066_/A mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A top_left_grid_pin_7_ vgnd vpwr scs8hd_diode_2
XFILLER_37_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_269 vgnd vpwr scs8hd_decap_8
XFILLER_5_137 vgnd vpwr scs8hd_decap_4
XFILLER_5_159 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_233 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_4_192 vgnd vpwr scs8hd_decap_4
XFILLER_4_74 vpwr vgnd scs8hd_fill_2
XFILLER_23_269 vgnd vpwr scs8hd_decap_8
XFILLER_23_39 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_247 vgnd vpwr scs8hd_decap_12
XFILLER_13_83 vpwr vgnd scs8hd_fill_2
XFILLER_1_162 vpwr vgnd scs8hd_fill_2
XFILLER_38_80 vgnd vpwr scs8hd_decap_12
Xmux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ _072_/Y mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_206 vgnd vpwr scs8hd_decap_6
XFILLER_9_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A bottom_left_grid_pin_5_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _066_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
XFILLER_11_217 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.INVTX1_1_.scs8hd_inv_1 top_left_grid_pin_11_ mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_6 vpwr vgnd scs8hd_fill_2
XFILLER_24_93 vgnd vpwr scs8hd_decap_4
XFILLER_6_210 vgnd vpwr scs8hd_decap_4
X_166_ chany_top_in[2] chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
X_097_ _076_/A _099_/B _097_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_243 vpwr vgnd scs8hd_fill_2
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
XFILLER_37_147 vgnd vpwr scs8hd_decap_12
XFILLER_1_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.LATCH_4_.latch_SLEEPB _113_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _072_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_29_38 vgnd vpwr scs8hd_decap_12
XFILLER_34_117 vgnd vpwr scs8hd_decap_12
X_149_ _149_/HI _149_/LO vgnd vpwr scs8hd_conb_1
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
XFILLER_25_117 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_191 vpwr vgnd scs8hd_fill_2
XFILLER_0_249 vgnd vpwr scs8hd_decap_6
XFILLER_0_238 vpwr vgnd scs8hd_fill_2
XFILLER_0_227 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_194 vpwr vgnd scs8hd_fill_2
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A bottom_left_grid_pin_9_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_30_164 vpwr vgnd scs8hd_fill_2
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_30_186 vgnd vpwr scs8hd_decap_12
XFILLER_7_74 vpwr vgnd scs8hd_fill_2
XFILLER_7_85 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _141_/HI mem_bottom_track_9.LATCH_2_.latch/Q
+ mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_21_175 vpwr vgnd scs8hd_fill_2
XFILLER_21_153 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_253 vpwr vgnd scs8hd_fill_2
XFILLER_29_242 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _061_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_168 vpwr vgnd scs8hd_fill_2
XFILLER_12_186 vpwr vgnd scs8hd_fill_2
XFILLER_35_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _068_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_26_212 vpwr vgnd scs8hd_fill_2
XFILLER_26_201 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_201 vpwr vgnd scs8hd_fill_2
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB _109_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_215 vgnd vpwr scs8hd_decap_6
XFILLER_14_259 vgnd vpwr scs8hd_decap_12
XFILLER_13_73 vpwr vgnd scs8hd_fill_2
XANTENNA__100__A _082_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_2_.scs8hd_inv_1 top_left_grid_pin_15_ mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_18 vgnd vpwr scs8hd_decap_12
Xmux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _059_/Y mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB _100_/Y vgnd vpwr scs8hd_diode_2
X_165_ _165_/A chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_40_93 vgnd vpwr scs8hd_decap_12
X_096_ address[5] address[6] _096_/C _099_/B vgnd vpwr scs8hd_or3_4
XFILLER_37_159 vgnd vpwr scs8hd_decap_12
XFILLER_1_10 vgnd vpwr scs8hd_decap_12
XFILLER_20_19 vgnd vpwr scs8hd_decap_12
Xmem_top_track_0.LATCH_1_.latch data_in mem_top_track_0.LATCH_1_.latch/Q _084_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_258 vpwr vgnd scs8hd_fill_2
XFILLER_3_236 vpwr vgnd scs8hd_fill_2
XFILLER_3_214 vgnd vpwr scs8hd_decap_3
XFILLER_10_85 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _063_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_83 vpwr vgnd scs8hd_fill_2
XFILLER_19_104 vpwr vgnd scs8hd_fill_2
XFILLER_19_115 vpwr vgnd scs8hd_fill_2
XFILLER_34_129 vgnd vpwr scs8hd_decap_12
X_148_ _148_/HI _148_/LO vgnd vpwr scs8hd_conb_1
XFILLER_25_3 vgnd vpwr scs8hd_decap_12
X_079_ _079_/A address[2] _135_/D _080_/B vgnd vpwr scs8hd_or3_4
XANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_33_184 vgnd vpwr scs8hd_decap_6
XFILLER_24_162 vpwr vgnd scs8hd_fill_2
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_62 vgnd vpwr scs8hd_decap_3
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_95 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB _078_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_154 vgnd vpwr scs8hd_fill_1
XFILLER_30_110 vgnd vpwr scs8hd_decap_4
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_30_198 vgnd vpwr scs8hd_decap_12
XFILLER_7_53 vpwr vgnd scs8hd_fill_2
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_110 vpwr vgnd scs8hd_fill_2
XFILLER_29_221 vpwr vgnd scs8hd_fill_2
XFILLER_8_114 vpwr vgnd scs8hd_fill_2
XFILLER_12_154 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB _123_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__103__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_35_257 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_track_17.LATCH_4_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_track_1.LATCH_3_.latch data_in mem_bottom_track_1.LATCH_3_.latch/Q _106_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_32_227 vgnd vpwr scs8hd_decap_12
Xmux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ _065_/Y mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_205 vpwr vgnd scs8hd_fill_2
XFILLER_14_205 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
Xmem_right_track_14.LATCH_0_.latch data_in _072_/A _138_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_120 vpwr vgnd scs8hd_fill_2
XFILLER_38_93 vgnd vpwr scs8hd_decap_12
XFILLER_1_197 vpwr vgnd scs8hd_fill_2
XFILLER_1_175 vpwr vgnd scs8hd_fill_2
XANTENNA__100__B _099_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_231 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_5_.scs8hd_inv_1 chanx_right_in[7] mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_84 vgnd vpwr scs8hd_decap_8
X_164_ chany_top_in[4] chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
X_095_ _110_/A address[3] _110_/C _096_/C vgnd vpwr scs8hd_or3_4
XFILLER_1_22 vgnd vpwr scs8hd_decap_4
XFILLER_1_66 vgnd vpwr scs8hd_fill_1
XFILLER_1_99 vpwr vgnd scs8hd_fill_2
XANTENNA__111__A address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_28_127 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_12.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_160 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_62 vgnd vpwr scs8hd_fill_1
XFILLER_19_138 vpwr vgnd scs8hd_fill_2
XFILLER_27_193 vpwr vgnd scs8hd_fill_2
X_078_ _080_/A _078_/B _078_/Y vgnd vpwr scs8hd_nor2_4
X_147_ _147_/HI _147_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__106__A _080_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_270 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_218 vpwr vgnd scs8hd_fill_2
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_74 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_16.LATCH_3_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_15_130 vpwr vgnd scs8hd_fill_2
XFILLER_30_144 vgnd vpwr scs8hd_decap_8
Xmux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ _062_/Y mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_2_.latch/Q mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_199 vpwr vgnd scs8hd_fill_2
XFILLER_12_144 vpwr vgnd scs8hd_fill_2
XANTENNA__103__B _138_/B vgnd vpwr scs8hd_diode_2
XFILLER_35_269 vgnd vpwr scs8hd_decap_8
XFILLER_5_118 vpwr vgnd scs8hd_fill_2
XFILLER_32_239 vgnd vpwr scs8hd_decap_12
XFILLER_27_62 vgnd vpwr scs8hd_decap_12
XFILLER_27_51 vgnd vpwr scs8hd_decap_8
XFILLER_40_250 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB _130_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_151 vpwr vgnd scs8hd_fill_2
XFILLER_4_88 vpwr vgnd scs8hd_fill_2
XFILLER_4_55 vpwr vgnd scs8hd_fill_2
XFILLER_4_44 vgnd vpwr scs8hd_decap_8
XANTENNA__114__A _080_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_132 vgnd vpwr scs8hd_decap_3
XANTENNA__109__A _094_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_254 vpwr vgnd scs8hd_fill_2
XFILLER_9_265 vpwr vgnd scs8hd_fill_2
XFILLER_24_74 vgnd vpwr scs8hd_fill_1
X_163_ chany_top_in[5] chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
X_094_ _094_/A _091_/B _094_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__111__B _138_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _151_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_78 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_2_.latch data_in mem_top_track_8.LATCH_2_.latch/Q _092_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _067_/Y vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ _068_/Y mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_10_32 vgnd vpwr scs8hd_decap_12
XFILLER_10_54 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_62 vgnd vpwr scs8hd_decap_12
XANTENNA__106__B _105_/B vgnd vpwr scs8hd_diode_2
X_077_ address[1] _052_/Y address[0] _078_/B vgnd vpwr scs8hd_or3_4
X_146_ _146_/HI _146_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__122__A _082_/B vgnd vpwr scs8hd_diode_2
XFILLER_33_197 vgnd vpwr scs8hd_decap_4
XFILLER_25_109 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB _127_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_208 vpwr vgnd scs8hd_fill_2
XFILLER_24_120 vgnd vpwr scs8hd_decap_6
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_31 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_164 vpwr vgnd scs8hd_fill_2
XFILLER_15_175 vpwr vgnd scs8hd_fill_2
XFILLER_30_123 vgnd vpwr scs8hd_decap_3
XANTENNA__117__A _094_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_197 vgnd vpwr scs8hd_decap_4
X_129_ _135_/A address[6] _138_/C _135_/D _129_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_21_123 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_track_9.LATCH_3_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_245 vgnd vpwr scs8hd_decap_8
XFILLER_29_234 vgnd vpwr scs8hd_decap_8
XFILLER_8_127 vpwr vgnd scs8hd_fill_2
XFILLER_12_123 vgnd vpwr scs8hd_decap_4
Xmux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_2_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__103__C _096_/C vgnd vpwr scs8hd_diode_2
XFILLER_26_226 vpwr vgnd scs8hd_fill_2
XFILLER_26_215 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_9.LATCH_4_.latch data_in mem_bottom_track_9.LATCH_4_.latch/Q _113_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _142_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_237 vpwr vgnd scs8hd_fill_2
XFILLER_40_262 vgnd vpwr scs8hd_decap_12
XFILLER_27_74 vgnd vpwr scs8hd_decap_12
XFILLER_17_248 vgnd vpwr scs8hd_decap_4
XFILLER_17_259 vpwr vgnd scs8hd_fill_2
XANTENNA__114__B _113_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_196 vgnd vpwr scs8hd_fill_1
XFILLER_4_174 vgnd vpwr scs8hd_decap_4
XFILLER_4_163 vpwr vgnd scs8hd_fill_2
XFILLER_4_78 vgnd vpwr scs8hd_decap_4
XANTENNA__130__A _135_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _071_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_87 vpwr vgnd scs8hd_fill_2
XANTENNA__109__B _105_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_200 vpwr vgnd scs8hd_fill_2
XFILLER_13_240 vgnd vpwr scs8hd_decap_4
XFILLER_13_262 vgnd vpwr scs8hd_decap_12
XANTENNA__125__A address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_6_.scs8hd_inv_1 bottom_left_grid_pin_9_ mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _064_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB _116_/Y vgnd vpwr scs8hd_diode_2
X_162_ chany_top_in[6] chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
X_093_ _101_/A _091_/B _093_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_247 vpwr vgnd scs8hd_fill_2
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
Xmem_top_track_16.LATCH_4_.latch data_in mem_top_track_16.LATCH_4_.latch/Q _098_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__111__C _132_/C vgnd vpwr scs8hd_diode_2
XFILLER_1_57 vpwr vgnd scs8hd_fill_2
Xmem_right_track_10.LATCH_0_.latch data_in _066_/A _132_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_44 vgnd vpwr scs8hd_decap_6
XFILLER_10_88 vpwr vgnd scs8hd_fill_2
XFILLER_19_31 vgnd vpwr scs8hd_decap_12
XFILLER_19_53 vgnd vpwr scs8hd_decap_6
XFILLER_35_74 vgnd vpwr scs8hd_decap_12
XFILLER_27_173 vgnd vpwr scs8hd_decap_4
XFILLER_27_140 vpwr vgnd scs8hd_fill_2
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
X_145_ _145_/HI _145_/LO vgnd vpwr scs8hd_conb_1
X_076_ _076_/A _080_/A _076_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__122__B _119_/B vgnd vpwr scs8hd_diode_2
XFILLER_33_110 vgnd vpwr scs8hd_decap_12
XFILLER_18_195 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_198 vgnd vpwr scs8hd_decap_4
XFILLER_24_154 vgnd vpwr scs8hd_fill_1
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_43 vgnd vpwr scs8hd_decap_12
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_143 vpwr vgnd scs8hd_fill_2
XFILLER_30_168 vpwr vgnd scs8hd_fill_2
XFILLER_7_78 vpwr vgnd scs8hd_fill_2
XFILLER_7_89 vpwr vgnd scs8hd_fill_2
XANTENNA__133__A address[5] vgnd vpwr scs8hd_diode_2
X_128_ _135_/A address[6] _075_/C address[0] _128_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__117__B _113_/B vgnd vpwr scs8hd_diode_2
XFILLER_38_202 vgnd vpwr scs8hd_decap_12
XFILLER_23_3 vgnd vpwr scs8hd_decap_12
X_059_ _059_/A _059_/Y vgnd vpwr scs8hd_inv_8
Xmux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_179 vpwr vgnd scs8hd_fill_2
XFILLER_21_157 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _062_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_257 vgnd vpwr scs8hd_decap_12
XFILLER_12_102 vpwr vgnd scs8hd_fill_2
XFILLER_16_32 vpwr vgnd scs8hd_fill_2
XFILLER_16_54 vpwr vgnd scs8hd_fill_2
XANTENNA__128__A _135_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_161 vpwr vgnd scs8hd_fill_2
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _070_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_5_.latch_SLEEPB _089_/Y vgnd vpwr scs8hd_diode_2
XFILLER_27_86 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_17_216 vpwr vgnd scs8hd_fill_2
XFILLER_40_274 vgnd vpwr scs8hd_fill_1
XFILLER_27_97 vpwr vgnd scs8hd_fill_2
XFILLER_4_131 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__130__B address[6] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_17.LATCH_4_.latch data_in mem_bottom_track_17.LATCH_4_.latch/Q _120_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_77 vgnd vpwr scs8hd_decap_4
Xmem_right_track_6.LATCH_0_.latch data_in _064_/A _130_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__125__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_13_274 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__051__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_39_171 vgnd vpwr scs8hd_decap_12
XFILLER_24_32 vgnd vpwr scs8hd_decap_12
X_161_ _161_/A chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_6_226 vpwr vgnd scs8hd_fill_2
XFILLER_10_233 vpwr vgnd scs8hd_fill_2
XFILLER_10_244 vpwr vgnd scs8hd_fill_2
XFILLER_10_255 vgnd vpwr scs8hd_decap_12
X_092_ _082_/B _091_/B _092_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_108 vgnd vpwr scs8hd_decap_12
XFILLER_1_36 vpwr vgnd scs8hd_fill_2
XANTENNA__136__A _135_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _064_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_141 vgnd vpwr scs8hd_decap_12
XFILLER_28_108 vpwr vgnd scs8hd_fill_2
XFILLER_19_43 vgnd vpwr scs8hd_decap_4
XFILLER_19_87 vpwr vgnd scs8hd_fill_2
XFILLER_19_119 vgnd vpwr scs8hd_decap_3
XFILLER_35_86 vgnd vpwr scs8hd_decap_12
Xmux_right_track_12.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[7] mux_right_track_12.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
X_144_ _144_/HI _144_/LO vgnd vpwr scs8hd_conb_1
Xmux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _151_/HI mem_top_track_8.LATCH_2_.latch/Q
+ mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_075_ address[5] address[6] _075_/C _080_/A vgnd vpwr scs8hd_or3_4
Xmux_right_track_2.tap_buf4_0_.scs8hd_inv_1 mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ _159_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_6 vgnd vpwr scs8hd_decap_12
XFILLER_18_130 vpwr vgnd scs8hd_fill_2
XFILLER_18_174 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB _084_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_177 vgnd vpwr scs8hd_decap_8
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_9.INVTX1_5_.scs8hd_inv_1 bottom_left_grid_pin_1_ mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_55 vgnd vpwr scs8hd_decap_4
XPHY_8 vgnd vpwr scs8hd_decap_3
X_127_ _135_/A address[6] _075_/C _135_/D _127_/Y vgnd vpwr scs8hd_nor4_4
X_058_ enable _110_/C vgnd vpwr scs8hd_inv_8
XANTENNA_mem_bottom_track_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_13 vgnd vpwr scs8hd_decap_12
XFILLER_7_57 vpwr vgnd scs8hd_fill_2
XANTENNA__133__B _138_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_3 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _169_/A vgnd vpwr scs8hd_inv_1
Xmux_top_track_16.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[2] mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_136 vpwr vgnd scs8hd_fill_2
XFILLER_21_114 vpwr vgnd scs8hd_fill_2
XFILLER_29_269 vgnd vpwr scs8hd_decap_8
XFILLER_12_169 vpwr vgnd scs8hd_fill_2
XFILLER_16_99 vpwr vgnd scs8hd_fill_2
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XANTENNA__128__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_7_195 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ _060_/Y mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__054__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_4_143 vpwr vgnd scs8hd_fill_2
XANTENNA__130__C _138_/C vgnd vpwr scs8hd_diode_2
XFILLER_31_220 vgnd vpwr scs8hd_decap_12
XFILLER_14_209 vgnd vpwr scs8hd_decap_4
Xmux_top_track_0.INVTX1_2_.scs8hd_inv_1 top_left_grid_pin_13_ mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_14.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_220 vpwr vgnd scs8hd_fill_2
XFILLER_13_231 vpwr vgnd scs8hd_fill_2
XANTENNA__125__C _132_/C vgnd vpwr scs8hd_diode_2
XFILLER_9_213 vpwr vgnd scs8hd_fill_2
XFILLER_9_235 vgnd vpwr scs8hd_decap_3
XFILLER_13_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
X_160_ right_top_grid_pin_10_ chanx_right_out[0] vgnd vpwr scs8hd_buf_2
X_091_ _080_/B _091_/B _091_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_44 vgnd vpwr scs8hd_decap_12
XFILLER_10_223 vgnd vpwr scs8hd_fill_1
XFILLER_10_267 vgnd vpwr scs8hd_decap_8
XFILLER_1_26 vgnd vpwr scs8hd_fill_1
XANTENNA__136__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_3_219 vpwr vgnd scs8hd_fill_2
XANTENNA__062__A _062_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_79 vgnd vpwr scs8hd_decap_6
XFILLER_27_153 vgnd vpwr scs8hd_decap_4
XFILLER_19_66 vpwr vgnd scs8hd_fill_2
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
XFILLER_35_98 vgnd vpwr scs8hd_decap_12
XFILLER_27_197 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_track_1.LATCH_5_.latch_SLEEPB _104_/Y vgnd vpwr scs8hd_diode_2
X_074_ address[4] address[3] _110_/C _075_/C vgnd vpwr scs8hd_or3_4
X_143_ _143_/HI _143_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_274 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_123 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_80 vpwr vgnd scs8hd_fill_2
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__057__A address[3] vgnd vpwr scs8hd_diode_2
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_78 vpwr vgnd scs8hd_fill_2
XPHY_9 vgnd vpwr scs8hd_decap_3
Xmux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ _066_/Y mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_15_101 vpwr vgnd scs8hd_fill_2
XFILLER_15_112 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_25 vgnd vpwr scs8hd_decap_6
XFILLER_7_36 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[5] mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_126_ address[5] address[6] _132_/C address[0] _126_/Y vgnd vpwr scs8hd_nor4_4
X_057_ address[3] _110_/B vgnd vpwr scs8hd_inv_8
XANTENNA__133__C _075_/C vgnd vpwr scs8hd_diode_2
XFILLER_38_215 vgnd vpwr scs8hd_decap_12
XFILLER_30_6 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A top_left_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_10.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[8] mux_right_track_10.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_32_44 vgnd vpwr scs8hd_decap_12
XFILLER_12_148 vpwr vgnd scs8hd_fill_2
XFILLER_20_192 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _072_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA__128__C _075_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_11_170 vpwr vgnd scs8hd_fill_2
XANTENNA__160__A right_top_grid_pin_10_ vgnd vpwr scs8hd_diode_2
X_109_ _094_/A _105_/B _109_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_34_251 vgnd vpwr scs8hd_decap_12
XANTENNA__070__A _070_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_188 vpwr vgnd scs8hd_fill_2
XFILLER_4_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__130__D address[0] vgnd vpwr scs8hd_diode_2
XANTENNA__155__A _155_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A bottom_left_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_22_243 vgnd vpwr scs8hd_decap_12
XANTENNA__065__A _065_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_57 vpwr vgnd scs8hd_fill_2
XFILLER_1_158 vpwr vgnd scs8hd_fill_2
XFILLER_1_114 vgnd vpwr scs8hd_decap_4
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XANTENNA__125__D _135_/D vgnd vpwr scs8hd_diode_2
XFILLER_9_258 vgnd vpwr scs8hd_decap_4
XFILLER_9_269 vgnd vpwr scs8hd_decap_8
XFILLER_5_80 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_184 vgnd vpwr scs8hd_decap_12
XFILLER_24_56 vgnd vpwr scs8hd_decap_12
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
X_090_ _078_/B _091_/B _090_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_206 vpwr vgnd scs8hd_fill_2
XFILLER_10_213 vgnd vpwr scs8hd_fill_1
Xmux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _068_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB _138_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__136__C _096_/C vgnd vpwr scs8hd_diode_2
XFILLER_39_3 vgnd vpwr scs8hd_decap_12
XFILLER_36_154 vgnd vpwr scs8hd_decap_12
Xmem_right_track_2.LATCH_0_.latch data_in _060_/A _126_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_58 vpwr vgnd scs8hd_fill_2
XFILLER_35_11 vgnd vpwr scs8hd_decap_12
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
X_142_ _142_/HI _142_/LO vgnd vpwr scs8hd_conb_1
X_073_ address[1] _052_/Y _135_/D _076_/A vgnd vpwr scs8hd_or3_4
XANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A bottom_left_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_33_135 vgnd vpwr scs8hd_decap_12
XFILLER_18_121 vgnd vpwr scs8hd_decap_3
XFILLER_18_143 vpwr vgnd scs8hd_fill_2
XFILLER_18_154 vpwr vgnd scs8hd_fill_2
XANTENNA__163__A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__073__A address[1] vgnd vpwr scs8hd_diode_2
X_125_ address[5] address[6] _132_/C _135_/D _125_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_15_179 vpwr vgnd scs8hd_fill_2
X_056_ address[4] _110_/A vgnd vpwr scs8hd_inv_8
XANTENNA__133__D _135_/D vgnd vpwr scs8hd_diode_2
XFILLER_38_238 vgnd vpwr scs8hd_decap_12
XFILLER_38_227 vgnd vpwr scs8hd_decap_8
XANTENNA__158__A _158_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_205 vgnd vpwr scs8hd_decap_12
XANTENNA__068__A _068_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_56 vgnd vpwr scs8hd_decap_12
Xmem_top_track_0.LATCH_2_.latch data_in mem_top_track_0.LATCH_2_.latch/Q _082_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_182 vgnd vpwr scs8hd_decap_8
XFILLER_12_127 vgnd vpwr scs8hd_fill_1
XFILLER_35_208 vgnd vpwr scs8hd_decap_12
XFILLER_28_271 vgnd vpwr scs8hd_decap_4
XANTENNA__128__D address[0] vgnd vpwr scs8hd_diode_2
X_108_ _101_/A _105_/B _108_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_153 vpwr vgnd scs8hd_fill_2
XFILLER_7_175 vpwr vgnd scs8hd_fill_2
XFILLER_21_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _063_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_8.tap_buf4_0_.scs8hd_inv_1 mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _174_/A vgnd vpwr scs8hd_inv_1
XFILLER_25_241 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_101 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _143_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_263 vgnd vpwr scs8hd_decap_12
XANTENNA__171__A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_22_255 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_3_.scs8hd_inv_1 chanx_right_in[5] mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_137 vpwr vgnd scs8hd_fill_2
XANTENNA__081__A _079_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_7 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
XANTENNA__166__A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_39_196 vgnd vpwr scs8hd_decap_12
XANTENNA__076__A _076_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_68 vgnd vpwr scs8hd_decap_6
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
XANTENNA__136__D address[0] vgnd vpwr scs8hd_diode_2
XFILLER_5_240 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_1.LATCH_4_.latch data_in mem_bottom_track_1.LATCH_4_.latch/Q _105_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_166 vgnd vpwr scs8hd_decap_12
XFILLER_42_125 vgnd vpwr scs8hd_decap_12
XFILLER_35_23 vgnd vpwr scs8hd_decap_12
X_141_ _141_/HI _141_/LO vgnd vpwr scs8hd_conb_1
X_072_ _072_/A _072_/Y vgnd vpwr scs8hd_inv_8
Xmux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_8.LATCH_3_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_147 vgnd vpwr scs8hd_decap_12
Xmem_right_track_14.LATCH_1_.latch data_in _071_/A _137_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _069_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_158 vpwr vgnd scs8hd_fill_2
XFILLER_24_147 vgnd vpwr scs8hd_decap_6
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__073__B _052_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_128 vgnd vpwr scs8hd_decap_3
XFILLER_15_147 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
X_055_ address[6] _138_/B vgnd vpwr scs8hd_inv_8
XANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
X_124_ _094_/A _119_/B _124_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_80 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_bottom_track_17.LATCH_5_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__174__A _174_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_180 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_217 vpwr vgnd scs8hd_fill_2
XFILLER_16_58 vgnd vpwr scs8hd_decap_4
XFILLER_32_68 vgnd vpwr scs8hd_decap_12
XANTENNA__084__A _080_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_2_.latch_SLEEPB _092_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_110 vpwr vgnd scs8hd_fill_2
XFILLER_7_132 vgnd vpwr scs8hd_decap_4
XFILLER_7_165 vgnd vpwr scs8hd_fill_1
X_107_ _082_/B _105_/B _107_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_194 vpwr vgnd scs8hd_fill_2
XFILLER_14_3 vgnd vpwr scs8hd_decap_12
XFILLER_26_209 vgnd vpwr scs8hd_fill_1
XANTENNA__169__A _169_/A vgnd vpwr scs8hd_diode_2
XANTENNA__079__A _079_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_4_157 vgnd vpwr scs8hd_decap_4
XFILLER_4_135 vpwr vgnd scs8hd_fill_2
XFILLER_16_220 vgnd vpwr scs8hd_decap_3
XFILLER_17_90 vpwr vgnd scs8hd_fill_2
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_267 vgnd vpwr scs8hd_decap_8
XFILLER_13_15 vgnd vpwr scs8hd_decap_12
XANTENNA__081__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_38_56 vgnd vpwr scs8hd_decap_12
XFILLER_13_201 vgnd vpwr scs8hd_decap_8
XFILLER_13_245 vgnd vpwr scs8hd_decap_8
XFILLER_0_182 vpwr vgnd scs8hd_fill_2
XFILLER_0_171 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr
+ scs8hd_diode_2
XFILLER_39_120 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__076__B _080_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_215 vpwr vgnd scs8hd_fill_2
XFILLER_10_237 vgnd vpwr scs8hd_decap_4
XFILLER_10_248 vpwr vgnd scs8hd_fill_2
XFILLER_40_68 vgnd vpwr scs8hd_decap_12
XANTENNA__092__A _082_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_29 vpwr vgnd scs8hd_fill_2
XFILLER_36_178 vgnd vpwr scs8hd_decap_12
XANTENNA__177__A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_10.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_27_101 vpwr vgnd scs8hd_fill_2
XFILLER_42_137 vgnd vpwr scs8hd_decap_12
XFILLER_35_35 vgnd vpwr scs8hd_decap_12
XFILLER_27_123 vpwr vgnd scs8hd_fill_2
XANTENNA__087__A address[4] vgnd vpwr scs8hd_diode_2
X_071_ _071_/A _071_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_140_ _140_/HI _140_/LO vgnd vpwr scs8hd_conb_1
Xmux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_top_track_16.LATCH_4_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_bottom_track_9.INVTX1_2_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_33_159 vgnd vpwr scs8hd_decap_12
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_50 vgnd vpwr scs8hd_decap_4
XANTENNA__073__C _135_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_3_.scs8hd_inv_1 chanx_right_in[0] mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_126 vpwr vgnd scs8hd_fill_2
X_054_ address[5] _135_/A vgnd vpwr scs8hd_inv_8
X_123_ _101_/A _119_/B _123_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_21_118 vpwr vgnd scs8hd_fill_2
XFILLER_37_262 vgnd vpwr scs8hd_decap_12
Xmem_top_track_8.LATCH_3_.latch data_in mem_top_track_8.LATCH_3_.latch/Q _091_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_16_15 vgnd vpwr scs8hd_decap_12
XFILLER_16_37 vgnd vpwr scs8hd_decap_8
XANTENNA__084__B _101_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_106_ _080_/B _105_/B _106_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_199 vpwr vgnd scs8hd_fill_2
XFILLER_11_184 vgnd vpwr scs8hd_fill_1
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XANTENNA__079__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_40_202 vgnd vpwr scs8hd_decap_12
XANTENNA__095__A _110_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_147 vpwr vgnd scs8hd_fill_2
XFILLER_4_114 vpwr vgnd scs8hd_fill_2
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_257 vgnd vpwr scs8hd_decap_12
XFILLER_22_213 vgnd vpwr scs8hd_fill_1
XFILLER_13_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__081__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_38_68 vgnd vpwr scs8hd_decap_12
XFILLER_13_224 vpwr vgnd scs8hd_fill_2
XFILLER_9_217 vgnd vpwr scs8hd_decap_3
XFILLER_13_235 vgnd vpwr scs8hd_decap_3
Xmux_right_track_8.INVTX1_0_.scs8hd_inv_1 chany_top_in[4] mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_272 vgnd vpwr scs8hd_decap_3
XFILLER_5_83 vgnd vpwr scs8hd_decap_3
XFILLER_24_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_205 vpwr vgnd scs8hd_fill_2
XANTENNA__092__B _091_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_9.LATCH_5_.latch data_in mem_bottom_track_9.LATCH_5_.latch/Q _112_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_track_1.LATCH_2_.latch_SLEEPB _107_/Y vgnd vpwr scs8hd_diode_2
XFILLER_42_149 vgnd vpwr scs8hd_decap_6
XFILLER_35_47 vgnd vpwr scs8hd_decap_12
XFILLER_27_179 vpwr vgnd scs8hd_fill_2
XFILLER_27_157 vgnd vpwr scs8hd_fill_1
XANTENNA__087__B _110_/B vgnd vpwr scs8hd_diode_2
X_070_ _070_/A _070_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _071_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_5_.scs8hd_inv_1 bottom_right_grid_pin_11_ mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_41_171 vgnd vpwr scs8hd_decap_12
XPHY_80 vgnd vpwr scs8hd_decap_3
XFILLER_26_190 vpwr vgnd scs8hd_fill_2
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _144_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_2_84 vpwr vgnd scs8hd_fill_2
XFILLER_24_116 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_track_9.LATCH_4_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_8.INVTX1_4_.scs8hd_inv_1 chanx_right_in[5] mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__098__A _078_/B vgnd vpwr scs8hd_diode_2
XFILLER_15_105 vpwr vgnd scs8hd_fill_2
XFILLER_15_116 vgnd vpwr scs8hd_decap_4
XFILLER_23_193 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_053_ address[0] _135_/D vgnd vpwr scs8hd_inv_8
X_122_ _082_/B _119_/B _122_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB _098_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_5_.latch data_in mem_top_track_16.LATCH_5_.latch/Q _097_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_37_274 vgnd vpwr scs8hd_decap_3
XFILLER_32_15 vgnd vpwr scs8hd_decap_12
Xmem_right_track_10.LATCH_1_.latch data_in _065_/A _131_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_16_27 vgnd vpwr scs8hd_decap_4
XFILLER_20_152 vgnd vpwr scs8hd_fill_1
XFILLER_28_241 vgnd vpwr scs8hd_decap_12
X_105_ _078_/B _105_/B _105_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_163 vpwr vgnd scs8hd_fill_2
XFILLER_11_174 vgnd vpwr scs8hd_decap_3
XFILLER_19_263 vgnd vpwr scs8hd_decap_12
XFILLER_19_252 vpwr vgnd scs8hd_fill_2
XFILLER_8_72 vpwr vgnd scs8hd_fill_2
XFILLER_27_59 vpwr vgnd scs8hd_fill_2
XFILLER_27_15 vgnd vpwr scs8hd_decap_12
XFILLER_25_233 vpwr vgnd scs8hd_fill_2
XANTENNA__079__C _135_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__095__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_4_19 vgnd vpwr scs8hd_decap_12
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_39 vgnd vpwr scs8hd_decap_12
XFILLER_13_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_151 vpwr vgnd scs8hd_fill_2
XFILLER_28_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_17.LATCH_3_.latch_SLEEPB _121_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_62 vgnd vpwr scs8hd_decap_3
XFILLER_24_27 vgnd vpwr scs8hd_decap_4
XFILLER_40_15 vgnd vpwr scs8hd_decap_12
XFILLER_6_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_221 vpwr vgnd scs8hd_fill_2
XFILLER_5_232 vpwr vgnd scs8hd_fill_2
XFILLER_5_254 vpwr vgnd scs8hd_fill_2
XFILLER_5_265 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _070_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_39_90 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_2_.latch/Q mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_track_17.LATCH_5_.latch data_in mem_bottom_track_17.LATCH_5_.latch/Q _119_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_27_136 vpwr vgnd scs8hd_fill_2
XFILLER_27_114 vpwr vgnd scs8hd_fill_2
Xmux_right_track_6.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__087__C _110_/C vgnd vpwr scs8hd_diode_2
XFILLER_19_49 vgnd vpwr scs8hd_fill_1
XFILLER_42_106 vgnd vpwr scs8hd_decap_12
XFILLER_35_59 vpwr vgnd scs8hd_fill_2
XFILLER_2_213 vgnd vpwr scs8hd_fill_1
XFILLER_2_246 vgnd vpwr scs8hd_decap_12
XFILLER_2_235 vgnd vpwr scs8hd_decap_8
XFILLER_2_224 vpwr vgnd scs8hd_fill_2
XFILLER_18_147 vgnd vpwr scs8hd_decap_6
XFILLER_18_158 vgnd vpwr scs8hd_decap_3
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XFILLER_25_92 vpwr vgnd scs8hd_fill_2
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _139_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_63 vpwr vgnd scs8hd_fill_2
XFILLER_24_139 vgnd vpwr scs8hd_decap_6
Xmux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_right_track_6.LATCH_1_.latch data_in _063_/A _129_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_track_0.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[4] mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__098__B _099_/B vgnd vpwr scs8hd_diode_2
XFILLER_23_150 vgnd vpwr scs8hd_decap_4
X_121_ _080_/B _119_/B _121_/Y vgnd vpwr scs8hd_nor2_4
X_052_ address[2] _052_/Y vgnd vpwr scs8hd_inv_8
XFILLER_36_80 vgnd vpwr scs8hd_decap_12
XFILLER_37_253 vpwr vgnd scs8hd_fill_2
XFILLER_37_220 vgnd vpwr scs8hd_decap_12
XFILLER_32_27 vgnd vpwr scs8hd_decap_4
XFILLER_28_220 vgnd vpwr scs8hd_decap_6
XFILLER_28_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _064_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB _135_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_104_ _076_/A _105_/B _104_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_157 vpwr vgnd scs8hd_fill_2
XFILLER_7_179 vpwr vgnd scs8hd_fill_2
XFILLER_21_7 vgnd vpwr scs8hd_decap_12
XFILLER_19_275 vpwr vgnd scs8hd_fill_2
XFILLER_19_242 vpwr vgnd scs8hd_fill_2
XFILLER_8_51 vpwr vgnd scs8hd_fill_2
XFILLER_27_27 vgnd vpwr scs8hd_decap_12
XFILLER_40_215 vgnd vpwr scs8hd_decap_12
XFILLER_25_245 vgnd vpwr scs8hd_decap_6
XANTENNA__095__C _110_/C vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_234 vgnd vpwr scs8hd_decap_8
XFILLER_17_71 vpwr vgnd scs8hd_fill_2
XFILLER_17_82 vpwr vgnd scs8hd_fill_2
XFILLER_3_193 vgnd vpwr scs8hd_decap_4
XFILLER_12_3 vgnd vpwr scs8hd_decap_12
XFILLER_22_226 vgnd vpwr scs8hd_decap_8
XFILLER_38_15 vgnd vpwr scs8hd_decap_12
XFILLER_21_270 vgnd vpwr scs8hd_decap_6
XFILLER_0_196 vgnd vpwr scs8hd_decap_4
XFILLER_39_123 vgnd vpwr scs8hd_decap_12
XFILLER_40_27 vgnd vpwr scs8hd_decap_4
XFILLER_30_93 vgnd vpwr scs8hd_fill_1
XFILLER_10_19 vgnd vpwr scs8hd_decap_12
XFILLER_42_118 vgnd vpwr scs8hd_decap_6
XFILLER_2_203 vpwr vgnd scs8hd_fill_2
Xmux_right_track_14.tap_buf4_0_.scs8hd_inv_1 mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ _153_/A vgnd vpwr scs8hd_inv_1
XFILLER_2_258 vgnd vpwr scs8hd_decap_12
XFILLER_18_104 vgnd vpwr scs8hd_decap_8
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_18_126 vpwr vgnd scs8hd_fill_2
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.tap_buf4_0_.scs8hd_inv_1 mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _170_/A vgnd vpwr scs8hd_inv_1
XFILLER_32_151 vpwr vgnd scs8hd_fill_2
XFILLER_23_162 vpwr vgnd scs8hd_fill_2
X_051_ address[1] _079_/A vgnd vpwr scs8hd_inv_8
X_120_ _078_/B _119_/B _120_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_4.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_62 vgnd vpwr scs8hd_fill_1
XFILLER_11_84 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_184 vpwr vgnd scs8hd_fill_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_243 vgnd vpwr scs8hd_fill_1
XFILLER_37_232 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_165 vpwr vgnd scs8hd_fill_2
XFILLER_20_154 vpwr vgnd scs8hd_fill_2
XFILLER_20_143 vgnd vpwr scs8hd_fill_1
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
XFILLER_7_114 vpwr vgnd scs8hd_fill_2
X_103_ address[5] _138_/B _096_/C _105_/B vgnd vpwr scs8hd_or3_4
XFILLER_11_198 vpwr vgnd scs8hd_fill_2
XFILLER_34_213 vgnd vpwr scs8hd_fill_1
XFILLER_19_210 vpwr vgnd scs8hd_fill_2
XFILLER_8_85 vgnd vpwr scs8hd_fill_1
XFILLER_27_39 vgnd vpwr scs8hd_decap_12
XFILLER_40_238 vgnd vpwr scs8hd_decap_12
XFILLER_40_227 vgnd vpwr scs8hd_decap_8
XFILLER_25_257 vgnd vpwr scs8hd_decap_12
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_205 vpwr vgnd scs8hd_fill_2
XFILLER_30_271 vgnd vpwr scs8hd_decap_4
XFILLER_38_27 vgnd vpwr scs8hd_decap_4
Xmux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_12.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_120 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_93 vgnd vpwr scs8hd_decap_6
XFILLER_8_253 vgnd vpwr scs8hd_decap_8
XFILLER_8_264 vgnd vpwr scs8hd_decap_8
XFILLER_12_260 vgnd vpwr scs8hd_decap_12
XFILLER_5_53 vpwr vgnd scs8hd_fill_2
XFILLER_5_97 vpwr vgnd scs8hd_fill_2
XFILLER_39_135 vgnd vpwr scs8hd_decap_12
XFILLER_10_219 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_190 vgnd vpwr scs8hd_decap_12
XFILLER_5_201 vpwr vgnd scs8hd_fill_2
XFILLER_14_73 vgnd vpwr scs8hd_decap_8
XFILLER_14_84 vgnd vpwr scs8hd_decap_8
Xmux_right_track_8.tap_buf4_0_.scs8hd_inv_1 mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _156_/A vgnd vpwr scs8hd_inv_1
XFILLER_30_72 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_2_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_70 vgnd vpwr scs8hd_decap_12
XFILLER_36_105 vgnd vpwr scs8hd_decap_12
XANTENNA__101__A _101_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XFILLER_26_160 vgnd vpwr scs8hd_decap_3
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_5_ mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_32 vgnd vpwr scs8hd_decap_4
XFILLER_24_108 vgnd vpwr scs8hd_decap_8
XFILLER_32_163 vgnd vpwr scs8hd_decap_12
XFILLER_21_19 vgnd vpwr scs8hd_decap_12
XFILLER_23_130 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _139_/HI mem_bottom_track_1.LATCH_2_.latch/Q
+ mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_9.LATCH_3_.latch_SLEEPB _114_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_93 vgnd vpwr scs8hd_decap_12
XFILLER_14_163 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_100 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_2.LATCH_1_.latch data_in _059_/A _125_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_133 vpwr vgnd scs8hd_fill_2
XFILLER_22_84 vgnd vpwr scs8hd_decap_8
X_102_ _094_/A _099_/B _102_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_2.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_170 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_214 vpwr vgnd scs8hd_fill_2
XFILLER_25_269 vgnd vpwr scs8hd_decap_8
XFILLER_4_118 vpwr vgnd scs8hd_fill_2
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__104__A _076_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_162 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_110 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_top_track_0.LATCH_3_.latch data_in mem_top_track_0.LATCH_3_.latch/Q _080_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
XFILLER_12_272 vgnd vpwr scs8hd_decap_3
XFILLER_5_76 vgnd vpwr scs8hd_decap_4
Xmem_bottom_track_9.LATCH_0_.latch data_in mem_bottom_track_9.LATCH_0_.latch/Q _117_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_147 vgnd vpwr scs8hd_decap_12
XFILLER_10_209 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_82 vgnd vpwr scs8hd_decap_4
XFILLER_36_117 vgnd vpwr scs8hd_decap_12
XFILLER_29_180 vgnd vpwr scs8hd_fill_1
XANTENNA__101__B _099_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_2_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_19 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_7 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.INVTX1_1_.scs8hd_inv_1 top_left_grid_pin_9_ mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XFILLER_26_183 vgnd vpwr scs8hd_fill_1
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_62 vgnd vpwr scs8hd_decap_12
XFILLER_25_51 vgnd vpwr scs8hd_decap_8
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
XFILLER_37_7 vpwr vgnd scs8hd_fill_2
XANTENNA__112__A _076_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_175 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB _101_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_197 vgnd vpwr scs8hd_decap_8
XFILLER_23_175 vpwr vgnd scs8hd_fill_2
XFILLER_23_142 vpwr vgnd scs8hd_fill_2
Xmem_top_track_16.LATCH_0_.latch data_in mem_top_track_16.LATCH_0_.latch/Q _102_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_53 vpwr vgnd scs8hd_fill_2
XANTENNA__107__A _082_/B vgnd vpwr scs8hd_diode_2
X_178_ _178_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_245 vgnd vpwr scs8hd_decap_8
XFILLER_28_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_5_.latch data_in mem_bottom_track_1.LATCH_5_.latch/Q _104_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_201 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_101_ _101_/A _099_/B _101_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_138 vpwr vgnd scs8hd_fill_2
XFILLER_11_123 vgnd vpwr scs8hd_fill_1
XFILLER_7_149 vpwr vgnd scs8hd_fill_2
XFILLER_19_234 vpwr vgnd scs8hd_fill_2
XFILLER_19_223 vpwr vgnd scs8hd_fill_2
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XFILLER_6_160 vgnd vpwr scs8hd_fill_1
XFILLER_8_32 vgnd vpwr scs8hd_decap_8
XFILLER_6_193 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_237 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB _080_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_7_.scs8hd_inv_1 bottom_left_grid_pin_13_ mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _069_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_215 vgnd vpwr scs8hd_decap_3
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_62 vgnd vpwr scs8hd_decap_12
XFILLER_33_51 vgnd vpwr scs8hd_decap_8
XANTENNA__104__B _105_/B vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _078_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_251 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_240 vpwr vgnd scs8hd_fill_2
XFILLER_5_33 vgnd vpwr scs8hd_decap_3
XANTENNA__115__A _082_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_159 vgnd vpwr scs8hd_decap_12
XFILLER_39_104 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_track_17.LATCH_0_.latch data_in mem_bottom_track_17.LATCH_0_.latch/Q _124_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_30_30 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_top_track_8.LATCH_4_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_5_225 vgnd vpwr scs8hd_decap_4
XFILLER_5_236 vpwr vgnd scs8hd_fill_2
XFILLER_5_258 vpwr vgnd scs8hd_fill_2
XFILLER_5_269 vgnd vpwr scs8hd_decap_8
XFILLER_39_94 vgnd vpwr scs8hd_decap_6
XFILLER_36_129 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_3_ vgnd vpwr scs8hd_diode_2
XFILLER_27_118 vpwr vgnd scs8hd_fill_2
XFILLER_35_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_228 vgnd vpwr scs8hd_decap_4
XFILLER_26_151 vpwr vgnd scs8hd_fill_2
XPHY_30 vgnd vpwr scs8hd_decap_3
Xmux_top_track_0.INVTX1_4_.scs8hd_inv_1 chanx_right_in[4] mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XFILLER_25_96 vpwr vgnd scs8hd_fill_2
XFILLER_25_74 vgnd vpwr scs8hd_decap_12
XPHY_41 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr
+ scs8hd_diode_2
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
XFILLER_2_67 vpwr vgnd scs8hd_fill_2
XANTENNA__112__B _113_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_143 vgnd vpwr scs8hd_decap_8
XFILLER_17_162 vpwr vgnd scs8hd_fill_2
XFILLER_17_184 vpwr vgnd scs8hd_fill_2
XFILLER_32_187 vgnd vpwr scs8hd_decap_12
XFILLER_23_110 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
X_177_ chany_bottom_in[0] chany_top_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA__107__B _105_/B vgnd vpwr scs8hd_diode_2
XANTENNA__123__A _101_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_124 vgnd vpwr scs8hd_fill_1
XFILLER_20_146 vgnd vpwr scs8hd_decap_6
XFILLER_28_213 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A bottom_left_grid_pin_1_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_64 vgnd vpwr scs8hd_fill_1
X_100_ _082_/B _099_/B _100_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_179 vpwr vgnd scs8hd_fill_2
XFILLER_34_205 vgnd vpwr scs8hd_decap_8
XFILLER_34_227 vgnd vpwr scs8hd_decap_12
XANTENNA__118__A _135_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_55 vpwr vgnd scs8hd_fill_2
XFILLER_8_88 vpwr vgnd scs8hd_fill_2
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XFILLER_17_31 vgnd vpwr scs8hd_decap_8
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_208 vgnd vpwr scs8hd_decap_12
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_53 vpwr vgnd scs8hd_fill_2
XFILLER_17_75 vpwr vgnd scs8hd_fill_2
XFILLER_17_86 vpwr vgnd scs8hd_fill_2
XFILLER_33_74 vgnd vpwr scs8hd_decap_12
XFILLER_3_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA__120__B _119_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_2_.latch/Q mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_178 vpwr vgnd scs8hd_fill_2
XFILLER_0_167 vpwr vgnd scs8hd_fill_2
XFILLER_0_134 vpwr vgnd scs8hd_fill_2
Xmem_top_track_8.LATCH_4_.latch data_in mem_top_track_8.LATCH_4_.latch/Q _090_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__115__B _113_/B vgnd vpwr scs8hd_diode_2
XANTENNA__131__A _135_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_32 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_track_16.LATCH_5_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_39_51 vgnd vpwr scs8hd_decap_8
XFILLER_29_193 vgnd vpwr scs8hd_decap_12
XANTENNA__126__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_35_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_207 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XPHY_75 vgnd vpwr scs8hd_decap_3
XFILLER_25_86 vgnd vpwr scs8hd_decap_3
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_46 vpwr vgnd scs8hd_fill_2
XFILLER_1_262 vgnd vpwr scs8hd_decap_12
XFILLER_32_199 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_99 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_track_1.LATCH_3_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_144 vpwr vgnd scs8hd_fill_2
XFILLER_14_188 vgnd vpwr scs8hd_decap_4
X_176_ chany_bottom_in[1] chany_top_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA__123__B _119_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_258 vpwr vgnd scs8hd_fill_2
XFILLER_20_169 vgnd vpwr scs8hd_decap_4
XFILLER_9_170 vgnd vpwr scs8hd_fill_1
XFILLER_11_114 vpwr vgnd scs8hd_fill_2
XFILLER_22_32 vgnd vpwr scs8hd_decap_12
XFILLER_7_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB _128_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
XFILLER_34_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_203 vgnd vpwr scs8hd_decap_4
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XANTENNA__118__B _138_/B vgnd vpwr scs8hd_diode_2
X_159_ _159_/A chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA__134__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_33_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_206 vgnd vpwr scs8hd_decap_8
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_86 vgnd vpwr scs8hd_decap_12
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_132 vgnd vpwr scs8hd_decap_3
XFILLER_22_209 vgnd vpwr scs8hd_decap_4
XANTENNA__129__A _135_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_202 vgnd vpwr scs8hd_fill_1
XFILLER_8_224 vgnd vpwr scs8hd_decap_3
XFILLER_5_13 vgnd vpwr scs8hd_decap_12
XFILLER_5_57 vpwr vgnd scs8hd_fill_2
XANTENNA__131__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_30_98 vgnd vpwr scs8hd_decap_12
XFILLER_30_32 vgnd vpwr scs8hd_decap_12
XFILLER_5_205 vgnd vpwr scs8hd_decap_3
XFILLER_29_172 vpwr vgnd scs8hd_fill_2
XFILLER_29_161 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__126__B address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_271 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_track_9.LATCH_5_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__052__A address[2] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_5_.scs8hd_inv_1 bottom_left_grid_pin_3_ mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XFILLER_26_186 vpwr vgnd scs8hd_fill_2
XPHY_54 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_10 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
Xmux_right_track_14.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[3] mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_274 vgnd vpwr scs8hd_decap_3
XFILLER_2_36 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB _117_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_17_153 vgnd vpwr scs8hd_fill_1
XFILLER_32_123 vgnd vpwr scs8hd_fill_1
XANTENNA__137__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_17_175 vpwr vgnd scs8hd_fill_2
XFILLER_17_197 vpwr vgnd scs8hd_fill_2
XFILLER_23_123 vgnd vpwr scs8hd_decap_4
XFILLER_11_45 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
X_175_ chany_bottom_in[2] chany_top_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_35_7 vpwr vgnd scs8hd_fill_2
XFILLER_37_237 vgnd vpwr scs8hd_decap_6
XFILLER_9_182 vgnd vpwr scs8hd_fill_1
XFILLER_20_104 vgnd vpwr scs8hd_decap_4
XFILLER_20_137 vgnd vpwr scs8hd_decap_6
XFILLER_28_259 vgnd vpwr scs8hd_decap_12
XFILLER_28_226 vgnd vpwr scs8hd_fill_1
XFILLER_28_215 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_104 vpwr vgnd scs8hd_fill_2
XFILLER_11_137 vgnd vpwr scs8hd_decap_3
XFILLER_22_44 vgnd vpwr scs8hd_decap_12
XFILLER_11_159 vpwr vgnd scs8hd_fill_2
XFILLER_19_259 vpwr vgnd scs8hd_fill_2
XFILLER_19_248 vpwr vgnd scs8hd_fill_2
Xmux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_2_.scs8hd_inv_1/Y
+ _064_/A mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
XFILLER_8_68 vpwr vgnd scs8hd_fill_2
XFILLER_8_79 vgnd vpwr scs8hd_decap_6
XANTENNA__118__C _075_/C vgnd vpwr scs8hd_diode_2
X_089_ _076_/A _091_/B _089_/Y vgnd vpwr scs8hd_nor2_4
X_158_ _158_/A chanx_right_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA__134__B _138_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_152 vgnd vpwr scs8hd_fill_1
XFILLER_6_174 vpwr vgnd scs8hd_fill_2
XFILLER_26_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_218 vpwr vgnd scs8hd_fill_2
XANTENNA__060__A _060_/A vgnd vpwr scs8hd_diode_2
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_98 vgnd vpwr scs8hd_decap_12
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_199 vpwr vgnd scs8hd_fill_2
XFILLER_30_210 vgnd vpwr scs8hd_decap_4
XANTENNA__129__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_254 vgnd vpwr scs8hd_decap_8
XANTENNA__055__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_28_32 vgnd vpwr scs8hd_decap_12
XFILLER_0_114 vgnd vpwr scs8hd_decap_4
XFILLER_0_147 vpwr vgnd scs8hd_fill_2
XFILLER_8_236 vgnd vpwr scs8hd_decap_8
XFILLER_12_243 vgnd vpwr scs8hd_decap_8
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
XFILLER_5_25 vgnd vpwr scs8hd_decap_8
XANTENNA__131__C _132_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_4_.latch_SLEEPB _090_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_77 vgnd vpwr scs8hd_decap_12
XFILLER_30_44 vgnd vpwr scs8hd_decap_12
XFILLER_39_86 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_151 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__126__C _132_/C vgnd vpwr scs8hd_diode_2
XFILLER_35_110 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _149_/HI mem_top_track_0.LATCH_2_.latch/Q
+ mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_26_110 vgnd vpwr scs8hd_decap_6
XFILLER_41_135 vgnd vpwr scs8hd_decap_12
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_165 vgnd vpwr scs8hd_decap_3
XFILLER_26_154 vpwr vgnd scs8hd_fill_2
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_231 vpwr vgnd scs8hd_fill_2
XFILLER_17_143 vpwr vgnd scs8hd_fill_2
XFILLER_40_190 vgnd vpwr scs8hd_decap_12
XFILLER_32_157 vgnd vpwr scs8hd_decap_4
XANTENNA__137__B _138_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__153__A _153_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_179 vpwr vgnd scs8hd_fill_2
XFILLER_23_146 vpwr vgnd scs8hd_fill_2
XFILLER_23_102 vpwr vgnd scs8hd_fill_2
XANTENNA__063__A _063_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_57 vpwr vgnd scs8hd_fill_2
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_1.LATCH_0_.latch data_in mem_bottom_track_1.LATCH_0_.latch/Q _109_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_102 vgnd vpwr scs8hd_decap_4
X_174_ _174_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
Xmux_right_track_12.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[1] mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_127 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_91 vpwr vgnd scs8hd_fill_2
XFILLER_3_80 vpwr vgnd scs8hd_fill_2
XANTENNA__058__A enable vgnd vpwr scs8hd_diode_2
XFILLER_22_67 vgnd vpwr scs8hd_decap_6
XFILLER_22_56 vgnd vpwr scs8hd_decap_8
XFILLER_19_238 vpwr vgnd scs8hd_fill_2
XFILLER_19_227 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB _086_/Y vgnd vpwr scs8hd_diode_2
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.INVTX1_4_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_157_ _157_/A chanx_right_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA__134__C _075_/C vgnd vpwr scs8hd_diode_2
XFILLER_6_131 vpwr vgnd scs8hd_fill_2
XFILLER_10_193 vgnd vpwr scs8hd_fill_1
X_088_ address[5] address[6] _138_/C _091_/B vgnd vpwr scs8hd_or3_4
XFILLER_19_3 vpwr vgnd scs8hd_fill_2
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_274 vgnd vpwr scs8hd_fill_1
Xmux_top_track_16.INVTX1_5_.scs8hd_inv_1 chanx_right_in[6] mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_112 vpwr vgnd scs8hd_fill_2
XANTENNA__129__C _138_/C vgnd vpwr scs8hd_diode_2
XFILLER_15_252 vpwr vgnd scs8hd_fill_2
XANTENNA__161__A _161_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_266 vpwr vgnd scs8hd_fill_2
XFILLER_21_222 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__071__A _071_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_44 vgnd vpwr scs8hd_decap_12
XFILLER_8_215 vgnd vpwr scs8hd_fill_1
XFILLER_39_108 vgnd vpwr scs8hd_decap_12
XANTENNA__131__D _135_/D vgnd vpwr scs8hd_diode_2
XFILLER_10_7 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__156__A _156_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_10.tap_buf4_0_.scs8hd_inv_1 mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ _155_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__066__A _066_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_56 vgnd vpwr scs8hd_decap_12
XFILLER_14_46 vgnd vpwr scs8hd_decap_12
XFILLER_30_89 vgnd vpwr scs8hd_decap_3
XANTENNA__126__D address[0] vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_1_.scs8hd_inv_1 top_left_grid_pin_7_ mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_41_147 vgnd vpwr scs8hd_decap_12
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XFILLER_1_210 vgnd vpwr scs8hd_decap_4
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
XFILLER_1_243 vgnd vpwr scs8hd_fill_1
XANTENNA__137__C _138_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _060_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_158 vpwr vgnd scs8hd_fill_2
XFILLER_23_114 vpwr vgnd scs8hd_fill_2
XFILLER_36_44 vgnd vpwr scs8hd_decap_12
XFILLER_14_125 vgnd vpwr scs8hd_decap_3
X_173_ chany_bottom_in[4] chany_top_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA__164__A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_4_.latch_SLEEPB _105_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_140 vpwr vgnd scs8hd_fill_2
XFILLER_9_162 vpwr vgnd scs8hd_fill_2
XFILLER_9_184 vgnd vpwr scs8hd_decap_3
XANTENNA__074__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
X_156_ _156_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
X_087_ address[4] _110_/B _110_/C _138_/C vgnd vpwr scs8hd_or3_4
Xmux_bottom_track_1.INVTX1_7_.scs8hd_inv_1 bottom_left_grid_pin_11_ mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__134__D address[0] vgnd vpwr scs8hd_diode_2
XFILLER_6_110 vpwr vgnd scs8hd_fill_2
XFILLER_6_154 vgnd vpwr scs8hd_decap_6
XANTENNA__159__A _159_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[1] mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__069__A _069_/A vgnd vpwr scs8hd_diode_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_242 vgnd vpwr scs8hd_decap_12
XFILLER_24_231 vgnd vpwr scs8hd_decap_8
XFILLER_17_57 vpwr vgnd scs8hd_fill_2
Xmux_right_track_10.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[2] mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_223 vpwr vgnd scs8hd_fill_2
XANTENNA__129__D _135_/D vgnd vpwr scs8hd_diode_2
X_139_ _139_/HI _139_/LO vgnd vpwr scs8hd_conb_1
Xmux_right_track_4.tap_buf4_0_.scs8hd_inv_1 mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ _158_/A vgnd vpwr scs8hd_inv_1
XFILLER_0_71 vpwr vgnd scs8hd_fill_2
XFILLER_0_138 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_10.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_56 vgnd vpwr scs8hd_decap_12
XFILLER_5_38 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__172__A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_69 vpwr vgnd scs8hd_fill_2
XFILLER_30_68 vgnd vpwr scs8hd_decap_4
XANTENNA__082__A _080_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_66 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_35_123 vgnd vpwr scs8hd_decap_12
XANTENNA__167__A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XPHY_46 vgnd vpwr scs8hd_decap_3
XANTENNA__077__A address[1] vgnd vpwr scs8hd_diode_2
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XFILLER_41_159 vgnd vpwr scs8hd_decap_12
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_9_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__137__D _135_/D vgnd vpwr scs8hd_diode_2
XFILLER_17_123 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_17.LATCH_5_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XFILLER_31_170 vgnd vpwr scs8hd_decap_12
Xmem_top_track_0.LATCH_4_.latch data_in mem_top_track_0.LATCH_4_.latch/Q _078_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_15 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_9.LATCH_1_.latch data_in mem_bottom_track_9.LATCH_1_.latch/Q _116_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _069_/A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_36_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_148 vgnd vpwr scs8hd_decap_3
X_172_ chany_bottom_in[5] chany_top_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_22_192 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _145_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_170 vpwr vgnd scs8hd_fill_2
XFILLER_20_118 vgnd vpwr scs8hd_decap_6
XFILLER_9_174 vpwr vgnd scs8hd_fill_2
XFILLER_9_196 vpwr vgnd scs8hd_fill_2
XFILLER_28_229 vgnd vpwr scs8hd_decap_3
XFILLER_36_251 vgnd vpwr scs8hd_decap_12
XANTENNA__074__B address[3] vgnd vpwr scs8hd_diode_2
Xmux_right_track_6.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[5] mux_right_track_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_118 vpwr vgnd scs8hd_fill_2
XANTENNA__090__A _078_/B vgnd vpwr scs8hd_diode_2
XFILLER_27_262 vpwr vgnd scs8hd_fill_2
XFILLER_27_240 vgnd vpwr scs8hd_decap_4
XFILLER_19_207 vgnd vpwr scs8hd_fill_1
X_155_ _155_/A chanx_right_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_6_144 vpwr vgnd scs8hd_fill_2
X_086_ _080_/A _094_/A _086_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_243 vgnd vpwr scs8hd_fill_1
XANTENNA__175__A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XFILLER_24_254 vgnd vpwr scs8hd_decap_12
XANTENNA__085__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_3_158 vpwr vgnd scs8hd_fill_2
Xmem_top_track_16.LATCH_1_.latch data_in mem_top_track_16.LATCH_1_.latch/Q _101_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_276 vgnd vpwr scs8hd_fill_1
X_138_ address[5] _138_/B _138_/C address[0] _138_/Y vgnd vpwr scs8hd_nor4_4
X_069_ _069_/A _069_/Y vgnd vpwr scs8hd_inv_8
XFILLER_24_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_17.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_94 vgnd vpwr scs8hd_fill_1
Xmux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_2_.scs8hd_inv_1/Y
+ _062_/A mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_92 vpwr vgnd scs8hd_fill_2
XFILLER_0_106 vpwr vgnd scs8hd_fill_2
XFILLER_28_68 vgnd vpwr scs8hd_decap_12
XFILLER_8_206 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB _134_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_213 vgnd vpwr scs8hd_fill_1
Xmem_right_track_12.LATCH_0_.latch data_in _068_/A _134_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_154 vgnd vpwr scs8hd_decap_12
XFILLER_38_121 vgnd vpwr scs8hd_decap_12
XFILLER_14_15 vgnd vpwr scs8hd_decap_12
XANTENNA__082__B _082_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_176 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_2_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_135 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_0.LATCH_3_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_6_93 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.tap_buf4_0_.scs8hd_inv_1 mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _178_/A vgnd vpwr scs8hd_inv_1
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_179 vgnd vpwr scs8hd_decap_4
XFILLER_26_135 vpwr vgnd scs8hd_fill_2
XPHY_47 vgnd vpwr scs8hd_decap_3
XANTENNA__077__B _052_/Y vgnd vpwr scs8hd_diode_2
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XFILLER_34_190 vgnd vpwr scs8hd_decap_8
XANTENNA__093__A _101_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_245 vpwr vgnd scs8hd_fill_2
XFILLER_32_127 vgnd vpwr scs8hd_decap_12
XFILLER_32_105 vgnd vpwr scs8hd_decap_12
XFILLER_17_179 vpwr vgnd scs8hd_fill_2
XANTENNA__178__A _178_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_127 vgnd vpwr scs8hd_fill_1
XFILLER_31_182 vgnd vpwr scs8hd_fill_1
XFILLER_11_27 vgnd vpwr scs8hd_decap_12
XFILLER_11_49 vpwr vgnd scs8hd_fill_2
XANTENNA__088__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_36_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_171_ chany_bottom_in[6] chany_top_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_37_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_17.LATCH_1_.latch data_in mem_bottom_track_17.LATCH_1_.latch/Q _123_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_193 vpwr vgnd scs8hd_fill_2
XFILLER_20_108 vgnd vpwr scs8hd_fill_1
XFILLER_36_263 vgnd vpwr scs8hd_decap_12
XFILLER_11_108 vgnd vpwr scs8hd_decap_3
XANTENNA__074__C _110_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__090__B _091_/B vgnd vpwr scs8hd_diode_2
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XFILLER_27_274 vgnd vpwr scs8hd_decap_3
Xmux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_2_.scs8hd_inv_1/Y
+ _068_/A mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_085_ address[1] address[2] address[0] _094_/A vgnd vpwr scs8hd_or3_4
XFILLER_6_189 vpwr vgnd scs8hd_fill_2
X_154_ _154_/A chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_10_185 vpwr vgnd scs8hd_fill_2
XFILLER_12_81 vgnd vpwr scs8hd_decap_8
Xmux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_211 vgnd vpwr scs8hd_decap_3
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_266 vgnd vpwr scs8hd_decap_8
XANTENNA__085__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_3_137 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[6] mux_right_track_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_right_track_8.LATCH_0_.latch data_in _070_/A _136_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_137_ address[5] _138_/B _138_/C _135_/D _137_/Y vgnd vpwr scs8hd_nor4_4
X_068_ _068_/A _068_/Y vgnd vpwr scs8hd_inv_8
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_2_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_3 vpwr vgnd scs8hd_fill_2
XFILLER_21_236 vpwr vgnd scs8hd_fill_2
XFILLER_21_203 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB _093_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_12_203 vpwr vgnd scs8hd_fill_2
XANTENNA__096__A address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _066_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_8.LATCH_5_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_18_80 vpwr vgnd scs8hd_fill_2
XFILLER_7_240 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A top_left_grid_pin_9_ vgnd vpwr scs8hd_diode_2
XFILLER_38_166 vgnd vpwr scs8hd_decap_12
XFILLER_38_133 vgnd vpwr scs8hd_decap_12
XFILLER_14_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_10.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XFILLER_35_147 vgnd vpwr scs8hd_decap_12
XFILLER_6_61 vgnd vpwr scs8hd_decap_3
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_25_59 vpwr vgnd scs8hd_fill_2
XFILLER_25_15 vgnd vpwr scs8hd_decap_12
XPHY_48 vgnd vpwr scs8hd_decap_3
XANTENNA__077__C address[0] vgnd vpwr scs8hd_diode_2
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XPHY_37 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__093__B _091_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_235 vpwr vgnd scs8hd_fill_2
XFILLER_17_114 vpwr vgnd scs8hd_fill_2
XFILLER_17_147 vgnd vpwr scs8hd_decap_6
XFILLER_17_158 vpwr vgnd scs8hd_fill_2
XFILLER_32_139 vgnd vpwr scs8hd_fill_1
XFILLER_32_117 vgnd vpwr scs8hd_decap_6
XFILLER_15_81 vgnd vpwr scs8hd_decap_4
Xmem_top_track_8.LATCH_5_.latch data_in mem_top_track_8.LATCH_5_.latch/Q _089_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_106 vpwr vgnd scs8hd_fill_2
XFILLER_16_191 vgnd vpwr scs8hd_decap_4
XFILLER_11_39 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A bottom_left_grid_pin_7_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA__088__B address[6] vgnd vpwr scs8hd_diode_2
X_170_ _170_/A chany_top_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_14_106 vgnd vpwr scs8hd_fill_1
XFILLER_14_139 vgnd vpwr scs8hd_decap_3
XFILLER_26_80 vgnd vpwr scs8hd_fill_1
XFILLER_9_132 vpwr vgnd scs8hd_fill_2
XFILLER_3_84 vgnd vpwr scs8hd_decap_4
XFILLER_3_62 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_9.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__099__A _080_/B vgnd vpwr scs8hd_diode_2
XFILLER_27_253 vpwr vgnd scs8hd_fill_2
X_153_ _153_/A chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_12_93 vpwr vgnd scs8hd_fill_2
X_084_ _080_/A _101_/A _084_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_18_231 vpwr vgnd scs8hd_fill_2
XFILLER_19_7 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.INVTX1_2_.scs8hd_inv_1 top_right_grid_pin_11_ mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_33_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr
+ scs8hd_diode_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_6.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_33_59 vpwr vgnd scs8hd_fill_2
XFILLER_33_15 vgnd vpwr scs8hd_decap_12
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__085__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_3_116 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_9.LATCH_5_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_215 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_201 vgnd vpwr scs8hd_fill_1
XFILLER_15_234 vpwr vgnd scs8hd_fill_2
XFILLER_15_256 vgnd vpwr scs8hd_decap_12
XFILLER_30_259 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_70 vpwr vgnd scs8hd_fill_2
X_136_ _135_/A address[6] _096_/C address[0] _136_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_2_182 vpwr vgnd scs8hd_fill_2
X_067_ _067_/A _067_/Y vgnd vpwr scs8hd_inv_8
XFILLER_0_41 vpwr vgnd scs8hd_fill_2
XFILLER_28_15 vgnd vpwr scs8hd_decap_12
XANTENNA__096__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_12_226 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _149_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_219 vgnd vpwr scs8hd_decap_3
XFILLER_34_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _059_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_7_263 vgnd vpwr scs8hd_decap_12
X_119_ _076_/A _119_/B _119_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_38_145 vgnd vpwr scs8hd_decap_8
Xmux_right_track_2.INVTX1_2_.scs8hd_inv_1 right_bottom_grid_pin_12_ mux_right_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_38_178 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_134 vpwr vgnd scs8hd_fill_2
XFILLER_29_123 vpwr vgnd scs8hd_fill_2
XFILLER_4_222 vpwr vgnd scs8hd_fill_2
XFILLER_4_244 vgnd vpwr scs8hd_fill_1
XFILLER_35_159 vgnd vpwr scs8hd_decap_12
XFILLER_29_91 vgnd vpwr scs8hd_fill_1
XFILLER_6_73 vpwr vgnd scs8hd_fill_2
XFILLER_6_84 vpwr vgnd scs8hd_fill_2
XFILLER_25_27 vgnd vpwr scs8hd_decap_12
XPHY_49 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_258 vpwr vgnd scs8hd_fill_2
XFILLER_1_214 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_track_1.LATCH_4_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_71 vpwr vgnd scs8hd_fill_2
XFILLER_23_118 vpwr vgnd scs8hd_fill_2
XFILLER_31_184 vgnd vpwr scs8hd_decap_12
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XANTENNA__088__C _138_/C vgnd vpwr scs8hd_diode_2
XFILLER_22_173 vpwr vgnd scs8hd_fill_2
XFILLER_22_140 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB _108_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_3 vgnd vpwr scs8hd_decap_3
XFILLER_9_111 vpwr vgnd scs8hd_fill_2
XFILLER_9_166 vpwr vgnd scs8hd_fill_2
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_1.INVTX1_4_.scs8hd_inv_1 chanx_right_in[7] mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__099__B _099_/B vgnd vpwr scs8hd_diode_2
X_083_ address[1] address[2] _135_/D _101_/A vgnd vpwr scs8hd_or3_4
XFILLER_6_114 vpwr vgnd scs8hd_fill_2
XFILLER_8_19 vgnd vpwr scs8hd_decap_12
X_152_ _152_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_10_154 vgnd vpwr scs8hd_decap_3
Xmux_top_track_8.INVTX1_3_.scs8hd_inv_1 chanx_right_in[2] mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
Xmux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _063_/A mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_257 vgnd vpwr scs8hd_decap_12
XFILLER_5_180 vgnd vpwr scs8hd_decap_3
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_202 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB _099_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_39 vgnd vpwr scs8hd_decap_3
XFILLER_33_27 vgnd vpwr scs8hd_decap_12
XFILLER_30_227 vgnd vpwr scs8hd_decap_12
XFILLER_15_268 vgnd vpwr scs8hd_decap_8
X_135_ _135_/A address[6] _096_/C _135_/D _135_/Y vgnd vpwr scs8hd_nor4_4
X_066_ _066_/A _066_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mem_top_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_31_7 vpwr vgnd scs8hd_fill_2
XFILLER_9_62 vgnd vpwr scs8hd_fill_1
XFILLER_28_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__096__C _096_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_7_231 vpwr vgnd scs8hd_fill_2
XFILLER_11_260 vpwr vgnd scs8hd_fill_2
XFILLER_7_275 vpwr vgnd scs8hd_fill_2
X_118_ _135_/A _138_/B _075_/C _119_/B vgnd vpwr scs8hd_or3_4
Xmem_right_track_4.LATCH_0_.latch data_in _062_/A _128_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_59 vpwr vgnd scs8hd_fill_2
XFILLER_39_15 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_2_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_157 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB _076_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ _060_/A mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_4_212 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_20_50 vgnd vpwr scs8hd_decap_12
XFILLER_29_70 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_9.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_190 vpwr vgnd scs8hd_fill_2
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XFILLER_25_39 vgnd vpwr scs8hd_decap_12
XPHY_39 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_17.LATCH_2_.latch_SLEEPB _122_/Y vgnd vpwr scs8hd_diode_2
XFILLER_25_193 vpwr vgnd scs8hd_fill_2
XFILLER_25_171 vpwr vgnd scs8hd_fill_2
XFILLER_17_105 vpwr vgnd scs8hd_fill_2
XFILLER_40_141 vgnd vpwr scs8hd_decap_12
XFILLER_16_171 vpwr vgnd scs8hd_fill_2
XFILLER_31_196 vgnd vpwr scs8hd_decap_12
XFILLER_39_252 vgnd vpwr scs8hd_decap_4
Xmux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _071_/A mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_39_263 vgnd vpwr scs8hd_decap_12
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
XFILLER_14_119 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_152 vgnd vpwr scs8hd_fill_1
Xmux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _147_/HI _064_/Y mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_26_93 vgnd vpwr scs8hd_decap_6
XFILLER_13_163 vpwr vgnd scs8hd_fill_2
XFILLER_13_174 vpwr vgnd scs8hd_fill_2
XFILLER_9_145 vpwr vgnd scs8hd_fill_2
XFILLER_9_178 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _146_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_266 vgnd vpwr scs8hd_decap_8
X_151_ _151_/HI _151_/LO vgnd vpwr scs8hd_conb_1
X_082_ _080_/A _082_/B _082_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_148 vpwr vgnd scs8hd_fill_2
XFILLER_10_133 vgnd vpwr scs8hd_decap_3
XFILLER_12_40 vgnd vpwr scs8hd_decap_3
Xmux_top_track_0.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[0] mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _150_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_203 vgnd vpwr scs8hd_decap_12
XFILLER_18_244 vpwr vgnd scs8hd_fill_2
XFILLER_18_255 vgnd vpwr scs8hd_decap_12
XFILLER_33_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_8.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_33_39 vgnd vpwr scs8hd_decap_12
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_83 vpwr vgnd scs8hd_fill_2
X_134_ address[5] _138_/B _075_/C address[0] _134_/Y vgnd vpwr scs8hd_nor4_4
X_065_ _065_/A _065_/Y vgnd vpwr scs8hd_inv_8
Xmem_bottom_track_1.LATCH_1_.latch data_in mem_bottom_track_1.LATCH_1_.latch/Q _108_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_2_.scs8hd_inv_1/Y
+ _066_/A mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_0_32 vpwr vgnd scs8hd_fill_2
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
XFILLER_9_74 vpwr vgnd scs8hd_fill_2
XFILLER_9_96 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB _136_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_93 vgnd vpwr scs8hd_decap_12
XFILLER_7_254 vpwr vgnd scs8hd_fill_2
X_117_ _094_/A _113_/B _117_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_15_3 vgnd vpwr scs8hd_decap_12
XFILLER_30_18 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ _070_/A mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_39_27 vgnd vpwr scs8hd_decap_12
XFILLER_29_114 vpwr vgnd scs8hd_fill_2
XFILLER_29_103 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_62 vpwr vgnd scs8hd_fill_2
XFILLER_20_84 vpwr vgnd scs8hd_fill_2
XFILLER_6_97 vpwr vgnd scs8hd_fill_2
XFILLER_26_139 vgnd vpwr scs8hd_decap_12
XFILLER_19_180 vgnd vpwr scs8hd_decap_3
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XFILLER_1_249 vgnd vpwr scs8hd_decap_6
XFILLER_1_227 vpwr vgnd scs8hd_fill_2
XFILLER_15_40 vpwr vgnd scs8hd_fill_2
XFILLER_17_128 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__102__A _094_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_153 vpwr vgnd scs8hd_fill_2
XFILLER_39_275 vpwr vgnd scs8hd_fill_2
XFILLER_39_220 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_109 vgnd vpwr scs8hd_fill_1
XFILLER_13_197 vpwr vgnd scs8hd_fill_2
XFILLER_22_19 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _065_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_245 vgnd vpwr scs8hd_decap_8
XFILLER_27_223 vpwr vgnd scs8hd_fill_2
X_150_ _150_/HI _150_/LO vgnd vpwr scs8hd_conb_1
X_081_ _079_/A address[2] address[0] _082_/B vgnd vpwr scs8hd_or3_4
XFILLER_6_127 vpwr vgnd scs8hd_fill_2
XFILLER_10_145 vpwr vgnd scs8hd_fill_2
XFILLER_10_189 vgnd vpwr scs8hd_decap_4
XFILLER_12_52 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_215 vgnd vpwr scs8hd_decap_12
XFILLER_18_267 vgnd vpwr scs8hd_decap_8
XFILLER_5_193 vpwr vgnd scs8hd_fill_2
XFILLER_17_19 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A top_left_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_215 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _060_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_215 vpwr vgnd scs8hd_fill_2
XFILLER_15_248 vpwr vgnd scs8hd_fill_2
XFILLER_23_62 vpwr vgnd scs8hd_fill_2
XFILLER_23_51 vgnd vpwr scs8hd_decap_8
X_133_ address[5] _138_/B _075_/C _135_/D _133_/Y vgnd vpwr scs8hd_nor4_4
X_064_ _064_/A _064_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__110__A _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_7 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_218 vpwr vgnd scs8hd_fill_2
XFILLER_0_88 vgnd vpwr scs8hd_decap_3
XFILLER_9_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_207 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_84 vgnd vpwr scs8hd_decap_6
XANTENNA__105__A _078_/B vgnd vpwr scs8hd_diode_2
X_116_ _101_/A _113_/B _116_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_240 vpwr vgnd scs8hd_fill_2
XFILLER_39_39 vgnd vpwr scs8hd_decap_12
XFILLER_4_247 vgnd vpwr scs8hd_decap_12
XFILLER_20_96 vpwr vgnd scs8hd_fill_2
XFILLER_29_50 vgnd vpwr scs8hd_decap_8
XFILLER_6_32 vgnd vpwr scs8hd_decap_4
XFILLER_6_43 vgnd vpwr scs8hd_fill_1
XFILLER_26_118 vgnd vpwr scs8hd_decap_8
XPHY_19 vgnd vpwr scs8hd_decap_3
Xmem_top_track_8.LATCH_0_.latch data_in mem_top_track_8.LATCH_0_.latch/Q _094_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_239 vgnd vpwr scs8hd_decap_4
XFILLER_1_217 vgnd vpwr scs8hd_fill_1
XFILLER_17_118 vgnd vpwr scs8hd_decap_4
XFILLER_40_154 vgnd vpwr scs8hd_decap_12
XFILLER_15_85 vgnd vpwr scs8hd_fill_1
XFILLER_31_62 vgnd vpwr scs8hd_decap_12
XANTENNA__102__B _099_/B vgnd vpwr scs8hd_diode_2
XFILLER_31_110 vgnd vpwr scs8hd_decap_8
XFILLER_16_151 vpwr vgnd scs8hd_fill_2
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_243 vgnd vpwr scs8hd_fill_1
XFILLER_39_232 vgnd vpwr scs8hd_decap_3
XFILLER_22_154 vpwr vgnd scs8hd_fill_2
XFILLER_22_121 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _062_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_84 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_94 vgnd vpwr scs8hd_decap_12
XFILLER_9_136 vpwr vgnd scs8hd_fill_2
XFILLER_13_132 vpwr vgnd scs8hd_fill_2
XANTENNA__113__A _078_/B vgnd vpwr scs8hd_diode_2
XFILLER_36_202 vgnd vpwr scs8hd_decap_12
XFILLER_3_88 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_2_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
X_080_ _080_/A _080_/B _080_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_102 vgnd vpwr scs8hd_decap_4
XFILLER_10_168 vgnd vpwr scs8hd_decap_8
XFILLER_5_3 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_17.INVTX1_7_.scs8hd_inv_1 bottom_left_grid_pin_15_ mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_202 vgnd vpwr scs8hd_decap_3
XFILLER_18_213 vgnd vpwr scs8hd_fill_1
XFILLER_33_227 vgnd vpwr scs8hd_decap_12
XANTENNA__108__A _101_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_2_.latch_SLEEPB _115_/Y vgnd vpwr scs8hd_diode_2
XFILLER_38_3 vgnd vpwr scs8hd_decap_12
XFILLER_24_205 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_219 vgnd vpwr scs8hd_fill_1
XFILLER_15_238 vgnd vpwr scs8hd_decap_4
Xmem_top_track_0.LATCH_5_.latch data_in mem_top_track_0.LATCH_5_.latch/Q _076_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_063_ _063_/A _063_/Y vgnd vpwr scs8hd_inv_8
X_132_ _135_/A address[6] _132_/C address[0] _132_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_2_186 vpwr vgnd scs8hd_fill_2
XFILLER_2_131 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_9.LATCH_2_.latch data_in mem_bottom_track_9.LATCH_2_.latch/Q _115_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_23 vpwr vgnd scs8hd_fill_2
XANTENNA__110__B _110_/B vgnd vpwr scs8hd_diode_2
XFILLER_0_67 vpwr vgnd scs8hd_fill_2
XFILLER_14_271 vgnd vpwr scs8hd_decap_4
Xmux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _061_/A mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _060_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_274 vgnd vpwr scs8hd_fill_1
XFILLER_20_230 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_30 vgnd vpwr scs8hd_fill_1
XFILLER_18_52 vpwr vgnd scs8hd_fill_2
XFILLER_18_63 vpwr vgnd scs8hd_fill_2
XFILLER_11_230 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA__105__B _105_/B vgnd vpwr scs8hd_diode_2
X_115_ _082_/B _113_/B _115_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_38_105 vgnd vpwr scs8hd_fill_1
XANTENNA__121__A _080_/B vgnd vpwr scs8hd_diode_2
XFILLER_29_138 vpwr vgnd scs8hd_fill_2
XFILLER_37_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_226 vgnd vpwr scs8hd_decap_3
XFILLER_29_62 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_4_259 vgnd vpwr scs8hd_decap_12
XFILLER_29_95 vpwr vgnd scs8hd_fill_2
XFILLER_28_160 vgnd vpwr scs8hd_fill_1
XANTENNA__116__A _101_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_11 vgnd vpwr scs8hd_decap_12
XFILLER_6_77 vgnd vpwr scs8hd_decap_4
XFILLER_6_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_2_.latch data_in mem_top_track_16.LATCH_2_.latch/Q _100_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_34_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _148_/HI _069_/Y mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_141 vpwr vgnd scs8hd_fill_2
XFILLER_40_166 vgnd vpwr scs8hd_decap_12
XFILLER_15_53 vpwr vgnd scs8hd_fill_2
XFILLER_15_75 vgnd vpwr scs8hd_decap_4
XFILLER_31_74 vgnd vpwr scs8hd_decap_12
XFILLER_16_130 vpwr vgnd scs8hd_fill_2
XFILLER_16_163 vpwr vgnd scs8hd_fill_2
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _141_/HI vgnd vpwr
+ scs8hd_diode_2
.ends

