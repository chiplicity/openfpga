magic
tech EFS8A
magscale 1 2
timestamp 1604336936
<< locali >>
rect 7297 23511 7331 23613
rect 15577 5083 15611 5185
<< viali >>
rect 13185 25449 13219 25483
rect 19349 25449 19383 25483
rect 10517 25381 10551 25415
rect 10333 25313 10367 25347
rect 13001 25313 13035 25347
rect 19165 25313 19199 25347
rect 19809 25313 19843 25347
rect 10609 25245 10643 25279
rect 15945 25245 15979 25279
rect 10057 25177 10091 25211
rect 11069 25109 11103 25143
rect 11437 25109 11471 25143
rect 14013 24905 14047 24939
rect 6929 24837 6963 24871
rect 9965 24837 9999 24871
rect 10333 24837 10367 24871
rect 10609 24837 10643 24871
rect 13093 24837 13127 24871
rect 19625 24837 19659 24871
rect 6561 24769 6595 24803
rect 7849 24769 7883 24803
rect 12265 24769 12299 24803
rect 19993 24769 20027 24803
rect 10885 24701 10919 24735
rect 11529 24701 11563 24735
rect 14565 24701 14599 24735
rect 15669 24701 15703 24735
rect 16773 24701 16807 24735
rect 17325 24701 17359 24735
rect 18429 24701 18463 24735
rect 18981 24701 19015 24735
rect 21097 24701 21131 24735
rect 21649 24701 21683 24735
rect 22201 24701 22235 24735
rect 22753 24701 22787 24735
rect 7205 24633 7239 24667
rect 7389 24633 7423 24667
rect 7481 24633 7515 24667
rect 11069 24633 11103 24667
rect 11161 24633 11195 24667
rect 13369 24633 13403 24667
rect 13645 24633 13679 24667
rect 18337 24633 18371 24667
rect 20177 24633 20211 24667
rect 6285 24565 6319 24599
rect 9689 24565 9723 24599
rect 12817 24565 12851 24599
rect 13553 24565 13587 24599
rect 14749 24565 14783 24599
rect 15209 24565 15243 24599
rect 15853 24565 15887 24599
rect 16313 24565 16347 24599
rect 16957 24565 16991 24599
rect 18613 24565 18647 24599
rect 19441 24565 19475 24599
rect 20085 24565 20119 24599
rect 20545 24565 20579 24599
rect 21281 24565 21315 24599
rect 22385 24565 22419 24599
rect 6929 24361 6963 24395
rect 7573 24361 7607 24395
rect 8309 24361 8343 24395
rect 13093 24361 13127 24395
rect 17049 24361 17083 24395
rect 18153 24361 18187 24395
rect 21557 24361 21591 24395
rect 22753 24361 22787 24395
rect 23857 24361 23891 24395
rect 24961 24361 24995 24395
rect 10762 24293 10796 24327
rect 13921 24293 13955 24327
rect 15853 24293 15887 24327
rect 19625 24293 19659 24327
rect 20085 24293 20119 24327
rect 7297 24225 7331 24259
rect 8401 24225 8435 24259
rect 13737 24225 13771 24259
rect 16865 24225 16899 24259
rect 17969 24225 18003 24259
rect 19717 24225 19751 24259
rect 22569 24225 22603 24259
rect 23673 24225 23707 24259
rect 24777 24225 24811 24259
rect 8217 24157 8251 24191
rect 10517 24157 10551 24191
rect 14013 24157 14047 24191
rect 15117 24157 15151 24191
rect 15761 24157 15795 24191
rect 15945 24157 15979 24191
rect 19533 24157 19567 24191
rect 21465 24157 21499 24191
rect 21649 24157 21683 24191
rect 18613 24089 18647 24123
rect 21097 24089 21131 24123
rect 7849 24021 7883 24055
rect 10425 24021 10459 24055
rect 11897 24021 11931 24055
rect 12449 24021 12483 24055
rect 13461 24021 13495 24055
rect 15393 24021 15427 24055
rect 16405 24021 16439 24055
rect 18889 24021 18923 24055
rect 19165 24021 19199 24055
rect 9873 23817 9907 23851
rect 11345 23817 11379 23851
rect 12265 23817 12299 23851
rect 12633 23817 12667 23851
rect 14933 23817 14967 23851
rect 15577 23817 15611 23851
rect 16497 23817 16531 23851
rect 21833 23817 21867 23851
rect 22569 23817 22603 23851
rect 23857 23817 23891 23851
rect 24961 23817 24995 23851
rect 10425 23749 10459 23783
rect 18337 23749 18371 23783
rect 22293 23749 22327 23783
rect 10977 23681 11011 23715
rect 13369 23681 13403 23715
rect 13553 23681 13587 23715
rect 16865 23681 16899 23715
rect 17509 23681 17543 23715
rect 18797 23681 18831 23715
rect 7297 23613 7331 23647
rect 7573 23613 7607 23647
rect 7829 23613 7863 23647
rect 10701 23613 10735 23647
rect 12449 23613 12483 23647
rect 15945 23613 15979 23647
rect 17049 23613 17083 23647
rect 19809 23613 19843 23647
rect 19901 23613 19935 23647
rect 22385 23613 22419 23647
rect 23673 23613 23707 23647
rect 24225 23613 24259 23647
rect 24777 23613 24811 23647
rect 7113 23545 7147 23579
rect 10885 23545 10919 23579
rect 13093 23545 13127 23579
rect 13820 23545 13854 23579
rect 16221 23545 16255 23579
rect 18889 23545 18923 23579
rect 20146 23545 20180 23579
rect 24593 23545 24627 23579
rect 7297 23477 7331 23511
rect 7389 23477 7423 23511
rect 8953 23477 8987 23511
rect 10149 23477 10183 23511
rect 11805 23477 11839 23511
rect 16957 23477 16991 23511
rect 17785 23477 17819 23511
rect 18797 23477 18831 23511
rect 19349 23477 19383 23511
rect 21281 23477 21315 23511
rect 23029 23477 23063 23511
rect 23489 23477 23523 23511
rect 25329 23477 25363 23511
rect 8401 23273 8435 23307
rect 11529 23273 11563 23307
rect 13185 23273 13219 23307
rect 14013 23273 14047 23307
rect 15117 23273 15151 23307
rect 20269 23273 20303 23307
rect 22937 23273 22971 23307
rect 24777 23273 24811 23307
rect 10416 23205 10450 23239
rect 13737 23205 13771 23239
rect 15568 23205 15602 23239
rect 21272 23205 21306 23239
rect 7277 23137 7311 23171
rect 13001 23137 13035 23171
rect 18041 23137 18075 23171
rect 21005 23137 21039 23171
rect 24593 23137 24627 23171
rect 7021 23069 7055 23103
rect 10149 23069 10183 23103
rect 13277 23069 13311 23103
rect 14197 23069 14231 23103
rect 15301 23069 15335 23103
rect 17785 23069 17819 23103
rect 12725 23001 12759 23035
rect 17601 23001 17635 23035
rect 10057 22933 10091 22967
rect 12081 22933 12115 22967
rect 12541 22933 12575 22967
rect 16681 22933 16715 22967
rect 17233 22933 17267 22967
rect 19165 22933 19199 22967
rect 19901 22933 19935 22967
rect 20729 22933 20763 22967
rect 22385 22933 22419 22967
rect 6653 22729 6687 22763
rect 11345 22729 11379 22763
rect 13461 22729 13495 22763
rect 14473 22729 14507 22763
rect 16957 22729 16991 22763
rect 20913 22729 20947 22763
rect 24777 22729 24811 22763
rect 10333 22661 10367 22695
rect 11805 22661 11839 22695
rect 12541 22661 12575 22695
rect 15117 22661 15151 22695
rect 21097 22661 21131 22695
rect 10885 22593 10919 22627
rect 13093 22593 13127 22627
rect 14933 22593 14967 22627
rect 15669 22593 15703 22627
rect 22385 22593 22419 22627
rect 7113 22525 7147 22559
rect 7757 22525 7791 22559
rect 8024 22525 8058 22559
rect 10609 22525 10643 22559
rect 12265 22525 12299 22559
rect 14197 22525 14231 22559
rect 15393 22525 15427 22559
rect 16773 22525 16807 22559
rect 17325 22525 17359 22559
rect 18521 22525 18555 22559
rect 20545 22525 20579 22559
rect 21649 22525 21683 22559
rect 24593 22525 24627 22559
rect 12817 22457 12851 22491
rect 13001 22457 13035 22491
rect 16037 22457 16071 22491
rect 17785 22457 17819 22491
rect 18337 22457 18371 22491
rect 18766 22457 18800 22491
rect 21373 22457 21407 22491
rect 21557 22457 21591 22491
rect 7665 22389 7699 22423
rect 9137 22389 9171 22423
rect 9689 22389 9723 22423
rect 10149 22389 10183 22423
rect 10793 22389 10827 22423
rect 15577 22389 15611 22423
rect 19901 22389 19935 22423
rect 22017 22389 22051 22423
rect 24409 22389 24443 22423
rect 25237 22389 25271 22423
rect 6653 22185 6687 22219
rect 8217 22185 8251 22219
rect 10241 22185 10275 22219
rect 11713 22185 11747 22219
rect 12449 22185 12483 22219
rect 16221 22185 16255 22219
rect 17785 22185 17819 22219
rect 21189 22185 21223 22219
rect 7573 22117 7607 22151
rect 8309 22117 8343 22151
rect 11805 22117 11839 22151
rect 14013 22117 14047 22151
rect 17877 22117 17911 22151
rect 18521 22117 18555 22151
rect 19349 22117 19383 22151
rect 22201 22117 22235 22151
rect 11529 22049 11563 22083
rect 15025 22049 15059 22083
rect 22293 22049 22327 22083
rect 23469 22049 23503 22083
rect 8125 21981 8159 22015
rect 12817 21981 12851 22015
rect 13921 21981 13955 22015
rect 14105 21981 14139 22015
rect 16221 21981 16255 22015
rect 16313 21981 16347 22015
rect 17785 21981 17819 22015
rect 19257 21981 19291 22015
rect 19441 21981 19475 22015
rect 21557 21981 21591 22015
rect 22201 21981 22235 22015
rect 23213 21981 23247 22015
rect 11253 21913 11287 21947
rect 13553 21913 13587 21947
rect 15761 21913 15795 21947
rect 17325 21913 17359 21947
rect 18889 21913 18923 21947
rect 19809 21913 19843 21947
rect 7757 21845 7791 21879
rect 10793 21845 10827 21879
rect 13185 21845 13219 21879
rect 15577 21845 15611 21879
rect 16681 21845 16715 21879
rect 20177 21845 20211 21879
rect 21741 21845 21775 21879
rect 24593 21845 24627 21879
rect 13829 21641 13863 21675
rect 14933 21641 14967 21675
rect 16497 21641 16531 21675
rect 17417 21641 17451 21675
rect 17785 21641 17819 21675
rect 19349 21641 19383 21675
rect 20361 21641 20395 21675
rect 10793 21573 10827 21607
rect 12817 21573 12851 21607
rect 14565 21573 14599 21607
rect 15209 21573 15243 21607
rect 21833 21573 21867 21607
rect 7941 21505 7975 21539
rect 8125 21505 8159 21539
rect 11161 21505 11195 21539
rect 11345 21505 11379 21539
rect 13277 21505 13311 21539
rect 15577 21505 15611 21539
rect 16865 21505 16899 21539
rect 18061 21505 18095 21539
rect 18797 21505 18831 21539
rect 19809 21505 19843 21539
rect 22201 21505 22235 21539
rect 24225 21505 24259 21539
rect 14197 21437 14231 21471
rect 16681 21437 16715 21471
rect 19901 21437 19935 21471
rect 21649 21437 21683 21471
rect 23949 21437 23983 21471
rect 24685 21437 24719 21471
rect 7297 21369 7331 21403
rect 7665 21369 7699 21403
rect 8370 21369 8404 21403
rect 11713 21369 11747 21403
rect 13277 21369 13311 21403
rect 13369 21369 13403 21403
rect 15761 21369 15795 21403
rect 22293 21369 22327 21403
rect 22385 21369 22419 21403
rect 23213 21369 23247 21403
rect 9505 21301 9539 21335
rect 10609 21301 10643 21335
rect 11253 21301 11287 21335
rect 12265 21301 12299 21335
rect 15669 21301 15703 21335
rect 16129 21301 16163 21335
rect 19165 21301 19199 21335
rect 19809 21301 19843 21335
rect 20821 21301 20855 21335
rect 21189 21301 21223 21335
rect 22937 21301 22971 21335
rect 7389 21097 7423 21131
rect 7757 21097 7791 21131
rect 9137 21097 9171 21131
rect 10793 21097 10827 21131
rect 11253 21097 11287 21131
rect 11621 21097 11655 21131
rect 14105 21097 14139 21131
rect 15117 21097 15151 21131
rect 17601 21097 17635 21131
rect 18337 21097 18371 21131
rect 19257 21097 19291 21131
rect 20729 21097 20763 21131
rect 22017 21097 22051 21131
rect 22293 21097 22327 21131
rect 23949 21097 23983 21131
rect 8401 21029 8435 21063
rect 8585 21029 8619 21063
rect 8677 21029 8711 21063
rect 11958 21029 11992 21063
rect 17325 21029 17359 21063
rect 18153 21029 18187 21063
rect 18889 21029 18923 21063
rect 19625 21029 19659 21063
rect 21465 21029 21499 21063
rect 21557 21029 21591 21063
rect 15568 20961 15602 20995
rect 19349 20961 19383 20995
rect 22825 20961 22859 20995
rect 9689 20893 9723 20927
rect 11713 20893 11747 20927
rect 14197 20893 14231 20927
rect 15301 20893 15335 20927
rect 18429 20893 18463 20927
rect 21465 20893 21499 20927
rect 22569 20893 22603 20927
rect 25053 20893 25087 20927
rect 21005 20825 21039 20859
rect 8125 20757 8159 20791
rect 13093 20757 13127 20791
rect 13645 20757 13679 20791
rect 16681 20757 16715 20791
rect 17877 20757 17911 20791
rect 20085 20757 20119 20791
rect 8125 20553 8159 20587
rect 12081 20553 12115 20587
rect 17509 20553 17543 20587
rect 20269 20553 20303 20587
rect 15485 20485 15519 20519
rect 25513 20485 25547 20519
rect 8769 20417 8803 20451
rect 20913 20417 20947 20451
rect 12817 20349 12851 20383
rect 12909 20349 12943 20383
rect 16037 20349 16071 20383
rect 17877 20349 17911 20383
rect 18061 20349 18095 20383
rect 20637 20349 20671 20383
rect 21097 20349 21131 20383
rect 23029 20349 23063 20383
rect 23949 20349 23983 20383
rect 24133 20349 24167 20383
rect 7757 20281 7791 20315
rect 9036 20281 9070 20315
rect 13176 20281 13210 20315
rect 15761 20281 15795 20315
rect 15945 20281 15979 20315
rect 16405 20281 16439 20315
rect 18328 20281 18362 20315
rect 21342 20281 21376 20315
rect 24378 20281 24412 20315
rect 8493 20213 8527 20247
rect 10149 20213 10183 20247
rect 11713 20213 11747 20247
rect 14289 20213 14323 20247
rect 14841 20213 14875 20247
rect 15301 20213 15335 20247
rect 16957 20213 16991 20247
rect 19441 20213 19475 20247
rect 22477 20213 22511 20247
rect 23397 20213 23431 20247
rect 8769 20009 8803 20043
rect 11897 20009 11931 20043
rect 13553 20009 13587 20043
rect 15853 20009 15887 20043
rect 19349 20009 19383 20043
rect 21741 20009 21775 20043
rect 22201 20009 22235 20043
rect 16129 19941 16163 19975
rect 19165 19941 19199 19975
rect 21557 19941 21591 19975
rect 23305 19941 23339 19975
rect 24869 19941 24903 19975
rect 10517 19873 10551 19907
rect 10784 19873 10818 19907
rect 13369 19873 13403 19907
rect 16580 19873 16614 19907
rect 21833 19873 21867 19907
rect 23397 19873 23431 19907
rect 24961 19873 24995 19907
rect 13645 19805 13679 19839
rect 15301 19805 15335 19839
rect 16313 19805 16347 19839
rect 18337 19805 18371 19839
rect 18705 19805 18739 19839
rect 19441 19805 19475 19839
rect 23305 19805 23339 19839
rect 24777 19805 24811 19839
rect 13093 19737 13127 19771
rect 17693 19737 17727 19771
rect 18889 19737 18923 19771
rect 20177 19737 20211 19771
rect 21281 19737 21315 19771
rect 24409 19737 24443 19771
rect 8125 19669 8159 19703
rect 12541 19669 12575 19703
rect 14105 19669 14139 19703
rect 19809 19669 19843 19703
rect 20729 19669 20763 19703
rect 22845 19669 22879 19703
rect 23857 19669 23891 19703
rect 24133 19669 24167 19703
rect 9413 19465 9447 19499
rect 13277 19465 13311 19499
rect 19165 19465 19199 19499
rect 21465 19465 21499 19499
rect 22845 19465 22879 19499
rect 23489 19465 23523 19499
rect 25513 19465 25547 19499
rect 23949 19397 23983 19431
rect 9597 19329 9631 19363
rect 18613 19329 18647 19363
rect 21189 19329 21223 19363
rect 24133 19329 24167 19363
rect 7941 19261 7975 19295
rect 8677 19261 8711 19295
rect 9864 19261 9898 19295
rect 12265 19261 12299 19295
rect 12449 19261 12483 19295
rect 12725 19261 12759 19295
rect 13829 19261 13863 19295
rect 14096 19261 14130 19295
rect 19441 19261 19475 19295
rect 19699 19261 19733 19295
rect 21741 19261 21775 19295
rect 8401 19193 8435 19227
rect 15761 19193 15795 19227
rect 16681 19193 16715 19227
rect 16957 19193 16991 19227
rect 17325 19193 17359 19227
rect 17877 19193 17911 19227
rect 18613 19193 18647 19227
rect 18705 19193 18739 19227
rect 19993 19193 20027 19227
rect 20269 19193 20303 19227
rect 22017 19193 22051 19227
rect 22385 19193 22419 19227
rect 24378 19193 24412 19227
rect 26065 19193 26099 19227
rect 8115 19125 8149 19159
rect 8585 19125 8619 19159
rect 9137 19125 9171 19159
rect 10977 19125 11011 19159
rect 11529 19125 11563 19159
rect 13645 19125 13679 19159
rect 15209 19125 15243 19159
rect 16129 19125 16163 19159
rect 16387 19125 16421 19159
rect 16865 19125 16899 19159
rect 18135 19125 18169 19159
rect 20177 19125 20211 19159
rect 20913 19125 20947 19159
rect 21925 19125 21959 19159
rect 9413 18921 9447 18955
rect 10241 18921 10275 18955
rect 10701 18921 10735 18955
rect 13553 18921 13587 18955
rect 14197 18921 14231 18955
rect 16681 18921 16715 18955
rect 19073 18921 19107 18955
rect 21189 18921 21223 18955
rect 21649 18921 21683 18955
rect 22937 18921 22971 18955
rect 24409 18921 24443 18955
rect 10333 18853 10367 18887
rect 12633 18853 12667 18887
rect 12725 18853 12759 18887
rect 15853 18853 15887 18887
rect 20729 18853 20763 18887
rect 22385 18853 22419 18887
rect 24501 18853 24535 18887
rect 24869 18853 24903 18887
rect 15669 18785 15703 18819
rect 17397 18785 17431 18819
rect 22201 18785 22235 18819
rect 23213 18785 23247 18819
rect 24225 18785 24259 18819
rect 25421 18785 25455 18819
rect 10241 18717 10275 18751
rect 12633 18717 12667 18751
rect 14105 18717 14139 18751
rect 14289 18717 14323 18751
rect 15945 18717 15979 18751
rect 16405 18717 16439 18751
rect 17141 18717 17175 18751
rect 19809 18717 19843 18751
rect 22477 18717 22511 18751
rect 8125 18649 8159 18683
rect 9781 18649 9815 18683
rect 12173 18649 12207 18683
rect 14657 18649 14691 18683
rect 20269 18649 20303 18683
rect 21925 18649 21959 18683
rect 23581 18649 23615 18683
rect 23949 18649 23983 18683
rect 25237 18649 25271 18683
rect 11897 18581 11931 18615
rect 13093 18581 13127 18615
rect 13737 18581 13771 18615
rect 15025 18581 15059 18615
rect 15393 18581 15427 18615
rect 18521 18581 18555 18615
rect 19717 18581 19751 18615
rect 9597 18377 9631 18411
rect 10609 18377 10643 18411
rect 11253 18377 11287 18411
rect 13829 18377 13863 18411
rect 15025 18377 15059 18411
rect 18153 18377 18187 18411
rect 23121 18377 23155 18411
rect 24409 18377 24443 18411
rect 19533 18309 19567 18343
rect 23489 18309 23523 18343
rect 8677 18241 8711 18275
rect 10149 18241 10183 18275
rect 12449 18241 12483 18275
rect 19625 18241 19659 18275
rect 22385 18241 22419 18275
rect 24961 18241 24995 18275
rect 25329 18241 25363 18275
rect 9045 18173 9079 18207
rect 9873 18173 9907 18207
rect 12173 18173 12207 18207
rect 15393 18173 15427 18207
rect 15485 18173 15519 18207
rect 17877 18173 17911 18207
rect 22109 18173 22143 18207
rect 24225 18173 24259 18207
rect 24685 18173 24719 18207
rect 25697 18173 25731 18207
rect 12716 18105 12750 18139
rect 15730 18105 15764 18139
rect 18429 18105 18463 18139
rect 18613 18105 18647 18139
rect 18705 18105 18739 18139
rect 19073 18105 19107 18139
rect 19870 18105 19904 18139
rect 24869 18105 24903 18139
rect 9321 18037 9355 18071
rect 10057 18037 10091 18071
rect 11345 18037 11379 18071
rect 14565 18037 14599 18071
rect 16865 18037 16899 18071
rect 17509 18037 17543 18071
rect 21005 18037 21039 18071
rect 21925 18037 21959 18071
rect 9505 17833 9539 17867
rect 13737 17833 13771 17867
rect 14473 17833 14507 17867
rect 15853 17833 15887 17867
rect 17325 17833 17359 17867
rect 18153 17833 18187 17867
rect 19717 17833 19751 17867
rect 20269 17833 20303 17867
rect 23213 17833 23247 17867
rect 25329 17833 25363 17867
rect 10333 17765 10367 17799
rect 15025 17765 15059 17799
rect 18582 17765 18616 17799
rect 11345 17697 11379 17731
rect 11601 17697 11635 17731
rect 15669 17697 15703 17731
rect 21180 17697 21214 17731
rect 24216 17697 24250 17731
rect 10333 17629 10367 17663
rect 10425 17629 10459 17663
rect 10885 17629 10919 17663
rect 15945 17629 15979 17663
rect 17141 17629 17175 17663
rect 18337 17629 18371 17663
rect 20913 17629 20947 17663
rect 23949 17629 23983 17663
rect 9873 17561 9907 17595
rect 15393 17561 15427 17595
rect 11253 17493 11287 17527
rect 12725 17493 12759 17527
rect 13277 17493 13311 17527
rect 14105 17493 14139 17527
rect 16405 17493 16439 17527
rect 22293 17493 22327 17527
rect 22845 17493 22879 17527
rect 23765 17493 23799 17527
rect 9505 17289 9539 17323
rect 10885 17289 10919 17323
rect 12265 17289 12299 17323
rect 12541 17289 12575 17323
rect 15393 17289 15427 17323
rect 15761 17289 15795 17323
rect 17877 17289 17911 17323
rect 18613 17289 18647 17323
rect 21741 17289 21775 17323
rect 22017 17289 22051 17323
rect 14105 17221 14139 17255
rect 16497 17221 16531 17255
rect 18337 17221 18371 17255
rect 19625 17221 19659 17255
rect 20177 17221 20211 17255
rect 10701 17153 10735 17187
rect 11345 17153 11379 17187
rect 13093 17153 13127 17187
rect 14565 17153 14599 17187
rect 17049 17153 17083 17187
rect 19073 17153 19107 17187
rect 19165 17153 19199 17187
rect 20637 17153 20671 17187
rect 20729 17153 20763 17187
rect 22385 17153 22419 17187
rect 11437 17085 11471 17119
rect 13553 17085 13587 17119
rect 14657 17085 14691 17119
rect 16773 17085 16807 17119
rect 17509 17085 17543 17119
rect 23673 17085 23707 17119
rect 9873 17017 9907 17051
rect 12817 17017 12851 17051
rect 13921 17017 13955 17051
rect 14565 17017 14599 17051
rect 19073 17017 19107 17051
rect 19993 17017 20027 17051
rect 22477 17017 22511 17051
rect 22569 17017 22603 17051
rect 23918 17017 23952 17051
rect 10149 16949 10183 16983
rect 11345 16949 11379 16983
rect 11897 16949 11931 16983
rect 13001 16949 13035 16983
rect 16313 16949 16347 16983
rect 16957 16949 16991 16983
rect 20637 16949 20671 16983
rect 21189 16949 21223 16983
rect 23029 16949 23063 16983
rect 23489 16949 23523 16983
rect 25053 16949 25087 16983
rect 9955 16745 9989 16779
rect 10977 16745 11011 16779
rect 12817 16745 12851 16779
rect 15375 16745 15409 16779
rect 16773 16745 16807 16779
rect 18419 16745 18453 16779
rect 19717 16745 19751 16779
rect 21189 16745 21223 16779
rect 23949 16745 23983 16779
rect 24317 16745 24351 16779
rect 24675 16745 24709 16779
rect 10241 16677 10275 16711
rect 10425 16677 10459 16711
rect 11253 16677 11287 16711
rect 11682 16677 11716 16711
rect 14197 16677 14231 16711
rect 14749 16677 14783 16711
rect 15853 16677 15887 16711
rect 17325 16677 17359 16711
rect 18245 16677 18279 16711
rect 18889 16677 18923 16711
rect 19441 16677 19475 16711
rect 22100 16677 22134 16711
rect 25145 16677 25179 16711
rect 11437 16609 11471 16643
rect 13921 16609 13955 16643
rect 15117 16609 15151 16643
rect 15669 16609 15703 16643
rect 16497 16609 16531 16643
rect 17049 16609 17083 16643
rect 18981 16609 19015 16643
rect 21833 16609 21867 16643
rect 25237 16609 25271 16643
rect 10517 16541 10551 16575
rect 15945 16541 15979 16575
rect 18797 16541 18831 16575
rect 25145 16541 25179 16575
rect 20177 16473 20211 16507
rect 13737 16405 13771 16439
rect 17877 16405 17911 16439
rect 20453 16405 20487 16439
rect 21465 16405 21499 16439
rect 23213 16405 23247 16439
rect 9597 16201 9631 16235
rect 9965 16201 9999 16235
rect 10885 16201 10919 16235
rect 12725 16201 12759 16235
rect 13185 16201 13219 16235
rect 15025 16201 15059 16235
rect 17509 16201 17543 16235
rect 18429 16201 18463 16235
rect 19717 16201 19751 16235
rect 22477 16201 22511 16235
rect 23489 16201 23523 16235
rect 25421 16201 25455 16235
rect 25973 16201 26007 16235
rect 16497 16133 16531 16167
rect 19993 16133 20027 16167
rect 21557 16133 21591 16167
rect 10333 16065 10367 16099
rect 11437 16065 11471 16099
rect 12265 16065 12299 16099
rect 21005 16065 21039 16099
rect 22109 16065 22143 16099
rect 13645 15997 13679 16031
rect 13912 15997 13946 16031
rect 15577 15997 15611 16031
rect 18981 15997 19015 16031
rect 24041 15997 24075 16031
rect 24297 15997 24331 16031
rect 11161 15929 11195 15963
rect 16773 15929 16807 15963
rect 16957 15929 16991 15963
rect 17049 15929 17083 15963
rect 17877 15929 17911 15963
rect 18705 15929 18739 15963
rect 20269 15929 20303 15963
rect 20545 15929 20579 15963
rect 21373 15929 21407 15963
rect 21833 15929 21867 15963
rect 22017 15929 22051 15963
rect 10701 15861 10735 15895
rect 11345 15861 11379 15895
rect 11897 15861 11931 15895
rect 13553 15861 13587 15895
rect 16313 15861 16347 15895
rect 18889 15861 18923 15895
rect 19441 15861 19475 15895
rect 20453 15861 20487 15895
rect 23949 15861 23983 15895
rect 9965 15657 9999 15691
rect 13921 15657 13955 15691
rect 15117 15657 15151 15691
rect 17601 15657 17635 15691
rect 19165 15657 19199 15691
rect 23029 15657 23063 15691
rect 24041 15657 24075 15691
rect 25421 15657 25455 15691
rect 12311 15589 12345 15623
rect 18052 15589 18086 15623
rect 21465 15589 21499 15623
rect 21925 15589 21959 15623
rect 22845 15589 22879 15623
rect 24685 15589 24719 15623
rect 24869 15589 24903 15623
rect 12173 15521 12207 15555
rect 12449 15521 12483 15555
rect 15568 15521 15602 15555
rect 21281 15521 21315 15555
rect 22293 15521 22327 15555
rect 13829 15453 13863 15487
rect 14013 15453 14047 15487
rect 15301 15453 15335 15487
rect 17785 15453 17819 15487
rect 20361 15453 20395 15487
rect 20729 15453 20763 15487
rect 21557 15453 21591 15487
rect 23121 15453 23155 15487
rect 24961 15453 24995 15487
rect 10793 15385 10827 15419
rect 11897 15385 11931 15419
rect 13277 15385 13311 15419
rect 22569 15385 22603 15419
rect 13461 15317 13495 15351
rect 14381 15317 14415 15351
rect 16681 15317 16715 15351
rect 17325 15317 17359 15351
rect 19993 15317 20027 15351
rect 21005 15317 21039 15351
rect 23765 15317 23799 15351
rect 24409 15317 24443 15351
rect 11529 15113 11563 15147
rect 11897 15113 11931 15147
rect 13093 15113 13127 15147
rect 15393 15113 15427 15147
rect 16773 15113 16807 15147
rect 18797 15113 18831 15147
rect 22845 15113 22879 15147
rect 23489 15113 23523 15147
rect 25145 15113 25179 15147
rect 13645 15045 13679 15079
rect 17417 15045 17451 15079
rect 22569 15045 22603 15079
rect 23765 15045 23799 15079
rect 12173 14977 12207 15011
rect 15945 14977 15979 15011
rect 19257 14977 19291 15011
rect 19809 14977 19843 15011
rect 24225 14977 24259 15011
rect 12725 14909 12759 14943
rect 13921 14909 13955 14943
rect 15669 14909 15703 14943
rect 20269 14909 20303 14943
rect 20536 14909 20570 14943
rect 24317 14909 24351 14943
rect 14105 14841 14139 14875
rect 14197 14841 14231 14875
rect 15209 14841 15243 14875
rect 15853 14841 15887 14875
rect 16405 14841 16439 14875
rect 16865 14841 16899 14875
rect 18613 14841 18647 14875
rect 19349 14841 19383 14875
rect 13369 14773 13403 14807
rect 14841 14773 14875 14807
rect 17785 14773 17819 14807
rect 19257 14773 19291 14807
rect 20177 14773 20211 14807
rect 21649 14773 21683 14807
rect 24225 14773 24259 14807
rect 24685 14773 24719 14807
rect 25237 14773 25271 14807
rect 12633 14569 12667 14603
rect 13461 14569 13495 14603
rect 15117 14569 15151 14603
rect 16497 14569 16531 14603
rect 17693 14569 17727 14603
rect 19809 14569 19843 14603
rect 22293 14569 22327 14603
rect 22937 14569 22971 14603
rect 23305 14569 23339 14603
rect 14013 14501 14047 14535
rect 14197 14501 14231 14535
rect 15853 14501 15887 14535
rect 18052 14501 18086 14535
rect 20545 14501 20579 14535
rect 21180 14501 21214 14535
rect 24032 14501 24066 14535
rect 12725 14433 12759 14467
rect 15945 14433 15979 14467
rect 20177 14433 20211 14467
rect 23765 14433 23799 14467
rect 12633 14365 12667 14399
rect 14289 14365 14323 14399
rect 15761 14365 15795 14399
rect 17785 14365 17819 14399
rect 20913 14365 20947 14399
rect 15393 14297 15427 14331
rect 12173 14229 12207 14263
rect 13737 14229 13771 14263
rect 19165 14229 19199 14263
rect 23581 14229 23615 14263
rect 25145 14229 25179 14263
rect 11805 14025 11839 14059
rect 12173 14025 12207 14059
rect 12725 14025 12759 14059
rect 13369 14025 13403 14059
rect 13737 14025 13771 14059
rect 15209 14025 15243 14059
rect 15761 14025 15795 14059
rect 16497 14025 16531 14059
rect 17509 14025 17543 14059
rect 18429 14025 18463 14059
rect 18981 14025 19015 14059
rect 20269 14025 20303 14059
rect 20545 14025 20579 14059
rect 21557 14025 21591 14059
rect 23121 14025 23155 14059
rect 25513 14025 25547 14059
rect 22109 13957 22143 13991
rect 12817 13889 12851 13923
rect 16957 13889 16991 13923
rect 17049 13889 17083 13923
rect 19533 13889 19567 13923
rect 19993 13889 20027 13923
rect 21097 13889 21131 13923
rect 21925 13889 21959 13923
rect 22661 13889 22695 13923
rect 23489 13889 23523 13923
rect 13829 13821 13863 13855
rect 16313 13821 16347 13855
rect 18797 13821 18831 13855
rect 19257 13821 19291 13855
rect 24041 13821 24075 13855
rect 24133 13821 24167 13855
rect 24389 13821 24423 13855
rect 14096 13753 14130 13787
rect 16957 13753 16991 13787
rect 19441 13753 19475 13787
rect 20821 13753 20855 13787
rect 21005 13753 21039 13787
rect 22385 13753 22419 13787
rect 17785 13685 17819 13719
rect 22569 13685 22603 13719
rect 12817 13481 12851 13515
rect 13921 13481 13955 13515
rect 15577 13481 15611 13515
rect 16497 13481 16531 13515
rect 18153 13481 18187 13515
rect 19441 13481 19475 13515
rect 20545 13481 20579 13515
rect 21465 13481 21499 13515
rect 22109 13481 22143 13515
rect 23121 13481 23155 13515
rect 24593 13481 24627 13515
rect 11704 13413 11738 13447
rect 17325 13413 17359 13447
rect 18889 13413 18923 13447
rect 23765 13413 23799 13447
rect 23857 13413 23891 13447
rect 25145 13413 25179 13447
rect 25329 13413 25363 13447
rect 25421 13413 25455 13447
rect 18981 13345 19015 13379
rect 23581 13345 23615 13379
rect 11437 13277 11471 13311
rect 15761 13277 15795 13311
rect 17233 13277 17267 13311
rect 17417 13277 17451 13311
rect 18889 13277 18923 13311
rect 21373 13277 21407 13311
rect 21557 13277 21591 13311
rect 22477 13277 22511 13311
rect 18429 13209 18463 13243
rect 23305 13209 23339 13243
rect 24869 13209 24903 13243
rect 14289 13141 14323 13175
rect 14657 13141 14691 13175
rect 15117 13141 15151 13175
rect 16865 13141 16899 13175
rect 19809 13141 19843 13175
rect 20177 13141 20211 13175
rect 21005 13141 21039 13175
rect 24225 13141 24259 13175
rect 11161 12937 11195 12971
rect 16405 12937 16439 12971
rect 17049 12937 17083 12971
rect 19073 12937 19107 12971
rect 22661 12937 22695 12971
rect 24869 12937 24903 12971
rect 25697 12937 25731 12971
rect 17509 12869 17543 12903
rect 17785 12869 17819 12903
rect 18153 12869 18187 12903
rect 20177 12869 20211 12903
rect 21189 12869 21223 12903
rect 23765 12869 23799 12903
rect 11897 12801 11931 12835
rect 21465 12801 21499 12835
rect 21649 12801 21683 12835
rect 24225 12801 24259 12835
rect 25237 12801 25271 12835
rect 11529 12733 11563 12767
rect 12265 12733 12299 12767
rect 12449 12733 12483 12767
rect 15025 12733 15059 12767
rect 18429 12733 18463 12767
rect 20453 12733 20487 12767
rect 12694 12665 12728 12699
rect 15292 12665 15326 12699
rect 18705 12665 18739 12699
rect 19533 12665 19567 12699
rect 19809 12665 19843 12699
rect 20729 12665 20763 12699
rect 24317 12665 24351 12699
rect 13829 12597 13863 12631
rect 14933 12597 14967 12631
rect 18613 12597 18647 12631
rect 20637 12597 20671 12631
rect 22201 12597 22235 12631
rect 23121 12597 23155 12631
rect 23489 12597 23523 12631
rect 24225 12597 24259 12631
rect 17417 12393 17451 12427
rect 17785 12393 17819 12427
rect 19257 12393 19291 12427
rect 23857 12393 23891 12427
rect 24869 12393 24903 12427
rect 12265 12325 12299 12359
rect 12357 12325 12391 12359
rect 13829 12325 13863 12359
rect 18144 12325 18178 12359
rect 21465 12325 21499 12359
rect 13921 12257 13955 12291
rect 15393 12257 15427 12291
rect 15660 12257 15694 12291
rect 17877 12257 17911 12291
rect 21281 12257 21315 12291
rect 22744 12257 22778 12291
rect 12173 12189 12207 12223
rect 13737 12189 13771 12223
rect 21557 12189 21591 12223
rect 22477 12189 22511 12223
rect 13001 12121 13035 12155
rect 21005 12121 21039 12155
rect 11805 12053 11839 12087
rect 13369 12053 13403 12087
rect 14289 12053 14323 12087
rect 14749 12053 14783 12087
rect 15117 12053 15151 12087
rect 16773 12053 16807 12087
rect 20177 12053 20211 12087
rect 20729 12053 20763 12087
rect 22017 12053 22051 12087
rect 24409 12053 24443 12087
rect 25145 12053 25179 12087
rect 11805 11849 11839 11883
rect 12173 11849 12207 11883
rect 12817 11849 12851 11883
rect 14289 11849 14323 11883
rect 16221 11849 16255 11883
rect 17509 11849 17543 11883
rect 20637 11849 20671 11883
rect 21005 11849 21039 11883
rect 22477 11849 22511 11883
rect 23489 11849 23523 11883
rect 25513 11849 25547 11883
rect 13001 11781 13035 11815
rect 14933 11781 14967 11815
rect 16497 11781 16531 11815
rect 18153 11781 18187 11815
rect 13369 11713 13403 11747
rect 13553 11713 13587 11747
rect 14657 11713 14691 11747
rect 15485 11713 15519 11747
rect 16865 11713 16899 11747
rect 17049 11713 17083 11747
rect 20085 11713 20119 11747
rect 15209 11645 15243 11679
rect 21097 11645 21131 11679
rect 23029 11645 23063 11679
rect 23949 11645 23983 11679
rect 24133 11645 24167 11679
rect 24389 11645 24423 11679
rect 13921 11577 13955 11611
rect 15393 11577 15427 11611
rect 16957 11577 16991 11611
rect 18429 11577 18463 11611
rect 18613 11577 18647 11611
rect 18705 11577 18739 11611
rect 21364 11577 21398 11611
rect 11437 11509 11471 11543
rect 13461 11509 13495 11543
rect 15945 11509 15979 11543
rect 17785 11509 17819 11543
rect 19165 11509 19199 11543
rect 19441 11509 19475 11543
rect 13829 11305 13863 11339
rect 14933 11305 14967 11339
rect 16037 11305 16071 11339
rect 16405 11305 16439 11339
rect 18613 11305 18647 11339
rect 22293 11305 22327 11339
rect 22845 11305 22879 11339
rect 11437 11237 11471 11271
rect 15577 11237 15611 11271
rect 17049 11237 17083 11271
rect 20729 11237 20763 11271
rect 21180 11237 21214 11271
rect 11253 11169 11287 11203
rect 12705 11169 12739 11203
rect 16865 11169 16899 11203
rect 18429 11169 18463 11203
rect 20913 11169 20947 11203
rect 23949 11169 23983 11203
rect 24205 11169 24239 11203
rect 11529 11101 11563 11135
rect 12449 11101 12483 11135
rect 17141 11101 17175 11135
rect 18705 11101 18739 11135
rect 19809 11101 19843 11135
rect 10977 11033 11011 11067
rect 12265 11033 12299 11067
rect 16589 11033 16623 11067
rect 18153 11033 18187 11067
rect 25329 11033 25363 11067
rect 17601 10965 17635 10999
rect 17969 10965 18003 10999
rect 19073 10965 19107 10999
rect 23673 10965 23707 10999
rect 17877 10761 17911 10795
rect 18705 10761 18739 10795
rect 21557 10761 21591 10795
rect 22477 10761 22511 10795
rect 23121 10761 23155 10795
rect 24777 10761 24811 10795
rect 16497 10693 16531 10727
rect 18337 10693 18371 10727
rect 20361 10693 20395 10727
rect 21281 10693 21315 10727
rect 23765 10693 23799 10727
rect 15945 10625 15979 10659
rect 17049 10625 17083 10659
rect 17417 10625 17451 10659
rect 18981 10625 19015 10659
rect 21925 10625 21959 10659
rect 23489 10625 23523 10659
rect 24133 10625 24167 10659
rect 10609 10557 10643 10591
rect 12725 10557 12759 10591
rect 13185 10557 13219 10591
rect 13277 10557 13311 10591
rect 13544 10557 13578 10591
rect 24317 10557 24351 10591
rect 25237 10557 25271 10591
rect 25789 10557 25823 10591
rect 11345 10489 11379 10523
rect 16313 10489 16347 10523
rect 16773 10489 16807 10523
rect 16957 10489 16991 10523
rect 19226 10489 19260 10523
rect 20913 10489 20947 10523
rect 22109 10489 22143 10523
rect 10977 10421 11011 10455
rect 12173 10421 12207 10455
rect 14657 10421 14691 10455
rect 15577 10421 15611 10455
rect 22017 10421 22051 10455
rect 24225 10421 24259 10455
rect 25421 10421 25455 10455
rect 10977 10217 11011 10251
rect 13553 10217 13587 10251
rect 15853 10217 15887 10251
rect 17325 10217 17359 10251
rect 18981 10217 19015 10251
rect 21465 10217 21499 10251
rect 23029 10217 23063 10251
rect 14013 10149 14047 10183
rect 18797 10149 18831 10183
rect 20729 10149 20763 10183
rect 21557 10149 21591 10183
rect 23673 10149 23707 10183
rect 24409 10149 24443 10183
rect 24593 10149 24627 10183
rect 16212 10081 16246 10115
rect 18245 10081 18279 10115
rect 19073 10081 19107 10115
rect 21925 10081 21959 10115
rect 22845 10081 22879 10115
rect 13553 10013 13587 10047
rect 13645 10013 13679 10047
rect 15945 10013 15979 10047
rect 21465 10013 21499 10047
rect 22385 10013 22419 10047
rect 23121 10013 23155 10047
rect 24685 10013 24719 10047
rect 18521 9945 18555 9979
rect 13093 9877 13127 9911
rect 19441 9877 19475 9911
rect 21005 9877 21039 9911
rect 22569 9877 22603 9911
rect 24133 9877 24167 9911
rect 25237 9877 25271 9911
rect 15853 9673 15887 9707
rect 16865 9673 16899 9707
rect 17417 9673 17451 9707
rect 19441 9673 19475 9707
rect 21557 9673 21591 9707
rect 23121 9673 23155 9707
rect 12725 9605 12759 9639
rect 13001 9605 13035 9639
rect 13921 9605 13955 9639
rect 16405 9605 16439 9639
rect 17785 9605 17819 9639
rect 19993 9605 20027 9639
rect 20545 9605 20579 9639
rect 21833 9605 21867 9639
rect 22109 9605 22143 9639
rect 23765 9605 23799 9639
rect 25789 9605 25823 9639
rect 13369 9537 13403 9571
rect 13553 9537 13587 9571
rect 16957 9537 16991 9571
rect 20821 9537 20855 9571
rect 22569 9537 22603 9571
rect 24685 9537 24719 9571
rect 12265 9469 12299 9503
rect 14381 9469 14415 9503
rect 14473 9469 14507 9503
rect 14740 9469 14774 9503
rect 18061 9469 18095 9503
rect 18317 9469 18351 9503
rect 24041 9469 24075 9503
rect 25237 9469 25271 9503
rect 13461 9401 13495 9435
rect 22569 9401 22603 9435
rect 22661 9401 22695 9435
rect 24317 9401 24351 9435
rect 25053 9401 25087 9435
rect 21005 9333 21039 9367
rect 23489 9333 23523 9367
rect 24225 9333 24259 9367
rect 25421 9333 25455 9367
rect 13369 9129 13403 9163
rect 13737 9129 13771 9163
rect 14565 9129 14599 9163
rect 16865 9129 16899 9163
rect 18061 9129 18095 9163
rect 20361 9129 20395 9163
rect 20729 9129 20763 9163
rect 22109 9129 22143 9163
rect 23765 9129 23799 9163
rect 24317 9129 24351 9163
rect 24685 9129 24719 9163
rect 25421 9129 25455 9163
rect 13093 9061 13127 9095
rect 16681 9061 16715 9095
rect 16957 9061 16991 9095
rect 18582 9061 18616 9095
rect 25237 9061 25271 9095
rect 21281 8993 21315 9027
rect 22385 8993 22419 9027
rect 22652 8993 22686 9027
rect 18337 8925 18371 8959
rect 25513 8925 25547 8959
rect 16405 8789 16439 8823
rect 19717 8789 19751 8823
rect 21189 8789 21223 8823
rect 21465 8789 21499 8823
rect 24961 8789 24995 8823
rect 16497 8585 16531 8619
rect 17417 8585 17451 8619
rect 17877 8585 17911 8619
rect 19073 8585 19107 8619
rect 22477 8585 22511 8619
rect 25973 8585 26007 8619
rect 15945 8517 15979 8551
rect 19349 8517 19383 8551
rect 19625 8517 19659 8551
rect 23029 8517 23063 8551
rect 23397 8517 23431 8551
rect 25697 8517 25731 8551
rect 15577 8449 15611 8483
rect 17049 8449 17083 8483
rect 18337 8449 18371 8483
rect 19993 8449 20027 8483
rect 23673 8449 23707 8483
rect 18521 8381 18555 8415
rect 21097 8381 21131 8415
rect 23929 8381 23963 8415
rect 16313 8313 16347 8347
rect 16773 8313 16807 8347
rect 16957 8313 16991 8347
rect 20085 8313 20119 8347
rect 20177 8313 20211 8347
rect 21342 8313 21376 8347
rect 26341 8313 26375 8347
rect 20637 8245 20671 8279
rect 20913 8245 20947 8279
rect 25053 8245 25087 8279
rect 16497 8041 16531 8075
rect 16865 8041 16899 8075
rect 22845 8041 22879 8075
rect 23765 8041 23799 8075
rect 19625 7973 19659 8007
rect 19809 7973 19843 8007
rect 23397 7973 23431 8007
rect 17969 7905 18003 7939
rect 18705 7905 18739 7939
rect 19901 7905 19935 7939
rect 21180 7905 21214 7939
rect 23949 7905 23983 7939
rect 24216 7905 24250 7939
rect 16957 7837 16991 7871
rect 18245 7837 18279 7871
rect 20913 7837 20947 7871
rect 14657 7701 14691 7735
rect 19349 7701 19383 7735
rect 20545 7701 20579 7735
rect 22293 7701 22327 7735
rect 25329 7701 25363 7735
rect 14381 7497 14415 7531
rect 15853 7497 15887 7531
rect 19441 7497 19475 7531
rect 21557 7497 21591 7531
rect 21925 7497 21959 7531
rect 23489 7497 23523 7531
rect 14657 7429 14691 7463
rect 16497 7429 16531 7463
rect 20637 7429 20671 7463
rect 24041 7429 24075 7463
rect 20453 7361 20487 7395
rect 21189 7361 21223 7395
rect 22569 7361 22603 7395
rect 24501 7361 24535 7395
rect 25053 7361 25087 7395
rect 14933 7293 14967 7327
rect 17877 7293 17911 7327
rect 18061 7293 18095 7327
rect 20913 7293 20947 7327
rect 22293 7293 22327 7327
rect 24593 7293 24627 7327
rect 25513 7293 25547 7327
rect 26065 7293 26099 7327
rect 15117 7225 15151 7259
rect 15209 7225 15243 7259
rect 16773 7225 16807 7259
rect 16957 7225 16991 7259
rect 17049 7225 17083 7259
rect 18306 7225 18340 7259
rect 21097 7225 21131 7259
rect 23121 7225 23155 7259
rect 16221 7157 16255 7191
rect 17509 7157 17543 7191
rect 20085 7157 20119 7191
rect 24501 7157 24535 7191
rect 25329 7157 25363 7191
rect 25697 7157 25731 7191
rect 14657 6953 14691 6987
rect 18153 6953 18187 6987
rect 19533 6953 19567 6987
rect 19993 6953 20027 6987
rect 23213 6953 23247 6987
rect 24685 6953 24719 6987
rect 19027 6885 19061 6919
rect 23857 6885 23891 6919
rect 25421 6885 25455 6919
rect 8033 6817 8067 6851
rect 16304 6817 16338 6851
rect 18889 6817 18923 6851
rect 20545 6817 20579 6851
rect 20913 6817 20947 6851
rect 21465 6817 21499 6851
rect 22017 6817 22051 6851
rect 22753 6817 22787 6851
rect 25237 6817 25271 6851
rect 16037 6749 16071 6783
rect 19165 6749 19199 6783
rect 22201 6749 22235 6783
rect 23765 6749 23799 6783
rect 23949 6749 23983 6783
rect 25513 6749 25547 6783
rect 8217 6681 8251 6715
rect 17417 6681 17451 6715
rect 18613 6681 18647 6715
rect 24961 6681 24995 6715
rect 21097 6613 21131 6647
rect 23397 6613 23431 6647
rect 24317 6613 24351 6647
rect 14565 6409 14599 6443
rect 16681 6409 16715 6443
rect 17877 6409 17911 6443
rect 19441 6409 19475 6443
rect 20085 6409 20119 6443
rect 21925 6409 21959 6443
rect 22937 6409 22971 6443
rect 23305 6409 23339 6443
rect 24041 6409 24075 6443
rect 26065 6409 26099 6443
rect 13645 6273 13679 6307
rect 14657 6273 14691 6307
rect 18061 6273 18095 6307
rect 24133 6273 24167 6307
rect 13369 6205 13403 6239
rect 20361 6205 20395 6239
rect 20545 6205 20579 6239
rect 22661 6205 22695 6239
rect 24400 6205 24434 6239
rect 14924 6137 14958 6171
rect 16957 6137 16991 6171
rect 18306 6137 18340 6171
rect 20812 6137 20846 6171
rect 8125 6069 8159 6103
rect 14197 6069 14231 6103
rect 16037 6069 16071 6103
rect 25513 6069 25547 6103
rect 18153 5865 18187 5899
rect 18521 5865 18555 5899
rect 19257 5865 19291 5899
rect 19901 5865 19935 5899
rect 20637 5865 20671 5899
rect 22293 5865 22327 5899
rect 25329 5865 25363 5899
rect 14197 5797 14231 5831
rect 15568 5797 15602 5831
rect 18981 5797 19015 5831
rect 14289 5729 14323 5763
rect 14657 5729 14691 5763
rect 19717 5729 19751 5763
rect 20913 5729 20947 5763
rect 21180 5729 21214 5763
rect 23397 5729 23431 5763
rect 23664 5729 23698 5763
rect 14197 5661 14231 5695
rect 15301 5661 15335 5695
rect 13737 5593 13771 5627
rect 15025 5593 15059 5627
rect 16681 5525 16715 5559
rect 24777 5525 24811 5559
rect 13277 5321 13311 5355
rect 14197 5321 14231 5355
rect 14473 5321 14507 5355
rect 15853 5321 15887 5355
rect 20545 5321 20579 5355
rect 23029 5321 23063 5355
rect 16037 5253 16071 5287
rect 19809 5253 19843 5287
rect 23489 5253 23523 5287
rect 23765 5253 23799 5287
rect 24685 5253 24719 5287
rect 13369 5185 13403 5219
rect 14841 5185 14875 5219
rect 15485 5185 15519 5219
rect 15577 5185 15611 5219
rect 16497 5185 16531 5219
rect 19349 5185 19383 5219
rect 21005 5185 21039 5219
rect 24225 5185 24259 5219
rect 25053 5185 25087 5219
rect 25421 5185 25455 5219
rect 18613 5117 18647 5151
rect 18889 5117 18923 5151
rect 20269 5117 20303 5151
rect 20729 5117 20763 5151
rect 22477 5117 22511 5151
rect 25237 5117 25271 5151
rect 25973 5117 26007 5151
rect 14933 5049 14967 5083
rect 15025 5049 15059 5083
rect 15577 5049 15611 5083
rect 16589 5049 16623 5083
rect 22293 5049 22327 5083
rect 24317 5049 24351 5083
rect 13921 4981 13955 5015
rect 16497 4981 16531 5015
rect 16957 4981 16991 5015
rect 21557 4981 21591 5015
rect 22661 4981 22695 5015
rect 24225 4981 24259 5015
rect 14841 4777 14875 4811
rect 16221 4777 16255 4811
rect 23857 4777 23891 4811
rect 24317 4777 24351 4811
rect 14473 4709 14507 4743
rect 15853 4709 15887 4743
rect 23949 4709 23983 4743
rect 13369 4641 13403 4675
rect 15301 4641 15335 4675
rect 19809 4641 19843 4675
rect 21833 4641 21867 4675
rect 23673 4641 23707 4675
rect 24869 4641 24903 4675
rect 23397 4505 23431 4539
rect 13553 4437 13587 4471
rect 15485 4437 15519 4471
rect 22017 4437 22051 4471
rect 25053 4437 25087 4471
rect 21833 4233 21867 4267
rect 23857 4233 23891 4267
rect 13277 4097 13311 4131
rect 15301 4097 15335 4131
rect 19349 4097 19383 4131
rect 23305 4097 23339 4131
rect 25973 4097 26007 4131
rect 13369 4029 13403 4063
rect 14749 4029 14783 4063
rect 15853 4029 15887 4063
rect 16589 4029 16623 4063
rect 18705 4029 18739 4063
rect 19809 4029 19843 4063
rect 20361 4029 20395 4063
rect 20913 4029 20947 4063
rect 21465 4029 21499 4063
rect 22385 4029 22419 4063
rect 22477 4029 22511 4063
rect 24317 4029 24351 4063
rect 24869 4029 24903 4063
rect 25237 4029 25271 4063
rect 25421 4029 25455 4063
rect 13645 3961 13679 3995
rect 16129 3961 16163 3995
rect 14105 3893 14139 3927
rect 14933 3893 14967 3927
rect 15669 3893 15703 3927
rect 18889 3893 18923 3927
rect 19993 3893 20027 3927
rect 21097 3893 21131 3927
rect 22661 3893 22695 3927
rect 24501 3893 24535 3927
rect 25605 3893 25639 3927
rect 18521 3689 18555 3723
rect 20453 3689 20487 3723
rect 23949 3689 23983 3723
rect 13645 3621 13679 3655
rect 10241 3553 10275 3587
rect 12265 3553 12299 3587
rect 13369 3553 13403 3587
rect 15945 3553 15979 3587
rect 17233 3553 17267 3587
rect 18337 3553 18371 3587
rect 19441 3553 19475 3587
rect 20913 3553 20947 3587
rect 22017 3553 22051 3587
rect 23121 3553 23155 3587
rect 23397 3553 23431 3587
rect 24593 3553 24627 3587
rect 10517 3485 10551 3519
rect 16129 3485 16163 3519
rect 19625 3485 19659 3519
rect 12449 3349 12483 3383
rect 17417 3349 17451 3383
rect 21097 3349 21131 3383
rect 22201 3349 22235 3383
rect 24777 3349 24811 3383
rect 10241 3145 10275 3179
rect 14013 3145 14047 3179
rect 16037 3145 16071 3179
rect 16681 3145 16715 3179
rect 17417 3145 17451 3179
rect 18337 3145 18371 3179
rect 18705 3145 18739 3179
rect 19441 3145 19475 3179
rect 20269 3145 20303 3179
rect 21189 3145 21223 3179
rect 23121 3145 23155 3179
rect 23397 3145 23431 3179
rect 24409 3145 24443 3179
rect 24777 3145 24811 3179
rect 13645 3077 13679 3111
rect 13185 3009 13219 3043
rect 22109 3009 22143 3043
rect 23857 3009 23891 3043
rect 8677 2941 8711 2975
rect 9413 2941 9447 2975
rect 10885 2941 10919 2975
rect 11621 2941 11655 2975
rect 12909 2941 12943 2975
rect 14841 2941 14875 2975
rect 15577 2941 15611 2975
rect 16865 2941 16899 2975
rect 18153 2941 18187 2975
rect 19257 2941 19291 2975
rect 19809 2941 19843 2975
rect 20361 2941 20395 2975
rect 22293 2941 22327 2975
rect 23673 2941 23707 2975
rect 24961 2941 24995 2975
rect 25513 2941 25547 2975
rect 8953 2873 8987 2907
rect 11161 2873 11195 2907
rect 12725 2873 12759 2907
rect 15117 2873 15151 2907
rect 17785 2873 17819 2907
rect 20637 2873 20671 2907
rect 22569 2873 22603 2907
rect 17049 2805 17083 2839
rect 25145 2805 25179 2839
rect 14933 2601 14967 2635
rect 16221 2601 16255 2635
rect 17785 2601 17819 2635
rect 18797 2601 18831 2635
rect 20269 2601 20303 2635
rect 22385 2601 22419 2635
rect 23029 2601 23063 2635
rect 11161 2465 11195 2499
rect 11713 2465 11747 2499
rect 12633 2465 12667 2499
rect 13185 2465 13219 2499
rect 14289 2465 14323 2499
rect 16037 2465 16071 2499
rect 16589 2465 16623 2499
rect 17141 2465 17175 2499
rect 18613 2465 18647 2499
rect 19165 2465 19199 2499
rect 19717 2465 19751 2499
rect 21741 2465 21775 2499
rect 22845 2465 22879 2499
rect 23397 2465 23431 2499
rect 24593 2465 24627 2499
rect 25145 2465 25179 2499
rect 12817 2329 12851 2363
rect 14473 2329 14507 2363
rect 17325 2329 17359 2363
rect 19901 2329 19935 2363
rect 11345 2261 11379 2295
rect 21925 2261 21959 2295
rect 24777 2261 24811 2295
<< metal1 >>
rect 12986 27412 12992 27464
rect 13044 27452 13050 27464
rect 13170 27452 13176 27464
rect 13044 27424 13176 27452
rect 13044 27412 13050 27424
rect 13170 27412 13176 27424
rect 13228 27412 13234 27464
rect 22186 26256 22192 26308
rect 22244 26296 22250 26308
rect 24578 26296 24584 26308
rect 22244 26268 24584 26296
rect 22244 26256 22250 26268
rect 24578 26256 24584 26268
rect 24636 26256 24642 26308
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 13173 25483 13231 25489
rect 13173 25449 13185 25483
rect 13219 25480 13231 25483
rect 15930 25480 15936 25492
rect 13219 25452 15936 25480
rect 13219 25449 13231 25452
rect 13173 25443 13231 25449
rect 15930 25440 15936 25452
rect 15988 25440 15994 25492
rect 19337 25483 19395 25489
rect 19337 25449 19349 25483
rect 19383 25480 19395 25483
rect 20070 25480 20076 25492
rect 19383 25452 20076 25480
rect 19383 25449 19395 25452
rect 19337 25443 19395 25449
rect 20070 25440 20076 25452
rect 20128 25440 20134 25492
rect 9950 25372 9956 25424
rect 10008 25412 10014 25424
rect 10505 25415 10563 25421
rect 10505 25412 10517 25415
rect 10008 25384 10517 25412
rect 10008 25372 10014 25384
rect 10505 25381 10517 25384
rect 10551 25381 10563 25415
rect 10505 25375 10563 25381
rect 10318 25344 10324 25356
rect 10279 25316 10324 25344
rect 10318 25304 10324 25316
rect 10376 25304 10382 25356
rect 12710 25304 12716 25356
rect 12768 25344 12774 25356
rect 12989 25347 13047 25353
rect 12989 25344 13001 25347
rect 12768 25316 13001 25344
rect 12768 25304 12774 25316
rect 12989 25313 13001 25316
rect 13035 25313 13047 25347
rect 19150 25344 19156 25356
rect 19111 25316 19156 25344
rect 12989 25307 13047 25313
rect 19150 25304 19156 25316
rect 19208 25304 19214 25356
rect 19797 25347 19855 25353
rect 19797 25313 19809 25347
rect 19843 25344 19855 25347
rect 19978 25344 19984 25356
rect 19843 25316 19984 25344
rect 19843 25313 19855 25316
rect 19797 25307 19855 25313
rect 19978 25304 19984 25316
rect 20036 25344 20042 25356
rect 24762 25344 24768 25356
rect 20036 25316 24768 25344
rect 20036 25304 20042 25316
rect 24762 25304 24768 25316
rect 24820 25304 24826 25356
rect 9858 25236 9864 25288
rect 9916 25276 9922 25288
rect 10597 25279 10655 25285
rect 10597 25276 10609 25279
rect 9916 25248 10609 25276
rect 9916 25236 9922 25248
rect 10597 25245 10609 25248
rect 10643 25245 10655 25279
rect 11054 25276 11060 25288
rect 10597 25239 10655 25245
rect 10796 25248 11060 25276
rect 10045 25211 10103 25217
rect 10045 25177 10057 25211
rect 10091 25208 10103 25211
rect 10796 25208 10824 25248
rect 11054 25236 11060 25248
rect 11112 25236 11118 25288
rect 15933 25279 15991 25285
rect 15933 25245 15945 25279
rect 15979 25276 15991 25279
rect 16206 25276 16212 25288
rect 15979 25248 16212 25276
rect 15979 25245 15991 25248
rect 15933 25239 15991 25245
rect 16206 25236 16212 25248
rect 16264 25236 16270 25288
rect 10091 25180 10824 25208
rect 10091 25177 10103 25180
rect 10045 25171 10103 25177
rect 10870 25168 10876 25220
rect 10928 25208 10934 25220
rect 10928 25180 11468 25208
rect 10928 25168 10934 25180
rect 11057 25143 11115 25149
rect 11057 25109 11069 25143
rect 11103 25140 11115 25143
rect 11238 25140 11244 25152
rect 11103 25112 11244 25140
rect 11103 25109 11115 25112
rect 11057 25103 11115 25109
rect 11238 25100 11244 25112
rect 11296 25100 11302 25152
rect 11440 25149 11468 25180
rect 11425 25143 11483 25149
rect 11425 25109 11437 25143
rect 11471 25140 11483 25143
rect 12434 25140 12440 25152
rect 11471 25112 12440 25140
rect 11471 25109 11483 25112
rect 11425 25103 11483 25109
rect 12434 25100 12440 25112
rect 12492 25100 12498 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 12710 24896 12716 24948
rect 12768 24936 12774 24948
rect 14001 24939 14059 24945
rect 14001 24936 14013 24939
rect 12768 24908 14013 24936
rect 12768 24896 12774 24908
rect 14001 24905 14013 24908
rect 14047 24905 14059 24939
rect 14001 24899 14059 24905
rect 6917 24871 6975 24877
rect 6917 24837 6929 24871
rect 6963 24837 6975 24871
rect 9950 24868 9956 24880
rect 9911 24840 9956 24868
rect 6917 24831 6975 24837
rect 5994 24760 6000 24812
rect 6052 24800 6058 24812
rect 6549 24803 6607 24809
rect 6549 24800 6561 24803
rect 6052 24772 6561 24800
rect 6052 24760 6058 24772
rect 6549 24769 6561 24772
rect 6595 24769 6607 24803
rect 6932 24800 6960 24831
rect 9950 24828 9956 24840
rect 10008 24828 10014 24880
rect 10318 24868 10324 24880
rect 10279 24840 10324 24868
rect 10318 24828 10324 24840
rect 10376 24828 10382 24880
rect 10597 24871 10655 24877
rect 10597 24837 10609 24871
rect 10643 24868 10655 24871
rect 10778 24868 10784 24880
rect 10643 24840 10784 24868
rect 10643 24837 10655 24840
rect 10597 24831 10655 24837
rect 10778 24828 10784 24840
rect 10836 24828 10842 24880
rect 13081 24871 13139 24877
rect 13081 24837 13093 24871
rect 13127 24837 13139 24871
rect 13081 24831 13139 24837
rect 19613 24871 19671 24877
rect 19613 24837 19625 24871
rect 19659 24837 19671 24871
rect 23566 24868 23572 24880
rect 19613 24831 19671 24837
rect 22112 24840 23572 24868
rect 7837 24803 7895 24809
rect 7837 24800 7849 24803
rect 6932 24772 7849 24800
rect 6549 24763 6607 24769
rect 7837 24769 7849 24772
rect 7883 24800 7895 24803
rect 8294 24800 8300 24812
rect 7883 24772 8300 24800
rect 7883 24769 7895 24772
rect 7837 24763 7895 24769
rect 6564 24732 6592 24763
rect 8294 24760 8300 24772
rect 8352 24760 8358 24812
rect 12253 24803 12311 24809
rect 12253 24769 12265 24803
rect 12299 24800 12311 24803
rect 13096 24800 13124 24831
rect 13998 24800 14004 24812
rect 12299 24772 13032 24800
rect 13096 24772 14004 24800
rect 12299 24769 12311 24772
rect 12253 24763 12311 24769
rect 10870 24732 10876 24744
rect 6564 24704 7420 24732
rect 10831 24704 10876 24732
rect 7190 24664 7196 24676
rect 7151 24636 7196 24664
rect 7190 24624 7196 24636
rect 7248 24624 7254 24676
rect 7392 24673 7420 24704
rect 10870 24692 10876 24704
rect 10928 24692 10934 24744
rect 11517 24735 11575 24741
rect 11517 24732 11529 24735
rect 11072 24704 11529 24732
rect 11072 24676 11100 24704
rect 11517 24701 11529 24704
rect 11563 24701 11575 24735
rect 13004 24732 13032 24772
rect 13998 24760 14004 24772
rect 14056 24760 14062 24812
rect 19518 24760 19524 24812
rect 19576 24800 19582 24812
rect 19628 24800 19656 24831
rect 19978 24800 19984 24812
rect 19576 24772 19656 24800
rect 19939 24772 19984 24800
rect 19576 24760 19582 24772
rect 19978 24760 19984 24772
rect 20036 24760 20042 24812
rect 21542 24760 21548 24812
rect 21600 24800 21606 24812
rect 22112 24800 22140 24840
rect 22480 24812 22508 24840
rect 23566 24828 23572 24840
rect 23624 24828 23630 24880
rect 21600 24772 22140 24800
rect 21600 24760 21606 24772
rect 22462 24760 22468 24812
rect 22520 24760 22526 24812
rect 14553 24735 14611 24741
rect 13004 24704 13492 24732
rect 11517 24695 11575 24701
rect 7377 24667 7435 24673
rect 7377 24633 7389 24667
rect 7423 24633 7435 24667
rect 7377 24627 7435 24633
rect 7469 24667 7527 24673
rect 7469 24633 7481 24667
rect 7515 24633 7527 24667
rect 11054 24664 11060 24676
rect 11015 24636 11060 24664
rect 7469 24627 7527 24633
rect 6273 24599 6331 24605
rect 6273 24565 6285 24599
rect 6319 24596 6331 24599
rect 7484 24596 7512 24627
rect 11054 24624 11060 24636
rect 11112 24624 11118 24676
rect 11149 24667 11207 24673
rect 11149 24633 11161 24667
rect 11195 24664 11207 24667
rect 11238 24664 11244 24676
rect 11195 24636 11244 24664
rect 11195 24633 11207 24636
rect 11149 24627 11207 24633
rect 11238 24624 11244 24636
rect 11296 24664 11302 24676
rect 11974 24664 11980 24676
rect 11296 24636 11980 24664
rect 11296 24624 11302 24636
rect 11974 24624 11980 24636
rect 12032 24624 12038 24676
rect 13078 24624 13084 24676
rect 13136 24664 13142 24676
rect 13357 24667 13415 24673
rect 13357 24664 13369 24667
rect 13136 24636 13369 24664
rect 13136 24624 13142 24636
rect 13357 24633 13369 24636
rect 13403 24633 13415 24667
rect 13464 24664 13492 24704
rect 14553 24701 14565 24735
rect 14599 24732 14611 24735
rect 15657 24735 15715 24741
rect 14599 24704 15240 24732
rect 14599 24701 14611 24704
rect 14553 24695 14611 24701
rect 13633 24667 13691 24673
rect 13633 24664 13645 24667
rect 13464 24636 13645 24664
rect 13357 24627 13415 24633
rect 13633 24633 13645 24636
rect 13679 24664 13691 24667
rect 14090 24664 14096 24676
rect 13679 24636 14096 24664
rect 13679 24633 13691 24636
rect 13633 24627 13691 24633
rect 14090 24624 14096 24636
rect 14148 24624 14154 24676
rect 7558 24596 7564 24608
rect 6319 24568 7564 24596
rect 6319 24565 6331 24568
rect 6273 24559 6331 24565
rect 7558 24556 7564 24568
rect 7616 24556 7622 24608
rect 9677 24599 9735 24605
rect 9677 24565 9689 24599
rect 9723 24596 9735 24599
rect 9858 24596 9864 24608
rect 9723 24568 9864 24596
rect 9723 24565 9735 24568
rect 9677 24559 9735 24565
rect 9858 24556 9864 24568
rect 9916 24556 9922 24608
rect 10042 24556 10048 24608
rect 10100 24596 10106 24608
rect 12805 24599 12863 24605
rect 12805 24596 12817 24599
rect 10100 24568 12817 24596
rect 10100 24556 10106 24568
rect 12805 24565 12817 24568
rect 12851 24596 12863 24599
rect 13541 24599 13599 24605
rect 13541 24596 13553 24599
rect 12851 24568 13553 24596
rect 12851 24565 12863 24568
rect 12805 24559 12863 24565
rect 13541 24565 13553 24568
rect 13587 24565 13599 24599
rect 13541 24559 13599 24565
rect 14550 24556 14556 24608
rect 14608 24596 14614 24608
rect 15212 24605 15240 24704
rect 15657 24701 15669 24735
rect 15703 24732 15715 24735
rect 16298 24732 16304 24744
rect 15703 24704 16304 24732
rect 15703 24701 15715 24704
rect 15657 24695 15715 24701
rect 16298 24692 16304 24704
rect 16356 24692 16362 24744
rect 16761 24735 16819 24741
rect 16761 24701 16773 24735
rect 16807 24732 16819 24735
rect 17313 24735 17371 24741
rect 17313 24732 17325 24735
rect 16807 24704 17325 24732
rect 16807 24701 16819 24704
rect 16761 24695 16819 24701
rect 17313 24701 17325 24704
rect 17359 24732 17371 24735
rect 17770 24732 17776 24744
rect 17359 24704 17776 24732
rect 17359 24701 17371 24704
rect 17313 24695 17371 24701
rect 17770 24692 17776 24704
rect 17828 24692 17834 24744
rect 18417 24735 18475 24741
rect 18417 24701 18429 24735
rect 18463 24732 18475 24735
rect 18506 24732 18512 24744
rect 18463 24704 18512 24732
rect 18463 24701 18475 24704
rect 18417 24695 18475 24701
rect 18506 24692 18512 24704
rect 18564 24732 18570 24744
rect 18969 24735 19027 24741
rect 18969 24732 18981 24735
rect 18564 24704 18981 24732
rect 18564 24692 18570 24704
rect 18969 24701 18981 24704
rect 19015 24701 19027 24735
rect 18969 24695 19027 24701
rect 20898 24692 20904 24744
rect 20956 24732 20962 24744
rect 21085 24735 21143 24741
rect 21085 24732 21097 24735
rect 20956 24704 21097 24732
rect 20956 24692 20962 24704
rect 21085 24701 21097 24704
rect 21131 24732 21143 24735
rect 21637 24735 21695 24741
rect 21637 24732 21649 24735
rect 21131 24704 21649 24732
rect 21131 24701 21143 24704
rect 21085 24695 21143 24701
rect 21637 24701 21649 24704
rect 21683 24701 21695 24735
rect 21637 24695 21695 24701
rect 22189 24735 22247 24741
rect 22189 24701 22201 24735
rect 22235 24732 22247 24735
rect 22278 24732 22284 24744
rect 22235 24704 22284 24732
rect 22235 24701 22247 24704
rect 22189 24695 22247 24701
rect 22278 24692 22284 24704
rect 22336 24732 22342 24744
rect 22741 24735 22799 24741
rect 22741 24732 22753 24735
rect 22336 24704 22753 24732
rect 22336 24692 22342 24704
rect 22741 24701 22753 24704
rect 22787 24701 22799 24735
rect 22741 24695 22799 24701
rect 16482 24664 16488 24676
rect 15856 24636 16488 24664
rect 14737 24599 14795 24605
rect 14737 24596 14749 24599
rect 14608 24568 14749 24596
rect 14608 24556 14614 24568
rect 14737 24565 14749 24568
rect 14783 24565 14795 24599
rect 14737 24559 14795 24565
rect 15197 24599 15255 24605
rect 15197 24565 15209 24599
rect 15243 24596 15255 24599
rect 15470 24596 15476 24608
rect 15243 24568 15476 24596
rect 15243 24565 15255 24568
rect 15197 24559 15255 24565
rect 15470 24556 15476 24568
rect 15528 24556 15534 24608
rect 15856 24605 15884 24636
rect 16482 24624 16488 24636
rect 16540 24624 16546 24676
rect 18325 24667 18383 24673
rect 18325 24633 18337 24667
rect 18371 24664 18383 24667
rect 19150 24664 19156 24676
rect 18371 24636 19156 24664
rect 18371 24633 18383 24636
rect 18325 24627 18383 24633
rect 19150 24624 19156 24636
rect 19208 24624 19214 24676
rect 20165 24667 20223 24673
rect 20165 24633 20177 24667
rect 20211 24664 20223 24667
rect 23382 24664 23388 24676
rect 20211 24636 20392 24664
rect 20211 24633 20223 24636
rect 20165 24627 20223 24633
rect 20364 24608 20392 24636
rect 22388 24636 23388 24664
rect 15841 24599 15899 24605
rect 15841 24565 15853 24599
rect 15887 24565 15899 24599
rect 16298 24596 16304 24608
rect 16259 24568 16304 24596
rect 15841 24559 15899 24565
rect 16298 24556 16304 24568
rect 16356 24556 16362 24608
rect 16945 24599 17003 24605
rect 16945 24565 16957 24599
rect 16991 24596 17003 24599
rect 17862 24596 17868 24608
rect 16991 24568 17868 24596
rect 16991 24565 17003 24568
rect 16945 24559 17003 24565
rect 17862 24556 17868 24568
rect 17920 24556 17926 24608
rect 18598 24596 18604 24608
rect 18559 24568 18604 24596
rect 18598 24556 18604 24568
rect 18656 24556 18662 24608
rect 19426 24596 19432 24608
rect 19339 24568 19432 24596
rect 19426 24556 19432 24568
rect 19484 24596 19490 24608
rect 20070 24596 20076 24608
rect 19484 24568 20076 24596
rect 19484 24556 19490 24568
rect 20070 24556 20076 24568
rect 20128 24556 20134 24608
rect 20346 24556 20352 24608
rect 20404 24596 20410 24608
rect 20533 24599 20591 24605
rect 20533 24596 20545 24599
rect 20404 24568 20545 24596
rect 20404 24556 20410 24568
rect 20533 24565 20545 24568
rect 20579 24565 20591 24599
rect 20533 24559 20591 24565
rect 21269 24599 21327 24605
rect 21269 24565 21281 24599
rect 21315 24596 21327 24599
rect 21358 24596 21364 24608
rect 21315 24568 21364 24596
rect 21315 24565 21327 24568
rect 21269 24559 21327 24565
rect 21358 24556 21364 24568
rect 21416 24556 21422 24608
rect 22388 24605 22416 24636
rect 23382 24624 23388 24636
rect 23440 24624 23446 24676
rect 22373 24599 22431 24605
rect 22373 24565 22385 24599
rect 22419 24565 22431 24599
rect 22373 24559 22431 24565
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 6362 24352 6368 24404
rect 6420 24392 6426 24404
rect 6917 24395 6975 24401
rect 6917 24392 6929 24395
rect 6420 24364 6929 24392
rect 6420 24352 6426 24364
rect 6917 24361 6929 24364
rect 6963 24392 6975 24395
rect 7190 24392 7196 24404
rect 6963 24364 7196 24392
rect 6963 24361 6975 24364
rect 6917 24355 6975 24361
rect 7190 24352 7196 24364
rect 7248 24352 7254 24404
rect 7558 24392 7564 24404
rect 7519 24364 7564 24392
rect 7558 24352 7564 24364
rect 7616 24352 7622 24404
rect 8294 24392 8300 24404
rect 8255 24364 8300 24392
rect 8294 24352 8300 24364
rect 8352 24352 8358 24404
rect 13078 24392 13084 24404
rect 13039 24364 13084 24392
rect 13078 24352 13084 24364
rect 13136 24352 13142 24404
rect 17037 24395 17095 24401
rect 17037 24361 17049 24395
rect 17083 24392 17095 24395
rect 17310 24392 17316 24404
rect 17083 24364 17316 24392
rect 17083 24361 17095 24364
rect 17037 24355 17095 24361
rect 17310 24352 17316 24364
rect 17368 24352 17374 24404
rect 18141 24395 18199 24401
rect 18141 24361 18153 24395
rect 18187 24392 18199 24395
rect 19242 24392 19248 24404
rect 18187 24364 19248 24392
rect 18187 24361 18199 24364
rect 18141 24355 18199 24361
rect 19242 24352 19248 24364
rect 19300 24352 19306 24404
rect 21542 24392 21548 24404
rect 21503 24364 21548 24392
rect 21542 24352 21548 24364
rect 21600 24352 21606 24404
rect 22738 24392 22744 24404
rect 22699 24364 22744 24392
rect 22738 24352 22744 24364
rect 22796 24352 22802 24404
rect 23845 24395 23903 24401
rect 23845 24361 23857 24395
rect 23891 24392 23903 24395
rect 24118 24392 24124 24404
rect 23891 24364 24124 24392
rect 23891 24361 23903 24364
rect 23845 24355 23903 24361
rect 24118 24352 24124 24364
rect 24176 24352 24182 24404
rect 24949 24395 25007 24401
rect 24949 24361 24961 24395
rect 24995 24392 25007 24395
rect 26878 24392 26884 24404
rect 24995 24364 26884 24392
rect 24995 24361 25007 24364
rect 24949 24355 25007 24361
rect 26878 24352 26884 24364
rect 26936 24352 26942 24404
rect 9858 24284 9864 24336
rect 9916 24324 9922 24336
rect 10750 24327 10808 24333
rect 10750 24324 10762 24327
rect 9916 24296 10762 24324
rect 9916 24284 9922 24296
rect 10750 24293 10762 24296
rect 10796 24324 10808 24327
rect 10870 24324 10876 24336
rect 10796 24296 10876 24324
rect 10796 24293 10808 24296
rect 10750 24287 10808 24293
rect 10870 24284 10876 24296
rect 10928 24284 10934 24336
rect 13909 24327 13967 24333
rect 13909 24293 13921 24327
rect 13955 24324 13967 24327
rect 13998 24324 14004 24336
rect 13955 24296 14004 24324
rect 13955 24293 13967 24296
rect 13909 24287 13967 24293
rect 13998 24284 14004 24296
rect 14056 24284 14062 24336
rect 15838 24324 15844 24336
rect 15799 24296 15844 24324
rect 15838 24284 15844 24296
rect 15896 24284 15902 24336
rect 19610 24324 19616 24336
rect 19571 24296 19616 24324
rect 19610 24284 19616 24296
rect 19668 24324 19674 24336
rect 20073 24327 20131 24333
rect 20073 24324 20085 24327
rect 19668 24296 20085 24324
rect 19668 24284 19674 24296
rect 20073 24293 20085 24296
rect 20119 24293 20131 24327
rect 20073 24287 20131 24293
rect 7285 24259 7343 24265
rect 7285 24225 7297 24259
rect 7331 24256 7343 24259
rect 8018 24256 8024 24268
rect 7331 24228 8024 24256
rect 7331 24225 7343 24228
rect 7285 24219 7343 24225
rect 8018 24216 8024 24228
rect 8076 24256 8082 24268
rect 8389 24259 8447 24265
rect 8389 24256 8401 24259
rect 8076 24228 8401 24256
rect 8076 24216 8082 24228
rect 8389 24225 8401 24228
rect 8435 24225 8447 24259
rect 8389 24219 8447 24225
rect 12250 24216 12256 24268
rect 12308 24256 12314 24268
rect 13538 24256 13544 24268
rect 12308 24228 13544 24256
rect 12308 24216 12314 24228
rect 13538 24216 13544 24228
rect 13596 24256 13602 24268
rect 13725 24259 13783 24265
rect 13725 24256 13737 24259
rect 13596 24228 13737 24256
rect 13596 24216 13602 24228
rect 13725 24225 13737 24228
rect 13771 24225 13783 24259
rect 16850 24256 16856 24268
rect 16811 24228 16856 24256
rect 13725 24219 13783 24225
rect 16850 24216 16856 24228
rect 16908 24216 16914 24268
rect 17586 24216 17592 24268
rect 17644 24256 17650 24268
rect 17957 24259 18015 24265
rect 17957 24256 17969 24259
rect 17644 24228 17969 24256
rect 17644 24216 17650 24228
rect 17957 24225 17969 24228
rect 18003 24225 18015 24259
rect 17957 24219 18015 24225
rect 19426 24216 19432 24268
rect 19484 24256 19490 24268
rect 19705 24259 19763 24265
rect 19705 24256 19717 24259
rect 19484 24228 19717 24256
rect 19484 24216 19490 24228
rect 19705 24225 19717 24228
rect 19751 24225 19763 24259
rect 22554 24256 22560 24268
rect 22515 24228 22560 24256
rect 19705 24219 19763 24225
rect 22554 24216 22560 24228
rect 22612 24216 22618 24268
rect 23661 24259 23719 24265
rect 23661 24225 23673 24259
rect 23707 24256 23719 24259
rect 24210 24256 24216 24268
rect 23707 24228 24216 24256
rect 23707 24225 23719 24228
rect 23661 24219 23719 24225
rect 24210 24216 24216 24228
rect 24268 24216 24274 24268
rect 24765 24259 24823 24265
rect 24765 24225 24777 24259
rect 24811 24256 24823 24259
rect 24854 24256 24860 24268
rect 24811 24228 24860 24256
rect 24811 24225 24823 24228
rect 24765 24219 24823 24225
rect 24854 24216 24860 24228
rect 24912 24216 24918 24268
rect 8110 24148 8116 24200
rect 8168 24188 8174 24200
rect 8205 24191 8263 24197
rect 8205 24188 8217 24191
rect 8168 24160 8217 24188
rect 8168 24148 8174 24160
rect 8205 24157 8217 24160
rect 8251 24157 8263 24191
rect 8205 24151 8263 24157
rect 9674 24148 9680 24200
rect 9732 24188 9738 24200
rect 10502 24188 10508 24200
rect 9732 24160 10508 24188
rect 9732 24148 9738 24160
rect 10502 24148 10508 24160
rect 10560 24148 10566 24200
rect 14001 24191 14059 24197
rect 14001 24157 14013 24191
rect 14047 24188 14059 24191
rect 14458 24188 14464 24200
rect 14047 24160 14464 24188
rect 14047 24157 14059 24160
rect 14001 24151 14059 24157
rect 14458 24148 14464 24160
rect 14516 24148 14522 24200
rect 15105 24191 15163 24197
rect 15105 24157 15117 24191
rect 15151 24188 15163 24191
rect 15746 24188 15752 24200
rect 15151 24160 15752 24188
rect 15151 24157 15163 24160
rect 15105 24151 15163 24157
rect 15746 24148 15752 24160
rect 15804 24148 15810 24200
rect 15930 24188 15936 24200
rect 15891 24160 15936 24188
rect 15930 24148 15936 24160
rect 15988 24148 15994 24200
rect 19518 24188 19524 24200
rect 19479 24160 19524 24188
rect 19518 24148 19524 24160
rect 19576 24148 19582 24200
rect 21450 24188 21456 24200
rect 21411 24160 21456 24188
rect 21450 24148 21456 24160
rect 21508 24148 21514 24200
rect 21634 24188 21640 24200
rect 21595 24160 21640 24188
rect 21634 24148 21640 24160
rect 21692 24148 21698 24200
rect 18601 24123 18659 24129
rect 18601 24089 18613 24123
rect 18647 24120 18659 24123
rect 19058 24120 19064 24132
rect 18647 24092 19064 24120
rect 18647 24089 18659 24092
rect 18601 24083 18659 24089
rect 19058 24080 19064 24092
rect 19116 24080 19122 24132
rect 21082 24120 21088 24132
rect 21043 24092 21088 24120
rect 21082 24080 21088 24092
rect 21140 24080 21146 24132
rect 7834 24052 7840 24064
rect 7795 24024 7840 24052
rect 7834 24012 7840 24024
rect 7892 24012 7898 24064
rect 10410 24052 10416 24064
rect 10371 24024 10416 24052
rect 10410 24012 10416 24024
rect 10468 24052 10474 24064
rect 10778 24052 10784 24064
rect 10468 24024 10784 24052
rect 10468 24012 10474 24024
rect 10778 24012 10784 24024
rect 10836 24012 10842 24064
rect 11885 24055 11943 24061
rect 11885 24021 11897 24055
rect 11931 24052 11943 24055
rect 11974 24052 11980 24064
rect 11931 24024 11980 24052
rect 11931 24021 11943 24024
rect 11885 24015 11943 24021
rect 11974 24012 11980 24024
rect 12032 24012 12038 24064
rect 12434 24012 12440 24064
rect 12492 24052 12498 24064
rect 13449 24055 13507 24061
rect 12492 24024 12537 24052
rect 12492 24012 12498 24024
rect 13449 24021 13461 24055
rect 13495 24052 13507 24055
rect 13814 24052 13820 24064
rect 13495 24024 13820 24052
rect 13495 24021 13507 24024
rect 13449 24015 13507 24021
rect 13814 24012 13820 24024
rect 13872 24012 13878 24064
rect 15378 24052 15384 24064
rect 15339 24024 15384 24052
rect 15378 24012 15384 24024
rect 15436 24012 15442 24064
rect 16390 24052 16396 24064
rect 16351 24024 16396 24052
rect 16390 24012 16396 24024
rect 16448 24012 16454 24064
rect 18874 24052 18880 24064
rect 18835 24024 18880 24052
rect 18874 24012 18880 24024
rect 18932 24012 18938 24064
rect 19150 24052 19156 24064
rect 19111 24024 19156 24052
rect 19150 24012 19156 24024
rect 19208 24012 19214 24064
rect 19334 24012 19340 24064
rect 19392 24052 19398 24064
rect 19978 24052 19984 24064
rect 19392 24024 19984 24052
rect 19392 24012 19398 24024
rect 19978 24012 19984 24024
rect 20036 24012 20042 24064
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 9858 23848 9864 23860
rect 9819 23820 9864 23848
rect 9858 23808 9864 23820
rect 9916 23808 9922 23860
rect 10502 23808 10508 23860
rect 10560 23848 10566 23860
rect 11333 23851 11391 23857
rect 11333 23848 11345 23851
rect 10560 23820 11345 23848
rect 10560 23808 10566 23820
rect 11333 23817 11345 23820
rect 11379 23817 11391 23851
rect 12250 23848 12256 23860
rect 12211 23820 12256 23848
rect 11333 23811 11391 23817
rect 10042 23740 10048 23792
rect 10100 23780 10106 23792
rect 10413 23783 10471 23789
rect 10413 23780 10425 23783
rect 10100 23752 10425 23780
rect 10100 23740 10106 23752
rect 10413 23749 10425 23752
rect 10459 23749 10471 23783
rect 10413 23743 10471 23749
rect 9858 23672 9864 23724
rect 9916 23712 9922 23724
rect 10134 23712 10140 23724
rect 9916 23684 10140 23712
rect 9916 23672 9922 23684
rect 10134 23672 10140 23684
rect 10192 23672 10198 23724
rect 10962 23712 10968 23724
rect 10244 23684 10968 23712
rect 7285 23647 7343 23653
rect 7285 23613 7297 23647
rect 7331 23644 7343 23647
rect 7561 23647 7619 23653
rect 7561 23644 7573 23647
rect 7331 23616 7573 23644
rect 7331 23613 7343 23616
rect 7285 23607 7343 23613
rect 7561 23613 7573 23616
rect 7607 23613 7619 23647
rect 7561 23607 7619 23613
rect 7650 23604 7656 23656
rect 7708 23644 7714 23656
rect 7817 23647 7875 23653
rect 7817 23644 7829 23647
rect 7708 23616 7829 23644
rect 7708 23604 7714 23616
rect 7817 23613 7829 23616
rect 7863 23644 7875 23647
rect 8294 23644 8300 23656
rect 7863 23616 8300 23644
rect 7863 23613 7875 23616
rect 7817 23607 7875 23613
rect 8294 23604 8300 23616
rect 8352 23604 8358 23656
rect 10244 23644 10272 23684
rect 10962 23672 10968 23684
rect 11020 23672 11026 23724
rect 11348 23712 11376 23811
rect 12250 23808 12256 23820
rect 12308 23808 12314 23860
rect 12618 23848 12624 23860
rect 12579 23820 12624 23848
rect 12618 23808 12624 23820
rect 12676 23808 12682 23860
rect 14458 23808 14464 23860
rect 14516 23848 14522 23860
rect 14921 23851 14979 23857
rect 14921 23848 14933 23851
rect 14516 23820 14933 23848
rect 14516 23808 14522 23820
rect 14921 23817 14933 23820
rect 14967 23848 14979 23851
rect 15565 23851 15623 23857
rect 15565 23848 15577 23851
rect 14967 23820 15577 23848
rect 14967 23817 14979 23820
rect 14921 23811 14979 23817
rect 15565 23817 15577 23820
rect 15611 23848 15623 23851
rect 15930 23848 15936 23860
rect 15611 23820 15936 23848
rect 15611 23817 15623 23820
rect 15565 23811 15623 23817
rect 15930 23808 15936 23820
rect 15988 23808 15994 23860
rect 16482 23848 16488 23860
rect 16443 23820 16488 23848
rect 16482 23808 16488 23820
rect 16540 23808 16546 23860
rect 21542 23808 21548 23860
rect 21600 23848 21606 23860
rect 21821 23851 21879 23857
rect 21821 23848 21833 23851
rect 21600 23820 21833 23848
rect 21600 23808 21606 23820
rect 21821 23817 21833 23820
rect 21867 23817 21879 23851
rect 21821 23811 21879 23817
rect 22094 23808 22100 23860
rect 22152 23848 22158 23860
rect 22557 23851 22615 23857
rect 22557 23848 22569 23851
rect 22152 23820 22569 23848
rect 22152 23808 22158 23820
rect 22557 23817 22569 23820
rect 22603 23817 22615 23851
rect 22557 23811 22615 23817
rect 23845 23851 23903 23857
rect 23845 23817 23857 23851
rect 23891 23848 23903 23851
rect 24670 23848 24676 23860
rect 23891 23820 24676 23848
rect 23891 23817 23903 23820
rect 23845 23811 23903 23817
rect 24670 23808 24676 23820
rect 24728 23808 24734 23860
rect 24946 23848 24952 23860
rect 24907 23820 24952 23848
rect 24946 23808 24952 23820
rect 25004 23808 25010 23860
rect 18322 23780 18328 23792
rect 18283 23752 18328 23780
rect 18322 23740 18328 23752
rect 18380 23740 18386 23792
rect 21450 23740 21456 23792
rect 21508 23780 21514 23792
rect 22281 23783 22339 23789
rect 22281 23780 22293 23783
rect 21508 23752 22293 23780
rect 21508 23740 21514 23752
rect 22281 23749 22293 23752
rect 22327 23780 22339 23783
rect 23290 23780 23296 23792
rect 22327 23752 23296 23780
rect 22327 23749 22339 23752
rect 22281 23743 22339 23749
rect 23290 23740 23296 23752
rect 23348 23740 23354 23792
rect 13357 23715 13415 23721
rect 13357 23712 13369 23715
rect 11348 23684 13369 23712
rect 13357 23681 13369 23684
rect 13403 23712 13415 23715
rect 13541 23715 13599 23721
rect 13541 23712 13553 23715
rect 13403 23684 13553 23712
rect 13403 23681 13415 23684
rect 13357 23675 13415 23681
rect 13541 23681 13553 23684
rect 13587 23681 13599 23715
rect 13541 23675 13599 23681
rect 16390 23672 16396 23724
rect 16448 23712 16454 23724
rect 16853 23715 16911 23721
rect 16853 23712 16865 23715
rect 16448 23684 16865 23712
rect 16448 23672 16454 23684
rect 16853 23681 16865 23684
rect 16899 23681 16911 23715
rect 16853 23675 16911 23681
rect 17497 23715 17555 23721
rect 17497 23681 17509 23715
rect 17543 23712 17555 23715
rect 18785 23715 18843 23721
rect 18785 23712 18797 23715
rect 17543 23684 18797 23712
rect 17543 23681 17555 23684
rect 17497 23675 17555 23681
rect 18785 23681 18797 23684
rect 18831 23712 18843 23715
rect 18966 23712 18972 23724
rect 18831 23684 18972 23712
rect 18831 23681 18843 23684
rect 18785 23675 18843 23681
rect 18966 23672 18972 23684
rect 19024 23672 19030 23724
rect 10152 23616 10272 23644
rect 10689 23647 10747 23653
rect 7101 23579 7159 23585
rect 7101 23545 7113 23579
rect 7147 23576 7159 23579
rect 8110 23576 8116 23588
rect 7147 23548 8116 23576
rect 7147 23545 7159 23548
rect 7101 23539 7159 23545
rect 8110 23536 8116 23548
rect 8168 23536 8174 23588
rect 10152 23520 10180 23616
rect 10689 23613 10701 23647
rect 10735 23644 10747 23647
rect 10735 23616 11836 23644
rect 10735 23613 10747 23616
rect 10689 23607 10747 23613
rect 10410 23536 10416 23588
rect 10468 23576 10474 23588
rect 10873 23579 10931 23585
rect 10873 23576 10885 23579
rect 10468 23548 10885 23576
rect 10468 23536 10474 23548
rect 10873 23545 10885 23548
rect 10919 23545 10931 23579
rect 10873 23539 10931 23545
rect 7006 23468 7012 23520
rect 7064 23508 7070 23520
rect 7285 23511 7343 23517
rect 7285 23508 7297 23511
rect 7064 23480 7297 23508
rect 7064 23468 7070 23480
rect 7285 23477 7297 23480
rect 7331 23508 7343 23511
rect 7377 23511 7435 23517
rect 7377 23508 7389 23511
rect 7331 23480 7389 23508
rect 7331 23477 7343 23480
rect 7285 23471 7343 23477
rect 7377 23477 7389 23480
rect 7423 23477 7435 23511
rect 7377 23471 7435 23477
rect 8018 23468 8024 23520
rect 8076 23508 8082 23520
rect 8941 23511 8999 23517
rect 8941 23508 8953 23511
rect 8076 23480 8953 23508
rect 8076 23468 8082 23480
rect 8941 23477 8953 23480
rect 8987 23508 8999 23511
rect 9582 23508 9588 23520
rect 8987 23480 9588 23508
rect 8987 23477 8999 23480
rect 8941 23471 8999 23477
rect 9582 23468 9588 23480
rect 9640 23468 9646 23520
rect 10134 23508 10140 23520
rect 10095 23480 10140 23508
rect 10134 23468 10140 23480
rect 10192 23468 10198 23520
rect 11808 23517 11836 23616
rect 12434 23604 12440 23656
rect 12492 23644 12498 23656
rect 13630 23644 13636 23656
rect 12492 23616 13636 23644
rect 12492 23604 12498 23616
rect 13630 23604 13636 23616
rect 13688 23604 13694 23656
rect 15933 23647 15991 23653
rect 15933 23613 15945 23647
rect 15979 23644 15991 23647
rect 17037 23647 17095 23653
rect 17037 23644 17049 23647
rect 15979 23616 17049 23644
rect 15979 23613 15991 23616
rect 15933 23607 15991 23613
rect 17037 23613 17049 23616
rect 17083 23644 17095 23647
rect 17862 23644 17868 23656
rect 17083 23616 17868 23644
rect 17083 23613 17095 23616
rect 17037 23607 17095 23613
rect 17862 23604 17868 23616
rect 17920 23604 17926 23656
rect 19797 23647 19855 23653
rect 19797 23613 19809 23647
rect 19843 23644 19855 23647
rect 19889 23647 19947 23653
rect 19889 23644 19901 23647
rect 19843 23616 19901 23644
rect 19843 23613 19855 23616
rect 19797 23607 19855 23613
rect 19889 23613 19901 23616
rect 19935 23644 19947 23647
rect 20990 23644 20996 23656
rect 19935 23616 20996 23644
rect 19935 23613 19947 23616
rect 19889 23607 19947 23613
rect 20990 23604 20996 23616
rect 21048 23604 21054 23656
rect 22373 23647 22431 23653
rect 22373 23613 22385 23647
rect 22419 23644 22431 23647
rect 23661 23647 23719 23653
rect 23661 23644 23673 23647
rect 22419 23616 23060 23644
rect 22419 23613 22431 23616
rect 22373 23607 22431 23613
rect 13081 23579 13139 23585
rect 13081 23545 13093 23579
rect 13127 23576 13139 23579
rect 13808 23579 13866 23585
rect 13808 23576 13820 23579
rect 13127 23548 13820 23576
rect 13127 23545 13139 23548
rect 13081 23539 13139 23545
rect 13808 23545 13820 23548
rect 13854 23576 13866 23579
rect 14090 23576 14096 23588
rect 13854 23548 14096 23576
rect 13854 23545 13866 23548
rect 13808 23539 13866 23545
rect 14090 23536 14096 23548
rect 14148 23536 14154 23588
rect 16114 23536 16120 23588
rect 16172 23576 16178 23588
rect 16209 23579 16267 23585
rect 16209 23576 16221 23579
rect 16172 23548 16221 23576
rect 16172 23536 16178 23548
rect 16209 23545 16221 23548
rect 16255 23545 16267 23579
rect 18874 23576 18880 23588
rect 18835 23548 18880 23576
rect 16209 23539 16267 23545
rect 11793 23511 11851 23517
rect 11793 23477 11805 23511
rect 11839 23508 11851 23511
rect 12342 23508 12348 23520
rect 11839 23480 12348 23508
rect 11839 23477 11851 23480
rect 11793 23471 11851 23477
rect 12342 23468 12348 23480
rect 12400 23468 12406 23520
rect 15102 23468 15108 23520
rect 15160 23508 15166 23520
rect 15838 23508 15844 23520
rect 15160 23480 15844 23508
rect 15160 23468 15166 23480
rect 15838 23468 15844 23480
rect 15896 23468 15902 23520
rect 16224 23508 16252 23539
rect 18874 23536 18880 23548
rect 18932 23536 18938 23588
rect 20134 23579 20192 23585
rect 20134 23576 20146 23579
rect 19444 23548 20146 23576
rect 19444 23520 19472 23548
rect 20134 23545 20146 23548
rect 20180 23545 20192 23579
rect 20134 23539 20192 23545
rect 16945 23511 17003 23517
rect 16945 23508 16957 23511
rect 16224 23480 16957 23508
rect 16945 23477 16957 23480
rect 16991 23477 17003 23511
rect 16945 23471 17003 23477
rect 17586 23468 17592 23520
rect 17644 23508 17650 23520
rect 17773 23511 17831 23517
rect 17773 23508 17785 23511
rect 17644 23480 17785 23508
rect 17644 23468 17650 23480
rect 17773 23477 17785 23480
rect 17819 23477 17831 23511
rect 17773 23471 17831 23477
rect 18785 23511 18843 23517
rect 18785 23477 18797 23511
rect 18831 23508 18843 23511
rect 19058 23508 19064 23520
rect 18831 23480 19064 23508
rect 18831 23477 18843 23480
rect 18785 23471 18843 23477
rect 19058 23468 19064 23480
rect 19116 23468 19122 23520
rect 19337 23511 19395 23517
rect 19337 23477 19349 23511
rect 19383 23508 19395 23511
rect 19426 23508 19432 23520
rect 19383 23480 19432 23508
rect 19383 23477 19395 23480
rect 19337 23471 19395 23477
rect 19426 23468 19432 23480
rect 19484 23468 19490 23520
rect 21266 23508 21272 23520
rect 21227 23480 21272 23508
rect 21266 23468 21272 23480
rect 21324 23468 21330 23520
rect 23032 23517 23060 23616
rect 23492 23616 23673 23644
rect 23492 23520 23520 23616
rect 23661 23613 23673 23616
rect 23707 23613 23719 23647
rect 24210 23644 24216 23656
rect 24171 23616 24216 23644
rect 23661 23607 23719 23613
rect 24210 23604 24216 23616
rect 24268 23604 24274 23656
rect 24765 23647 24823 23653
rect 24765 23613 24777 23647
rect 24811 23613 24823 23647
rect 24765 23607 24823 23613
rect 23934 23536 23940 23588
rect 23992 23576 23998 23588
rect 24581 23579 24639 23585
rect 24581 23576 24593 23579
rect 23992 23548 24593 23576
rect 23992 23536 23998 23548
rect 24581 23545 24593 23548
rect 24627 23576 24639 23579
rect 24780 23576 24808 23607
rect 24627 23548 24808 23576
rect 24627 23545 24639 23548
rect 24581 23539 24639 23545
rect 23017 23511 23075 23517
rect 23017 23477 23029 23511
rect 23063 23508 23075 23511
rect 23106 23508 23112 23520
rect 23063 23480 23112 23508
rect 23063 23477 23075 23480
rect 23017 23471 23075 23477
rect 23106 23468 23112 23480
rect 23164 23468 23170 23520
rect 23474 23508 23480 23520
rect 23435 23480 23480 23508
rect 23474 23468 23480 23480
rect 23532 23468 23538 23520
rect 23842 23468 23848 23520
rect 23900 23508 23906 23520
rect 24854 23508 24860 23520
rect 23900 23480 24860 23508
rect 23900 23468 23906 23480
rect 24854 23468 24860 23480
rect 24912 23508 24918 23520
rect 25317 23511 25375 23517
rect 25317 23508 25329 23511
rect 24912 23480 25329 23508
rect 24912 23468 24918 23480
rect 25317 23477 25329 23480
rect 25363 23477 25375 23511
rect 25317 23471 25375 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 8294 23264 8300 23316
rect 8352 23304 8358 23316
rect 8389 23307 8447 23313
rect 8389 23304 8401 23307
rect 8352 23276 8401 23304
rect 8352 23264 8358 23276
rect 8389 23273 8401 23276
rect 8435 23273 8447 23307
rect 8389 23267 8447 23273
rect 11054 23264 11060 23316
rect 11112 23304 11118 23316
rect 11517 23307 11575 23313
rect 11517 23304 11529 23307
rect 11112 23276 11529 23304
rect 11112 23264 11118 23276
rect 11517 23273 11529 23276
rect 11563 23273 11575 23307
rect 11517 23267 11575 23273
rect 12618 23264 12624 23316
rect 12676 23304 12682 23316
rect 13173 23307 13231 23313
rect 13173 23304 13185 23307
rect 12676 23276 13185 23304
rect 12676 23264 12682 23276
rect 13173 23273 13185 23276
rect 13219 23304 13231 23307
rect 13262 23304 13268 23316
rect 13219 23276 13268 23304
rect 13219 23273 13231 23276
rect 13173 23267 13231 23273
rect 13262 23264 13268 23276
rect 13320 23264 13326 23316
rect 13998 23304 14004 23316
rect 13959 23276 14004 23304
rect 13998 23264 14004 23276
rect 14056 23264 14062 23316
rect 15102 23304 15108 23316
rect 15063 23276 15108 23304
rect 15102 23264 15108 23276
rect 15160 23264 15166 23316
rect 19518 23264 19524 23316
rect 19576 23304 19582 23316
rect 20257 23307 20315 23313
rect 20257 23304 20269 23307
rect 19576 23276 20269 23304
rect 19576 23264 19582 23276
rect 20257 23273 20269 23276
rect 20303 23273 20315 23307
rect 20257 23267 20315 23273
rect 22554 23264 22560 23316
rect 22612 23304 22618 23316
rect 22830 23304 22836 23316
rect 22612 23276 22836 23304
rect 22612 23264 22618 23276
rect 22830 23264 22836 23276
rect 22888 23304 22894 23316
rect 22925 23307 22983 23313
rect 22925 23304 22937 23307
rect 22888 23276 22937 23304
rect 22888 23264 22894 23276
rect 22925 23273 22937 23276
rect 22971 23273 22983 23307
rect 24762 23304 24768 23316
rect 24723 23276 24768 23304
rect 22925 23267 22983 23273
rect 24762 23264 24768 23276
rect 24820 23264 24826 23316
rect 10404 23239 10462 23245
rect 10404 23205 10416 23239
rect 10450 23236 10462 23239
rect 11974 23236 11980 23248
rect 10450 23208 11980 23236
rect 10450 23205 10462 23208
rect 10404 23199 10462 23205
rect 11974 23196 11980 23208
rect 12032 23196 12038 23248
rect 13725 23239 13783 23245
rect 13725 23205 13737 23239
rect 13771 23236 13783 23239
rect 14458 23236 14464 23248
rect 13771 23208 14464 23236
rect 13771 23205 13783 23208
rect 13725 23199 13783 23205
rect 14458 23196 14464 23208
rect 14516 23196 14522 23248
rect 15556 23239 15614 23245
rect 15556 23205 15568 23239
rect 15602 23236 15614 23239
rect 15930 23236 15936 23248
rect 15602 23208 15936 23236
rect 15602 23205 15614 23208
rect 15556 23199 15614 23205
rect 15930 23196 15936 23208
rect 15988 23196 15994 23248
rect 21266 23245 21272 23248
rect 21260 23236 21272 23245
rect 21227 23208 21272 23236
rect 21260 23199 21272 23208
rect 21266 23196 21272 23199
rect 21324 23196 21330 23248
rect 6638 23128 6644 23180
rect 6696 23168 6702 23180
rect 7265 23171 7323 23177
rect 7265 23168 7277 23171
rect 6696 23140 7277 23168
rect 6696 23128 6702 23140
rect 7265 23137 7277 23140
rect 7311 23168 7323 23171
rect 8202 23168 8208 23180
rect 7311 23140 8208 23168
rect 7311 23137 7323 23140
rect 7265 23131 7323 23137
rect 8202 23128 8208 23140
rect 8260 23128 8266 23180
rect 12066 23128 12072 23180
rect 12124 23168 12130 23180
rect 12989 23171 13047 23177
rect 12989 23168 13001 23171
rect 12124 23140 13001 23168
rect 12124 23128 12130 23140
rect 12989 23137 13001 23140
rect 13035 23137 13047 23171
rect 18029 23171 18087 23177
rect 18029 23168 18041 23171
rect 12989 23131 13047 23137
rect 17604 23140 18041 23168
rect 7006 23100 7012 23112
rect 6967 23072 7012 23100
rect 7006 23060 7012 23072
rect 7064 23060 7070 23112
rect 9674 23060 9680 23112
rect 9732 23100 9738 23112
rect 10137 23103 10195 23109
rect 10137 23100 10149 23103
rect 9732 23072 10149 23100
rect 9732 23060 9738 23072
rect 10137 23069 10149 23072
rect 10183 23069 10195 23103
rect 10137 23063 10195 23069
rect 12434 23060 12440 23112
rect 12492 23100 12498 23112
rect 13262 23100 13268 23112
rect 12492 23072 12756 23100
rect 13223 23072 13268 23100
rect 12492 23060 12498 23072
rect 12728 23041 12756 23072
rect 13262 23060 13268 23072
rect 13320 23060 13326 23112
rect 14182 23100 14188 23112
rect 14143 23072 14188 23100
rect 14182 23060 14188 23072
rect 14240 23060 14246 23112
rect 15286 23100 15292 23112
rect 15247 23072 15292 23100
rect 15286 23060 15292 23072
rect 15344 23060 15350 23112
rect 17604 23041 17632 23140
rect 18029 23137 18041 23140
rect 18075 23137 18087 23171
rect 20990 23168 20996 23180
rect 20951 23140 20996 23168
rect 18029 23131 18087 23137
rect 20990 23128 20996 23140
rect 21048 23128 21054 23180
rect 24581 23171 24639 23177
rect 24581 23137 24593 23171
rect 24627 23168 24639 23171
rect 24854 23168 24860 23180
rect 24627 23140 24860 23168
rect 24627 23137 24639 23140
rect 24581 23131 24639 23137
rect 24854 23128 24860 23140
rect 24912 23128 24918 23180
rect 17678 23060 17684 23112
rect 17736 23100 17742 23112
rect 17773 23103 17831 23109
rect 17773 23100 17785 23103
rect 17736 23072 17785 23100
rect 17736 23060 17742 23072
rect 17773 23069 17785 23072
rect 17819 23069 17831 23103
rect 17773 23063 17831 23069
rect 12713 23035 12771 23041
rect 12713 23001 12725 23035
rect 12759 23001 12771 23035
rect 17589 23035 17647 23041
rect 17589 23032 17601 23035
rect 12713 22995 12771 23001
rect 16684 23004 17601 23032
rect 16684 22976 16712 23004
rect 17589 23001 17601 23004
rect 17635 23001 17647 23035
rect 17589 22995 17647 23001
rect 9582 22924 9588 22976
rect 9640 22964 9646 22976
rect 10045 22967 10103 22973
rect 10045 22964 10057 22967
rect 9640 22936 10057 22964
rect 9640 22924 9646 22936
rect 10045 22933 10057 22936
rect 10091 22964 10103 22967
rect 10870 22964 10876 22976
rect 10091 22936 10876 22964
rect 10091 22933 10103 22936
rect 10045 22927 10103 22933
rect 10870 22924 10876 22936
rect 10928 22924 10934 22976
rect 12066 22964 12072 22976
rect 12027 22936 12072 22964
rect 12066 22924 12072 22936
rect 12124 22924 12130 22976
rect 12529 22967 12587 22973
rect 12529 22933 12541 22967
rect 12575 22964 12587 22967
rect 12802 22964 12808 22976
rect 12575 22936 12808 22964
rect 12575 22933 12587 22936
rect 12529 22927 12587 22933
rect 12802 22924 12808 22936
rect 12860 22924 12866 22976
rect 16666 22964 16672 22976
rect 16627 22936 16672 22964
rect 16666 22924 16672 22936
rect 16724 22924 16730 22976
rect 16850 22924 16856 22976
rect 16908 22964 16914 22976
rect 17221 22967 17279 22973
rect 17221 22964 17233 22967
rect 16908 22936 17233 22964
rect 16908 22924 16914 22936
rect 17221 22933 17233 22936
rect 17267 22933 17279 22967
rect 17221 22927 17279 22933
rect 18874 22924 18880 22976
rect 18932 22964 18938 22976
rect 19153 22967 19211 22973
rect 19153 22964 19165 22967
rect 18932 22936 19165 22964
rect 18932 22924 18938 22936
rect 19153 22933 19165 22936
rect 19199 22933 19211 22967
rect 19153 22927 19211 22933
rect 19426 22924 19432 22976
rect 19484 22964 19490 22976
rect 19889 22967 19947 22973
rect 19889 22964 19901 22967
rect 19484 22936 19901 22964
rect 19484 22924 19490 22936
rect 19889 22933 19901 22936
rect 19935 22933 19947 22967
rect 20714 22964 20720 22976
rect 20675 22936 20720 22964
rect 19889 22927 19947 22933
rect 20714 22924 20720 22936
rect 20772 22964 20778 22976
rect 21634 22964 21640 22976
rect 20772 22936 21640 22964
rect 20772 22924 20778 22936
rect 21634 22924 21640 22936
rect 21692 22964 21698 22976
rect 22373 22967 22431 22973
rect 22373 22964 22385 22967
rect 21692 22936 22385 22964
rect 21692 22924 21698 22936
rect 22373 22933 22385 22936
rect 22419 22933 22431 22967
rect 22373 22927 22431 22933
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 6638 22760 6644 22772
rect 6599 22732 6644 22760
rect 6638 22720 6644 22732
rect 6696 22720 6702 22772
rect 11333 22763 11391 22769
rect 11333 22729 11345 22763
rect 11379 22760 11391 22763
rect 11974 22760 11980 22772
rect 11379 22732 11980 22760
rect 11379 22729 11391 22732
rect 11333 22723 11391 22729
rect 11974 22720 11980 22732
rect 12032 22760 12038 22772
rect 13262 22760 13268 22772
rect 12032 22732 13268 22760
rect 12032 22720 12038 22732
rect 13262 22720 13268 22732
rect 13320 22760 13326 22772
rect 13449 22763 13507 22769
rect 13449 22760 13461 22763
rect 13320 22732 13461 22760
rect 13320 22720 13326 22732
rect 13449 22729 13461 22732
rect 13495 22729 13507 22763
rect 14458 22760 14464 22772
rect 14419 22732 14464 22760
rect 13449 22723 13507 22729
rect 14458 22720 14464 22732
rect 14516 22720 14522 22772
rect 16942 22760 16948 22772
rect 16903 22732 16948 22760
rect 16942 22720 16948 22732
rect 17000 22720 17006 22772
rect 20901 22763 20959 22769
rect 20901 22729 20913 22763
rect 20947 22760 20959 22763
rect 20990 22760 20996 22772
rect 20947 22732 20996 22760
rect 20947 22729 20959 22732
rect 20901 22723 20959 22729
rect 20990 22720 20996 22732
rect 21048 22720 21054 22772
rect 24670 22720 24676 22772
rect 24728 22760 24734 22772
rect 24765 22763 24823 22769
rect 24765 22760 24777 22763
rect 24728 22732 24777 22760
rect 24728 22720 24734 22732
rect 24765 22729 24777 22732
rect 24811 22729 24823 22763
rect 24765 22723 24823 22729
rect 10318 22692 10324 22704
rect 10279 22664 10324 22692
rect 10318 22652 10324 22664
rect 10376 22652 10382 22704
rect 11054 22652 11060 22704
rect 11112 22692 11118 22704
rect 11790 22692 11796 22704
rect 11112 22664 11796 22692
rect 11112 22652 11118 22664
rect 11790 22652 11796 22664
rect 11848 22652 11854 22704
rect 12526 22692 12532 22704
rect 12487 22664 12532 22692
rect 12526 22652 12532 22664
rect 12584 22652 12590 22704
rect 14550 22652 14556 22704
rect 14608 22692 14614 22704
rect 15105 22695 15163 22701
rect 15105 22692 15117 22695
rect 14608 22664 15117 22692
rect 14608 22652 14614 22664
rect 15105 22661 15117 22664
rect 15151 22661 15163 22695
rect 15105 22655 15163 22661
rect 21085 22695 21143 22701
rect 21085 22661 21097 22695
rect 21131 22692 21143 22695
rect 21634 22692 21640 22704
rect 21131 22664 21640 22692
rect 21131 22661 21143 22664
rect 21085 22655 21143 22661
rect 21634 22652 21640 22664
rect 21692 22652 21698 22704
rect 10870 22624 10876 22636
rect 10831 22596 10876 22624
rect 10870 22584 10876 22596
rect 10928 22584 10934 22636
rect 11808 22624 11836 22652
rect 13078 22624 13084 22636
rect 11808 22596 13084 22624
rect 13078 22584 13084 22596
rect 13136 22584 13142 22636
rect 14921 22627 14979 22633
rect 14921 22593 14933 22627
rect 14967 22624 14979 22627
rect 15657 22627 15715 22633
rect 15657 22624 15669 22627
rect 14967 22596 15669 22624
rect 14967 22593 14979 22596
rect 14921 22587 14979 22593
rect 15657 22593 15669 22596
rect 15703 22624 15715 22627
rect 16666 22624 16672 22636
rect 15703 22596 16672 22624
rect 15703 22593 15715 22596
rect 15657 22587 15715 22593
rect 16666 22584 16672 22596
rect 16724 22584 16730 22636
rect 21358 22584 21364 22636
rect 21416 22624 21422 22636
rect 22373 22627 22431 22633
rect 22373 22624 22385 22627
rect 21416 22596 22385 22624
rect 21416 22584 21422 22596
rect 22373 22593 22385 22596
rect 22419 22593 22431 22627
rect 22373 22587 22431 22593
rect 7006 22516 7012 22568
rect 7064 22556 7070 22568
rect 8018 22565 8024 22568
rect 7101 22559 7159 22565
rect 7101 22556 7113 22559
rect 7064 22528 7113 22556
rect 7064 22516 7070 22528
rect 7101 22525 7113 22528
rect 7147 22556 7159 22559
rect 7745 22559 7803 22565
rect 7745 22556 7757 22559
rect 7147 22528 7757 22556
rect 7147 22525 7159 22528
rect 7101 22519 7159 22525
rect 7668 22432 7696 22528
rect 7745 22525 7757 22528
rect 7791 22525 7803 22559
rect 8012 22556 8024 22565
rect 7979 22528 8024 22556
rect 7745 22519 7803 22525
rect 8012 22519 8024 22528
rect 8018 22516 8024 22519
rect 8076 22516 8082 22568
rect 10134 22516 10140 22568
rect 10192 22556 10198 22568
rect 10597 22559 10655 22565
rect 10597 22556 10609 22559
rect 10192 22528 10609 22556
rect 10192 22516 10198 22528
rect 10597 22525 10609 22528
rect 10643 22525 10655 22559
rect 10597 22519 10655 22525
rect 12253 22559 12311 22565
rect 12253 22525 12265 22559
rect 12299 22556 12311 22559
rect 14185 22559 14243 22565
rect 12299 22528 13032 22556
rect 12299 22525 12311 22528
rect 12253 22519 12311 22525
rect 12802 22488 12808 22500
rect 12763 22460 12808 22488
rect 12802 22448 12808 22460
rect 12860 22448 12866 22500
rect 13004 22497 13032 22528
rect 14185 22525 14197 22559
rect 14231 22556 14243 22559
rect 15378 22556 15384 22568
rect 14231 22528 15384 22556
rect 14231 22525 14243 22528
rect 14185 22519 14243 22525
rect 15378 22516 15384 22528
rect 15436 22516 15442 22568
rect 16758 22556 16764 22568
rect 16671 22528 16764 22556
rect 16758 22516 16764 22528
rect 16816 22556 16822 22568
rect 17313 22559 17371 22565
rect 17313 22556 17325 22559
rect 16816 22528 17325 22556
rect 16816 22516 16822 22528
rect 17313 22525 17325 22528
rect 17359 22525 17371 22559
rect 17313 22519 17371 22525
rect 18509 22559 18567 22565
rect 18509 22525 18521 22559
rect 18555 22525 18567 22559
rect 18509 22519 18567 22525
rect 20533 22559 20591 22565
rect 20533 22525 20545 22559
rect 20579 22556 20591 22559
rect 21266 22556 21272 22568
rect 20579 22528 21272 22556
rect 20579 22525 20591 22528
rect 20533 22519 20591 22525
rect 12989 22491 13047 22497
rect 12989 22457 13001 22491
rect 13035 22488 13047 22491
rect 13446 22488 13452 22500
rect 13035 22460 13452 22488
rect 13035 22457 13047 22460
rect 12989 22451 13047 22457
rect 13446 22448 13452 22460
rect 13504 22448 13510 22500
rect 15286 22448 15292 22500
rect 15344 22488 15350 22500
rect 16025 22491 16083 22497
rect 16025 22488 16037 22491
rect 15344 22460 16037 22488
rect 15344 22448 15350 22460
rect 16025 22457 16037 22460
rect 16071 22488 16083 22491
rect 17678 22488 17684 22500
rect 16071 22460 17684 22488
rect 16071 22457 16083 22460
rect 16025 22451 16083 22457
rect 17678 22448 17684 22460
rect 17736 22488 17742 22500
rect 17773 22491 17831 22497
rect 17773 22488 17785 22491
rect 17736 22460 17785 22488
rect 17736 22448 17742 22460
rect 17773 22457 17785 22460
rect 17819 22488 17831 22491
rect 18325 22491 18383 22497
rect 18325 22488 18337 22491
rect 17819 22460 18337 22488
rect 17819 22457 17831 22460
rect 17773 22451 17831 22457
rect 18325 22457 18337 22460
rect 18371 22488 18383 22491
rect 18524 22488 18552 22519
rect 21266 22516 21272 22528
rect 21324 22556 21330 22568
rect 21637 22559 21695 22565
rect 21637 22556 21649 22559
rect 21324 22528 21649 22556
rect 21324 22516 21330 22528
rect 21637 22525 21649 22528
rect 21683 22525 21695 22559
rect 24581 22559 24639 22565
rect 24581 22556 24593 22559
rect 21637 22519 21695 22525
rect 24412 22528 24593 22556
rect 18371 22460 18552 22488
rect 18371 22457 18383 22460
rect 18325 22451 18383 22457
rect 18690 22448 18696 22500
rect 18748 22497 18754 22500
rect 18748 22491 18812 22497
rect 18748 22457 18766 22491
rect 18800 22457 18812 22491
rect 21358 22488 21364 22500
rect 21319 22460 21364 22488
rect 18748 22451 18812 22457
rect 18748 22448 18754 22451
rect 21358 22448 21364 22460
rect 21416 22448 21422 22500
rect 21542 22488 21548 22500
rect 21503 22460 21548 22488
rect 21542 22448 21548 22460
rect 21600 22448 21606 22500
rect 7650 22420 7656 22432
rect 7611 22392 7656 22420
rect 7650 22380 7656 22392
rect 7708 22380 7714 22432
rect 8294 22380 8300 22432
rect 8352 22420 8358 22432
rect 9125 22423 9183 22429
rect 9125 22420 9137 22423
rect 8352 22392 9137 22420
rect 8352 22380 8358 22392
rect 9125 22389 9137 22392
rect 9171 22389 9183 22423
rect 9674 22420 9680 22432
rect 9635 22392 9680 22420
rect 9125 22383 9183 22389
rect 9674 22380 9680 22392
rect 9732 22380 9738 22432
rect 10137 22423 10195 22429
rect 10137 22389 10149 22423
rect 10183 22420 10195 22423
rect 10778 22420 10784 22432
rect 10183 22392 10784 22420
rect 10183 22389 10195 22392
rect 10137 22383 10195 22389
rect 10778 22380 10784 22392
rect 10836 22380 10842 22432
rect 15102 22380 15108 22432
rect 15160 22420 15166 22432
rect 15565 22423 15623 22429
rect 15565 22420 15577 22423
rect 15160 22392 15577 22420
rect 15160 22380 15166 22392
rect 15565 22389 15577 22392
rect 15611 22389 15623 22423
rect 15565 22383 15623 22389
rect 19426 22380 19432 22432
rect 19484 22420 19490 22432
rect 19889 22423 19947 22429
rect 19889 22420 19901 22423
rect 19484 22392 19901 22420
rect 19484 22380 19490 22392
rect 19889 22389 19901 22392
rect 19935 22389 19947 22423
rect 21560 22420 21588 22448
rect 22005 22423 22063 22429
rect 22005 22420 22017 22423
rect 21560 22392 22017 22420
rect 19889 22383 19947 22389
rect 22005 22389 22017 22392
rect 22051 22389 22063 22423
rect 22005 22383 22063 22389
rect 24210 22380 24216 22432
rect 24268 22420 24274 22432
rect 24412 22429 24440 22528
rect 24581 22525 24593 22528
rect 24627 22525 24639 22559
rect 24581 22519 24639 22525
rect 24397 22423 24455 22429
rect 24397 22420 24409 22423
rect 24268 22392 24409 22420
rect 24268 22380 24274 22392
rect 24397 22389 24409 22392
rect 24443 22389 24455 22423
rect 24397 22383 24455 22389
rect 24854 22380 24860 22432
rect 24912 22420 24918 22432
rect 25225 22423 25283 22429
rect 25225 22420 25237 22423
rect 24912 22392 25237 22420
rect 24912 22380 24918 22392
rect 25225 22389 25237 22392
rect 25271 22420 25283 22423
rect 25774 22420 25780 22432
rect 25271 22392 25780 22420
rect 25271 22389 25283 22392
rect 25225 22383 25283 22389
rect 25774 22380 25780 22392
rect 25832 22380 25838 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 6638 22216 6644 22228
rect 6599 22188 6644 22216
rect 6638 22176 6644 22188
rect 6696 22176 6702 22228
rect 7834 22176 7840 22228
rect 7892 22216 7898 22228
rect 8205 22219 8263 22225
rect 8205 22216 8217 22219
rect 7892 22188 8217 22216
rect 7892 22176 7898 22188
rect 8205 22185 8217 22188
rect 8251 22185 8263 22219
rect 8205 22179 8263 22185
rect 10134 22176 10140 22228
rect 10192 22216 10198 22228
rect 10229 22219 10287 22225
rect 10229 22216 10241 22219
rect 10192 22188 10241 22216
rect 10192 22176 10198 22188
rect 10229 22185 10241 22188
rect 10275 22185 10287 22219
rect 10229 22179 10287 22185
rect 11701 22219 11759 22225
rect 11701 22185 11713 22219
rect 11747 22216 11759 22219
rect 11882 22216 11888 22228
rect 11747 22188 11888 22216
rect 11747 22185 11759 22188
rect 11701 22179 11759 22185
rect 11882 22176 11888 22188
rect 11940 22176 11946 22228
rect 12437 22219 12495 22225
rect 12437 22185 12449 22219
rect 12483 22216 12495 22219
rect 12618 22216 12624 22228
rect 12483 22188 12624 22216
rect 12483 22185 12495 22188
rect 12437 22179 12495 22185
rect 12618 22176 12624 22188
rect 12676 22176 12682 22228
rect 16209 22219 16267 22225
rect 16209 22185 16221 22219
rect 16255 22216 16267 22219
rect 16298 22216 16304 22228
rect 16255 22188 16304 22216
rect 16255 22185 16267 22188
rect 16209 22179 16267 22185
rect 16298 22176 16304 22188
rect 16356 22216 16362 22228
rect 16758 22216 16764 22228
rect 16356 22188 16764 22216
rect 16356 22176 16362 22188
rect 16758 22176 16764 22188
rect 16816 22176 16822 22228
rect 17218 22176 17224 22228
rect 17276 22216 17282 22228
rect 17770 22216 17776 22228
rect 17276 22188 17776 22216
rect 17276 22176 17282 22188
rect 17770 22176 17776 22188
rect 17828 22176 17834 22228
rect 19242 22216 19248 22228
rect 19168 22188 19248 22216
rect 7561 22151 7619 22157
rect 7561 22117 7573 22151
rect 7607 22148 7619 22151
rect 8018 22148 8024 22160
rect 7607 22120 8024 22148
rect 7607 22117 7619 22120
rect 7561 22111 7619 22117
rect 8018 22108 8024 22120
rect 8076 22108 8082 22160
rect 8294 22108 8300 22160
rect 8352 22148 8358 22160
rect 11790 22148 11796 22160
rect 8352 22120 8397 22148
rect 11751 22120 11796 22148
rect 8352 22108 8358 22120
rect 11790 22108 11796 22120
rect 11848 22108 11854 22160
rect 13998 22148 14004 22160
rect 13911 22120 14004 22148
rect 13998 22108 14004 22120
rect 14056 22148 14062 22160
rect 14642 22148 14648 22160
rect 14056 22120 14648 22148
rect 14056 22108 14062 22120
rect 14642 22108 14648 22120
rect 14700 22108 14706 22160
rect 17862 22148 17868 22160
rect 17823 22120 17868 22148
rect 17862 22108 17868 22120
rect 17920 22148 17926 22160
rect 18509 22151 18567 22157
rect 18509 22148 18521 22151
rect 17920 22120 18521 22148
rect 17920 22108 17926 22120
rect 18509 22117 18521 22120
rect 18555 22148 18567 22151
rect 18690 22148 18696 22160
rect 18555 22120 18696 22148
rect 18555 22117 18567 22120
rect 18509 22111 18567 22117
rect 18690 22108 18696 22120
rect 18748 22108 18754 22160
rect 19168 22092 19196 22188
rect 19242 22176 19248 22188
rect 19300 22176 19306 22228
rect 21177 22219 21235 22225
rect 21177 22185 21189 22219
rect 21223 22216 21235 22219
rect 21266 22216 21272 22228
rect 21223 22188 21272 22216
rect 21223 22185 21235 22188
rect 21177 22179 21235 22185
rect 21266 22176 21272 22188
rect 21324 22176 21330 22228
rect 19334 22148 19340 22160
rect 19295 22120 19340 22148
rect 19334 22108 19340 22120
rect 19392 22108 19398 22160
rect 22186 22148 22192 22160
rect 22147 22120 22192 22148
rect 22186 22108 22192 22120
rect 22244 22108 22250 22160
rect 11514 22080 11520 22092
rect 11475 22052 11520 22080
rect 11514 22040 11520 22052
rect 11572 22080 11578 22092
rect 11698 22080 11704 22092
rect 11572 22052 11704 22080
rect 11572 22040 11578 22052
rect 11698 22040 11704 22052
rect 11756 22040 11762 22092
rect 13814 22040 13820 22092
rect 13872 22080 13878 22092
rect 15013 22083 15071 22089
rect 15013 22080 15025 22083
rect 13872 22052 15025 22080
rect 13872 22040 13878 22052
rect 15013 22049 15025 22052
rect 15059 22080 15071 22083
rect 15102 22080 15108 22092
rect 15059 22052 15108 22080
rect 15059 22049 15071 22052
rect 15013 22043 15071 22049
rect 15102 22040 15108 22052
rect 15160 22040 15166 22092
rect 19150 22040 19156 22092
rect 19208 22040 19214 22092
rect 22281 22083 22339 22089
rect 22281 22049 22293 22083
rect 22327 22080 22339 22083
rect 23014 22080 23020 22092
rect 22327 22052 23020 22080
rect 22327 22049 22339 22052
rect 22281 22043 22339 22049
rect 23014 22040 23020 22052
rect 23072 22080 23078 22092
rect 23457 22083 23515 22089
rect 23457 22080 23469 22083
rect 23072 22052 23469 22080
rect 23072 22040 23078 22052
rect 23457 22049 23469 22052
rect 23503 22049 23515 22083
rect 23457 22043 23515 22049
rect 7374 21972 7380 22024
rect 7432 22012 7438 22024
rect 8113 22015 8171 22021
rect 8113 22012 8125 22015
rect 7432 21984 8125 22012
rect 7432 21972 7438 21984
rect 8113 21981 8125 21984
rect 8159 22012 8171 22015
rect 8202 22012 8208 22024
rect 8159 21984 8208 22012
rect 8159 21981 8171 21984
rect 8113 21975 8171 21981
rect 8202 21972 8208 21984
rect 8260 21972 8266 22024
rect 12805 22015 12863 22021
rect 12805 21981 12817 22015
rect 12851 22012 12863 22015
rect 13909 22015 13967 22021
rect 13909 22012 13921 22015
rect 12851 21984 13921 22012
rect 12851 21981 12863 21984
rect 12805 21975 12863 21981
rect 13909 21981 13921 21984
rect 13955 21981 13967 22015
rect 14090 22012 14096 22024
rect 14051 21984 14096 22012
rect 13909 21975 13967 21981
rect 11241 21947 11299 21953
rect 11241 21913 11253 21947
rect 11287 21944 11299 21947
rect 12066 21944 12072 21956
rect 11287 21916 12072 21944
rect 11287 21913 11299 21916
rect 11241 21907 11299 21913
rect 12066 21904 12072 21916
rect 12124 21904 12130 21956
rect 13538 21944 13544 21956
rect 13499 21916 13544 21944
rect 13538 21904 13544 21916
rect 13596 21904 13602 21956
rect 13924 21944 13952 21975
rect 14090 21972 14096 21984
rect 14148 21972 14154 22024
rect 16206 22012 16212 22024
rect 16167 21984 16212 22012
rect 16206 21972 16212 21984
rect 16264 21972 16270 22024
rect 16301 22015 16359 22021
rect 16301 21981 16313 22015
rect 16347 22012 16359 22015
rect 16390 22012 16396 22024
rect 16347 21984 16396 22012
rect 16347 21981 16359 21984
rect 16301 21975 16359 21981
rect 16390 21972 16396 21984
rect 16448 21972 16454 22024
rect 17770 22012 17776 22024
rect 17731 21984 17776 22012
rect 17770 21972 17776 21984
rect 17828 21972 17834 22024
rect 19245 22015 19303 22021
rect 19245 22012 19257 22015
rect 18769 21984 19257 22012
rect 14182 21944 14188 21956
rect 13924 21916 14188 21944
rect 14182 21904 14188 21916
rect 14240 21904 14246 21956
rect 15746 21944 15752 21956
rect 15707 21916 15752 21944
rect 15746 21904 15752 21916
rect 15804 21904 15810 21956
rect 17313 21947 17371 21953
rect 17313 21913 17325 21947
rect 17359 21944 17371 21947
rect 18769 21944 18797 21984
rect 19245 21981 19257 21984
rect 19291 21981 19303 22015
rect 19426 22012 19432 22024
rect 19387 21984 19432 22012
rect 19245 21975 19303 21981
rect 18874 21944 18880 21956
rect 17359 21916 18797 21944
rect 18835 21916 18880 21944
rect 17359 21913 17371 21916
rect 17313 21907 17371 21913
rect 18874 21904 18880 21916
rect 18932 21904 18938 21956
rect 19260 21944 19288 21975
rect 19426 21972 19432 21984
rect 19484 21972 19490 22024
rect 21545 22015 21603 22021
rect 21545 21981 21557 22015
rect 21591 22012 21603 22015
rect 22189 22015 22247 22021
rect 22189 22012 22201 22015
rect 21591 21984 22201 22012
rect 21591 21981 21603 21984
rect 21545 21975 21603 21981
rect 22189 21981 22201 21984
rect 22235 22012 22247 22015
rect 22370 22012 22376 22024
rect 22235 21984 22376 22012
rect 22235 21981 22247 21984
rect 22189 21975 22247 21981
rect 22370 21972 22376 21984
rect 22428 21972 22434 22024
rect 23198 22012 23204 22024
rect 23159 21984 23204 22012
rect 23198 21972 23204 21984
rect 23256 21972 23262 22024
rect 19797 21947 19855 21953
rect 19797 21944 19809 21947
rect 19260 21916 19809 21944
rect 19797 21913 19809 21916
rect 19843 21913 19855 21947
rect 19797 21907 19855 21913
rect 7742 21876 7748 21888
rect 7703 21848 7748 21876
rect 7742 21836 7748 21848
rect 7800 21836 7806 21888
rect 10781 21879 10839 21885
rect 10781 21845 10793 21879
rect 10827 21876 10839 21879
rect 11330 21876 11336 21888
rect 10827 21848 11336 21876
rect 10827 21845 10839 21848
rect 10781 21839 10839 21845
rect 11330 21836 11336 21848
rect 11388 21836 11394 21888
rect 13170 21876 13176 21888
rect 13131 21848 13176 21876
rect 13170 21836 13176 21848
rect 13228 21836 13234 21888
rect 15562 21876 15568 21888
rect 15523 21848 15568 21876
rect 15562 21836 15568 21848
rect 15620 21836 15626 21888
rect 16022 21836 16028 21888
rect 16080 21876 16086 21888
rect 16482 21876 16488 21888
rect 16080 21848 16488 21876
rect 16080 21836 16086 21848
rect 16482 21836 16488 21848
rect 16540 21836 16546 21888
rect 16666 21876 16672 21888
rect 16627 21848 16672 21876
rect 16666 21836 16672 21848
rect 16724 21836 16730 21888
rect 20162 21876 20168 21888
rect 20123 21848 20168 21876
rect 20162 21836 20168 21848
rect 20220 21836 20226 21888
rect 21542 21836 21548 21888
rect 21600 21876 21606 21888
rect 21729 21879 21787 21885
rect 21729 21876 21741 21879
rect 21600 21848 21741 21876
rect 21600 21836 21606 21848
rect 21729 21845 21741 21848
rect 21775 21845 21787 21879
rect 21729 21839 21787 21845
rect 23474 21836 23480 21888
rect 23532 21876 23538 21888
rect 24581 21879 24639 21885
rect 24581 21876 24593 21879
rect 23532 21848 24593 21876
rect 23532 21836 23538 21848
rect 24581 21845 24593 21848
rect 24627 21845 24639 21879
rect 24581 21839 24639 21845
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 13817 21675 13875 21681
rect 13817 21641 13829 21675
rect 13863 21672 13875 21675
rect 13998 21672 14004 21684
rect 13863 21644 14004 21672
rect 13863 21641 13875 21644
rect 13817 21635 13875 21641
rect 13998 21632 14004 21644
rect 14056 21632 14062 21684
rect 14734 21632 14740 21684
rect 14792 21672 14798 21684
rect 14921 21675 14979 21681
rect 14921 21672 14933 21675
rect 14792 21644 14933 21672
rect 14792 21632 14798 21644
rect 14921 21641 14933 21644
rect 14967 21641 14979 21675
rect 14921 21635 14979 21641
rect 16206 21632 16212 21684
rect 16264 21672 16270 21684
rect 16485 21675 16543 21681
rect 16485 21672 16497 21675
rect 16264 21644 16497 21672
rect 16264 21632 16270 21644
rect 16485 21641 16497 21644
rect 16531 21641 16543 21675
rect 16485 21635 16543 21641
rect 17218 21632 17224 21684
rect 17276 21672 17282 21684
rect 17405 21675 17463 21681
rect 17405 21672 17417 21675
rect 17276 21644 17417 21672
rect 17276 21632 17282 21644
rect 17405 21641 17417 21644
rect 17451 21641 17463 21675
rect 17770 21672 17776 21684
rect 17731 21644 17776 21672
rect 17405 21635 17463 21641
rect 17770 21632 17776 21644
rect 17828 21632 17834 21684
rect 19334 21672 19340 21684
rect 19295 21644 19340 21672
rect 19334 21632 19340 21644
rect 19392 21632 19398 21684
rect 20346 21672 20352 21684
rect 20307 21644 20352 21672
rect 20346 21632 20352 21644
rect 20404 21632 20410 21684
rect 10781 21607 10839 21613
rect 10781 21573 10793 21607
rect 10827 21573 10839 21607
rect 12802 21604 12808 21616
rect 12763 21576 12808 21604
rect 10781 21567 10839 21573
rect 7650 21496 7656 21548
rect 7708 21536 7714 21548
rect 7929 21539 7987 21545
rect 7929 21536 7941 21539
rect 7708 21508 7941 21536
rect 7708 21496 7714 21508
rect 7929 21505 7941 21508
rect 7975 21536 7987 21539
rect 8113 21539 8171 21545
rect 8113 21536 8125 21539
rect 7975 21508 8125 21536
rect 7975 21505 7987 21508
rect 7929 21499 7987 21505
rect 8113 21505 8125 21508
rect 8159 21505 8171 21539
rect 8113 21499 8171 21505
rect 10796 21468 10824 21567
rect 12802 21564 12808 21576
rect 12860 21564 12866 21616
rect 13906 21564 13912 21616
rect 13964 21604 13970 21616
rect 14553 21607 14611 21613
rect 14553 21604 14565 21607
rect 13964 21576 14565 21604
rect 13964 21564 13970 21576
rect 14553 21573 14565 21576
rect 14599 21573 14611 21607
rect 14553 21567 14611 21573
rect 15197 21607 15255 21613
rect 15197 21573 15209 21607
rect 15243 21604 15255 21607
rect 17586 21604 17592 21616
rect 15243 21576 17592 21604
rect 15243 21573 15255 21576
rect 15197 21567 15255 21573
rect 11146 21536 11152 21548
rect 11107 21508 11152 21536
rect 11146 21496 11152 21508
rect 11204 21496 11210 21548
rect 11330 21536 11336 21548
rect 11291 21508 11336 21536
rect 11330 21496 11336 21508
rect 11388 21496 11394 21548
rect 13265 21539 13323 21545
rect 13265 21505 13277 21539
rect 13311 21505 13323 21539
rect 14568 21536 14596 21567
rect 17586 21564 17592 21576
rect 17644 21564 17650 21616
rect 15565 21539 15623 21545
rect 15565 21536 15577 21539
rect 14568 21508 15577 21536
rect 13265 21499 13323 21505
rect 15565 21505 15577 21508
rect 15611 21505 15623 21539
rect 16850 21536 16856 21548
rect 16811 21508 16856 21536
rect 15565 21499 15623 21505
rect 13280 21468 13308 21499
rect 16850 21496 16856 21508
rect 16908 21496 16914 21548
rect 17788 21536 17816 21632
rect 21726 21564 21732 21616
rect 21784 21604 21790 21616
rect 21821 21607 21879 21613
rect 21821 21604 21833 21607
rect 21784 21576 21833 21604
rect 21784 21564 21790 21576
rect 21821 21573 21833 21576
rect 21867 21573 21879 21607
rect 21821 21567 21879 21573
rect 18049 21539 18107 21545
rect 18049 21536 18061 21539
rect 17788 21508 18061 21536
rect 18049 21505 18061 21508
rect 18095 21505 18107 21539
rect 18049 21499 18107 21505
rect 18785 21539 18843 21545
rect 18785 21505 18797 21539
rect 18831 21536 18843 21539
rect 18966 21536 18972 21548
rect 18831 21508 18972 21536
rect 18831 21505 18843 21508
rect 18785 21499 18843 21505
rect 18966 21496 18972 21508
rect 19024 21536 19030 21548
rect 19797 21539 19855 21545
rect 19797 21536 19809 21539
rect 19024 21508 19809 21536
rect 19024 21496 19030 21508
rect 19797 21505 19809 21508
rect 19843 21536 19855 21539
rect 19978 21536 19984 21548
rect 19843 21508 19984 21536
rect 19843 21505 19855 21508
rect 19797 21499 19855 21505
rect 19978 21496 19984 21508
rect 20036 21496 20042 21548
rect 21174 21496 21180 21548
rect 21232 21536 21238 21548
rect 22189 21539 22247 21545
rect 22189 21536 22201 21539
rect 21232 21508 22201 21536
rect 21232 21496 21238 21508
rect 22189 21505 22201 21508
rect 22235 21536 22247 21539
rect 22462 21536 22468 21548
rect 22235 21508 22468 21536
rect 22235 21505 22247 21508
rect 22189 21499 22247 21505
rect 22462 21496 22468 21508
rect 22520 21496 22526 21548
rect 24210 21536 24216 21548
rect 24171 21508 24216 21536
rect 24210 21496 24216 21508
rect 24268 21496 24274 21548
rect 14182 21468 14188 21480
rect 10796 21440 13216 21468
rect 13280 21440 14188 21468
rect 13188 21412 13216 21440
rect 14182 21428 14188 21440
rect 14240 21428 14246 21480
rect 16482 21428 16488 21480
rect 16540 21468 16546 21480
rect 16666 21468 16672 21480
rect 16540 21440 16672 21468
rect 16540 21428 16546 21440
rect 16666 21428 16672 21440
rect 16724 21428 16730 21480
rect 18690 21428 18696 21480
rect 18748 21468 18754 21480
rect 19889 21471 19947 21477
rect 19889 21468 19901 21471
rect 18748 21440 19901 21468
rect 18748 21428 18754 21440
rect 19889 21437 19901 21440
rect 19935 21468 19947 21471
rect 20346 21468 20352 21480
rect 19935 21440 20352 21468
rect 19935 21437 19947 21440
rect 19889 21431 19947 21437
rect 20346 21428 20352 21440
rect 20404 21428 20410 21480
rect 20714 21428 20720 21480
rect 20772 21468 20778 21480
rect 21637 21471 21695 21477
rect 21637 21468 21649 21471
rect 20772 21440 21649 21468
rect 20772 21428 20778 21440
rect 21637 21437 21649 21440
rect 21683 21468 21695 21471
rect 23750 21468 23756 21480
rect 21683 21440 23756 21468
rect 21683 21437 21695 21440
rect 21637 21431 21695 21437
rect 7285 21403 7343 21409
rect 7285 21369 7297 21403
rect 7331 21400 7343 21403
rect 7653 21403 7711 21409
rect 7653 21400 7665 21403
rect 7331 21372 7665 21400
rect 7331 21369 7343 21372
rect 7285 21363 7343 21369
rect 7653 21369 7665 21372
rect 7699 21400 7711 21403
rect 8294 21400 8300 21412
rect 7699 21372 8300 21400
rect 7699 21369 7711 21372
rect 7653 21363 7711 21369
rect 8294 21360 8300 21372
rect 8352 21409 8358 21412
rect 8352 21403 8416 21409
rect 8352 21369 8370 21403
rect 8404 21369 8416 21403
rect 8352 21363 8416 21369
rect 8352 21360 8358 21363
rect 11054 21360 11060 21412
rect 11112 21400 11118 21412
rect 11701 21403 11759 21409
rect 11701 21400 11713 21403
rect 11112 21372 11713 21400
rect 11112 21360 11118 21372
rect 11701 21369 11713 21372
rect 11747 21400 11759 21403
rect 11882 21400 11888 21412
rect 11747 21372 11888 21400
rect 11747 21369 11759 21372
rect 11701 21363 11759 21369
rect 11882 21360 11888 21372
rect 11940 21360 11946 21412
rect 13170 21360 13176 21412
rect 13228 21400 13234 21412
rect 13265 21403 13323 21409
rect 13265 21400 13277 21403
rect 13228 21372 13277 21400
rect 13228 21360 13234 21372
rect 13265 21369 13277 21372
rect 13311 21369 13323 21403
rect 13265 21363 13323 21369
rect 13357 21403 13415 21409
rect 13357 21369 13369 21403
rect 13403 21400 13415 21403
rect 13538 21400 13544 21412
rect 13403 21372 13544 21400
rect 13403 21369 13415 21372
rect 13357 21363 13415 21369
rect 13538 21360 13544 21372
rect 13596 21360 13602 21412
rect 15562 21360 15568 21412
rect 15620 21400 15626 21412
rect 15749 21403 15807 21409
rect 15749 21400 15761 21403
rect 15620 21372 15761 21400
rect 15620 21360 15626 21372
rect 15749 21369 15761 21372
rect 15795 21400 15807 21403
rect 16574 21400 16580 21412
rect 15795 21372 16580 21400
rect 15795 21369 15807 21372
rect 15749 21363 15807 21369
rect 16574 21360 16580 21372
rect 16632 21360 16638 21412
rect 22296 21409 22324 21440
rect 23750 21428 23756 21440
rect 23808 21428 23814 21480
rect 23937 21471 23995 21477
rect 23937 21437 23949 21471
rect 23983 21468 23995 21471
rect 24670 21468 24676 21480
rect 23983 21440 24676 21468
rect 23983 21437 23995 21440
rect 23937 21431 23995 21437
rect 24670 21428 24676 21440
rect 24728 21428 24734 21480
rect 22281 21403 22339 21409
rect 22281 21369 22293 21403
rect 22327 21369 22339 21403
rect 22281 21363 22339 21369
rect 22373 21403 22431 21409
rect 22373 21369 22385 21403
rect 22419 21400 22431 21403
rect 22554 21400 22560 21412
rect 22419 21372 22560 21400
rect 22419 21369 22431 21372
rect 22373 21363 22431 21369
rect 22554 21360 22560 21372
rect 22612 21360 22618 21412
rect 22738 21360 22744 21412
rect 22796 21400 22802 21412
rect 23198 21400 23204 21412
rect 22796 21372 23204 21400
rect 22796 21360 22802 21372
rect 23198 21360 23204 21372
rect 23256 21360 23262 21412
rect 9122 21292 9128 21344
rect 9180 21332 9186 21344
rect 9493 21335 9551 21341
rect 9493 21332 9505 21335
rect 9180 21304 9505 21332
rect 9180 21292 9186 21304
rect 9493 21301 9505 21304
rect 9539 21301 9551 21335
rect 9493 21295 9551 21301
rect 9766 21292 9772 21344
rect 9824 21332 9830 21344
rect 10597 21335 10655 21341
rect 10597 21332 10609 21335
rect 9824 21304 10609 21332
rect 9824 21292 9830 21304
rect 10597 21301 10609 21304
rect 10643 21332 10655 21335
rect 11241 21335 11299 21341
rect 11241 21332 11253 21335
rect 10643 21304 11253 21332
rect 10643 21301 10655 21304
rect 10597 21295 10655 21301
rect 11241 21301 11253 21304
rect 11287 21332 11299 21335
rect 11974 21332 11980 21344
rect 11287 21304 11980 21332
rect 11287 21301 11299 21304
rect 11241 21295 11299 21301
rect 11974 21292 11980 21304
rect 12032 21292 12038 21344
rect 12250 21332 12256 21344
rect 12211 21304 12256 21332
rect 12250 21292 12256 21304
rect 12308 21292 12314 21344
rect 14734 21292 14740 21344
rect 14792 21332 14798 21344
rect 15654 21332 15660 21344
rect 14792 21304 15660 21332
rect 14792 21292 14798 21304
rect 15654 21292 15660 21304
rect 15712 21292 15718 21344
rect 16114 21332 16120 21344
rect 16075 21304 16120 21332
rect 16114 21292 16120 21304
rect 16172 21292 16178 21344
rect 19058 21292 19064 21344
rect 19116 21332 19122 21344
rect 19153 21335 19211 21341
rect 19153 21332 19165 21335
rect 19116 21304 19165 21332
rect 19116 21292 19122 21304
rect 19153 21301 19165 21304
rect 19199 21332 19211 21335
rect 19797 21335 19855 21341
rect 19797 21332 19809 21335
rect 19199 21304 19809 21332
rect 19199 21301 19211 21304
rect 19153 21295 19211 21301
rect 19797 21301 19809 21304
rect 19843 21332 19855 21335
rect 20070 21332 20076 21344
rect 19843 21304 20076 21332
rect 19843 21301 19855 21304
rect 19797 21295 19855 21301
rect 20070 21292 20076 21304
rect 20128 21292 20134 21344
rect 20806 21332 20812 21344
rect 20767 21304 20812 21332
rect 20806 21292 20812 21304
rect 20864 21292 20870 21344
rect 21174 21332 21180 21344
rect 21135 21304 21180 21332
rect 21174 21292 21180 21304
rect 21232 21292 21238 21344
rect 22002 21292 22008 21344
rect 22060 21332 22066 21344
rect 22925 21335 22983 21341
rect 22925 21332 22937 21335
rect 22060 21304 22937 21332
rect 22060 21292 22066 21304
rect 22925 21301 22937 21304
rect 22971 21332 22983 21335
rect 23014 21332 23020 21344
rect 22971 21304 23020 21332
rect 22971 21301 22983 21304
rect 22925 21295 22983 21301
rect 23014 21292 23020 21304
rect 23072 21292 23078 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 7374 21128 7380 21140
rect 7335 21100 7380 21128
rect 7374 21088 7380 21100
rect 7432 21088 7438 21140
rect 7745 21131 7803 21137
rect 7745 21097 7757 21131
rect 7791 21128 7803 21131
rect 7834 21128 7840 21140
rect 7791 21100 7840 21128
rect 7791 21097 7803 21100
rect 7745 21091 7803 21097
rect 7834 21088 7840 21100
rect 7892 21088 7898 21140
rect 9122 21128 9128 21140
rect 8680 21100 9128 21128
rect 8386 21060 8392 21072
rect 8347 21032 8392 21060
rect 8386 21020 8392 21032
rect 8444 21020 8450 21072
rect 8478 21020 8484 21072
rect 8536 21060 8542 21072
rect 8680 21069 8708 21100
rect 9122 21088 9128 21100
rect 9180 21088 9186 21140
rect 10781 21131 10839 21137
rect 10781 21097 10793 21131
rect 10827 21128 10839 21131
rect 11146 21128 11152 21140
rect 10827 21100 11152 21128
rect 10827 21097 10839 21100
rect 10781 21091 10839 21097
rect 11146 21088 11152 21100
rect 11204 21088 11210 21140
rect 11241 21131 11299 21137
rect 11241 21097 11253 21131
rect 11287 21128 11299 21131
rect 11514 21128 11520 21140
rect 11287 21100 11520 21128
rect 11287 21097 11299 21100
rect 11241 21091 11299 21097
rect 11514 21088 11520 21100
rect 11572 21088 11578 21140
rect 11609 21131 11667 21137
rect 11609 21097 11621 21131
rect 11655 21128 11667 21131
rect 11790 21128 11796 21140
rect 11655 21100 11796 21128
rect 11655 21097 11667 21100
rect 11609 21091 11667 21097
rect 11790 21088 11796 21100
rect 11848 21088 11854 21140
rect 12250 21088 12256 21140
rect 12308 21128 12314 21140
rect 13538 21128 13544 21140
rect 12308 21100 13544 21128
rect 12308 21088 12314 21100
rect 13538 21088 13544 21100
rect 13596 21088 13602 21140
rect 14090 21128 14096 21140
rect 14003 21100 14096 21128
rect 14090 21088 14096 21100
rect 14148 21128 14154 21140
rect 15105 21131 15163 21137
rect 15105 21128 15117 21131
rect 14148 21100 15117 21128
rect 14148 21088 14154 21100
rect 15105 21097 15117 21100
rect 15151 21128 15163 21131
rect 16390 21128 16396 21140
rect 15151 21100 16396 21128
rect 15151 21097 15163 21100
rect 15105 21091 15163 21097
rect 16390 21088 16396 21100
rect 16448 21088 16454 21140
rect 17586 21128 17592 21140
rect 17547 21100 17592 21128
rect 17586 21088 17592 21100
rect 17644 21128 17650 21140
rect 18325 21131 18383 21137
rect 18325 21128 18337 21131
rect 17644 21100 18337 21128
rect 17644 21088 17650 21100
rect 18325 21097 18337 21100
rect 18371 21097 18383 21131
rect 18325 21091 18383 21097
rect 19245 21131 19303 21137
rect 19245 21097 19257 21131
rect 19291 21128 19303 21131
rect 19334 21128 19340 21140
rect 19291 21100 19340 21128
rect 19291 21097 19303 21100
rect 19245 21091 19303 21097
rect 19334 21088 19340 21100
rect 19392 21088 19398 21140
rect 20717 21131 20775 21137
rect 20717 21097 20729 21131
rect 20763 21128 20775 21131
rect 20806 21128 20812 21140
rect 20763 21100 20812 21128
rect 20763 21097 20775 21100
rect 20717 21091 20775 21097
rect 20806 21088 20812 21100
rect 20864 21128 20870 21140
rect 22002 21128 22008 21140
rect 20864 21100 21588 21128
rect 21963 21100 22008 21128
rect 20864 21088 20870 21100
rect 8573 21063 8631 21069
rect 8573 21060 8585 21063
rect 8536 21032 8585 21060
rect 8536 21020 8542 21032
rect 8573 21029 8585 21032
rect 8619 21029 8631 21063
rect 8573 21023 8631 21029
rect 8665 21063 8723 21069
rect 8665 21029 8677 21063
rect 8711 21029 8723 21063
rect 8665 21023 8723 21029
rect 11330 21020 11336 21072
rect 11388 21060 11394 21072
rect 11946 21063 12004 21069
rect 11946 21060 11958 21063
rect 11388 21032 11958 21060
rect 11388 21020 11394 21032
rect 11946 21029 11958 21032
rect 11992 21060 12004 21063
rect 12066 21060 12072 21072
rect 11992 21032 12072 21060
rect 11992 21029 12004 21032
rect 11946 21023 12004 21029
rect 12066 21020 12072 21032
rect 12124 21020 12130 21072
rect 15470 21020 15476 21072
rect 15528 21060 15534 21072
rect 16758 21060 16764 21072
rect 15528 21032 16764 21060
rect 15528 21020 15534 21032
rect 16758 21020 16764 21032
rect 16816 21020 16822 21072
rect 17313 21063 17371 21069
rect 17313 21029 17325 21063
rect 17359 21060 17371 21063
rect 17770 21060 17776 21072
rect 17359 21032 17776 21060
rect 17359 21029 17371 21032
rect 17313 21023 17371 21029
rect 17770 21020 17776 21032
rect 17828 21020 17834 21072
rect 17862 21020 17868 21072
rect 17920 21060 17926 21072
rect 18138 21060 18144 21072
rect 17920 21032 18144 21060
rect 17920 21020 17926 21032
rect 18138 21020 18144 21032
rect 18196 21020 18202 21072
rect 18877 21063 18935 21069
rect 18877 21029 18889 21063
rect 18923 21060 18935 21063
rect 19426 21060 19432 21072
rect 18923 21032 19432 21060
rect 18923 21029 18935 21032
rect 18877 21023 18935 21029
rect 19426 21020 19432 21032
rect 19484 21020 19490 21072
rect 19518 21020 19524 21072
rect 19576 21060 19582 21072
rect 21560 21069 21588 21100
rect 22002 21088 22008 21100
rect 22060 21088 22066 21140
rect 22186 21088 22192 21140
rect 22244 21128 22250 21140
rect 22281 21131 22339 21137
rect 22281 21128 22293 21131
rect 22244 21100 22293 21128
rect 22244 21088 22250 21100
rect 22281 21097 22293 21100
rect 22327 21097 22339 21131
rect 22554 21128 22560 21140
rect 22281 21091 22339 21097
rect 22388 21100 22560 21128
rect 19613 21063 19671 21069
rect 19613 21060 19625 21063
rect 19576 21032 19625 21060
rect 19576 21020 19582 21032
rect 19613 21029 19625 21032
rect 19659 21029 19671 21063
rect 19613 21023 19671 21029
rect 21453 21063 21511 21069
rect 21453 21029 21465 21063
rect 21499 21029 21511 21063
rect 21453 21023 21511 21029
rect 21545 21063 21603 21069
rect 21545 21029 21557 21063
rect 21591 21060 21603 21063
rect 21591 21032 22140 21060
rect 21591 21029 21603 21032
rect 21545 21023 21603 21029
rect 15556 20995 15614 21001
rect 15556 20961 15568 20995
rect 15602 20992 15614 20995
rect 15838 20992 15844 21004
rect 15602 20964 15844 20992
rect 15602 20961 15614 20964
rect 15556 20955 15614 20961
rect 15838 20952 15844 20964
rect 15896 20952 15902 21004
rect 19337 20995 19395 21001
rect 19337 20961 19349 20995
rect 19383 20992 19395 20995
rect 20162 20992 20168 21004
rect 19383 20964 20168 20992
rect 19383 20961 19395 20964
rect 19337 20955 19395 20961
rect 20162 20952 20168 20964
rect 20220 20952 20226 21004
rect 20806 20952 20812 21004
rect 20864 20992 20870 21004
rect 21468 20992 21496 21023
rect 20864 20964 21496 20992
rect 22112 20992 22140 21032
rect 22388 20992 22416 21100
rect 22554 21088 22560 21100
rect 22612 21088 22618 21140
rect 23014 21088 23020 21140
rect 23072 21128 23078 21140
rect 23937 21131 23995 21137
rect 23937 21128 23949 21131
rect 23072 21100 23949 21128
rect 23072 21088 23078 21100
rect 23937 21097 23949 21100
rect 23983 21097 23995 21131
rect 23937 21091 23995 21097
rect 22922 21020 22928 21072
rect 22980 21060 22986 21072
rect 23842 21060 23848 21072
rect 22980 21032 23848 21060
rect 22980 21020 22986 21032
rect 23842 21020 23848 21032
rect 23900 21020 23906 21072
rect 22112 20964 22416 20992
rect 20864 20952 20870 20964
rect 22462 20952 22468 21004
rect 22520 20992 22526 21004
rect 22813 20995 22871 21001
rect 22813 20992 22825 20995
rect 22520 20964 22825 20992
rect 22520 20952 22526 20964
rect 22813 20961 22825 20964
rect 22859 20961 22871 20995
rect 22813 20955 22871 20961
rect 9677 20927 9735 20933
rect 9677 20893 9689 20927
rect 9723 20924 9735 20927
rect 9858 20924 9864 20936
rect 9723 20896 9864 20924
rect 9723 20893 9735 20896
rect 9677 20887 9735 20893
rect 9858 20884 9864 20896
rect 9916 20884 9922 20936
rect 11698 20924 11704 20936
rect 11659 20896 11704 20924
rect 11698 20884 11704 20896
rect 11756 20884 11762 20936
rect 13814 20884 13820 20936
rect 13872 20924 13878 20936
rect 14185 20927 14243 20933
rect 14185 20924 14197 20927
rect 13872 20896 14197 20924
rect 13872 20884 13878 20896
rect 14185 20893 14197 20896
rect 14231 20893 14243 20927
rect 15286 20924 15292 20936
rect 15247 20896 15292 20924
rect 14185 20887 14243 20893
rect 15286 20884 15292 20896
rect 15344 20884 15350 20936
rect 18322 20884 18328 20936
rect 18380 20924 18386 20936
rect 18417 20927 18475 20933
rect 18417 20924 18429 20927
rect 18380 20896 18429 20924
rect 18380 20884 18386 20896
rect 18417 20893 18429 20896
rect 18463 20893 18475 20927
rect 18417 20887 18475 20893
rect 20714 20884 20720 20936
rect 20772 20924 20778 20936
rect 21453 20927 21511 20933
rect 21453 20924 21465 20927
rect 20772 20896 21465 20924
rect 20772 20884 20778 20896
rect 21453 20893 21465 20896
rect 21499 20924 21511 20927
rect 21910 20924 21916 20936
rect 21499 20896 21916 20924
rect 21499 20893 21511 20896
rect 21453 20887 21511 20893
rect 21910 20884 21916 20896
rect 21968 20884 21974 20936
rect 22557 20927 22615 20933
rect 22557 20893 22569 20927
rect 22603 20893 22615 20927
rect 22557 20887 22615 20893
rect 20993 20859 21051 20865
rect 20993 20825 21005 20859
rect 21039 20856 21051 20859
rect 22002 20856 22008 20868
rect 21039 20828 22008 20856
rect 21039 20825 21051 20828
rect 20993 20819 21051 20825
rect 22002 20816 22008 20828
rect 22060 20816 22066 20868
rect 8110 20788 8116 20800
rect 8071 20760 8116 20788
rect 8110 20748 8116 20760
rect 8168 20748 8174 20800
rect 13081 20791 13139 20797
rect 13081 20757 13093 20791
rect 13127 20788 13139 20791
rect 13538 20788 13544 20800
rect 13127 20760 13544 20788
rect 13127 20757 13139 20760
rect 13081 20751 13139 20757
rect 13538 20748 13544 20760
rect 13596 20788 13602 20800
rect 13633 20791 13691 20797
rect 13633 20788 13645 20791
rect 13596 20760 13645 20788
rect 13596 20748 13602 20760
rect 13633 20757 13645 20760
rect 13679 20757 13691 20791
rect 13633 20751 13691 20757
rect 16574 20748 16580 20800
rect 16632 20788 16638 20800
rect 16669 20791 16727 20797
rect 16669 20788 16681 20791
rect 16632 20760 16681 20788
rect 16632 20748 16638 20760
rect 16669 20757 16681 20760
rect 16715 20757 16727 20791
rect 16669 20751 16727 20757
rect 17865 20791 17923 20797
rect 17865 20757 17877 20791
rect 17911 20788 17923 20791
rect 17954 20788 17960 20800
rect 17911 20760 17960 20788
rect 17911 20757 17923 20760
rect 17865 20751 17923 20757
rect 17954 20748 17960 20760
rect 18012 20748 18018 20800
rect 19978 20748 19984 20800
rect 20036 20788 20042 20800
rect 20073 20791 20131 20797
rect 20073 20788 20085 20791
rect 20036 20760 20085 20788
rect 20036 20748 20042 20760
rect 20073 20757 20085 20760
rect 20119 20757 20131 20791
rect 20073 20751 20131 20757
rect 21450 20748 21456 20800
rect 21508 20788 21514 20800
rect 22186 20788 22192 20800
rect 21508 20760 22192 20788
rect 21508 20748 21514 20760
rect 22186 20748 22192 20760
rect 22244 20748 22250 20800
rect 22572 20788 22600 20887
rect 24854 20884 24860 20936
rect 24912 20924 24918 20936
rect 25041 20927 25099 20933
rect 25041 20924 25053 20927
rect 24912 20896 25053 20924
rect 24912 20884 24918 20896
rect 25041 20893 25053 20896
rect 25087 20893 25099 20927
rect 25041 20887 25099 20893
rect 22738 20788 22744 20800
rect 22572 20760 22744 20788
rect 22738 20748 22744 20760
rect 22796 20748 22802 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 8113 20587 8171 20593
rect 8113 20553 8125 20587
rect 8159 20584 8171 20587
rect 8202 20584 8208 20596
rect 8159 20556 8208 20584
rect 8159 20553 8171 20556
rect 8113 20547 8171 20553
rect 8202 20544 8208 20556
rect 8260 20544 8266 20596
rect 12066 20584 12072 20596
rect 12027 20556 12072 20584
rect 12066 20544 12072 20556
rect 12124 20544 12130 20596
rect 17497 20587 17555 20593
rect 17497 20553 17509 20587
rect 17543 20584 17555 20587
rect 17862 20584 17868 20596
rect 17543 20556 17868 20584
rect 17543 20553 17555 20556
rect 17497 20547 17555 20553
rect 17862 20544 17868 20556
rect 17920 20544 17926 20596
rect 20257 20587 20315 20593
rect 20257 20553 20269 20587
rect 20303 20584 20315 20587
rect 20622 20584 20628 20596
rect 20303 20556 20628 20584
rect 20303 20553 20315 20556
rect 20257 20547 20315 20553
rect 20622 20544 20628 20556
rect 20680 20544 20686 20596
rect 15470 20516 15476 20528
rect 15431 20488 15476 20516
rect 15470 20476 15476 20488
rect 15528 20476 15534 20528
rect 25498 20516 25504 20528
rect 25459 20488 25504 20516
rect 25498 20476 25504 20488
rect 25556 20476 25562 20528
rect 8754 20448 8760 20460
rect 8715 20420 8760 20448
rect 8754 20408 8760 20420
rect 8812 20408 8818 20460
rect 20806 20408 20812 20460
rect 20864 20448 20870 20460
rect 20901 20451 20959 20457
rect 20901 20448 20913 20451
rect 20864 20420 20913 20448
rect 20864 20408 20870 20420
rect 20901 20417 20913 20420
rect 20947 20417 20959 20451
rect 20901 20411 20959 20417
rect 11698 20340 11704 20392
rect 11756 20380 11762 20392
rect 12805 20383 12863 20389
rect 12805 20380 12817 20383
rect 11756 20352 12817 20380
rect 11756 20340 11762 20352
rect 12805 20349 12817 20352
rect 12851 20380 12863 20383
rect 12897 20383 12955 20389
rect 12897 20380 12909 20383
rect 12851 20352 12909 20380
rect 12851 20349 12863 20352
rect 12805 20343 12863 20349
rect 12897 20349 12909 20352
rect 12943 20380 12955 20383
rect 12986 20380 12992 20392
rect 12943 20352 12992 20380
rect 12943 20349 12955 20352
rect 12897 20343 12955 20349
rect 12986 20340 12992 20352
rect 13044 20340 13050 20392
rect 15838 20380 15844 20392
rect 14844 20352 15844 20380
rect 7745 20315 7803 20321
rect 7745 20281 7757 20315
rect 7791 20312 7803 20315
rect 9024 20315 9082 20321
rect 9024 20312 9036 20315
rect 7791 20284 9036 20312
rect 7791 20281 7803 20284
rect 7745 20275 7803 20281
rect 9024 20281 9036 20284
rect 9070 20312 9082 20315
rect 9122 20312 9128 20324
rect 9070 20284 9128 20312
rect 9070 20281 9082 20284
rect 9024 20275 9082 20281
rect 9122 20272 9128 20284
rect 9180 20272 9186 20324
rect 13164 20315 13222 20321
rect 13164 20281 13176 20315
rect 13210 20312 13222 20315
rect 13538 20312 13544 20324
rect 13210 20284 13544 20312
rect 13210 20281 13222 20284
rect 13164 20275 13222 20281
rect 13538 20272 13544 20284
rect 13596 20272 13602 20324
rect 8478 20244 8484 20256
rect 8439 20216 8484 20244
rect 8478 20204 8484 20216
rect 8536 20204 8542 20256
rect 10134 20244 10140 20256
rect 10095 20216 10140 20244
rect 10134 20204 10140 20216
rect 10192 20204 10198 20256
rect 10686 20204 10692 20256
rect 10744 20244 10750 20256
rect 11698 20244 11704 20256
rect 10744 20216 11704 20244
rect 10744 20204 10750 20216
rect 11698 20204 11704 20216
rect 11756 20204 11762 20256
rect 14844 20253 14872 20352
rect 15838 20340 15844 20352
rect 15896 20380 15902 20392
rect 16025 20383 16083 20389
rect 16025 20380 16037 20383
rect 15896 20352 16037 20380
rect 15896 20340 15902 20352
rect 16025 20349 16037 20352
rect 16071 20349 16083 20383
rect 16025 20343 16083 20349
rect 17494 20340 17500 20392
rect 17552 20380 17558 20392
rect 17865 20383 17923 20389
rect 17865 20380 17877 20383
rect 17552 20352 17877 20380
rect 17552 20340 17558 20352
rect 17865 20349 17877 20352
rect 17911 20380 17923 20383
rect 18049 20383 18107 20389
rect 18049 20380 18061 20383
rect 17911 20352 18061 20380
rect 17911 20349 17923 20352
rect 17865 20343 17923 20349
rect 18049 20349 18061 20352
rect 18095 20380 18107 20383
rect 19518 20380 19524 20392
rect 18095 20352 19524 20380
rect 18095 20349 18107 20352
rect 18049 20343 18107 20349
rect 19518 20340 19524 20352
rect 19576 20380 19582 20392
rect 20625 20383 20683 20389
rect 20625 20380 20637 20383
rect 19576 20352 20637 20380
rect 19576 20340 19582 20352
rect 20625 20349 20637 20352
rect 20671 20380 20683 20383
rect 20990 20380 20996 20392
rect 20671 20352 20996 20380
rect 20671 20349 20683 20352
rect 20625 20343 20683 20349
rect 20990 20340 20996 20352
rect 21048 20380 21054 20392
rect 21085 20383 21143 20389
rect 21085 20380 21097 20383
rect 21048 20352 21097 20380
rect 21048 20340 21054 20352
rect 21085 20349 21097 20352
rect 21131 20380 21143 20383
rect 22738 20380 22744 20392
rect 21131 20352 22744 20380
rect 21131 20349 21143 20352
rect 21085 20343 21143 20349
rect 22738 20340 22744 20352
rect 22796 20380 22802 20392
rect 23017 20383 23075 20389
rect 23017 20380 23029 20383
rect 22796 20352 23029 20380
rect 22796 20340 22802 20352
rect 23017 20349 23029 20352
rect 23063 20380 23075 20383
rect 23934 20380 23940 20392
rect 23063 20352 23940 20380
rect 23063 20349 23075 20352
rect 23017 20343 23075 20349
rect 23934 20340 23940 20352
rect 23992 20380 23998 20392
rect 24121 20383 24179 20389
rect 24121 20380 24133 20383
rect 23992 20352 24133 20380
rect 23992 20340 23998 20352
rect 24121 20349 24133 20352
rect 24167 20349 24179 20383
rect 24121 20343 24179 20349
rect 15746 20312 15752 20324
rect 15707 20284 15752 20312
rect 15746 20272 15752 20284
rect 15804 20272 15810 20324
rect 15930 20312 15936 20324
rect 15891 20284 15936 20312
rect 15930 20272 15936 20284
rect 15988 20312 15994 20324
rect 18322 20321 18328 20324
rect 16393 20315 16451 20321
rect 16393 20312 16405 20315
rect 15988 20284 16405 20312
rect 15988 20272 15994 20284
rect 16393 20281 16405 20284
rect 16439 20281 16451 20315
rect 18316 20312 18328 20321
rect 18283 20284 18328 20312
rect 16393 20275 16451 20281
rect 18316 20275 18328 20284
rect 18322 20272 18328 20275
rect 18380 20272 18386 20324
rect 21174 20272 21180 20324
rect 21232 20312 21238 20324
rect 21330 20315 21388 20321
rect 21330 20312 21342 20315
rect 21232 20284 21342 20312
rect 21232 20272 21238 20284
rect 21330 20281 21342 20284
rect 21376 20281 21388 20315
rect 24366 20315 24424 20321
rect 24366 20312 24378 20315
rect 21330 20275 21388 20281
rect 24136 20284 24378 20312
rect 24136 20256 24164 20284
rect 24366 20281 24378 20284
rect 24412 20281 24424 20315
rect 24366 20275 24424 20281
rect 14277 20247 14335 20253
rect 14277 20213 14289 20247
rect 14323 20244 14335 20247
rect 14829 20247 14887 20253
rect 14829 20244 14841 20247
rect 14323 20216 14841 20244
rect 14323 20213 14335 20216
rect 14277 20207 14335 20213
rect 14829 20213 14841 20216
rect 14875 20213 14887 20247
rect 15286 20244 15292 20256
rect 15199 20216 15292 20244
rect 14829 20207 14887 20213
rect 15286 20204 15292 20216
rect 15344 20244 15350 20256
rect 16298 20244 16304 20256
rect 15344 20216 16304 20244
rect 15344 20204 15350 20216
rect 16298 20204 16304 20216
rect 16356 20204 16362 20256
rect 16942 20244 16948 20256
rect 16903 20216 16948 20244
rect 16942 20204 16948 20216
rect 17000 20204 17006 20256
rect 19426 20244 19432 20256
rect 19387 20216 19432 20244
rect 19426 20204 19432 20216
rect 19484 20204 19490 20256
rect 22462 20244 22468 20256
rect 22423 20216 22468 20244
rect 22462 20204 22468 20216
rect 22520 20204 22526 20256
rect 23382 20244 23388 20256
rect 23343 20216 23388 20244
rect 23382 20204 23388 20216
rect 23440 20204 23446 20256
rect 24118 20204 24124 20256
rect 24176 20204 24182 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 8754 20040 8760 20052
rect 8715 20012 8760 20040
rect 8754 20000 8760 20012
rect 8812 20000 8818 20052
rect 11885 20043 11943 20049
rect 11885 20009 11897 20043
rect 11931 20040 11943 20043
rect 12066 20040 12072 20052
rect 11931 20012 12072 20040
rect 11931 20009 11943 20012
rect 11885 20003 11943 20009
rect 12066 20000 12072 20012
rect 12124 20000 12130 20052
rect 13354 20000 13360 20052
rect 13412 20040 13418 20052
rect 13541 20043 13599 20049
rect 13541 20040 13553 20043
rect 13412 20012 13553 20040
rect 13412 20000 13418 20012
rect 13541 20009 13553 20012
rect 13587 20040 13599 20043
rect 13722 20040 13728 20052
rect 13587 20012 13728 20040
rect 13587 20009 13599 20012
rect 13541 20003 13599 20009
rect 13722 20000 13728 20012
rect 13780 20000 13786 20052
rect 15838 20040 15844 20052
rect 15799 20012 15844 20040
rect 15838 20000 15844 20012
rect 15896 20000 15902 20052
rect 19334 20040 19340 20052
rect 19295 20012 19340 20040
rect 19334 20000 19340 20012
rect 19392 20000 19398 20052
rect 21358 20000 21364 20052
rect 21416 20040 21422 20052
rect 21729 20043 21787 20049
rect 21729 20040 21741 20043
rect 21416 20012 21741 20040
rect 21416 20000 21422 20012
rect 21729 20009 21741 20012
rect 21775 20009 21787 20043
rect 21729 20003 21787 20009
rect 22094 20000 22100 20052
rect 22152 20040 22158 20052
rect 22189 20043 22247 20049
rect 22189 20040 22201 20043
rect 22152 20012 22201 20040
rect 22152 20000 22158 20012
rect 22189 20009 22201 20012
rect 22235 20009 22247 20043
rect 22189 20003 22247 20009
rect 22738 20000 22744 20052
rect 22796 20040 22802 20052
rect 23474 20040 23480 20052
rect 22796 20012 23480 20040
rect 22796 20000 22802 20012
rect 23474 20000 23480 20012
rect 23532 20000 23538 20052
rect 15746 19932 15752 19984
rect 15804 19972 15810 19984
rect 16117 19975 16175 19981
rect 16117 19972 16129 19975
rect 15804 19944 16129 19972
rect 15804 19932 15810 19944
rect 16117 19941 16129 19944
rect 16163 19941 16175 19975
rect 16117 19935 16175 19941
rect 16942 19932 16948 19984
rect 17000 19972 17006 19984
rect 19153 19975 19211 19981
rect 19153 19972 19165 19975
rect 17000 19944 19165 19972
rect 17000 19932 17006 19944
rect 19153 19941 19165 19944
rect 19199 19972 19211 19975
rect 19242 19972 19248 19984
rect 19199 19944 19248 19972
rect 19199 19941 19211 19944
rect 19153 19935 19211 19941
rect 19242 19932 19248 19944
rect 19300 19932 19306 19984
rect 20530 19932 20536 19984
rect 20588 19972 20594 19984
rect 21545 19975 21603 19981
rect 21545 19972 21557 19975
rect 20588 19944 21557 19972
rect 20588 19932 20594 19944
rect 21545 19941 21557 19944
rect 21591 19941 21603 19975
rect 22554 19972 22560 19984
rect 21545 19935 21603 19941
rect 21836 19944 22560 19972
rect 8754 19864 8760 19916
rect 8812 19904 8818 19916
rect 10505 19907 10563 19913
rect 10505 19904 10517 19907
rect 8812 19876 10517 19904
rect 8812 19864 8818 19876
rect 10505 19873 10517 19876
rect 10551 19904 10563 19907
rect 10594 19904 10600 19916
rect 10551 19876 10600 19904
rect 10551 19873 10563 19876
rect 10505 19867 10563 19873
rect 10594 19864 10600 19876
rect 10652 19864 10658 19916
rect 10778 19913 10784 19916
rect 10772 19904 10784 19913
rect 10739 19876 10784 19904
rect 10772 19867 10784 19876
rect 10778 19864 10784 19867
rect 10836 19864 10842 19916
rect 12342 19864 12348 19916
rect 12400 19904 12406 19916
rect 13357 19907 13415 19913
rect 13357 19904 13369 19907
rect 12400 19876 13369 19904
rect 12400 19864 12406 19876
rect 13357 19873 13369 19876
rect 13403 19904 13415 19907
rect 13722 19904 13728 19916
rect 13403 19876 13728 19904
rect 13403 19873 13415 19876
rect 13357 19867 13415 19873
rect 13722 19864 13728 19876
rect 13780 19864 13786 19916
rect 16574 19913 16580 19916
rect 16568 19904 16580 19913
rect 16535 19876 16580 19904
rect 16568 19867 16580 19876
rect 16574 19864 16580 19867
rect 16632 19864 16638 19916
rect 21174 19864 21180 19916
rect 21232 19904 21238 19916
rect 21836 19913 21864 19944
rect 22554 19932 22560 19944
rect 22612 19932 22618 19984
rect 22922 19932 22928 19984
rect 22980 19972 22986 19984
rect 23293 19975 23351 19981
rect 23293 19972 23305 19975
rect 22980 19944 23305 19972
rect 22980 19932 22986 19944
rect 23293 19941 23305 19944
rect 23339 19941 23351 19975
rect 24854 19972 24860 19984
rect 24815 19944 24860 19972
rect 23293 19935 23351 19941
rect 24854 19932 24860 19944
rect 24912 19932 24918 19984
rect 21821 19907 21879 19913
rect 21821 19904 21833 19907
rect 21232 19876 21833 19904
rect 21232 19864 21238 19876
rect 21821 19873 21833 19876
rect 21867 19873 21879 19907
rect 21821 19867 21879 19873
rect 22462 19864 22468 19916
rect 22520 19904 22526 19916
rect 23382 19904 23388 19916
rect 22520 19876 23388 19904
rect 22520 19864 22526 19876
rect 23382 19864 23388 19876
rect 23440 19864 23446 19916
rect 24118 19864 24124 19916
rect 24176 19904 24182 19916
rect 24949 19907 25007 19913
rect 24949 19904 24961 19907
rect 24176 19876 24961 19904
rect 24176 19864 24182 19876
rect 24949 19873 24961 19876
rect 24995 19873 25007 19907
rect 24949 19867 25007 19873
rect 13538 19796 13544 19848
rect 13596 19836 13602 19848
rect 13633 19839 13691 19845
rect 13633 19836 13645 19839
rect 13596 19808 13645 19836
rect 13596 19796 13602 19808
rect 13633 19805 13645 19808
rect 13679 19805 13691 19839
rect 13633 19799 13691 19805
rect 15289 19839 15347 19845
rect 15289 19805 15301 19839
rect 15335 19836 15347 19839
rect 15654 19836 15660 19848
rect 15335 19808 15660 19836
rect 15335 19805 15347 19808
rect 15289 19799 15347 19805
rect 15654 19796 15660 19808
rect 15712 19796 15718 19848
rect 16298 19836 16304 19848
rect 16259 19808 16304 19836
rect 16298 19796 16304 19808
rect 16356 19796 16362 19848
rect 18322 19836 18328 19848
rect 18235 19808 18328 19836
rect 18322 19796 18328 19808
rect 18380 19836 18386 19848
rect 18693 19839 18751 19845
rect 18693 19836 18705 19839
rect 18380 19808 18705 19836
rect 18380 19796 18386 19808
rect 18693 19805 18705 19808
rect 18739 19836 18751 19839
rect 19058 19836 19064 19848
rect 18739 19808 19064 19836
rect 18739 19805 18751 19808
rect 18693 19799 18751 19805
rect 19058 19796 19064 19808
rect 19116 19836 19122 19848
rect 19429 19839 19487 19845
rect 19429 19836 19441 19839
rect 19116 19808 19441 19836
rect 19116 19796 19122 19808
rect 19429 19805 19441 19808
rect 19475 19805 19487 19839
rect 23290 19836 23296 19848
rect 23251 19808 23296 19836
rect 19429 19799 19487 19805
rect 23290 19796 23296 19808
rect 23348 19796 23354 19848
rect 24762 19836 24768 19848
rect 24723 19808 24768 19836
rect 24762 19796 24768 19808
rect 24820 19796 24826 19848
rect 13078 19768 13084 19780
rect 13039 19740 13084 19768
rect 13078 19728 13084 19740
rect 13136 19728 13142 19780
rect 17681 19771 17739 19777
rect 17681 19737 17693 19771
rect 17727 19768 17739 19771
rect 18340 19768 18368 19796
rect 18874 19768 18880 19780
rect 17727 19740 18368 19768
rect 18787 19740 18880 19768
rect 17727 19737 17739 19740
rect 17681 19731 17739 19737
rect 18874 19728 18880 19740
rect 18932 19768 18938 19780
rect 20165 19771 20223 19777
rect 20165 19768 20177 19771
rect 18932 19740 20177 19768
rect 18932 19728 18938 19740
rect 20165 19737 20177 19740
rect 20211 19737 20223 19771
rect 20165 19731 20223 19737
rect 21269 19771 21327 19777
rect 21269 19737 21281 19771
rect 21315 19768 21327 19771
rect 22922 19768 22928 19780
rect 21315 19740 22928 19768
rect 21315 19737 21327 19740
rect 21269 19731 21327 19737
rect 22922 19728 22928 19740
rect 22980 19728 22986 19780
rect 24397 19771 24455 19777
rect 24397 19737 24409 19771
rect 24443 19768 24455 19771
rect 24670 19768 24676 19780
rect 24443 19740 24676 19768
rect 24443 19737 24455 19740
rect 24397 19731 24455 19737
rect 24670 19728 24676 19740
rect 24728 19728 24734 19780
rect 8113 19703 8171 19709
rect 8113 19669 8125 19703
rect 8159 19700 8171 19703
rect 8202 19700 8208 19712
rect 8159 19672 8208 19700
rect 8159 19669 8171 19672
rect 8113 19663 8171 19669
rect 8202 19660 8208 19672
rect 8260 19660 8266 19712
rect 12526 19700 12532 19712
rect 12487 19672 12532 19700
rect 12526 19660 12532 19672
rect 12584 19660 12590 19712
rect 14090 19700 14096 19712
rect 14051 19672 14096 19700
rect 14090 19660 14096 19672
rect 14148 19660 14154 19712
rect 19794 19700 19800 19712
rect 19755 19672 19800 19700
rect 19794 19660 19800 19672
rect 19852 19660 19858 19712
rect 20717 19703 20775 19709
rect 20717 19669 20729 19703
rect 20763 19700 20775 19703
rect 21174 19700 21180 19712
rect 20763 19672 21180 19700
rect 20763 19669 20775 19672
rect 20717 19663 20775 19669
rect 21174 19660 21180 19672
rect 21232 19660 21238 19712
rect 22370 19660 22376 19712
rect 22428 19700 22434 19712
rect 22833 19703 22891 19709
rect 22833 19700 22845 19703
rect 22428 19672 22845 19700
rect 22428 19660 22434 19672
rect 22833 19669 22845 19672
rect 22879 19669 22891 19703
rect 23842 19700 23848 19712
rect 23803 19672 23848 19700
rect 22833 19663 22891 19669
rect 23842 19660 23848 19672
rect 23900 19660 23906 19712
rect 24118 19700 24124 19712
rect 24079 19672 24124 19700
rect 24118 19660 24124 19672
rect 24176 19660 24182 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 8754 19456 8760 19508
rect 8812 19496 8818 19508
rect 9401 19499 9459 19505
rect 9401 19496 9413 19499
rect 8812 19468 9413 19496
rect 8812 19456 8818 19468
rect 9401 19465 9413 19468
rect 9447 19465 9459 19499
rect 9401 19459 9459 19465
rect 9416 19360 9444 19459
rect 12802 19456 12808 19508
rect 12860 19496 12866 19508
rect 13265 19499 13323 19505
rect 13265 19496 13277 19499
rect 12860 19468 13277 19496
rect 12860 19456 12866 19468
rect 13265 19465 13277 19468
rect 13311 19496 13323 19499
rect 13354 19496 13360 19508
rect 13311 19468 13360 19496
rect 13311 19465 13323 19468
rect 13265 19459 13323 19465
rect 13354 19456 13360 19468
rect 13412 19456 13418 19508
rect 19153 19499 19211 19505
rect 19153 19465 19165 19499
rect 19199 19496 19211 19499
rect 19334 19496 19340 19508
rect 19199 19468 19340 19496
rect 19199 19465 19211 19468
rect 19153 19459 19211 19465
rect 19334 19456 19340 19468
rect 19392 19496 19398 19508
rect 20254 19496 20260 19508
rect 19392 19468 20260 19496
rect 19392 19456 19398 19468
rect 20254 19456 20260 19468
rect 20312 19456 20318 19508
rect 21450 19496 21456 19508
rect 21411 19468 21456 19496
rect 21450 19456 21456 19468
rect 21508 19456 21514 19508
rect 22833 19499 22891 19505
rect 22833 19465 22845 19499
rect 22879 19496 22891 19499
rect 23290 19496 23296 19508
rect 22879 19468 23296 19496
rect 22879 19465 22891 19468
rect 22833 19459 22891 19465
rect 23290 19456 23296 19468
rect 23348 19456 23354 19508
rect 23477 19499 23535 19505
rect 23477 19465 23489 19499
rect 23523 19496 23535 19499
rect 24118 19496 24124 19508
rect 23523 19468 24124 19496
rect 23523 19465 23535 19468
rect 23477 19459 23535 19465
rect 24118 19456 24124 19468
rect 24176 19496 24182 19508
rect 25501 19499 25559 19505
rect 25501 19496 25513 19499
rect 24176 19468 25513 19496
rect 24176 19456 24182 19468
rect 25501 19465 25513 19468
rect 25547 19465 25559 19499
rect 25501 19459 25559 19465
rect 13170 19388 13176 19440
rect 13228 19428 13234 19440
rect 23934 19428 23940 19440
rect 13228 19400 13308 19428
rect 23895 19400 23940 19428
rect 13228 19388 13234 19400
rect 13280 19372 13308 19400
rect 23934 19388 23940 19400
rect 23992 19428 23998 19440
rect 23992 19400 24164 19428
rect 23992 19388 23998 19400
rect 9585 19363 9643 19369
rect 9585 19360 9597 19363
rect 9416 19332 9597 19360
rect 9585 19329 9597 19332
rect 9631 19329 9643 19363
rect 9585 19323 9643 19329
rect 13262 19320 13268 19372
rect 13320 19320 13326 19372
rect 18601 19363 18659 19369
rect 18601 19329 18613 19363
rect 18647 19360 18659 19363
rect 18874 19360 18880 19372
rect 18647 19332 18880 19360
rect 18647 19329 18659 19332
rect 18601 19323 18659 19329
rect 18874 19320 18880 19332
rect 18932 19320 18938 19372
rect 19794 19360 19800 19372
rect 19260 19332 19800 19360
rect 7929 19295 7987 19301
rect 7929 19261 7941 19295
rect 7975 19292 7987 19295
rect 8665 19295 8723 19301
rect 8665 19292 8677 19295
rect 7975 19264 8677 19292
rect 7975 19261 7987 19264
rect 7929 19255 7987 19261
rect 8665 19261 8677 19264
rect 8711 19261 8723 19295
rect 8665 19255 8723 19261
rect 8386 19224 8392 19236
rect 8347 19196 8392 19224
rect 8386 19184 8392 19196
rect 8444 19184 8450 19236
rect 8680 19224 8708 19255
rect 9674 19252 9680 19304
rect 9732 19292 9738 19304
rect 9852 19295 9910 19301
rect 9852 19292 9864 19295
rect 9732 19264 9864 19292
rect 9732 19252 9738 19264
rect 9852 19261 9864 19264
rect 9898 19292 9910 19295
rect 10134 19292 10140 19304
rect 9898 19264 10140 19292
rect 9898 19261 9910 19264
rect 9852 19255 9910 19261
rect 10134 19252 10140 19264
rect 10192 19252 10198 19304
rect 12253 19295 12311 19301
rect 12253 19261 12265 19295
rect 12299 19292 12311 19295
rect 12342 19292 12348 19304
rect 12299 19264 12348 19292
rect 12299 19261 12311 19264
rect 12253 19255 12311 19261
rect 12342 19252 12348 19264
rect 12400 19252 12406 19304
rect 12437 19295 12495 19301
rect 12437 19261 12449 19295
rect 12483 19292 12495 19295
rect 12526 19292 12532 19304
rect 12483 19264 12532 19292
rect 12483 19261 12495 19264
rect 12437 19255 12495 19261
rect 12526 19252 12532 19264
rect 12584 19252 12590 19304
rect 12710 19292 12716 19304
rect 12671 19264 12716 19292
rect 12710 19252 12716 19264
rect 12768 19252 12774 19304
rect 14090 19301 14096 19304
rect 13817 19295 13875 19301
rect 13817 19292 13829 19295
rect 13648 19264 13829 19292
rect 13648 19224 13676 19264
rect 13817 19261 13829 19264
rect 13863 19261 13875 19295
rect 14084 19292 14096 19301
rect 14003 19264 14096 19292
rect 13817 19255 13875 19261
rect 14084 19255 14096 19264
rect 14148 19292 14154 19304
rect 14148 19264 16988 19292
rect 14090 19252 14096 19255
rect 14148 19252 14154 19264
rect 15286 19224 15292 19236
rect 8680 19196 9812 19224
rect 8110 19165 8116 19168
rect 8103 19159 8116 19165
rect 8103 19125 8115 19159
rect 8168 19156 8174 19168
rect 8570 19156 8576 19168
rect 8168 19128 8203 19156
rect 8531 19128 8576 19156
rect 8103 19119 8116 19125
rect 8110 19116 8116 19119
rect 8168 19116 8174 19128
rect 8570 19116 8576 19128
rect 8628 19116 8634 19168
rect 9125 19159 9183 19165
rect 9125 19125 9137 19159
rect 9171 19156 9183 19159
rect 9674 19156 9680 19168
rect 9171 19128 9680 19156
rect 9171 19125 9183 19128
rect 9125 19119 9183 19125
rect 9674 19116 9680 19128
rect 9732 19116 9738 19168
rect 9784 19156 9812 19196
rect 13648 19196 15292 19224
rect 10778 19156 10784 19168
rect 9784 19128 10784 19156
rect 10778 19116 10784 19128
rect 10836 19156 10842 19168
rect 10965 19159 11023 19165
rect 10965 19156 10977 19159
rect 10836 19128 10977 19156
rect 10836 19116 10842 19128
rect 10965 19125 10977 19128
rect 11011 19156 11023 19159
rect 11517 19159 11575 19165
rect 11517 19156 11529 19159
rect 11011 19128 11529 19156
rect 11011 19125 11023 19128
rect 10965 19119 11023 19125
rect 11517 19125 11529 19128
rect 11563 19125 11575 19159
rect 11517 19119 11575 19125
rect 12986 19116 12992 19168
rect 13044 19156 13050 19168
rect 13354 19156 13360 19168
rect 13044 19128 13360 19156
rect 13044 19116 13050 19128
rect 13354 19116 13360 19128
rect 13412 19156 13418 19168
rect 13648 19165 13676 19196
rect 15286 19184 15292 19196
rect 15344 19184 15350 19236
rect 15746 19224 15752 19236
rect 15707 19196 15752 19224
rect 15746 19184 15752 19196
rect 15804 19224 15810 19236
rect 15804 19196 16620 19224
rect 15804 19184 15810 19196
rect 13633 19159 13691 19165
rect 13633 19156 13645 19159
rect 13412 19128 13645 19156
rect 13412 19116 13418 19128
rect 13633 19125 13645 19128
rect 13679 19125 13691 19159
rect 13633 19119 13691 19125
rect 14274 19116 14280 19168
rect 14332 19156 14338 19168
rect 15197 19159 15255 19165
rect 15197 19156 15209 19159
rect 14332 19128 15209 19156
rect 14332 19116 14338 19128
rect 15197 19125 15209 19128
rect 15243 19125 15255 19159
rect 15197 19119 15255 19125
rect 15838 19116 15844 19168
rect 15896 19156 15902 19168
rect 16117 19159 16175 19165
rect 16117 19156 16129 19159
rect 15896 19128 16129 19156
rect 15896 19116 15902 19128
rect 16117 19125 16129 19128
rect 16163 19125 16175 19159
rect 16117 19119 16175 19125
rect 16206 19116 16212 19168
rect 16264 19156 16270 19168
rect 16375 19159 16433 19165
rect 16375 19156 16387 19159
rect 16264 19128 16387 19156
rect 16264 19116 16270 19128
rect 16375 19125 16387 19128
rect 16421 19125 16433 19159
rect 16592 19156 16620 19196
rect 16666 19184 16672 19236
rect 16724 19224 16730 19236
rect 16960 19233 16988 19264
rect 17954 19252 17960 19304
rect 18012 19292 18018 19304
rect 19260 19292 19288 19332
rect 19794 19320 19800 19332
rect 19852 19320 19858 19372
rect 20530 19320 20536 19372
rect 20588 19360 20594 19372
rect 20990 19360 20996 19372
rect 20588 19332 20996 19360
rect 20588 19320 20594 19332
rect 20990 19320 20996 19332
rect 21048 19360 21054 19372
rect 24136 19369 24164 19400
rect 21177 19363 21235 19369
rect 21177 19360 21189 19363
rect 21048 19332 21189 19360
rect 21048 19320 21054 19332
rect 21177 19329 21189 19332
rect 21223 19329 21235 19363
rect 21177 19323 21235 19329
rect 24121 19363 24179 19369
rect 24121 19329 24133 19363
rect 24167 19329 24179 19363
rect 24121 19323 24179 19329
rect 18012 19264 19288 19292
rect 18012 19252 18018 19264
rect 18616 19233 18644 19264
rect 19334 19252 19340 19304
rect 19392 19292 19398 19304
rect 19429 19295 19487 19301
rect 19429 19292 19441 19295
rect 19392 19264 19441 19292
rect 19392 19252 19398 19264
rect 19429 19261 19441 19264
rect 19475 19261 19487 19295
rect 19429 19255 19487 19261
rect 19687 19295 19745 19301
rect 19687 19261 19699 19295
rect 19733 19292 19745 19295
rect 20162 19292 20168 19304
rect 19733 19264 20168 19292
rect 19733 19261 19745 19264
rect 19687 19255 19745 19261
rect 20162 19252 20168 19264
rect 20220 19252 20226 19304
rect 21726 19292 21732 19304
rect 21687 19264 21732 19292
rect 21726 19252 21732 19264
rect 21784 19252 21790 19304
rect 16945 19227 17003 19233
rect 16724 19196 16769 19224
rect 16724 19184 16730 19196
rect 16945 19193 16957 19227
rect 16991 19224 17003 19227
rect 17313 19227 17371 19233
rect 17313 19224 17325 19227
rect 16991 19196 17325 19224
rect 16991 19193 17003 19196
rect 16945 19187 17003 19193
rect 17313 19193 17325 19196
rect 17359 19193 17371 19227
rect 17313 19187 17371 19193
rect 17865 19227 17923 19233
rect 17865 19193 17877 19227
rect 17911 19224 17923 19227
rect 18601 19227 18659 19233
rect 17911 19196 18552 19224
rect 17911 19193 17923 19196
rect 17865 19187 17923 19193
rect 16853 19159 16911 19165
rect 16853 19156 16865 19159
rect 16592 19128 16865 19156
rect 16375 19119 16433 19125
rect 16853 19125 16865 19128
rect 16899 19156 16911 19159
rect 17770 19156 17776 19168
rect 16899 19128 17776 19156
rect 16899 19125 16911 19128
rect 16853 19119 16911 19125
rect 17770 19116 17776 19128
rect 17828 19116 17834 19168
rect 17954 19116 17960 19168
rect 18012 19156 18018 19168
rect 18123 19159 18181 19165
rect 18123 19156 18135 19159
rect 18012 19128 18135 19156
rect 18012 19116 18018 19128
rect 18123 19125 18135 19128
rect 18169 19125 18181 19159
rect 18524 19156 18552 19196
rect 18601 19193 18613 19227
rect 18647 19193 18659 19227
rect 18601 19187 18659 19193
rect 18693 19227 18751 19233
rect 18693 19193 18705 19227
rect 18739 19224 18751 19227
rect 18874 19224 18880 19236
rect 18739 19196 18880 19224
rect 18739 19193 18751 19196
rect 18693 19187 18751 19193
rect 18708 19156 18736 19187
rect 18874 19184 18880 19196
rect 18932 19184 18938 19236
rect 19978 19224 19984 19236
rect 19939 19196 19984 19224
rect 19978 19184 19984 19196
rect 20036 19184 20042 19236
rect 20257 19227 20315 19233
rect 20257 19193 20269 19227
rect 20303 19224 20315 19227
rect 20346 19224 20352 19236
rect 20303 19196 20352 19224
rect 20303 19193 20315 19196
rect 20257 19187 20315 19193
rect 20346 19184 20352 19196
rect 20404 19184 20410 19236
rect 22002 19224 22008 19236
rect 21963 19196 22008 19224
rect 22002 19184 22008 19196
rect 22060 19224 22066 19236
rect 22373 19227 22431 19233
rect 22373 19224 22385 19227
rect 22060 19196 22385 19224
rect 22060 19184 22066 19196
rect 22373 19193 22385 19196
rect 22419 19224 22431 19227
rect 22462 19224 22468 19236
rect 22419 19196 22468 19224
rect 22419 19193 22431 19196
rect 22373 19187 22431 19193
rect 22462 19184 22468 19196
rect 22520 19184 22526 19236
rect 23842 19184 23848 19236
rect 23900 19224 23906 19236
rect 24366 19227 24424 19233
rect 24366 19224 24378 19227
rect 23900 19196 24378 19224
rect 23900 19184 23906 19196
rect 24366 19193 24378 19196
rect 24412 19224 24424 19227
rect 24486 19224 24492 19236
rect 24412 19196 24492 19224
rect 24412 19193 24424 19196
rect 24366 19187 24424 19193
rect 24486 19184 24492 19196
rect 24544 19184 24550 19236
rect 24854 19184 24860 19236
rect 24912 19224 24918 19236
rect 26053 19227 26111 19233
rect 26053 19224 26065 19227
rect 24912 19196 26065 19224
rect 24912 19184 24918 19196
rect 26053 19193 26065 19196
rect 26099 19193 26111 19227
rect 26053 19187 26111 19193
rect 19426 19156 19432 19168
rect 18524 19128 19432 19156
rect 18123 19119 18181 19125
rect 19426 19116 19432 19128
rect 19484 19116 19490 19168
rect 20162 19156 20168 19168
rect 20123 19128 20168 19156
rect 20162 19116 20168 19128
rect 20220 19116 20226 19168
rect 20901 19159 20959 19165
rect 20901 19125 20913 19159
rect 20947 19156 20959 19159
rect 21358 19156 21364 19168
rect 20947 19128 21364 19156
rect 20947 19125 20959 19128
rect 20901 19119 20959 19125
rect 21358 19116 21364 19128
rect 21416 19116 21422 19168
rect 21910 19156 21916 19168
rect 21871 19128 21916 19156
rect 21910 19116 21916 19128
rect 21968 19116 21974 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 8294 18912 8300 18964
rect 8352 18952 8358 18964
rect 9401 18955 9459 18961
rect 9401 18952 9413 18955
rect 8352 18924 9413 18952
rect 8352 18912 8358 18924
rect 9401 18921 9413 18924
rect 9447 18952 9459 18955
rect 10229 18955 10287 18961
rect 10229 18952 10241 18955
rect 9447 18924 10241 18952
rect 9447 18921 9459 18924
rect 9401 18915 9459 18921
rect 10229 18921 10241 18924
rect 10275 18921 10287 18955
rect 10686 18952 10692 18964
rect 10647 18924 10692 18952
rect 10229 18915 10287 18921
rect 10686 18912 10692 18924
rect 10744 18912 10750 18964
rect 13538 18952 13544 18964
rect 13499 18924 13544 18952
rect 13538 18912 13544 18924
rect 13596 18912 13602 18964
rect 14185 18955 14243 18961
rect 14185 18921 14197 18955
rect 14231 18952 14243 18955
rect 14458 18952 14464 18964
rect 14231 18924 14464 18952
rect 14231 18921 14243 18924
rect 14185 18915 14243 18921
rect 14458 18912 14464 18924
rect 14516 18952 14522 18964
rect 16206 18952 16212 18964
rect 14516 18924 16212 18952
rect 14516 18912 14522 18924
rect 16206 18912 16212 18924
rect 16264 18912 16270 18964
rect 16574 18912 16580 18964
rect 16632 18952 16638 18964
rect 16669 18955 16727 18961
rect 16669 18952 16681 18955
rect 16632 18924 16681 18952
rect 16632 18912 16638 18924
rect 16669 18921 16681 18924
rect 16715 18921 16727 18955
rect 19058 18952 19064 18964
rect 19019 18924 19064 18952
rect 16669 18915 16727 18921
rect 19058 18912 19064 18924
rect 19116 18912 19122 18964
rect 21174 18952 21180 18964
rect 21135 18924 21180 18952
rect 21174 18912 21180 18924
rect 21232 18912 21238 18964
rect 21637 18955 21695 18961
rect 21637 18921 21649 18955
rect 21683 18952 21695 18955
rect 22002 18952 22008 18964
rect 21683 18924 22008 18952
rect 21683 18921 21695 18924
rect 21637 18915 21695 18921
rect 22002 18912 22008 18924
rect 22060 18912 22066 18964
rect 22922 18952 22928 18964
rect 22883 18924 22928 18952
rect 22922 18912 22928 18924
rect 22980 18912 22986 18964
rect 23474 18912 23480 18964
rect 23532 18952 23538 18964
rect 24397 18955 24455 18961
rect 24397 18952 24409 18955
rect 23532 18924 24409 18952
rect 23532 18912 23538 18924
rect 24397 18921 24409 18924
rect 24443 18921 24455 18955
rect 24397 18915 24455 18921
rect 10134 18844 10140 18896
rect 10192 18884 10198 18896
rect 10321 18887 10379 18893
rect 10321 18884 10333 18887
rect 10192 18856 10333 18884
rect 10192 18844 10198 18856
rect 10321 18853 10333 18856
rect 10367 18853 10379 18887
rect 10321 18847 10379 18853
rect 12158 18844 12164 18896
rect 12216 18884 12222 18896
rect 12621 18887 12679 18893
rect 12621 18884 12633 18887
rect 12216 18856 12633 18884
rect 12216 18844 12222 18856
rect 12621 18853 12633 18856
rect 12667 18853 12679 18887
rect 12621 18847 12679 18853
rect 12713 18887 12771 18893
rect 12713 18853 12725 18887
rect 12759 18884 12771 18887
rect 14090 18884 14096 18896
rect 12759 18856 14096 18884
rect 12759 18853 12771 18856
rect 12713 18847 12771 18853
rect 12728 18816 12756 18847
rect 14090 18844 14096 18856
rect 14148 18844 14154 18896
rect 15841 18887 15899 18893
rect 15841 18884 15853 18887
rect 15028 18856 15853 18884
rect 11900 18788 12756 18816
rect 10229 18751 10287 18757
rect 10229 18717 10241 18751
rect 10275 18748 10287 18751
rect 10594 18748 10600 18760
rect 10275 18720 10600 18748
rect 10275 18717 10287 18720
rect 10229 18711 10287 18717
rect 10594 18708 10600 18720
rect 10652 18708 10658 18760
rect 8113 18683 8171 18689
rect 8113 18649 8125 18683
rect 8159 18680 8171 18683
rect 8570 18680 8576 18692
rect 8159 18652 8576 18680
rect 8159 18649 8171 18652
rect 8113 18643 8171 18649
rect 8570 18640 8576 18652
rect 8628 18680 8634 18692
rect 9769 18683 9827 18689
rect 9769 18680 9781 18683
rect 8628 18652 9781 18680
rect 8628 18640 8634 18652
rect 9769 18649 9781 18652
rect 9815 18649 9827 18683
rect 9769 18643 9827 18649
rect 10778 18572 10784 18624
rect 10836 18612 10842 18624
rect 11900 18621 11928 18788
rect 12618 18748 12624 18760
rect 12579 18720 12624 18748
rect 12618 18708 12624 18720
rect 12676 18708 12682 18760
rect 14093 18751 14151 18757
rect 14093 18717 14105 18751
rect 14139 18717 14151 18751
rect 14274 18748 14280 18760
rect 14235 18720 14280 18748
rect 14093 18711 14151 18717
rect 12161 18683 12219 18689
rect 12161 18649 12173 18683
rect 12207 18680 12219 18683
rect 14108 18680 14136 18711
rect 14274 18708 14280 18720
rect 14332 18708 14338 18760
rect 14645 18683 14703 18689
rect 14645 18680 14657 18683
rect 12207 18652 14657 18680
rect 12207 18649 12219 18652
rect 12161 18643 12219 18649
rect 14645 18649 14657 18652
rect 14691 18649 14703 18683
rect 14645 18643 14703 18649
rect 11885 18615 11943 18621
rect 11885 18612 11897 18615
rect 10836 18584 11897 18612
rect 10836 18572 10842 18584
rect 11885 18581 11897 18584
rect 11931 18581 11943 18615
rect 11885 18575 11943 18581
rect 12434 18572 12440 18624
rect 12492 18612 12498 18624
rect 13081 18615 13139 18621
rect 13081 18612 13093 18615
rect 12492 18584 13093 18612
rect 12492 18572 12498 18584
rect 13081 18581 13093 18584
rect 13127 18612 13139 18615
rect 13354 18612 13360 18624
rect 13127 18584 13360 18612
rect 13127 18581 13139 18584
rect 13081 18575 13139 18581
rect 13354 18572 13360 18584
rect 13412 18572 13418 18624
rect 13722 18612 13728 18624
rect 13683 18584 13728 18612
rect 13722 18572 13728 18584
rect 13780 18572 13786 18624
rect 14826 18572 14832 18624
rect 14884 18612 14890 18624
rect 15028 18621 15056 18856
rect 15841 18853 15853 18856
rect 15887 18853 15899 18887
rect 15841 18847 15899 18853
rect 20717 18887 20775 18893
rect 20717 18853 20729 18887
rect 20763 18884 20775 18887
rect 21726 18884 21732 18896
rect 20763 18856 21732 18884
rect 20763 18853 20775 18856
rect 20717 18847 20775 18853
rect 21726 18844 21732 18856
rect 21784 18844 21790 18896
rect 22370 18884 22376 18896
rect 22331 18856 22376 18884
rect 22370 18844 22376 18856
rect 22428 18844 22434 18896
rect 24486 18884 24492 18896
rect 24447 18856 24492 18884
rect 24486 18844 24492 18856
rect 24544 18884 24550 18896
rect 24857 18887 24915 18893
rect 24857 18884 24869 18887
rect 24544 18856 24869 18884
rect 24544 18844 24550 18856
rect 24857 18853 24869 18856
rect 24903 18884 24915 18887
rect 24946 18884 24952 18896
rect 24903 18856 24952 18884
rect 24903 18853 24915 18856
rect 24857 18847 24915 18853
rect 24946 18844 24952 18856
rect 25004 18844 25010 18896
rect 15654 18816 15660 18828
rect 15615 18788 15660 18816
rect 15654 18776 15660 18788
rect 15712 18776 15718 18828
rect 16758 18776 16764 18828
rect 16816 18816 16822 18828
rect 17385 18819 17443 18825
rect 17385 18816 17397 18819
rect 16816 18788 17397 18816
rect 16816 18776 16822 18788
rect 17385 18785 17397 18788
rect 17431 18785 17443 18819
rect 22186 18816 22192 18828
rect 22147 18788 22192 18816
rect 17385 18779 17443 18785
rect 22186 18776 22192 18788
rect 22244 18816 22250 18828
rect 23201 18819 23259 18825
rect 23201 18816 23213 18819
rect 22244 18788 23213 18816
rect 22244 18776 22250 18788
rect 23201 18785 23213 18788
rect 23247 18785 23259 18819
rect 24210 18816 24216 18828
rect 24171 18788 24216 18816
rect 23201 18779 23259 18785
rect 24210 18776 24216 18788
rect 24268 18816 24274 18828
rect 25409 18819 25467 18825
rect 25409 18816 25421 18819
rect 24268 18788 25421 18816
rect 24268 18776 24274 18788
rect 25409 18785 25421 18788
rect 25455 18785 25467 18819
rect 25409 18779 25467 18785
rect 15930 18748 15936 18760
rect 15891 18720 15936 18748
rect 15930 18708 15936 18720
rect 15988 18708 15994 18760
rect 16298 18708 16304 18760
rect 16356 18748 16362 18760
rect 16393 18751 16451 18757
rect 16393 18748 16405 18751
rect 16356 18720 16405 18748
rect 16356 18708 16362 18720
rect 16393 18717 16405 18720
rect 16439 18748 16451 18751
rect 17126 18748 17132 18760
rect 16439 18720 17132 18748
rect 16439 18717 16451 18720
rect 16393 18711 16451 18717
rect 17126 18708 17132 18720
rect 17184 18708 17190 18760
rect 19797 18751 19855 18757
rect 19797 18717 19809 18751
rect 19843 18748 19855 18751
rect 20622 18748 20628 18760
rect 19843 18720 20628 18748
rect 19843 18717 19855 18720
rect 19797 18711 19855 18717
rect 20622 18708 20628 18720
rect 20680 18708 20686 18760
rect 22462 18748 22468 18760
rect 22423 18720 22468 18748
rect 22462 18708 22468 18720
rect 22520 18708 22526 18760
rect 24578 18708 24584 18760
rect 24636 18748 24642 18760
rect 25038 18748 25044 18760
rect 24636 18720 25044 18748
rect 24636 18708 24642 18720
rect 25038 18708 25044 18720
rect 25096 18708 25102 18760
rect 19334 18640 19340 18692
rect 19392 18680 19398 18692
rect 20162 18680 20168 18692
rect 19392 18652 20168 18680
rect 19392 18640 19398 18652
rect 20162 18640 20168 18652
rect 20220 18680 20226 18692
rect 20257 18683 20315 18689
rect 20257 18680 20269 18683
rect 20220 18652 20269 18680
rect 20220 18640 20226 18652
rect 20257 18649 20269 18652
rect 20303 18649 20315 18683
rect 20257 18643 20315 18649
rect 21913 18683 21971 18689
rect 21913 18649 21925 18683
rect 21959 18680 21971 18683
rect 22094 18680 22100 18692
rect 21959 18652 22100 18680
rect 21959 18649 21971 18652
rect 21913 18643 21971 18649
rect 22094 18640 22100 18652
rect 22152 18680 22158 18692
rect 23569 18683 23627 18689
rect 23569 18680 23581 18683
rect 22152 18652 23581 18680
rect 22152 18640 22158 18652
rect 23569 18649 23581 18652
rect 23615 18649 23627 18683
rect 23569 18643 23627 18649
rect 23937 18683 23995 18689
rect 23937 18649 23949 18683
rect 23983 18680 23995 18683
rect 24762 18680 24768 18692
rect 23983 18652 24768 18680
rect 23983 18649 23995 18652
rect 23937 18643 23995 18649
rect 24762 18640 24768 18652
rect 24820 18680 24826 18692
rect 25225 18683 25283 18689
rect 25225 18680 25237 18683
rect 24820 18652 25237 18680
rect 24820 18640 24826 18652
rect 25225 18649 25237 18652
rect 25271 18649 25283 18683
rect 25225 18643 25283 18649
rect 15013 18615 15071 18621
rect 15013 18612 15025 18615
rect 14884 18584 15025 18612
rect 14884 18572 14890 18584
rect 15013 18581 15025 18584
rect 15059 18581 15071 18615
rect 15378 18612 15384 18624
rect 15339 18584 15384 18612
rect 15013 18575 15071 18581
rect 15378 18572 15384 18584
rect 15436 18572 15442 18624
rect 18506 18612 18512 18624
rect 18467 18584 18512 18612
rect 18506 18572 18512 18584
rect 18564 18572 18570 18624
rect 19705 18615 19763 18621
rect 19705 18581 19717 18615
rect 19751 18612 19763 18615
rect 20346 18612 20352 18624
rect 19751 18584 20352 18612
rect 19751 18581 19763 18584
rect 19705 18575 19763 18581
rect 20346 18572 20352 18584
rect 20404 18612 20410 18624
rect 21174 18612 21180 18624
rect 20404 18584 21180 18612
rect 20404 18572 20410 18584
rect 21174 18572 21180 18584
rect 21232 18572 21238 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 8386 18368 8392 18420
rect 8444 18408 8450 18420
rect 9585 18411 9643 18417
rect 9585 18408 9597 18411
rect 8444 18380 9597 18408
rect 8444 18368 8450 18380
rect 9585 18377 9597 18380
rect 9631 18377 9643 18411
rect 10594 18408 10600 18420
rect 10555 18380 10600 18408
rect 9585 18371 9643 18377
rect 10594 18368 10600 18380
rect 10652 18368 10658 18420
rect 11241 18411 11299 18417
rect 11241 18377 11253 18411
rect 11287 18408 11299 18411
rect 12710 18408 12716 18420
rect 11287 18380 12716 18408
rect 11287 18377 11299 18380
rect 11241 18371 11299 18377
rect 12710 18368 12716 18380
rect 12768 18368 12774 18420
rect 13817 18411 13875 18417
rect 13817 18377 13829 18411
rect 13863 18408 13875 18411
rect 14090 18408 14096 18420
rect 13863 18380 14096 18408
rect 13863 18377 13875 18380
rect 13817 18371 13875 18377
rect 14090 18368 14096 18380
rect 14148 18368 14154 18420
rect 15013 18411 15071 18417
rect 15013 18377 15025 18411
rect 15059 18408 15071 18411
rect 15654 18408 15660 18420
rect 15059 18380 15660 18408
rect 15059 18377 15071 18380
rect 15013 18371 15071 18377
rect 15654 18368 15660 18380
rect 15712 18368 15718 18420
rect 18141 18411 18199 18417
rect 18141 18377 18153 18411
rect 18187 18408 18199 18411
rect 19978 18408 19984 18420
rect 18187 18380 19984 18408
rect 18187 18377 18199 18380
rect 18141 18371 18199 18377
rect 19978 18368 19984 18380
rect 20036 18368 20042 18420
rect 23109 18411 23167 18417
rect 23109 18377 23121 18411
rect 23155 18408 23167 18411
rect 24210 18408 24216 18420
rect 23155 18380 24216 18408
rect 23155 18377 23167 18380
rect 23109 18371 23167 18377
rect 24210 18368 24216 18380
rect 24268 18368 24274 18420
rect 24397 18411 24455 18417
rect 24397 18377 24409 18411
rect 24443 18408 24455 18411
rect 24854 18408 24860 18420
rect 24443 18380 24860 18408
rect 24443 18377 24455 18380
rect 24397 18371 24455 18377
rect 24854 18368 24860 18380
rect 24912 18368 24918 18420
rect 19518 18340 19524 18352
rect 19479 18312 19524 18340
rect 19518 18300 19524 18312
rect 19576 18340 19582 18352
rect 23474 18340 23480 18352
rect 19576 18312 19656 18340
rect 23435 18312 23480 18340
rect 19576 18300 19582 18312
rect 8665 18275 8723 18281
rect 8665 18241 8677 18275
rect 8711 18272 8723 18275
rect 9490 18272 9496 18284
rect 8711 18244 9496 18272
rect 8711 18241 8723 18244
rect 8665 18235 8723 18241
rect 9490 18232 9496 18244
rect 9548 18272 9554 18284
rect 10134 18272 10140 18284
rect 9548 18244 10140 18272
rect 9548 18232 9554 18244
rect 10134 18232 10140 18244
rect 10192 18232 10198 18284
rect 11514 18232 11520 18284
rect 11572 18272 11578 18284
rect 12434 18272 12440 18284
rect 11572 18244 12440 18272
rect 11572 18232 11578 18244
rect 12434 18232 12440 18244
rect 12492 18232 12498 18284
rect 19628 18281 19656 18312
rect 23474 18300 23480 18312
rect 23532 18300 23538 18352
rect 19613 18275 19671 18281
rect 19613 18241 19625 18275
rect 19659 18241 19671 18275
rect 19613 18235 19671 18241
rect 22373 18275 22431 18281
rect 22373 18241 22385 18275
rect 22419 18272 22431 18275
rect 22830 18272 22836 18284
rect 22419 18244 22836 18272
rect 22419 18241 22431 18244
rect 22373 18235 22431 18241
rect 22830 18232 22836 18244
rect 22888 18232 22894 18284
rect 24946 18272 24952 18284
rect 24907 18244 24952 18272
rect 24946 18232 24952 18244
rect 25004 18272 25010 18284
rect 25314 18272 25320 18284
rect 25004 18244 25320 18272
rect 25004 18232 25010 18244
rect 25314 18232 25320 18244
rect 25372 18232 25378 18284
rect 9033 18207 9091 18213
rect 9033 18173 9045 18207
rect 9079 18204 9091 18207
rect 9858 18204 9864 18216
rect 9079 18176 9864 18204
rect 9079 18173 9091 18176
rect 9033 18167 9091 18173
rect 9858 18164 9864 18176
rect 9916 18164 9922 18216
rect 12158 18204 12164 18216
rect 12119 18176 12164 18204
rect 12158 18164 12164 18176
rect 12216 18164 12222 18216
rect 15381 18207 15439 18213
rect 15381 18173 15393 18207
rect 15427 18204 15439 18207
rect 15473 18207 15531 18213
rect 15473 18204 15485 18207
rect 15427 18176 15485 18204
rect 15427 18173 15439 18176
rect 15381 18167 15439 18173
rect 15473 18173 15485 18176
rect 15519 18204 15531 18207
rect 16298 18204 16304 18216
rect 15519 18176 16304 18204
rect 15519 18173 15531 18176
rect 15473 18167 15531 18173
rect 16298 18164 16304 18176
rect 16356 18164 16362 18216
rect 17865 18207 17923 18213
rect 17865 18173 17877 18207
rect 17911 18204 17923 18207
rect 17911 18176 18644 18204
rect 17911 18173 17923 18176
rect 17865 18167 17923 18173
rect 18616 18148 18644 18176
rect 22094 18164 22100 18216
rect 22152 18204 22158 18216
rect 22152 18176 22197 18204
rect 22152 18164 22158 18176
rect 24026 18164 24032 18216
rect 24084 18204 24090 18216
rect 24213 18207 24271 18213
rect 24213 18204 24225 18207
rect 24084 18176 24225 18204
rect 24084 18164 24090 18176
rect 24213 18173 24225 18176
rect 24259 18204 24271 18207
rect 24670 18204 24676 18216
rect 24259 18176 24676 18204
rect 24259 18173 24271 18176
rect 24213 18167 24271 18173
rect 24670 18164 24676 18176
rect 24728 18164 24734 18216
rect 25685 18207 25743 18213
rect 25685 18204 25697 18207
rect 24872 18176 25697 18204
rect 12710 18145 12716 18148
rect 12704 18136 12716 18145
rect 12671 18108 12716 18136
rect 12704 18099 12716 18108
rect 12710 18096 12716 18099
rect 12768 18096 12774 18148
rect 15718 18139 15776 18145
rect 15718 18136 15730 18139
rect 14568 18108 15730 18136
rect 9306 18068 9312 18080
rect 9267 18040 9312 18068
rect 9306 18028 9312 18040
rect 9364 18068 9370 18080
rect 10045 18071 10103 18077
rect 10045 18068 10057 18071
rect 9364 18040 10057 18068
rect 9364 18028 9370 18040
rect 10045 18037 10057 18040
rect 10091 18068 10103 18071
rect 10686 18068 10692 18080
rect 10091 18040 10692 18068
rect 10091 18037 10103 18040
rect 10045 18031 10103 18037
rect 10686 18028 10692 18040
rect 10744 18028 10750 18080
rect 11330 18068 11336 18080
rect 11291 18040 11336 18068
rect 11330 18028 11336 18040
rect 11388 18028 11394 18080
rect 14274 18028 14280 18080
rect 14332 18068 14338 18080
rect 14568 18077 14596 18108
rect 15718 18105 15730 18108
rect 15764 18136 15776 18139
rect 15930 18136 15936 18148
rect 15764 18108 15936 18136
rect 15764 18105 15776 18108
rect 15718 18099 15776 18105
rect 15930 18096 15936 18108
rect 15988 18096 15994 18148
rect 18138 18096 18144 18148
rect 18196 18136 18202 18148
rect 18417 18139 18475 18145
rect 18417 18136 18429 18139
rect 18196 18108 18429 18136
rect 18196 18096 18202 18108
rect 18417 18105 18429 18108
rect 18463 18105 18475 18139
rect 18598 18136 18604 18148
rect 18559 18108 18604 18136
rect 18417 18099 18475 18105
rect 18598 18096 18604 18108
rect 18656 18096 18662 18148
rect 18693 18139 18751 18145
rect 18693 18105 18705 18139
rect 18739 18136 18751 18139
rect 19061 18139 19119 18145
rect 19061 18136 19073 18139
rect 18739 18108 19073 18136
rect 18739 18105 18751 18108
rect 18693 18099 18751 18105
rect 19061 18105 19073 18108
rect 19107 18136 19119 18139
rect 19518 18136 19524 18148
rect 19107 18108 19524 18136
rect 19107 18105 19119 18108
rect 19061 18099 19119 18105
rect 19518 18096 19524 18108
rect 19576 18136 19582 18148
rect 19858 18139 19916 18145
rect 19858 18136 19870 18139
rect 19576 18108 19870 18136
rect 19576 18096 19582 18108
rect 19858 18105 19870 18108
rect 19904 18105 19916 18139
rect 23474 18136 23480 18148
rect 19858 18099 19916 18105
rect 22480 18108 23480 18136
rect 22480 18080 22508 18108
rect 23474 18096 23480 18108
rect 23532 18096 23538 18148
rect 24762 18096 24768 18148
rect 24820 18136 24826 18148
rect 24872 18145 24900 18176
rect 25685 18173 25697 18176
rect 25731 18173 25743 18207
rect 25685 18167 25743 18173
rect 24857 18139 24915 18145
rect 24857 18136 24869 18139
rect 24820 18108 24869 18136
rect 24820 18096 24826 18108
rect 24857 18105 24869 18108
rect 24903 18105 24915 18139
rect 24857 18099 24915 18105
rect 14553 18071 14611 18077
rect 14553 18068 14565 18071
rect 14332 18040 14565 18068
rect 14332 18028 14338 18040
rect 14553 18037 14565 18040
rect 14599 18037 14611 18071
rect 14553 18031 14611 18037
rect 16758 18028 16764 18080
rect 16816 18068 16822 18080
rect 16853 18071 16911 18077
rect 16853 18068 16865 18071
rect 16816 18040 16865 18068
rect 16816 18028 16822 18040
rect 16853 18037 16865 18040
rect 16899 18037 16911 18071
rect 16853 18031 16911 18037
rect 17126 18028 17132 18080
rect 17184 18068 17190 18080
rect 17494 18068 17500 18080
rect 17184 18040 17500 18068
rect 17184 18028 17190 18040
rect 17494 18028 17500 18040
rect 17552 18068 17558 18080
rect 18322 18068 18328 18080
rect 17552 18040 18328 18068
rect 17552 18028 17558 18040
rect 18322 18028 18328 18040
rect 18380 18028 18386 18080
rect 20993 18071 21051 18077
rect 20993 18037 21005 18071
rect 21039 18068 21051 18071
rect 21174 18068 21180 18080
rect 21039 18040 21180 18068
rect 21039 18037 21051 18040
rect 20993 18031 21051 18037
rect 21174 18028 21180 18040
rect 21232 18028 21238 18080
rect 21913 18071 21971 18077
rect 21913 18037 21925 18071
rect 21959 18068 21971 18071
rect 22462 18068 22468 18080
rect 21959 18040 22468 18068
rect 21959 18037 21971 18040
rect 21913 18031 21971 18037
rect 22462 18028 22468 18040
rect 22520 18028 22526 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 9490 17864 9496 17876
rect 9451 17836 9496 17864
rect 9490 17824 9496 17836
rect 9548 17824 9554 17876
rect 11514 17864 11520 17876
rect 11348 17836 11520 17864
rect 9766 17756 9772 17808
rect 9824 17796 9830 17808
rect 10321 17799 10379 17805
rect 10321 17796 10333 17799
rect 9824 17768 10333 17796
rect 9824 17756 9830 17768
rect 10321 17765 10333 17768
rect 10367 17796 10379 17799
rect 11054 17796 11060 17808
rect 10367 17768 11060 17796
rect 10367 17765 10379 17768
rect 10321 17759 10379 17765
rect 11054 17756 11060 17768
rect 11112 17756 11118 17808
rect 11348 17737 11376 17836
rect 11514 17824 11520 17836
rect 11572 17824 11578 17876
rect 13725 17867 13783 17873
rect 13725 17833 13737 17867
rect 13771 17864 13783 17867
rect 14274 17864 14280 17876
rect 13771 17836 14280 17864
rect 13771 17833 13783 17836
rect 13725 17827 13783 17833
rect 14274 17824 14280 17836
rect 14332 17824 14338 17876
rect 14458 17864 14464 17876
rect 14419 17836 14464 17864
rect 14458 17824 14464 17836
rect 14516 17824 14522 17876
rect 15838 17864 15844 17876
rect 15799 17836 15844 17864
rect 15838 17824 15844 17836
rect 15896 17824 15902 17876
rect 17313 17867 17371 17873
rect 17313 17833 17325 17867
rect 17359 17864 17371 17867
rect 18138 17864 18144 17876
rect 17359 17836 18144 17864
rect 17359 17833 17371 17836
rect 17313 17827 17371 17833
rect 18138 17824 18144 17836
rect 18196 17824 18202 17876
rect 19518 17824 19524 17876
rect 19576 17864 19582 17876
rect 19705 17867 19763 17873
rect 19705 17864 19717 17867
rect 19576 17836 19717 17864
rect 19576 17824 19582 17836
rect 19705 17833 19717 17836
rect 19751 17864 19763 17867
rect 20257 17867 20315 17873
rect 20257 17864 20269 17867
rect 19751 17836 20269 17864
rect 19751 17833 19763 17836
rect 19705 17827 19763 17833
rect 20257 17833 20269 17836
rect 20303 17833 20315 17867
rect 20257 17827 20315 17833
rect 22370 17824 22376 17876
rect 22428 17864 22434 17876
rect 23201 17867 23259 17873
rect 23201 17864 23213 17867
rect 22428 17836 23213 17864
rect 22428 17824 22434 17836
rect 23201 17833 23213 17836
rect 23247 17833 23259 17867
rect 23201 17827 23259 17833
rect 23566 17824 23572 17876
rect 23624 17864 23630 17876
rect 23842 17864 23848 17876
rect 23624 17836 23848 17864
rect 23624 17824 23630 17836
rect 23842 17824 23848 17836
rect 23900 17824 23906 17876
rect 25314 17864 25320 17876
rect 25275 17836 25320 17864
rect 25314 17824 25320 17836
rect 25372 17824 25378 17876
rect 14292 17796 14320 17824
rect 15013 17799 15071 17805
rect 15013 17796 15025 17799
rect 14292 17768 15025 17796
rect 15013 17765 15025 17768
rect 15059 17765 15071 17799
rect 15013 17759 15071 17765
rect 18506 17756 18512 17808
rect 18564 17805 18570 17808
rect 18564 17799 18628 17805
rect 18564 17765 18582 17799
rect 18616 17765 18628 17799
rect 18564 17759 18628 17765
rect 18564 17756 18570 17759
rect 11333 17731 11391 17737
rect 11333 17697 11345 17731
rect 11379 17697 11391 17731
rect 11589 17731 11647 17737
rect 11589 17728 11601 17731
rect 11333 17691 11391 17697
rect 11440 17700 11601 17728
rect 10318 17660 10324 17672
rect 10279 17632 10324 17660
rect 10318 17620 10324 17632
rect 10376 17620 10382 17672
rect 10410 17620 10416 17672
rect 10468 17660 10474 17672
rect 10778 17660 10784 17672
rect 10468 17632 10784 17660
rect 10468 17620 10474 17632
rect 10778 17620 10784 17632
rect 10836 17620 10842 17672
rect 10873 17663 10931 17669
rect 10873 17629 10885 17663
rect 10919 17660 10931 17663
rect 11146 17660 11152 17672
rect 10919 17632 11152 17660
rect 10919 17629 10931 17632
rect 10873 17623 10931 17629
rect 11146 17620 11152 17632
rect 11204 17660 11210 17672
rect 11440 17660 11468 17700
rect 11589 17697 11601 17700
rect 11635 17697 11647 17731
rect 11589 17691 11647 17697
rect 14734 17688 14740 17740
rect 14792 17728 14798 17740
rect 15378 17728 15384 17740
rect 14792 17700 15384 17728
rect 14792 17688 14798 17700
rect 15378 17688 15384 17700
rect 15436 17728 15442 17740
rect 21174 17737 21180 17740
rect 15657 17731 15715 17737
rect 15657 17728 15669 17731
rect 15436 17700 15669 17728
rect 15436 17688 15442 17700
rect 15657 17697 15669 17700
rect 15703 17697 15715 17731
rect 21168 17728 21180 17737
rect 21135 17700 21180 17728
rect 15657 17691 15715 17697
rect 21168 17691 21180 17700
rect 21174 17688 21180 17691
rect 21232 17688 21238 17740
rect 24210 17737 24216 17740
rect 24204 17691 24216 17737
rect 24268 17728 24274 17740
rect 24268 17700 24304 17728
rect 24210 17688 24216 17691
rect 24268 17688 24274 17700
rect 11204 17632 11468 17660
rect 11204 17620 11210 17632
rect 15562 17620 15568 17672
rect 15620 17660 15626 17672
rect 15933 17663 15991 17669
rect 15933 17660 15945 17663
rect 15620 17632 15945 17660
rect 15620 17620 15626 17632
rect 15933 17629 15945 17632
rect 15979 17660 15991 17663
rect 16758 17660 16764 17672
rect 15979 17632 16764 17660
rect 15979 17629 15991 17632
rect 15933 17623 15991 17629
rect 16758 17620 16764 17632
rect 16816 17660 16822 17672
rect 17129 17663 17187 17669
rect 17129 17660 17141 17663
rect 16816 17632 17141 17660
rect 16816 17620 16822 17632
rect 17129 17629 17141 17632
rect 17175 17629 17187 17663
rect 18322 17660 18328 17672
rect 18283 17632 18328 17660
rect 17129 17623 17187 17629
rect 18322 17620 18328 17632
rect 18380 17620 18386 17672
rect 20898 17660 20904 17672
rect 20859 17632 20904 17660
rect 20898 17620 20904 17632
rect 20956 17620 20962 17672
rect 23658 17620 23664 17672
rect 23716 17660 23722 17672
rect 23937 17663 23995 17669
rect 23937 17660 23949 17663
rect 23716 17632 23949 17660
rect 23716 17620 23722 17632
rect 23937 17629 23949 17632
rect 23983 17629 23995 17663
rect 23937 17623 23995 17629
rect 9861 17595 9919 17601
rect 9861 17561 9873 17595
rect 9907 17592 9919 17595
rect 10962 17592 10968 17604
rect 9907 17564 10968 17592
rect 9907 17561 9919 17564
rect 9861 17555 9919 17561
rect 10962 17552 10968 17564
rect 11020 17552 11026 17604
rect 15381 17595 15439 17601
rect 15381 17561 15393 17595
rect 15427 17592 15439 17595
rect 16482 17592 16488 17604
rect 15427 17564 16488 17592
rect 15427 17561 15439 17564
rect 15381 17555 15439 17561
rect 16482 17552 16488 17564
rect 16540 17552 16546 17604
rect 11241 17527 11299 17533
rect 11241 17493 11253 17527
rect 11287 17524 11299 17527
rect 11698 17524 11704 17536
rect 11287 17496 11704 17524
rect 11287 17493 11299 17496
rect 11241 17487 11299 17493
rect 11698 17484 11704 17496
rect 11756 17484 11762 17536
rect 12250 17484 12256 17536
rect 12308 17524 12314 17536
rect 12710 17524 12716 17536
rect 12308 17496 12716 17524
rect 12308 17484 12314 17496
rect 12710 17484 12716 17496
rect 12768 17524 12774 17536
rect 13078 17524 13084 17536
rect 12768 17496 13084 17524
rect 12768 17484 12774 17496
rect 13078 17484 13084 17496
rect 13136 17524 13142 17536
rect 13265 17527 13323 17533
rect 13265 17524 13277 17527
rect 13136 17496 13277 17524
rect 13136 17484 13142 17496
rect 13265 17493 13277 17496
rect 13311 17493 13323 17527
rect 13265 17487 13323 17493
rect 14093 17527 14151 17533
rect 14093 17493 14105 17527
rect 14139 17524 14151 17527
rect 14826 17524 14832 17536
rect 14139 17496 14832 17524
rect 14139 17493 14151 17496
rect 14093 17487 14151 17493
rect 14826 17484 14832 17496
rect 14884 17484 14890 17536
rect 16393 17527 16451 17533
rect 16393 17493 16405 17527
rect 16439 17524 16451 17527
rect 17034 17524 17040 17536
rect 16439 17496 17040 17524
rect 16439 17493 16451 17496
rect 16393 17487 16451 17493
rect 17034 17484 17040 17496
rect 17092 17484 17098 17536
rect 22278 17524 22284 17536
rect 22239 17496 22284 17524
rect 22278 17484 22284 17496
rect 22336 17484 22342 17536
rect 22462 17484 22468 17536
rect 22520 17524 22526 17536
rect 22833 17527 22891 17533
rect 22833 17524 22845 17527
rect 22520 17496 22845 17524
rect 22520 17484 22526 17496
rect 22833 17493 22845 17496
rect 22879 17493 22891 17527
rect 23750 17524 23756 17536
rect 23711 17496 23756 17524
rect 22833 17487 22891 17493
rect 23750 17484 23756 17496
rect 23808 17484 23814 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 9493 17323 9551 17329
rect 9493 17289 9505 17323
rect 9539 17320 9551 17323
rect 10410 17320 10416 17332
rect 9539 17292 10416 17320
rect 9539 17289 9551 17292
rect 9493 17283 9551 17289
rect 10410 17280 10416 17292
rect 10468 17280 10474 17332
rect 10873 17323 10931 17329
rect 10873 17289 10885 17323
rect 10919 17320 10931 17323
rect 11790 17320 11796 17332
rect 10919 17292 11796 17320
rect 10919 17289 10931 17292
rect 10873 17283 10931 17289
rect 11790 17280 11796 17292
rect 11848 17280 11854 17332
rect 12250 17320 12256 17332
rect 12211 17292 12256 17320
rect 12250 17280 12256 17292
rect 12308 17280 12314 17332
rect 12526 17320 12532 17332
rect 12487 17292 12532 17320
rect 12526 17280 12532 17292
rect 12584 17280 12590 17332
rect 15381 17323 15439 17329
rect 15381 17289 15393 17323
rect 15427 17320 15439 17323
rect 15562 17320 15568 17332
rect 15427 17292 15568 17320
rect 15427 17289 15439 17292
rect 15381 17283 15439 17289
rect 15562 17280 15568 17292
rect 15620 17280 15626 17332
rect 15749 17323 15807 17329
rect 15749 17289 15761 17323
rect 15795 17320 15807 17323
rect 15838 17320 15844 17332
rect 15795 17292 15844 17320
rect 15795 17289 15807 17292
rect 15749 17283 15807 17289
rect 15838 17280 15844 17292
rect 15896 17280 15902 17332
rect 17865 17323 17923 17329
rect 17865 17289 17877 17323
rect 17911 17320 17923 17323
rect 18506 17320 18512 17332
rect 17911 17292 18512 17320
rect 17911 17289 17923 17292
rect 17865 17283 17923 17289
rect 18506 17280 18512 17292
rect 18564 17280 18570 17332
rect 18601 17323 18659 17329
rect 18601 17289 18613 17323
rect 18647 17320 18659 17323
rect 19334 17320 19340 17332
rect 18647 17292 19340 17320
rect 18647 17289 18659 17292
rect 18601 17283 18659 17289
rect 19334 17280 19340 17292
rect 19392 17280 19398 17332
rect 21726 17320 21732 17332
rect 19628 17292 20760 17320
rect 21687 17292 21732 17320
rect 14090 17252 14096 17264
rect 14051 17224 14096 17252
rect 14090 17212 14096 17224
rect 14148 17212 14154 17264
rect 16482 17252 16488 17264
rect 16443 17224 16488 17252
rect 16482 17212 16488 17224
rect 16540 17212 16546 17264
rect 18322 17252 18328 17264
rect 18283 17224 18328 17252
rect 18322 17212 18328 17224
rect 18380 17212 18386 17264
rect 18524 17252 18552 17280
rect 19628 17261 19656 17292
rect 19613 17255 19671 17261
rect 19613 17252 19625 17255
rect 18524 17224 19625 17252
rect 19613 17221 19625 17224
rect 19659 17221 19671 17255
rect 19613 17215 19671 17221
rect 20165 17255 20223 17261
rect 20165 17221 20177 17255
rect 20211 17221 20223 17255
rect 20165 17215 20223 17221
rect 10689 17187 10747 17193
rect 10689 17153 10701 17187
rect 10735 17184 10747 17187
rect 11330 17184 11336 17196
rect 10735 17156 11336 17184
rect 10735 17153 10747 17156
rect 10689 17147 10747 17153
rect 11330 17144 11336 17156
rect 11388 17144 11394 17196
rect 13078 17184 13084 17196
rect 13039 17156 13084 17184
rect 13078 17144 13084 17156
rect 13136 17144 13142 17196
rect 14458 17144 14464 17196
rect 14516 17184 14522 17196
rect 14553 17187 14611 17193
rect 14553 17184 14565 17187
rect 14516 17156 14565 17184
rect 14516 17144 14522 17156
rect 14553 17153 14565 17156
rect 14599 17184 14611 17187
rect 14826 17184 14832 17196
rect 14599 17156 14832 17184
rect 14599 17153 14611 17156
rect 14553 17147 14611 17153
rect 14826 17144 14832 17156
rect 14884 17144 14890 17196
rect 17034 17184 17040 17196
rect 16995 17156 17040 17184
rect 17034 17144 17040 17156
rect 17092 17144 17098 17196
rect 19058 17184 19064 17196
rect 19019 17156 19064 17184
rect 19058 17144 19064 17156
rect 19116 17144 19122 17196
rect 19153 17187 19211 17193
rect 19153 17153 19165 17187
rect 19199 17184 19211 17187
rect 19518 17184 19524 17196
rect 19199 17156 19524 17184
rect 19199 17153 19211 17156
rect 19153 17147 19211 17153
rect 19518 17144 19524 17156
rect 19576 17144 19582 17196
rect 11146 17076 11152 17128
rect 11204 17116 11210 17128
rect 11425 17119 11483 17125
rect 11425 17116 11437 17119
rect 11204 17088 11437 17116
rect 11204 17076 11210 17088
rect 11425 17085 11437 17088
rect 11471 17085 11483 17119
rect 11425 17079 11483 17085
rect 13541 17119 13599 17125
rect 13541 17085 13553 17119
rect 13587 17116 13599 17119
rect 14645 17119 14703 17125
rect 14645 17116 14657 17119
rect 13587 17088 14657 17116
rect 13587 17085 13599 17088
rect 13541 17079 13599 17085
rect 14645 17085 14657 17088
rect 14691 17085 14703 17119
rect 16758 17116 16764 17128
rect 16719 17088 16764 17116
rect 14645 17079 14703 17085
rect 9861 17051 9919 17057
rect 9861 17017 9873 17051
rect 9907 17048 9919 17051
rect 10318 17048 10324 17060
rect 9907 17020 10324 17048
rect 9907 17017 9919 17020
rect 9861 17011 9919 17017
rect 10318 17008 10324 17020
rect 10376 17048 10382 17060
rect 11238 17048 11244 17060
rect 10376 17020 11244 17048
rect 10376 17008 10382 17020
rect 11238 17008 11244 17020
rect 11296 17008 11302 17060
rect 11790 17008 11796 17060
rect 11848 17048 11854 17060
rect 12805 17051 12863 17057
rect 12805 17048 12817 17051
rect 11848 17020 12817 17048
rect 11848 17008 11854 17020
rect 12805 17017 12817 17020
rect 12851 17017 12863 17051
rect 12805 17011 12863 17017
rect 13814 17008 13820 17060
rect 13872 17048 13878 17060
rect 13909 17051 13967 17057
rect 13909 17048 13921 17051
rect 13872 17020 13921 17048
rect 13872 17008 13878 17020
rect 13909 17017 13921 17020
rect 13955 17048 13967 17051
rect 14366 17048 14372 17060
rect 13955 17020 14372 17048
rect 13955 17017 13967 17020
rect 13909 17011 13967 17017
rect 14366 17008 14372 17020
rect 14424 17048 14430 17060
rect 14553 17051 14611 17057
rect 14553 17048 14565 17051
rect 14424 17020 14565 17048
rect 14424 17008 14430 17020
rect 14553 17017 14565 17020
rect 14599 17017 14611 17051
rect 14660 17048 14688 17079
rect 16758 17076 16764 17088
rect 16816 17076 16822 17128
rect 17497 17119 17555 17125
rect 17497 17085 17509 17119
rect 17543 17116 17555 17119
rect 20180 17116 20208 17215
rect 20622 17184 20628 17196
rect 20583 17156 20628 17184
rect 20622 17144 20628 17156
rect 20680 17144 20686 17196
rect 20732 17193 20760 17292
rect 21726 17280 21732 17292
rect 21784 17280 21790 17332
rect 22005 17323 22063 17329
rect 22005 17289 22017 17323
rect 22051 17320 22063 17323
rect 22370 17320 22376 17332
rect 22051 17292 22376 17320
rect 22051 17289 22063 17292
rect 22005 17283 22063 17289
rect 22370 17280 22376 17292
rect 22428 17280 22434 17332
rect 20717 17187 20775 17193
rect 20717 17153 20729 17187
rect 20763 17153 20775 17187
rect 21744 17184 21772 17280
rect 22373 17187 22431 17193
rect 22373 17184 22385 17187
rect 21744 17156 22385 17184
rect 20717 17147 20775 17153
rect 22373 17153 22385 17156
rect 22419 17153 22431 17187
rect 22373 17147 22431 17153
rect 17543 17088 20208 17116
rect 17543 17085 17555 17088
rect 17497 17079 17555 17085
rect 14826 17048 14832 17060
rect 14660 17020 14832 17048
rect 14553 17011 14611 17017
rect 14826 17008 14832 17020
rect 14884 17008 14890 17060
rect 19076 17057 19104 17088
rect 19061 17051 19119 17057
rect 19061 17017 19073 17051
rect 19107 17017 19119 17051
rect 19061 17011 19119 17017
rect 19150 17008 19156 17060
rect 19208 17048 19214 17060
rect 19981 17051 20039 17057
rect 19981 17048 19993 17051
rect 19208 17020 19993 17048
rect 19208 17008 19214 17020
rect 19981 17017 19993 17020
rect 20027 17048 20039 17051
rect 20640 17048 20668 17144
rect 23658 17116 23664 17128
rect 23619 17088 23664 17116
rect 23658 17076 23664 17088
rect 23716 17076 23722 17128
rect 22462 17048 22468 17060
rect 20027 17020 20668 17048
rect 22423 17020 22468 17048
rect 20027 17017 20039 17020
rect 19981 17011 20039 17017
rect 22462 17008 22468 17020
rect 22520 17008 22526 17060
rect 22557 17051 22615 17057
rect 22557 17017 22569 17051
rect 22603 17017 22615 17051
rect 23750 17048 23756 17060
rect 22557 17011 22615 17017
rect 23124 17020 23756 17048
rect 9766 16940 9772 16992
rect 9824 16980 9830 16992
rect 10137 16983 10195 16989
rect 10137 16980 10149 16983
rect 9824 16952 10149 16980
rect 9824 16940 9830 16952
rect 10137 16949 10149 16952
rect 10183 16949 10195 16983
rect 10137 16943 10195 16949
rect 10962 16940 10968 16992
rect 11020 16980 11026 16992
rect 11333 16983 11391 16989
rect 11333 16980 11345 16983
rect 11020 16952 11345 16980
rect 11020 16940 11026 16952
rect 11333 16949 11345 16952
rect 11379 16949 11391 16983
rect 11333 16943 11391 16949
rect 11514 16940 11520 16992
rect 11572 16980 11578 16992
rect 11885 16983 11943 16989
rect 11885 16980 11897 16983
rect 11572 16952 11897 16980
rect 11572 16940 11578 16952
rect 11885 16949 11897 16952
rect 11931 16949 11943 16983
rect 12986 16980 12992 16992
rect 12947 16952 12992 16980
rect 11885 16943 11943 16949
rect 12986 16940 12992 16952
rect 13044 16940 13050 16992
rect 16301 16983 16359 16989
rect 16301 16949 16313 16983
rect 16347 16980 16359 16983
rect 16942 16980 16948 16992
rect 16347 16952 16948 16980
rect 16347 16949 16359 16952
rect 16301 16943 16359 16949
rect 16942 16940 16948 16952
rect 17000 16940 17006 16992
rect 20622 16980 20628 16992
rect 20583 16952 20628 16980
rect 20622 16940 20628 16952
rect 20680 16940 20686 16992
rect 20898 16940 20904 16992
rect 20956 16980 20962 16992
rect 21177 16983 21235 16989
rect 21177 16980 21189 16983
rect 20956 16952 21189 16980
rect 20956 16940 20962 16952
rect 21177 16949 21189 16952
rect 21223 16980 21235 16983
rect 21910 16980 21916 16992
rect 21223 16952 21916 16980
rect 21223 16949 21235 16952
rect 21177 16943 21235 16949
rect 21910 16940 21916 16952
rect 21968 16940 21974 16992
rect 22572 16980 22600 17011
rect 23124 16992 23152 17020
rect 23750 17008 23756 17020
rect 23808 17048 23814 17060
rect 23906 17051 23964 17057
rect 23906 17048 23918 17051
rect 23808 17020 23918 17048
rect 23808 17008 23814 17020
rect 23906 17017 23918 17020
rect 23952 17017 23964 17051
rect 23906 17011 23964 17017
rect 23017 16983 23075 16989
rect 23017 16980 23029 16983
rect 22572 16952 23029 16980
rect 23017 16949 23029 16952
rect 23063 16980 23075 16983
rect 23106 16980 23112 16992
rect 23063 16952 23112 16980
rect 23063 16949 23075 16952
rect 23017 16943 23075 16949
rect 23106 16940 23112 16952
rect 23164 16940 23170 16992
rect 23290 16940 23296 16992
rect 23348 16980 23354 16992
rect 23477 16983 23535 16989
rect 23477 16980 23489 16983
rect 23348 16952 23489 16980
rect 23348 16940 23354 16952
rect 23477 16949 23489 16952
rect 23523 16980 23535 16983
rect 23658 16980 23664 16992
rect 23523 16952 23664 16980
rect 23523 16949 23535 16952
rect 23477 16943 23535 16949
rect 23658 16940 23664 16952
rect 23716 16940 23722 16992
rect 24670 16940 24676 16992
rect 24728 16980 24734 16992
rect 25041 16983 25099 16989
rect 25041 16980 25053 16983
rect 24728 16952 25053 16980
rect 24728 16940 24734 16952
rect 25041 16949 25053 16952
rect 25087 16949 25099 16983
rect 25041 16943 25099 16949
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 9943 16779 10001 16785
rect 9943 16745 9955 16779
rect 9989 16776 10001 16779
rect 10778 16776 10784 16788
rect 9989 16748 10784 16776
rect 9989 16745 10001 16748
rect 9943 16739 10001 16745
rect 10778 16736 10784 16748
rect 10836 16736 10842 16788
rect 10962 16776 10968 16788
rect 10923 16748 10968 16776
rect 10962 16736 10968 16748
rect 11020 16736 11026 16788
rect 12805 16779 12863 16785
rect 12805 16776 12817 16779
rect 11256 16748 12817 16776
rect 10134 16668 10140 16720
rect 10192 16708 10198 16720
rect 10229 16711 10287 16717
rect 10229 16708 10241 16711
rect 10192 16680 10241 16708
rect 10192 16668 10198 16680
rect 10229 16677 10241 16680
rect 10275 16677 10287 16711
rect 10229 16671 10287 16677
rect 10413 16711 10471 16717
rect 10413 16677 10425 16711
rect 10459 16677 10471 16711
rect 10413 16671 10471 16677
rect 10428 16640 10456 16671
rect 10502 16668 10508 16720
rect 10560 16708 10566 16720
rect 11146 16708 11152 16720
rect 10560 16680 11152 16708
rect 10560 16668 10566 16680
rect 11146 16668 11152 16680
rect 11204 16708 11210 16720
rect 11256 16717 11284 16748
rect 12805 16745 12817 16748
rect 12851 16745 12863 16779
rect 15363 16779 15421 16785
rect 15363 16776 15375 16779
rect 12805 16739 12863 16745
rect 13924 16748 15375 16776
rect 11241 16711 11299 16717
rect 11241 16708 11253 16711
rect 11204 16680 11253 16708
rect 11204 16668 11210 16680
rect 11241 16677 11253 16680
rect 11287 16677 11299 16711
rect 11241 16671 11299 16677
rect 11606 16668 11612 16720
rect 11664 16717 11670 16720
rect 11664 16711 11728 16717
rect 11664 16677 11682 16711
rect 11716 16677 11728 16711
rect 11664 16671 11728 16677
rect 11664 16668 11670 16671
rect 11425 16643 11483 16649
rect 9600 16612 11100 16640
rect 9600 16584 9628 16612
rect 11072 16584 11100 16612
rect 11425 16609 11437 16643
rect 11471 16640 11483 16643
rect 11514 16640 11520 16652
rect 11471 16612 11520 16640
rect 11471 16609 11483 16612
rect 11425 16603 11483 16609
rect 11514 16600 11520 16612
rect 11572 16600 11578 16652
rect 13924 16649 13952 16748
rect 15363 16745 15375 16748
rect 15409 16745 15421 16779
rect 15363 16739 15421 16745
rect 16482 16736 16488 16788
rect 16540 16776 16546 16788
rect 16761 16779 16819 16785
rect 16761 16776 16773 16779
rect 16540 16748 16773 16776
rect 16540 16736 16546 16748
rect 16761 16745 16773 16748
rect 16807 16776 16819 16779
rect 16942 16776 16948 16788
rect 16807 16748 16948 16776
rect 16807 16745 16819 16748
rect 16761 16739 16819 16745
rect 16942 16736 16948 16748
rect 17000 16736 17006 16788
rect 18407 16779 18465 16785
rect 18407 16745 18419 16779
rect 18453 16776 18465 16779
rect 19058 16776 19064 16788
rect 18453 16748 19064 16776
rect 18453 16745 18465 16748
rect 18407 16739 18465 16745
rect 19058 16736 19064 16748
rect 19116 16776 19122 16788
rect 19705 16779 19763 16785
rect 19705 16776 19717 16779
rect 19116 16748 19717 16776
rect 19116 16736 19122 16748
rect 19705 16745 19717 16748
rect 19751 16745 19763 16779
rect 21174 16776 21180 16788
rect 21135 16748 21180 16776
rect 19705 16739 19763 16745
rect 21174 16736 21180 16748
rect 21232 16736 21238 16788
rect 23658 16736 23664 16788
rect 23716 16776 23722 16788
rect 23937 16779 23995 16785
rect 23937 16776 23949 16779
rect 23716 16748 23949 16776
rect 23716 16736 23722 16748
rect 23937 16745 23949 16748
rect 23983 16745 23995 16779
rect 23937 16739 23995 16745
rect 24210 16736 24216 16788
rect 24268 16776 24274 16788
rect 24305 16779 24363 16785
rect 24305 16776 24317 16779
rect 24268 16748 24317 16776
rect 24268 16736 24274 16748
rect 24305 16745 24317 16748
rect 24351 16745 24363 16779
rect 24305 16739 24363 16745
rect 24663 16779 24721 16785
rect 24663 16745 24675 16779
rect 24709 16776 24721 16779
rect 24762 16776 24768 16788
rect 24709 16748 24768 16776
rect 24709 16745 24721 16748
rect 24663 16739 24721 16745
rect 13998 16668 14004 16720
rect 14056 16708 14062 16720
rect 14185 16711 14243 16717
rect 14185 16708 14197 16711
rect 14056 16680 14197 16708
rect 14056 16668 14062 16680
rect 14185 16677 14197 16680
rect 14231 16677 14243 16711
rect 14734 16708 14740 16720
rect 14695 16680 14740 16708
rect 14185 16671 14243 16677
rect 14734 16668 14740 16680
rect 14792 16668 14798 16720
rect 15838 16708 15844 16720
rect 15799 16680 15844 16708
rect 15838 16668 15844 16680
rect 15896 16668 15902 16720
rect 16850 16668 16856 16720
rect 16908 16708 16914 16720
rect 17313 16711 17371 16717
rect 17313 16708 17325 16711
rect 16908 16680 17325 16708
rect 16908 16668 16914 16680
rect 17313 16677 17325 16680
rect 17359 16677 17371 16711
rect 17313 16671 17371 16677
rect 18233 16711 18291 16717
rect 18233 16677 18245 16711
rect 18279 16708 18291 16711
rect 18506 16708 18512 16720
rect 18279 16680 18512 16708
rect 18279 16677 18291 16680
rect 18233 16671 18291 16677
rect 18506 16668 18512 16680
rect 18564 16668 18570 16720
rect 18877 16711 18935 16717
rect 18877 16677 18889 16711
rect 18923 16708 18935 16711
rect 19242 16708 19248 16720
rect 18923 16680 19248 16708
rect 18923 16677 18935 16680
rect 18877 16671 18935 16677
rect 19242 16668 19248 16680
rect 19300 16668 19306 16720
rect 19429 16711 19487 16717
rect 19429 16677 19441 16711
rect 19475 16708 19487 16711
rect 19518 16708 19524 16720
rect 19475 16680 19524 16708
rect 19475 16677 19487 16680
rect 19429 16671 19487 16677
rect 19518 16668 19524 16680
rect 19576 16668 19582 16720
rect 22088 16711 22146 16717
rect 22088 16677 22100 16711
rect 22134 16708 22146 16711
rect 22278 16708 22284 16720
rect 22134 16680 22284 16708
rect 22134 16677 22146 16680
rect 22088 16671 22146 16677
rect 22278 16668 22284 16680
rect 22336 16668 22342 16720
rect 13909 16643 13967 16649
rect 13909 16640 13921 16643
rect 13832 16612 13921 16640
rect 9582 16532 9588 16584
rect 9640 16532 9646 16584
rect 10502 16572 10508 16584
rect 10463 16544 10508 16572
rect 10502 16532 10508 16544
rect 10560 16532 10566 16584
rect 11054 16532 11060 16584
rect 11112 16532 11118 16584
rect 13170 16532 13176 16584
rect 13228 16572 13234 16584
rect 13832 16572 13860 16612
rect 13909 16609 13921 16612
rect 13955 16609 13967 16643
rect 13909 16603 13967 16609
rect 15105 16643 15163 16649
rect 15105 16609 15117 16643
rect 15151 16640 15163 16643
rect 15378 16640 15384 16652
rect 15151 16612 15384 16640
rect 15151 16609 15163 16612
rect 15105 16603 15163 16609
rect 15378 16600 15384 16612
rect 15436 16640 15442 16652
rect 15657 16643 15715 16649
rect 15657 16640 15669 16643
rect 15436 16612 15669 16640
rect 15436 16600 15442 16612
rect 15657 16609 15669 16612
rect 15703 16609 15715 16643
rect 15657 16603 15715 16609
rect 16485 16643 16543 16649
rect 16485 16609 16497 16643
rect 16531 16640 16543 16643
rect 16758 16640 16764 16652
rect 16531 16612 16764 16640
rect 16531 16609 16543 16612
rect 16485 16603 16543 16609
rect 16758 16600 16764 16612
rect 16816 16600 16822 16652
rect 17034 16640 17040 16652
rect 16995 16612 17040 16640
rect 17034 16600 17040 16612
rect 17092 16600 17098 16652
rect 18524 16640 18552 16668
rect 18969 16643 19027 16649
rect 18969 16640 18981 16643
rect 18524 16612 18981 16640
rect 18969 16609 18981 16612
rect 19015 16609 19027 16643
rect 18969 16603 19027 16609
rect 21821 16643 21879 16649
rect 21821 16609 21833 16643
rect 21867 16640 21879 16643
rect 21910 16640 21916 16652
rect 21867 16612 21916 16640
rect 21867 16609 21879 16612
rect 21821 16603 21879 16609
rect 21910 16600 21916 16612
rect 21968 16600 21974 16652
rect 24320 16640 24348 16739
rect 24762 16736 24768 16748
rect 24820 16736 24826 16788
rect 24854 16668 24860 16720
rect 24912 16708 24918 16720
rect 25133 16711 25191 16717
rect 25133 16708 25145 16711
rect 24912 16680 25145 16708
rect 24912 16668 24918 16680
rect 25133 16677 25145 16680
rect 25179 16677 25191 16711
rect 25133 16671 25191 16677
rect 25225 16643 25283 16649
rect 25225 16640 25237 16643
rect 24320 16612 25237 16640
rect 25225 16609 25237 16612
rect 25271 16640 25283 16643
rect 25406 16640 25412 16652
rect 25271 16612 25412 16640
rect 25271 16609 25283 16612
rect 25225 16603 25283 16609
rect 25406 16600 25412 16612
rect 25464 16600 25470 16652
rect 15930 16572 15936 16584
rect 13228 16544 13860 16572
rect 15891 16544 15936 16572
rect 13228 16532 13234 16544
rect 15930 16532 15936 16544
rect 15988 16532 15994 16584
rect 18598 16532 18604 16584
rect 18656 16572 18662 16584
rect 18785 16575 18843 16581
rect 18785 16572 18797 16575
rect 18656 16544 18797 16572
rect 18656 16532 18662 16544
rect 18785 16541 18797 16544
rect 18831 16541 18843 16575
rect 18785 16535 18843 16541
rect 19978 16532 19984 16584
rect 20036 16572 20042 16584
rect 20438 16572 20444 16584
rect 20036 16544 20444 16572
rect 20036 16532 20042 16544
rect 20438 16532 20444 16544
rect 20496 16532 20502 16584
rect 25133 16575 25191 16581
rect 25133 16541 25145 16575
rect 25179 16572 25191 16575
rect 25314 16572 25320 16584
rect 25179 16544 25320 16572
rect 25179 16541 25191 16544
rect 25133 16535 25191 16541
rect 25314 16532 25320 16544
rect 25372 16532 25378 16584
rect 20165 16507 20223 16513
rect 20165 16473 20177 16507
rect 20211 16504 20223 16507
rect 20622 16504 20628 16516
rect 20211 16476 20628 16504
rect 20211 16473 20223 16476
rect 20165 16467 20223 16473
rect 20622 16464 20628 16476
rect 20680 16464 20686 16516
rect 13725 16439 13783 16445
rect 13725 16405 13737 16439
rect 13771 16436 13783 16439
rect 13906 16436 13912 16448
rect 13771 16408 13912 16436
rect 13771 16405 13783 16408
rect 13725 16399 13783 16405
rect 13906 16396 13912 16408
rect 13964 16396 13970 16448
rect 17865 16439 17923 16445
rect 17865 16405 17877 16439
rect 17911 16436 17923 16439
rect 18966 16436 18972 16448
rect 17911 16408 18972 16436
rect 17911 16405 17923 16408
rect 17865 16399 17923 16405
rect 18966 16396 18972 16408
rect 19024 16396 19030 16448
rect 20438 16436 20444 16448
rect 20399 16408 20444 16436
rect 20438 16396 20444 16408
rect 20496 16396 20502 16448
rect 21266 16396 21272 16448
rect 21324 16436 21330 16448
rect 21453 16439 21511 16445
rect 21453 16436 21465 16439
rect 21324 16408 21465 16436
rect 21324 16396 21330 16408
rect 21453 16405 21465 16408
rect 21499 16405 21511 16439
rect 21453 16399 21511 16405
rect 23106 16396 23112 16448
rect 23164 16436 23170 16448
rect 23201 16439 23259 16445
rect 23201 16436 23213 16439
rect 23164 16408 23213 16436
rect 23164 16396 23170 16408
rect 23201 16405 23213 16408
rect 23247 16405 23259 16439
rect 23201 16399 23259 16405
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 9582 16232 9588 16244
rect 9543 16204 9588 16232
rect 9582 16192 9588 16204
rect 9640 16192 9646 16244
rect 9953 16235 10011 16241
rect 9953 16201 9965 16235
rect 9999 16232 10011 16235
rect 10502 16232 10508 16244
rect 9999 16204 10508 16232
rect 9999 16201 10011 16204
rect 9953 16195 10011 16201
rect 10502 16192 10508 16204
rect 10560 16192 10566 16244
rect 10873 16235 10931 16241
rect 10873 16201 10885 16235
rect 10919 16232 10931 16235
rect 10962 16232 10968 16244
rect 10919 16204 10968 16232
rect 10919 16201 10931 16204
rect 10873 16195 10931 16201
rect 10962 16192 10968 16204
rect 11020 16192 11026 16244
rect 12713 16235 12771 16241
rect 12713 16201 12725 16235
rect 12759 16232 12771 16235
rect 12986 16232 12992 16244
rect 12759 16204 12992 16232
rect 12759 16201 12771 16204
rect 12713 16195 12771 16201
rect 12986 16192 12992 16204
rect 13044 16192 13050 16244
rect 13170 16232 13176 16244
rect 13131 16204 13176 16232
rect 13170 16192 13176 16204
rect 13228 16192 13234 16244
rect 14826 16232 14832 16244
rect 13648 16204 14832 16232
rect 10321 16099 10379 16105
rect 10321 16065 10333 16099
rect 10367 16096 10379 16099
rect 11425 16099 11483 16105
rect 11425 16096 11437 16099
rect 10367 16068 11437 16096
rect 10367 16065 10379 16068
rect 10321 16059 10379 16065
rect 11425 16065 11437 16068
rect 11471 16096 11483 16099
rect 11606 16096 11612 16108
rect 11471 16068 11612 16096
rect 11471 16065 11483 16068
rect 11425 16059 11483 16065
rect 11606 16056 11612 16068
rect 11664 16096 11670 16108
rect 12253 16099 12311 16105
rect 12253 16096 12265 16099
rect 11664 16068 12265 16096
rect 11664 16056 11670 16068
rect 12253 16065 12265 16068
rect 12299 16096 12311 16099
rect 12434 16096 12440 16108
rect 12299 16068 12440 16096
rect 12299 16065 12311 16068
rect 12253 16059 12311 16065
rect 12434 16056 12440 16068
rect 12492 16096 12498 16108
rect 13648 16096 13676 16204
rect 14826 16192 14832 16204
rect 14884 16232 14890 16244
rect 15013 16235 15071 16241
rect 15013 16232 15025 16235
rect 14884 16204 15025 16232
rect 14884 16192 14890 16204
rect 15013 16201 15025 16204
rect 15059 16201 15071 16235
rect 17494 16232 17500 16244
rect 17455 16204 17500 16232
rect 15013 16195 15071 16201
rect 17494 16192 17500 16204
rect 17552 16192 17558 16244
rect 18414 16232 18420 16244
rect 18375 16204 18420 16232
rect 18414 16192 18420 16204
rect 18472 16192 18478 16244
rect 18598 16192 18604 16244
rect 18656 16232 18662 16244
rect 19705 16235 19763 16241
rect 19705 16232 19717 16235
rect 18656 16204 19717 16232
rect 18656 16192 18662 16204
rect 19705 16201 19717 16204
rect 19751 16201 19763 16235
rect 19705 16195 19763 16201
rect 22094 16192 22100 16244
rect 22152 16232 22158 16244
rect 22465 16235 22523 16241
rect 22465 16232 22477 16235
rect 22152 16204 22477 16232
rect 22152 16192 22158 16204
rect 22465 16201 22477 16204
rect 22511 16232 22523 16235
rect 23290 16232 23296 16244
rect 22511 16204 23296 16232
rect 22511 16201 22523 16204
rect 22465 16195 22523 16201
rect 23290 16192 23296 16204
rect 23348 16192 23354 16244
rect 23474 16232 23480 16244
rect 23435 16204 23480 16232
rect 23474 16192 23480 16204
rect 23532 16192 23538 16244
rect 25406 16232 25412 16244
rect 25367 16204 25412 16232
rect 25406 16192 25412 16204
rect 25464 16232 25470 16244
rect 25961 16235 26019 16241
rect 25961 16232 25973 16235
rect 25464 16204 25973 16232
rect 25464 16192 25470 16204
rect 25961 16201 25973 16204
rect 26007 16201 26019 16235
rect 25961 16195 26019 16201
rect 15102 16124 15108 16176
rect 15160 16164 15166 16176
rect 15838 16164 15844 16176
rect 15160 16136 15844 16164
rect 15160 16124 15166 16136
rect 15838 16124 15844 16136
rect 15896 16164 15902 16176
rect 16485 16167 16543 16173
rect 16485 16164 16497 16167
rect 15896 16136 16497 16164
rect 15896 16124 15902 16136
rect 16485 16133 16497 16136
rect 16531 16133 16543 16167
rect 16485 16127 16543 16133
rect 19334 16124 19340 16176
rect 19392 16164 19398 16176
rect 19981 16167 20039 16173
rect 19981 16164 19993 16167
rect 19392 16136 19993 16164
rect 19392 16124 19398 16136
rect 19981 16133 19993 16136
rect 20027 16133 20039 16167
rect 21542 16164 21548 16176
rect 21503 16136 21548 16164
rect 19981 16127 20039 16133
rect 21542 16124 21548 16136
rect 21600 16124 21606 16176
rect 12492 16068 13676 16096
rect 20993 16099 21051 16105
rect 12492 16056 12498 16068
rect 20993 16065 21005 16099
rect 21039 16096 21051 16099
rect 21174 16096 21180 16108
rect 21039 16068 21180 16096
rect 21039 16065 21051 16068
rect 20993 16059 21051 16065
rect 21174 16056 21180 16068
rect 21232 16096 21238 16108
rect 22097 16099 22155 16105
rect 22097 16096 22109 16099
rect 21232 16068 22109 16096
rect 21232 16056 21238 16068
rect 22097 16065 22109 16068
rect 22143 16065 22155 16099
rect 23492 16096 23520 16192
rect 23492 16068 24164 16096
rect 22097 16059 22155 16065
rect 13906 16037 13912 16040
rect 13633 16031 13691 16037
rect 13633 15997 13645 16031
rect 13679 15997 13691 16031
rect 13900 16028 13912 16037
rect 13867 16000 13912 16028
rect 13633 15991 13691 15997
rect 13900 15991 13912 16000
rect 13964 16028 13970 16040
rect 15565 16031 15623 16037
rect 15565 16028 15577 16031
rect 13964 16000 15577 16028
rect 11146 15960 11152 15972
rect 11059 15932 11152 15960
rect 11146 15920 11152 15932
rect 11204 15920 11210 15972
rect 10686 15892 10692 15904
rect 10647 15864 10692 15892
rect 10686 15852 10692 15864
rect 10744 15892 10750 15904
rect 11164 15892 11192 15920
rect 10744 15864 11192 15892
rect 11333 15895 11391 15901
rect 10744 15852 10750 15864
rect 11333 15861 11345 15895
rect 11379 15892 11391 15895
rect 11422 15892 11428 15904
rect 11379 15864 11428 15892
rect 11379 15861 11391 15864
rect 11333 15855 11391 15861
rect 11422 15852 11428 15864
rect 11480 15852 11486 15904
rect 11514 15852 11520 15904
rect 11572 15892 11578 15904
rect 11885 15895 11943 15901
rect 11885 15892 11897 15895
rect 11572 15864 11897 15892
rect 11572 15852 11578 15864
rect 11885 15861 11897 15864
rect 11931 15892 11943 15895
rect 13541 15895 13599 15901
rect 13541 15892 13553 15895
rect 11931 15864 13553 15892
rect 11931 15861 11943 15864
rect 11885 15855 11943 15861
rect 13541 15861 13553 15864
rect 13587 15892 13599 15895
rect 13648 15892 13676 15991
rect 13906 15988 13912 15991
rect 13964 15988 13970 16000
rect 15565 15997 15577 16000
rect 15611 16028 15623 16031
rect 15930 16028 15936 16040
rect 15611 16000 15936 16028
rect 15611 15997 15623 16000
rect 15565 15991 15623 15997
rect 15930 15988 15936 16000
rect 15988 15988 15994 16040
rect 18966 16028 18972 16040
rect 18927 16000 18972 16028
rect 18966 15988 18972 16000
rect 19024 15988 19030 16040
rect 21266 15988 21272 16040
rect 21324 16028 21330 16040
rect 21324 16000 22048 16028
rect 21324 15988 21330 16000
rect 16574 15920 16580 15972
rect 16632 15960 16638 15972
rect 16761 15963 16819 15969
rect 16761 15960 16773 15963
rect 16632 15932 16773 15960
rect 16632 15920 16638 15932
rect 16761 15929 16773 15932
rect 16807 15929 16819 15963
rect 16942 15960 16948 15972
rect 16903 15932 16948 15960
rect 16761 15923 16819 15929
rect 16942 15920 16948 15932
rect 17000 15920 17006 15972
rect 17037 15963 17095 15969
rect 17037 15929 17049 15963
rect 17083 15960 17095 15963
rect 17678 15960 17684 15972
rect 17083 15932 17684 15960
rect 17083 15929 17095 15932
rect 17037 15923 17095 15929
rect 14826 15892 14832 15904
rect 13587 15864 14832 15892
rect 13587 15861 13599 15864
rect 13541 15855 13599 15861
rect 14826 15852 14832 15864
rect 14884 15852 14890 15904
rect 16301 15895 16359 15901
rect 16301 15861 16313 15895
rect 16347 15892 16359 15895
rect 17052 15892 17080 15923
rect 17678 15920 17684 15932
rect 17736 15920 17742 15972
rect 17865 15963 17923 15969
rect 17865 15929 17877 15963
rect 17911 15960 17923 15963
rect 18690 15960 18696 15972
rect 17911 15932 18696 15960
rect 17911 15929 17923 15932
rect 17865 15923 17923 15929
rect 18690 15920 18696 15932
rect 18748 15920 18754 15972
rect 20257 15963 20315 15969
rect 20257 15929 20269 15963
rect 20303 15960 20315 15963
rect 20346 15960 20352 15972
rect 20303 15932 20352 15960
rect 20303 15929 20315 15932
rect 20257 15923 20315 15929
rect 20346 15920 20352 15932
rect 20404 15920 20410 15972
rect 20530 15960 20536 15972
rect 20491 15932 20536 15960
rect 20530 15920 20536 15932
rect 20588 15920 20594 15972
rect 21361 15963 21419 15969
rect 21361 15929 21373 15963
rect 21407 15960 21419 15963
rect 21818 15960 21824 15972
rect 21407 15932 21824 15960
rect 21407 15929 21419 15932
rect 21361 15923 21419 15929
rect 21818 15920 21824 15932
rect 21876 15920 21882 15972
rect 22020 15969 22048 16000
rect 23290 15988 23296 16040
rect 23348 16028 23354 16040
rect 24026 16028 24032 16040
rect 23348 16000 24032 16028
rect 23348 15988 23354 16000
rect 24026 15988 24032 16000
rect 24084 15988 24090 16040
rect 24136 16028 24164 16068
rect 24285 16031 24343 16037
rect 24285 16028 24297 16031
rect 24136 16000 24297 16028
rect 24285 15997 24297 16000
rect 24331 16028 24343 16031
rect 24670 16028 24676 16040
rect 24331 16000 24676 16028
rect 24331 15997 24343 16000
rect 24285 15991 24343 15997
rect 24670 15988 24676 16000
rect 24728 15988 24734 16040
rect 22005 15963 22063 15969
rect 22005 15929 22017 15963
rect 22051 15929 22063 15963
rect 22005 15923 22063 15929
rect 16347 15864 17080 15892
rect 18877 15895 18935 15901
rect 16347 15861 16359 15864
rect 16301 15855 16359 15861
rect 18877 15861 18889 15895
rect 18923 15892 18935 15895
rect 19426 15892 19432 15904
rect 18923 15864 19432 15892
rect 18923 15861 18935 15864
rect 18877 15855 18935 15861
rect 19426 15852 19432 15864
rect 19484 15852 19490 15904
rect 20438 15892 20444 15904
rect 20399 15864 20444 15892
rect 20438 15852 20444 15864
rect 20496 15852 20502 15904
rect 23937 15895 23995 15901
rect 23937 15861 23949 15895
rect 23983 15892 23995 15895
rect 24670 15892 24676 15904
rect 23983 15864 24676 15892
rect 23983 15861 23995 15864
rect 23937 15855 23995 15861
rect 24670 15852 24676 15864
rect 24728 15852 24734 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 9953 15691 10011 15697
rect 9953 15657 9965 15691
rect 9999 15688 10011 15691
rect 10134 15688 10140 15700
rect 9999 15660 10140 15688
rect 9999 15657 10011 15660
rect 9953 15651 10011 15657
rect 10134 15648 10140 15660
rect 10192 15648 10198 15700
rect 13814 15648 13820 15700
rect 13872 15688 13878 15700
rect 13909 15691 13967 15697
rect 13909 15688 13921 15691
rect 13872 15660 13921 15688
rect 13872 15648 13878 15660
rect 13909 15657 13921 15660
rect 13955 15657 13967 15691
rect 15102 15688 15108 15700
rect 15063 15660 15108 15688
rect 13909 15651 13967 15657
rect 15102 15648 15108 15660
rect 15160 15648 15166 15700
rect 16574 15648 16580 15700
rect 16632 15688 16638 15700
rect 17589 15691 17647 15697
rect 17589 15688 17601 15691
rect 16632 15660 17601 15688
rect 16632 15648 16638 15660
rect 17589 15657 17601 15660
rect 17635 15657 17647 15691
rect 17589 15651 17647 15657
rect 17678 15648 17684 15700
rect 17736 15688 17742 15700
rect 19153 15691 19211 15697
rect 19153 15688 19165 15691
rect 17736 15660 19165 15688
rect 17736 15648 17742 15660
rect 19153 15657 19165 15660
rect 19199 15657 19211 15691
rect 19153 15651 19211 15657
rect 23017 15691 23075 15697
rect 23017 15657 23029 15691
rect 23063 15688 23075 15691
rect 23382 15688 23388 15700
rect 23063 15660 23388 15688
rect 23063 15657 23075 15660
rect 23017 15651 23075 15657
rect 23382 15648 23388 15660
rect 23440 15648 23446 15700
rect 24026 15688 24032 15700
rect 23987 15660 24032 15688
rect 24026 15648 24032 15660
rect 24084 15648 24090 15700
rect 25406 15688 25412 15700
rect 24688 15660 25412 15688
rect 12066 15580 12072 15632
rect 12124 15620 12130 15632
rect 12299 15623 12357 15629
rect 12299 15620 12311 15623
rect 12124 15592 12311 15620
rect 12124 15580 12130 15592
rect 12299 15589 12311 15592
rect 12345 15589 12357 15623
rect 12299 15583 12357 15589
rect 14182 15580 14188 15632
rect 14240 15620 14246 15632
rect 14734 15620 14740 15632
rect 14240 15592 14740 15620
rect 14240 15580 14246 15592
rect 14734 15580 14740 15592
rect 14792 15580 14798 15632
rect 18040 15623 18098 15629
rect 18040 15589 18052 15623
rect 18086 15620 18098 15623
rect 18138 15620 18144 15632
rect 18086 15592 18144 15620
rect 18086 15589 18098 15592
rect 18040 15583 18098 15589
rect 18138 15580 18144 15592
rect 18196 15580 18202 15632
rect 18322 15580 18328 15632
rect 18380 15620 18386 15632
rect 18874 15620 18880 15632
rect 18380 15592 18880 15620
rect 18380 15580 18386 15592
rect 18874 15580 18880 15592
rect 18932 15580 18938 15632
rect 20806 15580 20812 15632
rect 20864 15620 20870 15632
rect 21453 15623 21511 15629
rect 21453 15620 21465 15623
rect 20864 15592 21465 15620
rect 20864 15580 20870 15592
rect 21453 15589 21465 15592
rect 21499 15589 21511 15623
rect 21453 15583 21511 15589
rect 21542 15580 21548 15632
rect 21600 15580 21606 15632
rect 21726 15580 21732 15632
rect 21784 15620 21790 15632
rect 21913 15623 21971 15629
rect 21913 15620 21925 15623
rect 21784 15592 21925 15620
rect 21784 15580 21790 15592
rect 21913 15589 21925 15592
rect 21959 15589 21971 15623
rect 22830 15620 22836 15632
rect 22791 15592 22836 15620
rect 21913 15583 21971 15589
rect 22830 15580 22836 15592
rect 22888 15580 22894 15632
rect 24688 15629 24716 15660
rect 25406 15648 25412 15660
rect 25464 15648 25470 15700
rect 24673 15623 24731 15629
rect 24673 15589 24685 15623
rect 24719 15589 24731 15623
rect 24673 15583 24731 15589
rect 24762 15580 24768 15632
rect 24820 15620 24826 15632
rect 24857 15623 24915 15629
rect 24857 15620 24869 15623
rect 24820 15592 24869 15620
rect 24820 15580 24826 15592
rect 24857 15589 24869 15592
rect 24903 15589 24915 15623
rect 24857 15583 24915 15589
rect 12158 15552 12164 15564
rect 12119 15524 12164 15552
rect 12158 15512 12164 15524
rect 12216 15512 12222 15564
rect 12434 15512 12440 15564
rect 12492 15552 12498 15564
rect 15562 15561 15568 15564
rect 15556 15552 15568 15561
rect 12492 15524 12537 15552
rect 15523 15524 15568 15552
rect 12492 15512 12498 15524
rect 15556 15515 15568 15524
rect 15562 15512 15568 15515
rect 15620 15512 15626 15564
rect 21269 15555 21327 15561
rect 21269 15521 21281 15555
rect 21315 15552 21327 15555
rect 21560 15552 21588 15580
rect 22281 15555 22339 15561
rect 22281 15552 22293 15555
rect 21315 15524 22293 15552
rect 21315 15521 21327 15524
rect 21269 15515 21327 15521
rect 22281 15521 22293 15524
rect 22327 15521 22339 15555
rect 22281 15515 22339 15521
rect 11422 15484 11428 15496
rect 10796 15456 11428 15484
rect 10796 15428 10824 15456
rect 11422 15444 11428 15456
rect 11480 15444 11486 15496
rect 13814 15484 13820 15496
rect 13775 15456 13820 15484
rect 13814 15444 13820 15456
rect 13872 15444 13878 15496
rect 14001 15487 14059 15493
rect 14001 15453 14013 15487
rect 14047 15484 14059 15487
rect 14182 15484 14188 15496
rect 14047 15456 14188 15484
rect 14047 15453 14059 15456
rect 14001 15447 14059 15453
rect 14182 15444 14188 15456
rect 14240 15444 14246 15496
rect 14826 15444 14832 15496
rect 14884 15484 14890 15496
rect 15289 15487 15347 15493
rect 15289 15484 15301 15487
rect 14884 15456 15301 15484
rect 14884 15444 14890 15456
rect 15289 15453 15301 15456
rect 15335 15453 15347 15487
rect 17770 15484 17776 15496
rect 17731 15456 17776 15484
rect 15289 15447 15347 15453
rect 17770 15444 17776 15456
rect 17828 15444 17834 15496
rect 20349 15487 20407 15493
rect 20349 15453 20361 15487
rect 20395 15484 20407 15487
rect 20530 15484 20536 15496
rect 20395 15456 20536 15484
rect 20395 15453 20407 15456
rect 20349 15447 20407 15453
rect 20530 15444 20536 15456
rect 20588 15484 20594 15496
rect 20717 15487 20775 15493
rect 20717 15484 20729 15487
rect 20588 15456 20729 15484
rect 20588 15444 20594 15456
rect 20717 15453 20729 15456
rect 20763 15484 20775 15487
rect 21545 15487 21603 15493
rect 21545 15484 21557 15487
rect 20763 15456 21557 15484
rect 20763 15453 20775 15456
rect 20717 15447 20775 15453
rect 21545 15453 21557 15456
rect 21591 15484 21603 15487
rect 22002 15484 22008 15496
rect 21591 15456 22008 15484
rect 21591 15453 21603 15456
rect 21545 15447 21603 15453
rect 22002 15444 22008 15456
rect 22060 15444 22066 15496
rect 23106 15484 23112 15496
rect 23067 15456 23112 15484
rect 23106 15444 23112 15456
rect 23164 15444 23170 15496
rect 24854 15444 24860 15496
rect 24912 15484 24918 15496
rect 24949 15487 25007 15493
rect 24949 15484 24961 15487
rect 24912 15456 24961 15484
rect 24912 15444 24918 15456
rect 24949 15453 24961 15456
rect 24995 15453 25007 15487
rect 24949 15447 25007 15453
rect 10778 15416 10784 15428
rect 10739 15388 10784 15416
rect 10778 15376 10784 15388
rect 10836 15376 10842 15428
rect 11054 15376 11060 15428
rect 11112 15416 11118 15428
rect 11885 15419 11943 15425
rect 11885 15416 11897 15419
rect 11112 15388 11897 15416
rect 11112 15376 11118 15388
rect 11885 15385 11897 15388
rect 11931 15385 11943 15419
rect 11885 15379 11943 15385
rect 13265 15419 13323 15425
rect 13265 15385 13277 15419
rect 13311 15416 13323 15419
rect 13630 15416 13636 15428
rect 13311 15388 13636 15416
rect 13311 15385 13323 15388
rect 13265 15379 13323 15385
rect 13630 15376 13636 15388
rect 13688 15376 13694 15428
rect 22186 15376 22192 15428
rect 22244 15416 22250 15428
rect 22557 15419 22615 15425
rect 22557 15416 22569 15419
rect 22244 15388 22569 15416
rect 22244 15376 22250 15388
rect 22557 15385 22569 15388
rect 22603 15385 22615 15419
rect 22557 15379 22615 15385
rect 13446 15348 13452 15360
rect 13407 15320 13452 15348
rect 13446 15308 13452 15320
rect 13504 15308 13510 15360
rect 14090 15308 14096 15360
rect 14148 15348 14154 15360
rect 14369 15351 14427 15357
rect 14369 15348 14381 15351
rect 14148 15320 14381 15348
rect 14148 15308 14154 15320
rect 14369 15317 14381 15320
rect 14415 15317 14427 15351
rect 14369 15311 14427 15317
rect 15930 15308 15936 15360
rect 15988 15348 15994 15360
rect 16669 15351 16727 15357
rect 16669 15348 16681 15351
rect 15988 15320 16681 15348
rect 15988 15308 15994 15320
rect 16669 15317 16681 15320
rect 16715 15317 16727 15351
rect 16669 15311 16727 15317
rect 17034 15308 17040 15360
rect 17092 15348 17098 15360
rect 17313 15351 17371 15357
rect 17313 15348 17325 15351
rect 17092 15320 17325 15348
rect 17092 15308 17098 15320
rect 17313 15317 17325 15320
rect 17359 15348 17371 15351
rect 18046 15348 18052 15360
rect 17359 15320 18052 15348
rect 17359 15317 17371 15320
rect 17313 15311 17371 15317
rect 18046 15308 18052 15320
rect 18104 15308 18110 15360
rect 19981 15351 20039 15357
rect 19981 15317 19993 15351
rect 20027 15348 20039 15351
rect 20346 15348 20352 15360
rect 20027 15320 20352 15348
rect 20027 15317 20039 15320
rect 19981 15311 20039 15317
rect 20346 15308 20352 15320
rect 20404 15308 20410 15360
rect 20714 15308 20720 15360
rect 20772 15348 20778 15360
rect 20993 15351 21051 15357
rect 20993 15348 21005 15351
rect 20772 15320 21005 15348
rect 20772 15308 20778 15320
rect 20993 15317 21005 15320
rect 21039 15317 21051 15351
rect 20993 15311 21051 15317
rect 23753 15351 23811 15357
rect 23753 15317 23765 15351
rect 23799 15348 23811 15351
rect 23934 15348 23940 15360
rect 23799 15320 23940 15348
rect 23799 15317 23811 15320
rect 23753 15311 23811 15317
rect 23934 15308 23940 15320
rect 23992 15308 23998 15360
rect 24210 15308 24216 15360
rect 24268 15348 24274 15360
rect 24397 15351 24455 15357
rect 24397 15348 24409 15351
rect 24268 15320 24409 15348
rect 24268 15308 24274 15320
rect 24397 15317 24409 15320
rect 24443 15317 24455 15351
rect 24397 15311 24455 15317
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 11517 15147 11575 15153
rect 11517 15113 11529 15147
rect 11563 15144 11575 15147
rect 11606 15144 11612 15156
rect 11563 15116 11612 15144
rect 11563 15113 11575 15116
rect 11517 15107 11575 15113
rect 11606 15104 11612 15116
rect 11664 15104 11670 15156
rect 11885 15147 11943 15153
rect 11885 15113 11897 15147
rect 11931 15144 11943 15147
rect 12158 15144 12164 15156
rect 11931 15116 12164 15144
rect 11931 15113 11943 15116
rect 11885 15107 11943 15113
rect 12158 15104 12164 15116
rect 12216 15104 12222 15156
rect 12802 15104 12808 15156
rect 12860 15144 12866 15156
rect 13081 15147 13139 15153
rect 13081 15144 13093 15147
rect 12860 15116 13093 15144
rect 12860 15104 12866 15116
rect 13081 15113 13093 15116
rect 13127 15144 13139 15147
rect 13722 15144 13728 15156
rect 13127 15116 13728 15144
rect 13127 15113 13139 15116
rect 13081 15107 13139 15113
rect 13722 15104 13728 15116
rect 13780 15104 13786 15156
rect 15378 15144 15384 15156
rect 15339 15116 15384 15144
rect 15378 15104 15384 15116
rect 15436 15104 15442 15156
rect 15562 15104 15568 15156
rect 15620 15144 15626 15156
rect 16761 15147 16819 15153
rect 16761 15144 16773 15147
rect 15620 15116 16773 15144
rect 15620 15104 15626 15116
rect 12710 15036 12716 15088
rect 12768 15076 12774 15088
rect 13633 15079 13691 15085
rect 13633 15076 13645 15079
rect 12768 15048 13645 15076
rect 12768 15036 12774 15048
rect 13633 15045 13645 15048
rect 13679 15045 13691 15079
rect 13633 15039 13691 15045
rect 12066 14968 12072 15020
rect 12124 15008 12130 15020
rect 15948 15017 15976 15116
rect 16761 15113 16773 15116
rect 16807 15144 16819 15147
rect 17678 15144 17684 15156
rect 16807 15116 17684 15144
rect 16807 15113 16819 15116
rect 16761 15107 16819 15113
rect 17678 15104 17684 15116
rect 17736 15104 17742 15156
rect 18046 15104 18052 15156
rect 18104 15144 18110 15156
rect 18785 15147 18843 15153
rect 18785 15144 18797 15147
rect 18104 15116 18797 15144
rect 18104 15104 18110 15116
rect 18785 15113 18797 15116
rect 18831 15113 18843 15147
rect 22830 15144 22836 15156
rect 22791 15116 22836 15144
rect 18785 15107 18843 15113
rect 22830 15104 22836 15116
rect 22888 15104 22894 15156
rect 23477 15147 23535 15153
rect 23477 15113 23489 15147
rect 23523 15144 23535 15147
rect 24026 15144 24032 15156
rect 23523 15116 24032 15144
rect 23523 15113 23535 15116
rect 23477 15107 23535 15113
rect 24026 15104 24032 15116
rect 24084 15144 24090 15156
rect 24762 15144 24768 15156
rect 24084 15116 24768 15144
rect 24084 15104 24090 15116
rect 24762 15104 24768 15116
rect 24820 15104 24826 15156
rect 25133 15147 25191 15153
rect 25133 15113 25145 15147
rect 25179 15144 25191 15147
rect 25406 15144 25412 15156
rect 25179 15116 25412 15144
rect 25179 15113 25191 15116
rect 25133 15107 25191 15113
rect 25406 15104 25412 15116
rect 25464 15104 25470 15156
rect 17126 15036 17132 15088
rect 17184 15076 17190 15088
rect 17405 15079 17463 15085
rect 17405 15076 17417 15079
rect 17184 15048 17417 15076
rect 17184 15036 17190 15048
rect 17405 15045 17417 15048
rect 17451 15076 17463 15079
rect 18138 15076 18144 15088
rect 17451 15048 18144 15076
rect 17451 15045 17463 15048
rect 17405 15039 17463 15045
rect 18138 15036 18144 15048
rect 18196 15036 18202 15088
rect 22554 15076 22560 15088
rect 22467 15048 22560 15076
rect 22554 15036 22560 15048
rect 22612 15076 22618 15088
rect 23382 15076 23388 15088
rect 22612 15048 23388 15076
rect 22612 15036 22618 15048
rect 23382 15036 23388 15048
rect 23440 15036 23446 15088
rect 23750 15076 23756 15088
rect 23711 15048 23756 15076
rect 23750 15036 23756 15048
rect 23808 15036 23814 15088
rect 12161 15011 12219 15017
rect 12161 15008 12173 15011
rect 12124 14980 12173 15008
rect 12124 14968 12130 14980
rect 12161 14977 12173 14980
rect 12207 14977 12219 15011
rect 12161 14971 12219 14977
rect 15933 15011 15991 15017
rect 15933 14977 15945 15011
rect 15979 14977 15991 15011
rect 19242 15008 19248 15020
rect 19203 14980 19248 15008
rect 15933 14971 15991 14977
rect 19242 14968 19248 14980
rect 19300 14968 19306 15020
rect 19797 15011 19855 15017
rect 19797 14977 19809 15011
rect 19843 15008 19855 15011
rect 24210 15008 24216 15020
rect 19843 14980 20392 15008
rect 24171 14980 24216 15008
rect 19843 14977 19855 14980
rect 19797 14971 19855 14977
rect 12434 14900 12440 14952
rect 12492 14940 12498 14952
rect 12713 14943 12771 14949
rect 12713 14940 12725 14943
rect 12492 14912 12725 14940
rect 12492 14900 12498 14912
rect 12713 14909 12725 14912
rect 12759 14940 12771 14943
rect 13354 14940 13360 14952
rect 12759 14912 13360 14940
rect 12759 14909 12771 14912
rect 12713 14903 12771 14909
rect 13354 14900 13360 14912
rect 13412 14900 13418 14952
rect 13814 14900 13820 14952
rect 13872 14940 13878 14952
rect 13909 14943 13967 14949
rect 13909 14940 13921 14943
rect 13872 14912 13921 14940
rect 13872 14900 13878 14912
rect 13909 14909 13921 14912
rect 13955 14909 13967 14943
rect 13909 14903 13967 14909
rect 15657 14943 15715 14949
rect 15657 14909 15669 14943
rect 15703 14940 15715 14943
rect 20254 14940 20260 14952
rect 15703 14912 16436 14940
rect 20215 14912 20260 14940
rect 15703 14909 15715 14912
rect 15657 14903 15715 14909
rect 14090 14872 14096 14884
rect 14051 14844 14096 14872
rect 14090 14832 14096 14844
rect 14148 14832 14154 14884
rect 14182 14832 14188 14884
rect 14240 14872 14246 14884
rect 15197 14875 15255 14881
rect 14240 14844 14285 14872
rect 14240 14832 14246 14844
rect 15197 14841 15209 14875
rect 15243 14872 15255 14875
rect 15841 14875 15899 14881
rect 15841 14872 15853 14875
rect 15243 14844 15853 14872
rect 15243 14841 15255 14844
rect 15197 14835 15255 14841
rect 15841 14841 15853 14844
rect 15887 14872 15899 14875
rect 15930 14872 15936 14884
rect 15887 14844 15936 14872
rect 15887 14841 15899 14844
rect 15841 14835 15899 14841
rect 15930 14832 15936 14844
rect 15988 14832 15994 14884
rect 16408 14881 16436 14912
rect 20254 14900 20260 14912
rect 20312 14900 20318 14952
rect 20364 14940 20392 14980
rect 24210 14968 24216 14980
rect 24268 14968 24274 15020
rect 20530 14949 20536 14952
rect 20524 14940 20536 14949
rect 20364 14912 20536 14940
rect 20524 14903 20536 14912
rect 20530 14900 20536 14903
rect 20588 14900 20594 14952
rect 23934 14900 23940 14952
rect 23992 14940 23998 14952
rect 24305 14943 24363 14949
rect 24305 14940 24317 14943
rect 23992 14912 24317 14940
rect 23992 14900 23998 14912
rect 24305 14909 24317 14912
rect 24351 14909 24363 14943
rect 24305 14903 24363 14909
rect 16393 14875 16451 14881
rect 16393 14841 16405 14875
rect 16439 14872 16451 14875
rect 16853 14875 16911 14881
rect 16853 14872 16865 14875
rect 16439 14844 16865 14872
rect 16439 14841 16451 14844
rect 16393 14835 16451 14841
rect 16853 14841 16865 14844
rect 16899 14841 16911 14875
rect 18598 14872 18604 14884
rect 18511 14844 18604 14872
rect 16853 14835 16911 14841
rect 18598 14832 18604 14844
rect 18656 14872 18662 14884
rect 19337 14875 19395 14881
rect 19337 14872 19349 14875
rect 18656 14844 19349 14872
rect 18656 14832 18662 14844
rect 19337 14841 19349 14844
rect 19383 14872 19395 14875
rect 19383 14844 21680 14872
rect 19383 14841 19395 14844
rect 19337 14835 19395 14841
rect 13262 14764 13268 14816
rect 13320 14804 13326 14816
rect 13357 14807 13415 14813
rect 13357 14804 13369 14807
rect 13320 14776 13369 14804
rect 13320 14764 13326 14776
rect 13357 14773 13369 14776
rect 13403 14773 13415 14807
rect 14826 14804 14832 14816
rect 14787 14776 14832 14804
rect 13357 14767 13415 14773
rect 14826 14764 14832 14776
rect 14884 14764 14890 14816
rect 17770 14804 17776 14816
rect 17731 14776 17776 14804
rect 17770 14764 17776 14776
rect 17828 14764 17834 14816
rect 19242 14804 19248 14816
rect 19203 14776 19248 14804
rect 19242 14764 19248 14776
rect 19300 14764 19306 14816
rect 20165 14807 20223 14813
rect 20165 14773 20177 14807
rect 20211 14804 20223 14807
rect 20254 14804 20260 14816
rect 20211 14776 20260 14804
rect 20211 14773 20223 14776
rect 20165 14767 20223 14773
rect 20254 14764 20260 14776
rect 20312 14804 20318 14816
rect 20898 14804 20904 14816
rect 20312 14776 20904 14804
rect 20312 14764 20318 14776
rect 20898 14764 20904 14776
rect 20956 14764 20962 14816
rect 21652 14813 21680 14844
rect 21637 14807 21695 14813
rect 21637 14773 21649 14807
rect 21683 14773 21695 14807
rect 21637 14767 21695 14773
rect 23474 14764 23480 14816
rect 23532 14804 23538 14816
rect 24213 14807 24271 14813
rect 24213 14804 24225 14807
rect 23532 14776 24225 14804
rect 23532 14764 23538 14776
rect 24213 14773 24225 14776
rect 24259 14773 24271 14807
rect 24670 14804 24676 14816
rect 24631 14776 24676 14804
rect 24213 14767 24271 14773
rect 24670 14764 24676 14776
rect 24728 14764 24734 14816
rect 25222 14804 25228 14816
rect 25183 14776 25228 14804
rect 25222 14764 25228 14776
rect 25280 14764 25286 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 12621 14603 12679 14609
rect 12621 14569 12633 14603
rect 12667 14600 12679 14603
rect 12710 14600 12716 14612
rect 12667 14572 12716 14600
rect 12667 14569 12679 14572
rect 12621 14563 12679 14569
rect 12710 14560 12716 14572
rect 12768 14560 12774 14612
rect 13354 14560 13360 14612
rect 13412 14600 13418 14612
rect 13449 14603 13507 14609
rect 13449 14600 13461 14603
rect 13412 14572 13461 14600
rect 13412 14560 13418 14572
rect 13449 14569 13461 14572
rect 13495 14600 13507 14603
rect 14274 14600 14280 14612
rect 13495 14572 14280 14600
rect 13495 14569 13507 14572
rect 13449 14563 13507 14569
rect 14274 14560 14280 14572
rect 14332 14560 14338 14612
rect 15105 14603 15163 14609
rect 15105 14569 15117 14603
rect 15151 14600 15163 14603
rect 15562 14600 15568 14612
rect 15151 14572 15568 14600
rect 15151 14569 15163 14572
rect 15105 14563 15163 14569
rect 15562 14560 15568 14572
rect 15620 14560 15626 14612
rect 16485 14603 16543 14609
rect 16485 14569 16497 14603
rect 16531 14600 16543 14603
rect 17126 14600 17132 14612
rect 16531 14572 17132 14600
rect 16531 14569 16543 14572
rect 16485 14563 16543 14569
rect 17126 14560 17132 14572
rect 17184 14560 17190 14612
rect 17681 14603 17739 14609
rect 17681 14569 17693 14603
rect 17727 14600 17739 14603
rect 19150 14600 19156 14612
rect 17727 14572 19156 14600
rect 17727 14569 17739 14572
rect 17681 14563 17739 14569
rect 19150 14560 19156 14572
rect 19208 14560 19214 14612
rect 19242 14560 19248 14612
rect 19300 14600 19306 14612
rect 19797 14603 19855 14609
rect 19797 14600 19809 14603
rect 19300 14572 19809 14600
rect 19300 14560 19306 14572
rect 19797 14569 19809 14572
rect 19843 14600 19855 14603
rect 20622 14600 20628 14612
rect 19843 14572 20628 14600
rect 19843 14569 19855 14572
rect 19797 14563 19855 14569
rect 20622 14560 20628 14572
rect 20680 14560 20686 14612
rect 22094 14560 22100 14612
rect 22152 14600 22158 14612
rect 22281 14603 22339 14609
rect 22281 14600 22293 14603
rect 22152 14572 22293 14600
rect 22152 14560 22158 14572
rect 22281 14569 22293 14572
rect 22327 14569 22339 14603
rect 22281 14563 22339 14569
rect 22925 14603 22983 14609
rect 22925 14569 22937 14603
rect 22971 14600 22983 14603
rect 23106 14600 23112 14612
rect 22971 14572 23112 14600
rect 22971 14569 22983 14572
rect 22925 14563 22983 14569
rect 23106 14560 23112 14572
rect 23164 14560 23170 14612
rect 23293 14603 23351 14609
rect 23293 14569 23305 14603
rect 23339 14600 23351 14603
rect 24210 14600 24216 14612
rect 23339 14572 24216 14600
rect 23339 14569 23351 14572
rect 23293 14563 23351 14569
rect 24210 14560 24216 14572
rect 24268 14560 24274 14612
rect 13998 14532 14004 14544
rect 13959 14504 14004 14532
rect 13998 14492 14004 14504
rect 14056 14492 14062 14544
rect 14185 14535 14243 14541
rect 14185 14501 14197 14535
rect 14231 14532 14243 14535
rect 14366 14532 14372 14544
rect 14231 14504 14372 14532
rect 14231 14501 14243 14504
rect 14185 14495 14243 14501
rect 12158 14424 12164 14476
rect 12216 14464 12222 14476
rect 12713 14467 12771 14473
rect 12713 14464 12725 14467
rect 12216 14436 12725 14464
rect 12216 14424 12222 14436
rect 12713 14433 12725 14436
rect 12759 14433 12771 14467
rect 12713 14427 12771 14433
rect 13354 14424 13360 14476
rect 13412 14464 13418 14476
rect 14200 14464 14228 14495
rect 14366 14492 14372 14504
rect 14424 14492 14430 14544
rect 15838 14532 15844 14544
rect 15799 14504 15844 14532
rect 15838 14492 15844 14504
rect 15896 14492 15902 14544
rect 17494 14492 17500 14544
rect 17552 14532 17558 14544
rect 18040 14535 18098 14541
rect 18040 14532 18052 14535
rect 17552 14504 18052 14532
rect 17552 14492 17558 14504
rect 18040 14501 18052 14504
rect 18086 14532 18098 14535
rect 18598 14532 18604 14544
rect 18086 14504 18604 14532
rect 18086 14501 18098 14504
rect 18040 14495 18098 14501
rect 18598 14492 18604 14504
rect 18656 14492 18662 14544
rect 21174 14541 21180 14544
rect 20533 14535 20591 14541
rect 20533 14501 20545 14535
rect 20579 14532 20591 14535
rect 21168 14532 21180 14541
rect 20579 14504 21180 14532
rect 20579 14501 20591 14504
rect 20533 14495 20591 14501
rect 21168 14495 21180 14504
rect 21174 14492 21180 14495
rect 21232 14492 21238 14544
rect 24026 14541 24032 14544
rect 24020 14532 24032 14541
rect 23987 14504 24032 14532
rect 24020 14495 24032 14504
rect 24026 14492 24032 14495
rect 24084 14492 24090 14544
rect 15933 14467 15991 14473
rect 15933 14464 15945 14467
rect 13412 14436 14228 14464
rect 14292 14436 15945 14464
rect 13412 14424 13418 14436
rect 14292 14408 14320 14436
rect 15933 14433 15945 14436
rect 15979 14433 15991 14467
rect 15933 14427 15991 14433
rect 18966 14424 18972 14476
rect 19024 14464 19030 14476
rect 20165 14467 20223 14473
rect 20165 14464 20177 14467
rect 19024 14436 20177 14464
rect 19024 14424 19030 14436
rect 20165 14433 20177 14436
rect 20211 14464 20223 14467
rect 20622 14464 20628 14476
rect 20211 14436 20628 14464
rect 20211 14433 20223 14436
rect 20165 14427 20223 14433
rect 20622 14424 20628 14436
rect 20680 14424 20686 14476
rect 23753 14467 23811 14473
rect 23753 14433 23765 14467
rect 23799 14464 23811 14467
rect 23842 14464 23848 14476
rect 23799 14436 23848 14464
rect 23799 14433 23811 14436
rect 23753 14427 23811 14433
rect 23842 14424 23848 14436
rect 23900 14424 23906 14476
rect 11790 14356 11796 14408
rect 11848 14396 11854 14408
rect 12621 14399 12679 14405
rect 12621 14396 12633 14399
rect 11848 14368 12633 14396
rect 11848 14356 11854 14368
rect 12621 14365 12633 14368
rect 12667 14396 12679 14399
rect 13446 14396 13452 14408
rect 12667 14368 13452 14396
rect 12667 14365 12679 14368
rect 12621 14359 12679 14365
rect 13446 14356 13452 14368
rect 13504 14356 13510 14408
rect 14274 14396 14280 14408
rect 14235 14368 14280 14396
rect 14274 14356 14280 14368
rect 14332 14356 14338 14408
rect 15746 14396 15752 14408
rect 15707 14368 15752 14396
rect 15746 14356 15752 14368
rect 15804 14356 15810 14408
rect 17770 14396 17776 14408
rect 17731 14368 17776 14396
rect 17770 14356 17776 14368
rect 17828 14356 17834 14408
rect 20898 14396 20904 14408
rect 20859 14368 20904 14396
rect 20898 14356 20904 14368
rect 20956 14356 20962 14408
rect 13814 14288 13820 14340
rect 13872 14328 13878 14340
rect 15381 14331 15439 14337
rect 15381 14328 15393 14331
rect 13872 14300 15393 14328
rect 13872 14288 13878 14300
rect 15381 14297 15393 14300
rect 15427 14297 15439 14331
rect 15381 14291 15439 14297
rect 12161 14263 12219 14269
rect 12161 14229 12173 14263
rect 12207 14260 12219 14263
rect 13262 14260 13268 14272
rect 12207 14232 13268 14260
rect 12207 14229 12219 14232
rect 12161 14223 12219 14229
rect 13262 14220 13268 14232
rect 13320 14220 13326 14272
rect 13725 14263 13783 14269
rect 13725 14229 13737 14263
rect 13771 14260 13783 14263
rect 14090 14260 14096 14272
rect 13771 14232 14096 14260
rect 13771 14229 13783 14232
rect 13725 14223 13783 14229
rect 14090 14220 14096 14232
rect 14148 14220 14154 14272
rect 18138 14220 18144 14272
rect 18196 14260 18202 14272
rect 19153 14263 19211 14269
rect 19153 14260 19165 14263
rect 18196 14232 19165 14260
rect 18196 14220 18202 14232
rect 19153 14229 19165 14232
rect 19199 14229 19211 14263
rect 19153 14223 19211 14229
rect 23474 14220 23480 14272
rect 23532 14260 23538 14272
rect 23569 14263 23627 14269
rect 23569 14260 23581 14263
rect 23532 14232 23581 14260
rect 23532 14220 23538 14232
rect 23569 14229 23581 14232
rect 23615 14229 23627 14263
rect 23569 14223 23627 14229
rect 23934 14220 23940 14272
rect 23992 14260 23998 14272
rect 25133 14263 25191 14269
rect 25133 14260 25145 14263
rect 23992 14232 25145 14260
rect 23992 14220 23998 14232
rect 25133 14229 25145 14232
rect 25179 14229 25191 14263
rect 25133 14223 25191 14229
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 11790 14056 11796 14068
rect 11751 14028 11796 14056
rect 11790 14016 11796 14028
rect 11848 14016 11854 14068
rect 12158 14056 12164 14068
rect 12119 14028 12164 14056
rect 12158 14016 12164 14028
rect 12216 14016 12222 14068
rect 12710 14056 12716 14068
rect 12671 14028 12716 14056
rect 12710 14016 12716 14028
rect 12768 14016 12774 14068
rect 13354 14056 13360 14068
rect 13315 14028 13360 14056
rect 13354 14016 13360 14028
rect 13412 14016 13418 14068
rect 13725 14059 13783 14065
rect 13725 14025 13737 14059
rect 13771 14056 13783 14059
rect 13998 14056 14004 14068
rect 13771 14028 14004 14056
rect 13771 14025 13783 14028
rect 13725 14019 13783 14025
rect 13998 14016 14004 14028
rect 14056 14016 14062 14068
rect 14182 14016 14188 14068
rect 14240 14056 14246 14068
rect 15197 14059 15255 14065
rect 15197 14056 15209 14059
rect 14240 14028 15209 14056
rect 14240 14016 14246 14028
rect 15197 14025 15209 14028
rect 15243 14025 15255 14059
rect 15746 14056 15752 14068
rect 15707 14028 15752 14056
rect 15197 14019 15255 14025
rect 15746 14016 15752 14028
rect 15804 14016 15810 14068
rect 16482 14056 16488 14068
rect 16443 14028 16488 14056
rect 16482 14016 16488 14028
rect 16540 14016 16546 14068
rect 17494 14056 17500 14068
rect 17455 14028 17500 14056
rect 17494 14016 17500 14028
rect 17552 14016 17558 14068
rect 18414 14056 18420 14068
rect 18375 14028 18420 14056
rect 18414 14016 18420 14028
rect 18472 14016 18478 14068
rect 18966 14056 18972 14068
rect 18927 14028 18972 14056
rect 18966 14016 18972 14028
rect 19024 14016 19030 14068
rect 20162 14016 20168 14068
rect 20220 14056 20226 14068
rect 20257 14059 20315 14065
rect 20257 14056 20269 14059
rect 20220 14028 20269 14056
rect 20220 14016 20226 14028
rect 20257 14025 20269 14028
rect 20303 14025 20315 14059
rect 20257 14019 20315 14025
rect 20438 14016 20444 14068
rect 20496 14056 20502 14068
rect 20533 14059 20591 14065
rect 20533 14056 20545 14059
rect 20496 14028 20545 14056
rect 20496 14016 20502 14028
rect 20533 14025 20545 14028
rect 20579 14025 20591 14059
rect 20533 14019 20591 14025
rect 20898 14016 20904 14068
rect 20956 14056 20962 14068
rect 21545 14059 21603 14065
rect 21545 14056 21557 14059
rect 20956 14028 21557 14056
rect 20956 14016 20962 14028
rect 21545 14025 21557 14028
rect 21591 14056 21603 14059
rect 21910 14056 21916 14068
rect 21591 14028 21916 14056
rect 21591 14025 21603 14028
rect 21545 14019 21603 14025
rect 21910 14016 21916 14028
rect 21968 14016 21974 14068
rect 23106 14056 23112 14068
rect 23019 14028 23112 14056
rect 23106 14016 23112 14028
rect 23164 14056 23170 14068
rect 24026 14056 24032 14068
rect 23164 14028 24032 14056
rect 23164 14016 23170 14028
rect 24026 14016 24032 14028
rect 24084 14016 24090 14068
rect 25501 14059 25559 14065
rect 25501 14056 25513 14059
rect 24136 14028 25513 14056
rect 17218 13988 17224 14000
rect 16960 13960 17224 13988
rect 12802 13920 12808 13932
rect 12763 13892 12808 13920
rect 12802 13880 12808 13892
rect 12860 13880 12866 13932
rect 16574 13880 16580 13932
rect 16632 13920 16638 13932
rect 16960 13929 16988 13960
rect 17218 13948 17224 13960
rect 17276 13948 17282 14000
rect 18432 13988 18460 14016
rect 19242 13988 19248 14000
rect 18432 13960 19248 13988
rect 19242 13948 19248 13960
rect 19300 13948 19306 14000
rect 22097 13991 22155 13997
rect 22097 13957 22109 13991
rect 22143 13988 22155 13991
rect 23198 13988 23204 14000
rect 22143 13960 23204 13988
rect 22143 13957 22155 13960
rect 22097 13951 22155 13957
rect 23198 13948 23204 13960
rect 23256 13948 23262 14000
rect 23566 13988 23572 14000
rect 23400 13960 23572 13988
rect 16945 13923 17003 13929
rect 16945 13920 16957 13923
rect 16632 13892 16957 13920
rect 16632 13880 16638 13892
rect 16945 13889 16957 13892
rect 16991 13889 17003 13923
rect 16945 13883 17003 13889
rect 17037 13923 17095 13929
rect 17037 13889 17049 13923
rect 17083 13920 17095 13923
rect 17126 13920 17132 13932
rect 17083 13892 17132 13920
rect 17083 13889 17095 13892
rect 17037 13883 17095 13889
rect 17126 13880 17132 13892
rect 17184 13880 17190 13932
rect 19426 13880 19432 13932
rect 19484 13920 19490 13932
rect 19521 13923 19579 13929
rect 19521 13920 19533 13923
rect 19484 13892 19533 13920
rect 19484 13880 19490 13892
rect 19521 13889 19533 13892
rect 19567 13920 19579 13923
rect 19981 13923 20039 13929
rect 19981 13920 19993 13923
rect 19567 13892 19993 13920
rect 19567 13889 19579 13892
rect 19521 13883 19579 13889
rect 19981 13889 19993 13892
rect 20027 13920 20039 13923
rect 21085 13923 21143 13929
rect 21085 13920 21097 13923
rect 20027 13892 21097 13920
rect 20027 13889 20039 13892
rect 19981 13883 20039 13889
rect 21085 13889 21097 13892
rect 21131 13920 21143 13923
rect 21174 13920 21180 13932
rect 21131 13892 21180 13920
rect 21131 13889 21143 13892
rect 21085 13883 21143 13889
rect 21174 13880 21180 13892
rect 21232 13880 21238 13932
rect 21913 13923 21971 13929
rect 21913 13889 21925 13923
rect 21959 13920 21971 13923
rect 22649 13923 22707 13929
rect 22649 13920 22661 13923
rect 21959 13892 22661 13920
rect 21959 13889 21971 13892
rect 21913 13883 21971 13889
rect 22649 13889 22661 13892
rect 22695 13920 22707 13923
rect 23400 13920 23428 13960
rect 23566 13948 23572 13960
rect 23624 13988 23630 14000
rect 24136 13988 24164 14028
rect 25501 14025 25513 14028
rect 25547 14025 25559 14059
rect 25501 14019 25559 14025
rect 23624 13960 24164 13988
rect 23624 13948 23630 13960
rect 22695 13892 23428 13920
rect 23477 13923 23535 13929
rect 22695 13889 22707 13892
rect 22649 13883 22707 13889
rect 23477 13889 23489 13923
rect 23523 13920 23535 13923
rect 23842 13920 23848 13932
rect 23523 13892 23848 13920
rect 23523 13889 23535 13892
rect 23477 13883 23535 13889
rect 23842 13880 23848 13892
rect 23900 13880 23906 13932
rect 23934 13880 23940 13932
rect 23992 13920 23998 13932
rect 23992 13892 24256 13920
rect 23992 13880 23998 13892
rect 13814 13852 13820 13864
rect 13775 13824 13820 13852
rect 13814 13812 13820 13824
rect 13872 13812 13878 13864
rect 16301 13855 16359 13861
rect 16301 13821 16313 13855
rect 16347 13852 16359 13855
rect 18785 13855 18843 13861
rect 16347 13824 16528 13852
rect 16347 13821 16359 13824
rect 16301 13815 16359 13821
rect 14084 13787 14142 13793
rect 14084 13753 14096 13787
rect 14130 13784 14142 13787
rect 14274 13784 14280 13796
rect 14130 13756 14280 13784
rect 14130 13753 14142 13756
rect 14084 13747 14142 13753
rect 14274 13744 14280 13756
rect 14332 13744 14338 13796
rect 16500 13784 16528 13824
rect 18785 13821 18797 13855
rect 18831 13852 18843 13855
rect 19245 13855 19303 13861
rect 19245 13852 19257 13855
rect 18831 13824 19257 13852
rect 18831 13821 18843 13824
rect 18785 13815 18843 13821
rect 19245 13821 19257 13824
rect 19291 13852 19303 13855
rect 20530 13852 20536 13864
rect 19291 13824 20536 13852
rect 19291 13821 19303 13824
rect 19245 13815 19303 13821
rect 20530 13812 20536 13824
rect 20588 13812 20594 13864
rect 21192 13852 21220 13880
rect 22278 13852 22284 13864
rect 21192 13824 22284 13852
rect 22278 13812 22284 13824
rect 22336 13812 22342 13864
rect 23750 13852 23756 13864
rect 23400 13824 23756 13852
rect 16945 13787 17003 13793
rect 16945 13784 16957 13787
rect 16500 13756 16957 13784
rect 16945 13753 16957 13756
rect 16991 13784 17003 13787
rect 18230 13784 18236 13796
rect 16991 13756 18236 13784
rect 16991 13753 17003 13756
rect 16945 13747 17003 13753
rect 18230 13744 18236 13756
rect 18288 13744 18294 13796
rect 19334 13744 19340 13796
rect 19392 13784 19398 13796
rect 19429 13787 19487 13793
rect 19429 13784 19441 13787
rect 19392 13756 19441 13784
rect 19392 13744 19398 13756
rect 19429 13753 19441 13756
rect 19475 13753 19487 13787
rect 19429 13747 19487 13753
rect 20162 13744 20168 13796
rect 20220 13784 20226 13796
rect 20809 13787 20867 13793
rect 20809 13784 20821 13787
rect 20220 13756 20821 13784
rect 20220 13744 20226 13756
rect 20809 13753 20821 13756
rect 20855 13753 20867 13787
rect 20990 13784 20996 13796
rect 20951 13756 20996 13784
rect 20809 13747 20867 13753
rect 20990 13744 20996 13756
rect 21048 13744 21054 13796
rect 22373 13787 22431 13793
rect 22373 13753 22385 13787
rect 22419 13784 22431 13787
rect 22462 13784 22468 13796
rect 22419 13756 22468 13784
rect 22419 13753 22431 13756
rect 22373 13747 22431 13753
rect 22462 13744 22468 13756
rect 22520 13744 22526 13796
rect 23400 13784 23428 13824
rect 23750 13812 23756 13824
rect 23808 13812 23814 13864
rect 23860 13852 23888 13880
rect 24029 13855 24087 13861
rect 24029 13852 24041 13855
rect 23860 13824 24041 13852
rect 24029 13821 24041 13824
rect 24075 13852 24087 13855
rect 24121 13855 24179 13861
rect 24121 13852 24133 13855
rect 24075 13824 24133 13852
rect 24075 13821 24087 13824
rect 24029 13815 24087 13821
rect 24121 13821 24133 13824
rect 24167 13821 24179 13855
rect 24228 13852 24256 13892
rect 24394 13861 24400 13864
rect 24377 13855 24400 13861
rect 24377 13852 24389 13855
rect 24228 13824 24389 13852
rect 24121 13815 24179 13821
rect 24377 13821 24389 13824
rect 24452 13852 24458 13864
rect 24452 13824 24525 13852
rect 24377 13815 24400 13821
rect 24394 13812 24400 13815
rect 24452 13812 24458 13824
rect 22848 13756 23428 13784
rect 17126 13676 17132 13728
rect 17184 13716 17190 13728
rect 17770 13716 17776 13728
rect 17184 13688 17776 13716
rect 17184 13676 17190 13688
rect 17770 13676 17776 13688
rect 17828 13676 17834 13728
rect 22094 13676 22100 13728
rect 22152 13716 22158 13728
rect 22557 13719 22615 13725
rect 22557 13716 22569 13719
rect 22152 13688 22569 13716
rect 22152 13676 22158 13688
rect 22557 13685 22569 13688
rect 22603 13716 22615 13719
rect 22848 13716 22876 13756
rect 22603 13688 22876 13716
rect 22603 13685 22615 13688
rect 22557 13679 22615 13685
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 12158 13472 12164 13524
rect 12216 13512 12222 13524
rect 12434 13512 12440 13524
rect 12216 13484 12440 13512
rect 12216 13472 12222 13484
rect 12434 13472 12440 13484
rect 12492 13512 12498 13524
rect 12805 13515 12863 13521
rect 12805 13512 12817 13515
rect 12492 13484 12817 13512
rect 12492 13472 12498 13484
rect 12805 13481 12817 13484
rect 12851 13481 12863 13515
rect 12805 13475 12863 13481
rect 13814 13472 13820 13524
rect 13872 13512 13878 13524
rect 13909 13515 13967 13521
rect 13909 13512 13921 13515
rect 13872 13484 13921 13512
rect 13872 13472 13878 13484
rect 13909 13481 13921 13484
rect 13955 13512 13967 13515
rect 14826 13512 14832 13524
rect 13955 13484 14832 13512
rect 13955 13481 13967 13484
rect 13909 13475 13967 13481
rect 14826 13472 14832 13484
rect 14884 13472 14890 13524
rect 15565 13515 15623 13521
rect 15565 13481 15577 13515
rect 15611 13512 15623 13515
rect 15838 13512 15844 13524
rect 15611 13484 15844 13512
rect 15611 13481 15623 13484
rect 15565 13475 15623 13481
rect 15838 13472 15844 13484
rect 15896 13472 15902 13524
rect 16206 13472 16212 13524
rect 16264 13512 16270 13524
rect 16482 13512 16488 13524
rect 16264 13484 16488 13512
rect 16264 13472 16270 13484
rect 16482 13472 16488 13484
rect 16540 13472 16546 13524
rect 17402 13472 17408 13524
rect 17460 13512 17466 13524
rect 17678 13512 17684 13524
rect 17460 13484 17684 13512
rect 17460 13472 17466 13484
rect 17678 13472 17684 13484
rect 17736 13472 17742 13524
rect 17862 13472 17868 13524
rect 17920 13512 17926 13524
rect 18141 13515 18199 13521
rect 18141 13512 18153 13515
rect 17920 13484 18153 13512
rect 17920 13472 17926 13484
rect 18141 13481 18153 13484
rect 18187 13512 18199 13515
rect 18414 13512 18420 13524
rect 18187 13484 18420 13512
rect 18187 13481 18199 13484
rect 18141 13475 18199 13481
rect 18414 13472 18420 13484
rect 18472 13472 18478 13524
rect 19426 13512 19432 13524
rect 19387 13484 19432 13512
rect 19426 13472 19432 13484
rect 19484 13472 19490 13524
rect 20438 13512 20444 13524
rect 19536 13484 20444 13512
rect 11146 13404 11152 13456
rect 11204 13444 11210 13456
rect 11692 13447 11750 13453
rect 11692 13444 11704 13447
rect 11204 13416 11704 13444
rect 11204 13404 11210 13416
rect 11692 13413 11704 13416
rect 11738 13444 11750 13447
rect 12342 13444 12348 13456
rect 11738 13416 12348 13444
rect 11738 13413 11750 13416
rect 11692 13407 11750 13413
rect 12342 13404 12348 13416
rect 12400 13404 12406 13456
rect 17310 13444 17316 13456
rect 17271 13416 17316 13444
rect 17310 13404 17316 13416
rect 17368 13404 17374 13456
rect 18046 13404 18052 13456
rect 18104 13444 18110 13456
rect 18877 13447 18935 13453
rect 18877 13444 18889 13447
rect 18104 13416 18889 13444
rect 18104 13404 18110 13416
rect 18877 13413 18889 13416
rect 18923 13444 18935 13447
rect 19536 13444 19564 13484
rect 20438 13472 20444 13484
rect 20496 13472 20502 13524
rect 20533 13515 20591 13521
rect 20533 13481 20545 13515
rect 20579 13512 20591 13515
rect 20990 13512 20996 13524
rect 20579 13484 20996 13512
rect 20579 13481 20591 13484
rect 20533 13475 20591 13481
rect 20990 13472 20996 13484
rect 21048 13472 21054 13524
rect 21174 13472 21180 13524
rect 21232 13512 21238 13524
rect 21453 13515 21511 13521
rect 21453 13512 21465 13515
rect 21232 13484 21465 13512
rect 21232 13472 21238 13484
rect 21453 13481 21465 13484
rect 21499 13512 21511 13515
rect 21818 13512 21824 13524
rect 21499 13484 21824 13512
rect 21499 13481 21511 13484
rect 21453 13475 21511 13481
rect 21818 13472 21824 13484
rect 21876 13472 21882 13524
rect 22094 13472 22100 13524
rect 22152 13512 22158 13524
rect 23106 13512 23112 13524
rect 22152 13484 22197 13512
rect 23067 13484 23112 13512
rect 22152 13472 22158 13484
rect 23106 13472 23112 13484
rect 23164 13512 23170 13524
rect 23164 13484 23888 13512
rect 23164 13472 23170 13484
rect 23860 13456 23888 13484
rect 24394 13472 24400 13524
rect 24452 13512 24458 13524
rect 24581 13515 24639 13521
rect 24581 13512 24593 13515
rect 24452 13484 24593 13512
rect 24452 13472 24458 13484
rect 24581 13481 24593 13484
rect 24627 13512 24639 13515
rect 24627 13484 25452 13512
rect 24627 13481 24639 13484
rect 24581 13475 24639 13481
rect 18923 13416 19564 13444
rect 18923 13413 18935 13416
rect 18877 13407 18935 13413
rect 19610 13404 19616 13456
rect 19668 13444 19674 13456
rect 20070 13444 20076 13456
rect 19668 13416 20076 13444
rect 19668 13404 19674 13416
rect 20070 13404 20076 13416
rect 20128 13404 20134 13456
rect 22646 13404 22652 13456
rect 22704 13444 22710 13456
rect 23753 13447 23811 13453
rect 23753 13444 23765 13447
rect 22704 13416 23765 13444
rect 22704 13404 22710 13416
rect 23753 13413 23765 13416
rect 23799 13413 23811 13447
rect 23753 13407 23811 13413
rect 23842 13404 23848 13456
rect 23900 13444 23906 13456
rect 25133 13447 25191 13453
rect 23900 13416 23993 13444
rect 23900 13404 23906 13416
rect 25133 13413 25145 13447
rect 25179 13444 25191 13447
rect 25222 13444 25228 13456
rect 25179 13416 25228 13444
rect 25179 13413 25191 13416
rect 25133 13407 25191 13413
rect 25222 13404 25228 13416
rect 25280 13404 25286 13456
rect 25424 13453 25452 13484
rect 25317 13447 25375 13453
rect 25317 13413 25329 13447
rect 25363 13413 25375 13447
rect 25317 13407 25375 13413
rect 25409 13447 25467 13453
rect 25409 13413 25421 13447
rect 25455 13444 25467 13447
rect 25682 13444 25688 13456
rect 25455 13416 25688 13444
rect 25455 13413 25467 13416
rect 25409 13407 25467 13413
rect 18690 13336 18696 13388
rect 18748 13376 18754 13388
rect 18969 13379 19027 13385
rect 18969 13376 18981 13379
rect 18748 13348 18981 13376
rect 18748 13336 18754 13348
rect 18969 13345 18981 13348
rect 19015 13345 19027 13379
rect 18969 13339 19027 13345
rect 23106 13336 23112 13388
rect 23164 13376 23170 13388
rect 23569 13379 23627 13385
rect 23569 13376 23581 13379
rect 23164 13348 23581 13376
rect 23164 13336 23170 13348
rect 23569 13345 23581 13348
rect 23615 13345 23627 13379
rect 23569 13339 23627 13345
rect 24118 13336 24124 13388
rect 24176 13376 24182 13388
rect 24854 13376 24860 13388
rect 24176 13348 24860 13376
rect 24176 13336 24182 13348
rect 24854 13336 24860 13348
rect 24912 13376 24918 13388
rect 25332 13376 25360 13407
rect 25682 13404 25688 13416
rect 25740 13404 25746 13456
rect 24912 13348 25360 13376
rect 24912 13336 24918 13348
rect 11422 13308 11428 13320
rect 11383 13280 11428 13308
rect 11422 13268 11428 13280
rect 11480 13268 11486 13320
rect 15746 13308 15752 13320
rect 15707 13280 15752 13308
rect 15746 13268 15752 13280
rect 15804 13268 15810 13320
rect 17221 13311 17279 13317
rect 17221 13277 17233 13311
rect 17267 13277 17279 13311
rect 17402 13308 17408 13320
rect 17363 13280 17408 13308
rect 17221 13271 17279 13277
rect 17236 13240 17264 13271
rect 17402 13268 17408 13280
rect 17460 13268 17466 13320
rect 18877 13311 18935 13317
rect 18877 13277 18889 13311
rect 18923 13308 18935 13311
rect 19058 13308 19064 13320
rect 18923 13280 19064 13308
rect 18923 13277 18935 13280
rect 18877 13271 18935 13277
rect 19058 13268 19064 13280
rect 19116 13268 19122 13320
rect 21358 13308 21364 13320
rect 21319 13280 21364 13308
rect 21358 13268 21364 13280
rect 21416 13268 21422 13320
rect 21545 13311 21603 13317
rect 21545 13277 21557 13311
rect 21591 13308 21603 13311
rect 22278 13308 22284 13320
rect 21591 13280 22284 13308
rect 21591 13277 21603 13280
rect 21545 13271 21603 13277
rect 22278 13268 22284 13280
rect 22336 13268 22342 13320
rect 22462 13308 22468 13320
rect 22375 13280 22468 13308
rect 22462 13268 22468 13280
rect 22520 13308 22526 13320
rect 22520 13280 23612 13308
rect 22520 13268 22526 13280
rect 17770 13240 17776 13252
rect 17236 13212 17776 13240
rect 17770 13200 17776 13212
rect 17828 13240 17834 13252
rect 18417 13243 18475 13249
rect 18417 13240 18429 13243
rect 17828 13212 18429 13240
rect 17828 13200 17834 13212
rect 18417 13209 18429 13212
rect 18463 13209 18475 13243
rect 18417 13203 18475 13209
rect 23293 13243 23351 13249
rect 23293 13209 23305 13243
rect 23339 13240 23351 13243
rect 23474 13240 23480 13252
rect 23339 13212 23480 13240
rect 23339 13209 23351 13212
rect 23293 13203 23351 13209
rect 23474 13200 23480 13212
rect 23532 13200 23538 13252
rect 23584 13240 23612 13280
rect 24857 13243 24915 13249
rect 24857 13240 24869 13243
rect 23584 13212 24869 13240
rect 24857 13209 24869 13212
rect 24903 13209 24915 13243
rect 24857 13203 24915 13209
rect 14274 13172 14280 13184
rect 14187 13144 14280 13172
rect 14274 13132 14280 13144
rect 14332 13172 14338 13184
rect 14645 13175 14703 13181
rect 14645 13172 14657 13175
rect 14332 13144 14657 13172
rect 14332 13132 14338 13144
rect 14645 13141 14657 13144
rect 14691 13172 14703 13175
rect 15105 13175 15163 13181
rect 15105 13172 15117 13175
rect 14691 13144 15117 13172
rect 14691 13141 14703 13144
rect 14645 13135 14703 13141
rect 15105 13141 15117 13144
rect 15151 13172 15163 13175
rect 15286 13172 15292 13184
rect 15151 13144 15292 13172
rect 15151 13141 15163 13144
rect 15105 13135 15163 13141
rect 15286 13132 15292 13144
rect 15344 13132 15350 13184
rect 15562 13132 15568 13184
rect 15620 13172 15626 13184
rect 16853 13175 16911 13181
rect 16853 13172 16865 13175
rect 15620 13144 16865 13172
rect 15620 13132 15626 13144
rect 16853 13141 16865 13144
rect 16899 13141 16911 13175
rect 16853 13135 16911 13141
rect 19797 13175 19855 13181
rect 19797 13141 19809 13175
rect 19843 13172 19855 13175
rect 19978 13172 19984 13184
rect 19843 13144 19984 13172
rect 19843 13141 19855 13144
rect 19797 13135 19855 13141
rect 19978 13132 19984 13144
rect 20036 13132 20042 13184
rect 20162 13172 20168 13184
rect 20123 13144 20168 13172
rect 20162 13132 20168 13144
rect 20220 13132 20226 13184
rect 20993 13175 21051 13181
rect 20993 13141 21005 13175
rect 21039 13172 21051 13175
rect 21726 13172 21732 13184
rect 21039 13144 21732 13172
rect 21039 13141 21051 13144
rect 20993 13135 21051 13141
rect 21726 13132 21732 13144
rect 21784 13132 21790 13184
rect 24210 13172 24216 13184
rect 24171 13144 24216 13172
rect 24210 13132 24216 13144
rect 24268 13132 24274 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 11146 12968 11152 12980
rect 11107 12940 11152 12968
rect 11146 12928 11152 12940
rect 11204 12928 11210 12980
rect 15286 12928 15292 12980
rect 15344 12968 15350 12980
rect 16393 12971 16451 12977
rect 16393 12968 16405 12971
rect 15344 12940 16405 12968
rect 15344 12928 15350 12940
rect 16393 12937 16405 12940
rect 16439 12937 16451 12971
rect 17034 12968 17040 12980
rect 16947 12940 17040 12968
rect 16393 12931 16451 12937
rect 17034 12928 17040 12940
rect 17092 12968 17098 12980
rect 17402 12968 17408 12980
rect 17092 12940 17408 12968
rect 17092 12928 17098 12940
rect 17402 12928 17408 12940
rect 17460 12968 17466 12980
rect 17862 12968 17868 12980
rect 17460 12940 17868 12968
rect 17460 12928 17466 12940
rect 17862 12928 17868 12940
rect 17920 12928 17926 12980
rect 19058 12968 19064 12980
rect 19019 12940 19064 12968
rect 19058 12928 19064 12940
rect 19116 12928 19122 12980
rect 20346 12928 20352 12980
rect 20404 12968 20410 12980
rect 22646 12968 22652 12980
rect 20404 12940 21680 12968
rect 22607 12940 22652 12968
rect 20404 12928 20410 12940
rect 12434 12860 12440 12912
rect 12492 12860 12498 12912
rect 17497 12903 17555 12909
rect 17497 12869 17509 12903
rect 17543 12900 17555 12903
rect 17678 12900 17684 12912
rect 17543 12872 17684 12900
rect 17543 12869 17555 12872
rect 17497 12863 17555 12869
rect 17678 12860 17684 12872
rect 17736 12860 17742 12912
rect 17773 12903 17831 12909
rect 17773 12869 17785 12903
rect 17819 12900 17831 12903
rect 18046 12900 18052 12912
rect 17819 12872 18052 12900
rect 17819 12869 17831 12872
rect 17773 12863 17831 12869
rect 18046 12860 18052 12872
rect 18104 12860 18110 12912
rect 18141 12903 18199 12909
rect 18141 12869 18153 12903
rect 18187 12869 18199 12903
rect 18141 12863 18199 12869
rect 20165 12903 20223 12909
rect 20165 12869 20177 12903
rect 20211 12900 20223 12903
rect 20438 12900 20444 12912
rect 20211 12872 20444 12900
rect 20211 12869 20223 12872
rect 20165 12863 20223 12869
rect 11885 12835 11943 12841
rect 11885 12801 11897 12835
rect 11931 12832 11943 12835
rect 12452 12832 12480 12860
rect 11931 12804 12480 12832
rect 11931 12801 11943 12804
rect 11885 12795 11943 12801
rect 17402 12792 17408 12844
rect 17460 12832 17466 12844
rect 18156 12832 18184 12863
rect 20438 12860 20444 12872
rect 20496 12860 20502 12912
rect 21174 12900 21180 12912
rect 21135 12872 21180 12900
rect 21174 12860 21180 12872
rect 21232 12860 21238 12912
rect 17460 12804 18184 12832
rect 17460 12792 17466 12804
rect 20714 12792 20720 12844
rect 20772 12832 20778 12844
rect 21358 12832 21364 12844
rect 20772 12804 21364 12832
rect 20772 12792 20778 12804
rect 21358 12792 21364 12804
rect 21416 12832 21422 12844
rect 21652 12841 21680 12940
rect 22646 12928 22652 12940
rect 22704 12928 22710 12980
rect 24854 12968 24860 12980
rect 24815 12940 24860 12968
rect 24854 12928 24860 12940
rect 24912 12928 24918 12980
rect 25682 12968 25688 12980
rect 25643 12940 25688 12968
rect 25682 12928 25688 12940
rect 25740 12928 25746 12980
rect 23750 12900 23756 12912
rect 23711 12872 23756 12900
rect 23750 12860 23756 12872
rect 23808 12860 23814 12912
rect 21453 12835 21511 12841
rect 21453 12832 21465 12835
rect 21416 12804 21465 12832
rect 21416 12792 21422 12804
rect 21453 12801 21465 12804
rect 21499 12801 21511 12835
rect 21453 12795 21511 12801
rect 21637 12835 21695 12841
rect 21637 12801 21649 12835
rect 21683 12801 21695 12835
rect 24210 12832 24216 12844
rect 24171 12804 24216 12832
rect 21637 12795 21695 12801
rect 24210 12792 24216 12804
rect 24268 12832 24274 12844
rect 25225 12835 25283 12841
rect 25225 12832 25237 12835
rect 24268 12804 25237 12832
rect 24268 12792 24274 12804
rect 25225 12801 25237 12804
rect 25271 12801 25283 12835
rect 25225 12795 25283 12801
rect 11422 12724 11428 12776
rect 11480 12764 11486 12776
rect 11517 12767 11575 12773
rect 11517 12764 11529 12767
rect 11480 12736 11529 12764
rect 11480 12724 11486 12736
rect 11517 12733 11529 12736
rect 11563 12764 11575 12767
rect 12253 12767 12311 12773
rect 12253 12764 12265 12767
rect 11563 12736 12265 12764
rect 11563 12733 11575 12736
rect 11517 12727 11575 12733
rect 12253 12733 12265 12736
rect 12299 12764 12311 12767
rect 12434 12764 12440 12776
rect 12299 12736 12440 12764
rect 12299 12733 12311 12736
rect 12253 12727 12311 12733
rect 12434 12724 12440 12736
rect 12492 12724 12498 12776
rect 15013 12767 15071 12773
rect 15013 12764 15025 12767
rect 14936 12736 15025 12764
rect 12526 12656 12532 12708
rect 12584 12696 12590 12708
rect 12682 12699 12740 12705
rect 12682 12696 12694 12699
rect 12584 12668 12694 12696
rect 12584 12656 12590 12668
rect 12682 12665 12694 12668
rect 12728 12665 12740 12699
rect 12682 12659 12740 12665
rect 14936 12640 14964 12736
rect 15013 12733 15025 12736
rect 15059 12733 15071 12767
rect 18414 12764 18420 12776
rect 18375 12736 18420 12764
rect 15013 12727 15071 12733
rect 18414 12724 18420 12736
rect 18472 12764 18478 12776
rect 18598 12764 18604 12776
rect 18472 12736 18604 12764
rect 18472 12724 18478 12736
rect 18598 12724 18604 12736
rect 18656 12724 18662 12776
rect 19978 12724 19984 12776
rect 20036 12764 20042 12776
rect 20441 12767 20499 12773
rect 20441 12764 20453 12767
rect 20036 12736 20453 12764
rect 20036 12724 20042 12736
rect 20441 12733 20453 12736
rect 20487 12764 20499 12767
rect 20806 12764 20812 12776
rect 20487 12736 20812 12764
rect 20487 12733 20499 12736
rect 20441 12727 20499 12733
rect 20806 12724 20812 12736
rect 20864 12724 20870 12776
rect 15280 12699 15338 12705
rect 15280 12665 15292 12699
rect 15326 12696 15338 12699
rect 15378 12696 15384 12708
rect 15326 12668 15384 12696
rect 15326 12665 15338 12668
rect 15280 12659 15338 12665
rect 15378 12656 15384 12668
rect 15436 12656 15442 12708
rect 18690 12696 18696 12708
rect 18603 12668 18696 12696
rect 18690 12656 18696 12668
rect 18748 12696 18754 12708
rect 19334 12696 19340 12708
rect 18748 12668 19340 12696
rect 18748 12656 18754 12668
rect 19334 12656 19340 12668
rect 19392 12696 19398 12708
rect 19521 12699 19579 12705
rect 19521 12696 19533 12699
rect 19392 12668 19533 12696
rect 19392 12656 19398 12668
rect 19521 12665 19533 12668
rect 19567 12696 19579 12699
rect 19797 12699 19855 12705
rect 19797 12696 19809 12699
rect 19567 12668 19809 12696
rect 19567 12665 19579 12668
rect 19521 12659 19579 12665
rect 19797 12665 19809 12668
rect 19843 12665 19855 12699
rect 20714 12696 20720 12708
rect 20675 12668 20720 12696
rect 19797 12659 19855 12665
rect 20714 12656 20720 12668
rect 20772 12656 20778 12708
rect 21082 12656 21088 12708
rect 21140 12696 21146 12708
rect 21358 12696 21364 12708
rect 21140 12668 21364 12696
rect 21140 12656 21146 12668
rect 21358 12656 21364 12668
rect 21416 12656 21422 12708
rect 24302 12696 24308 12708
rect 24263 12668 24308 12696
rect 24302 12656 24308 12668
rect 24360 12656 24366 12708
rect 12342 12588 12348 12640
rect 12400 12628 12406 12640
rect 13817 12631 13875 12637
rect 13817 12628 13829 12631
rect 12400 12600 13829 12628
rect 12400 12588 12406 12600
rect 13817 12597 13829 12600
rect 13863 12628 13875 12631
rect 13906 12628 13912 12640
rect 13863 12600 13912 12628
rect 13863 12597 13875 12600
rect 13817 12591 13875 12597
rect 13906 12588 13912 12600
rect 13964 12588 13970 12640
rect 14918 12628 14924 12640
rect 14879 12600 14924 12628
rect 14918 12588 14924 12600
rect 14976 12588 14982 12640
rect 17678 12588 17684 12640
rect 17736 12628 17742 12640
rect 18601 12631 18659 12637
rect 18601 12628 18613 12631
rect 17736 12600 18613 12628
rect 17736 12588 17742 12600
rect 18601 12597 18613 12600
rect 18647 12597 18659 12631
rect 18601 12591 18659 12597
rect 20162 12588 20168 12640
rect 20220 12628 20226 12640
rect 20530 12628 20536 12640
rect 20220 12600 20536 12628
rect 20220 12588 20226 12600
rect 20530 12588 20536 12600
rect 20588 12628 20594 12640
rect 20625 12631 20683 12637
rect 20625 12628 20637 12631
rect 20588 12600 20637 12628
rect 20588 12588 20594 12600
rect 20625 12597 20637 12600
rect 20671 12597 20683 12631
rect 20625 12591 20683 12597
rect 22189 12631 22247 12637
rect 22189 12597 22201 12631
rect 22235 12628 22247 12631
rect 22278 12628 22284 12640
rect 22235 12600 22284 12628
rect 22235 12597 22247 12600
rect 22189 12591 22247 12597
rect 22278 12588 22284 12600
rect 22336 12588 22342 12640
rect 23106 12628 23112 12640
rect 23067 12600 23112 12628
rect 23106 12588 23112 12600
rect 23164 12588 23170 12640
rect 23477 12631 23535 12637
rect 23477 12597 23489 12631
rect 23523 12628 23535 12631
rect 24213 12631 24271 12637
rect 24213 12628 24225 12631
rect 23523 12600 24225 12628
rect 23523 12597 23535 12600
rect 23477 12591 23535 12597
rect 24213 12597 24225 12600
rect 24259 12628 24271 12631
rect 25038 12628 25044 12640
rect 24259 12600 25044 12628
rect 24259 12597 24271 12600
rect 24213 12591 24271 12597
rect 25038 12588 25044 12600
rect 25096 12588 25102 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 17402 12424 17408 12436
rect 17363 12396 17408 12424
rect 17402 12384 17408 12396
rect 17460 12384 17466 12436
rect 17770 12424 17776 12436
rect 17731 12396 17776 12424
rect 17770 12384 17776 12396
rect 17828 12384 17834 12436
rect 17862 12384 17868 12436
rect 17920 12424 17926 12436
rect 19245 12427 19303 12433
rect 19245 12424 19257 12427
rect 17920 12396 19257 12424
rect 17920 12384 17926 12396
rect 19245 12393 19257 12396
rect 19291 12393 19303 12427
rect 19245 12387 19303 12393
rect 20714 12384 20720 12436
rect 20772 12424 20778 12436
rect 21174 12424 21180 12436
rect 20772 12396 21180 12424
rect 20772 12384 20778 12396
rect 21174 12384 21180 12396
rect 21232 12384 21238 12436
rect 23842 12424 23848 12436
rect 23803 12396 23848 12424
rect 23842 12384 23848 12396
rect 23900 12384 23906 12436
rect 24857 12427 24915 12433
rect 24857 12393 24869 12427
rect 24903 12424 24915 12427
rect 25222 12424 25228 12436
rect 24903 12396 25228 12424
rect 24903 12393 24915 12396
rect 24857 12387 24915 12393
rect 25222 12384 25228 12396
rect 25280 12384 25286 12436
rect 12250 12356 12256 12368
rect 12211 12328 12256 12356
rect 12250 12316 12256 12328
rect 12308 12316 12314 12368
rect 12342 12316 12348 12368
rect 12400 12356 12406 12368
rect 13814 12356 13820 12368
rect 12400 12328 12445 12356
rect 13775 12328 13820 12356
rect 12400 12316 12406 12328
rect 13814 12316 13820 12328
rect 13872 12356 13878 12368
rect 14182 12356 14188 12368
rect 13872 12328 14188 12356
rect 13872 12316 13878 12328
rect 14182 12316 14188 12328
rect 14240 12316 14246 12368
rect 14918 12316 14924 12368
rect 14976 12356 14982 12368
rect 15930 12356 15936 12368
rect 14976 12328 15936 12356
rect 14976 12316 14982 12328
rect 13906 12248 13912 12300
rect 13964 12288 13970 12300
rect 15396 12297 15424 12328
rect 15930 12316 15936 12328
rect 15988 12316 15994 12368
rect 18132 12359 18190 12365
rect 18132 12325 18144 12359
rect 18178 12356 18190 12359
rect 18690 12356 18696 12368
rect 18178 12328 18696 12356
rect 18178 12325 18190 12328
rect 18132 12319 18190 12325
rect 18690 12316 18696 12328
rect 18748 12316 18754 12368
rect 19426 12316 19432 12368
rect 19484 12356 19490 12368
rect 20070 12356 20076 12368
rect 19484 12328 20076 12356
rect 19484 12316 19490 12328
rect 20070 12316 20076 12328
rect 20128 12316 20134 12368
rect 20990 12316 20996 12368
rect 21048 12356 21054 12368
rect 21453 12359 21511 12365
rect 21453 12356 21465 12359
rect 21048 12328 21465 12356
rect 21048 12316 21054 12328
rect 21453 12325 21465 12328
rect 21499 12356 21511 12359
rect 21542 12356 21548 12368
rect 21499 12328 21548 12356
rect 21499 12325 21511 12328
rect 21453 12319 21511 12325
rect 21542 12316 21548 12328
rect 21600 12316 21606 12368
rect 15381 12291 15439 12297
rect 13964 12260 14009 12288
rect 13964 12248 13970 12260
rect 15381 12257 15393 12291
rect 15427 12257 15439 12291
rect 15381 12251 15439 12257
rect 15648 12291 15706 12297
rect 15648 12257 15660 12291
rect 15694 12288 15706 12291
rect 17034 12288 17040 12300
rect 15694 12260 17040 12288
rect 15694 12257 15706 12260
rect 15648 12251 15706 12257
rect 17034 12248 17040 12260
rect 17092 12248 17098 12300
rect 17126 12248 17132 12300
rect 17184 12288 17190 12300
rect 17865 12291 17923 12297
rect 17865 12288 17877 12291
rect 17184 12260 17877 12288
rect 17184 12248 17190 12260
rect 17865 12257 17877 12260
rect 17911 12288 17923 12291
rect 17954 12288 17960 12300
rect 17911 12260 17960 12288
rect 17911 12257 17923 12260
rect 17865 12251 17923 12257
rect 17954 12248 17960 12260
rect 18012 12248 18018 12300
rect 20714 12248 20720 12300
rect 20772 12288 20778 12300
rect 21266 12288 21272 12300
rect 20772 12260 21272 12288
rect 20772 12248 20778 12260
rect 21266 12248 21272 12260
rect 21324 12248 21330 12300
rect 22738 12297 22744 12300
rect 22732 12251 22744 12297
rect 22796 12288 22802 12300
rect 22796 12260 22832 12288
rect 22738 12248 22744 12251
rect 22796 12248 22802 12260
rect 12158 12220 12164 12232
rect 12119 12192 12164 12220
rect 12158 12180 12164 12192
rect 12216 12180 12222 12232
rect 13722 12220 13728 12232
rect 13683 12192 13728 12220
rect 13722 12180 13728 12192
rect 13780 12180 13786 12232
rect 20254 12180 20260 12232
rect 20312 12220 20318 12232
rect 20898 12220 20904 12232
rect 20312 12192 20904 12220
rect 20312 12180 20318 12192
rect 20898 12180 20904 12192
rect 20956 12180 20962 12232
rect 21542 12220 21548 12232
rect 21503 12192 21548 12220
rect 21542 12180 21548 12192
rect 21600 12180 21606 12232
rect 22465 12223 22523 12229
rect 22465 12189 22477 12223
rect 22511 12189 22523 12223
rect 22465 12183 22523 12189
rect 12989 12155 13047 12161
rect 12989 12121 13001 12155
rect 13035 12152 13047 12155
rect 13538 12152 13544 12164
rect 13035 12124 13544 12152
rect 13035 12121 13047 12124
rect 12989 12115 13047 12121
rect 13538 12112 13544 12124
rect 13596 12112 13602 12164
rect 20806 12112 20812 12164
rect 20864 12152 20870 12164
rect 20993 12155 21051 12161
rect 20993 12152 21005 12155
rect 20864 12124 21005 12152
rect 20864 12112 20870 12124
rect 20993 12121 21005 12124
rect 21039 12121 21051 12155
rect 20993 12115 21051 12121
rect 11790 12084 11796 12096
rect 11751 12056 11796 12084
rect 11790 12044 11796 12056
rect 11848 12044 11854 12096
rect 13354 12084 13360 12096
rect 13315 12056 13360 12084
rect 13354 12044 13360 12056
rect 13412 12044 13418 12096
rect 13446 12044 13452 12096
rect 13504 12084 13510 12096
rect 14277 12087 14335 12093
rect 14277 12084 14289 12087
rect 13504 12056 14289 12084
rect 13504 12044 13510 12056
rect 14277 12053 14289 12056
rect 14323 12053 14335 12087
rect 14734 12084 14740 12096
rect 14695 12056 14740 12084
rect 14277 12047 14335 12053
rect 14734 12044 14740 12056
rect 14792 12044 14798 12096
rect 15105 12087 15163 12093
rect 15105 12053 15117 12087
rect 15151 12084 15163 12087
rect 15378 12084 15384 12096
rect 15151 12056 15384 12084
rect 15151 12053 15163 12056
rect 15105 12047 15163 12053
rect 15378 12044 15384 12056
rect 15436 12084 15442 12096
rect 16761 12087 16819 12093
rect 16761 12084 16773 12087
rect 15436 12056 16773 12084
rect 15436 12044 15442 12056
rect 16761 12053 16773 12056
rect 16807 12053 16819 12087
rect 16761 12047 16819 12053
rect 20165 12087 20223 12093
rect 20165 12053 20177 12087
rect 20211 12084 20223 12087
rect 20717 12087 20775 12093
rect 20717 12084 20729 12087
rect 20211 12056 20729 12084
rect 20211 12053 20223 12056
rect 20165 12047 20223 12053
rect 20717 12053 20729 12056
rect 20763 12084 20775 12087
rect 21174 12084 21180 12096
rect 20763 12056 21180 12084
rect 20763 12053 20775 12056
rect 20717 12047 20775 12053
rect 21174 12044 21180 12056
rect 21232 12044 21238 12096
rect 21910 12044 21916 12096
rect 21968 12084 21974 12096
rect 22005 12087 22063 12093
rect 22005 12084 22017 12087
rect 21968 12056 22017 12084
rect 21968 12044 21974 12056
rect 22005 12053 22017 12056
rect 22051 12084 22063 12087
rect 22480 12084 22508 12183
rect 24302 12112 24308 12164
rect 24360 12112 24366 12164
rect 22051 12056 22508 12084
rect 22051 12053 22063 12056
rect 22005 12047 22063 12053
rect 23658 12044 23664 12096
rect 23716 12084 23722 12096
rect 24320 12084 24348 12112
rect 24397 12087 24455 12093
rect 24397 12084 24409 12087
rect 23716 12056 24409 12084
rect 23716 12044 23722 12056
rect 24397 12053 24409 12056
rect 24443 12084 24455 12087
rect 24854 12084 24860 12096
rect 24443 12056 24860 12084
rect 24443 12053 24455 12056
rect 24397 12047 24455 12053
rect 24854 12044 24860 12056
rect 24912 12044 24918 12096
rect 25130 12084 25136 12096
rect 25091 12056 25136 12084
rect 25130 12044 25136 12056
rect 25188 12044 25194 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 11793 11883 11851 11889
rect 11793 11849 11805 11883
rect 11839 11880 11851 11883
rect 12066 11880 12072 11892
rect 11839 11852 12072 11880
rect 11839 11849 11851 11852
rect 11793 11843 11851 11849
rect 12066 11840 12072 11852
rect 12124 11840 12130 11892
rect 12161 11883 12219 11889
rect 12161 11849 12173 11883
rect 12207 11880 12219 11883
rect 12250 11880 12256 11892
rect 12207 11852 12256 11880
rect 12207 11849 12219 11852
rect 12161 11843 12219 11849
rect 12250 11840 12256 11852
rect 12308 11840 12314 11892
rect 12805 11883 12863 11889
rect 12805 11849 12817 11883
rect 12851 11880 12863 11883
rect 13814 11880 13820 11892
rect 12851 11852 13820 11880
rect 12851 11849 12863 11852
rect 12805 11843 12863 11849
rect 13814 11840 13820 11852
rect 13872 11840 13878 11892
rect 13906 11840 13912 11892
rect 13964 11880 13970 11892
rect 14277 11883 14335 11889
rect 14277 11880 14289 11883
rect 13964 11852 14289 11880
rect 13964 11840 13970 11852
rect 14277 11849 14289 11852
rect 14323 11849 14335 11883
rect 14277 11843 14335 11849
rect 15746 11840 15752 11892
rect 15804 11880 15810 11892
rect 16209 11883 16267 11889
rect 16209 11880 16221 11883
rect 15804 11852 16221 11880
rect 15804 11840 15810 11852
rect 16209 11849 16221 11852
rect 16255 11880 16267 11883
rect 17497 11883 17555 11889
rect 16255 11852 16896 11880
rect 16255 11849 16267 11852
rect 16209 11843 16267 11849
rect 12986 11812 12992 11824
rect 12947 11784 12992 11812
rect 12986 11772 12992 11784
rect 13044 11772 13050 11824
rect 14826 11772 14832 11824
rect 14884 11812 14890 11824
rect 14921 11815 14979 11821
rect 14921 11812 14933 11815
rect 14884 11784 14933 11812
rect 14884 11772 14890 11784
rect 14921 11781 14933 11784
rect 14967 11781 14979 11815
rect 14921 11775 14979 11781
rect 16485 11815 16543 11821
rect 16485 11781 16497 11815
rect 16531 11781 16543 11815
rect 16485 11775 16543 11781
rect 11790 11704 11796 11756
rect 11848 11744 11854 11756
rect 13357 11747 13415 11753
rect 13357 11744 13369 11747
rect 11848 11716 13369 11744
rect 11848 11704 11854 11716
rect 13357 11713 13369 11716
rect 13403 11744 13415 11747
rect 13446 11744 13452 11756
rect 13403 11716 13452 11744
rect 13403 11713 13415 11716
rect 13357 11707 13415 11713
rect 13446 11704 13452 11716
rect 13504 11704 13510 11756
rect 13538 11704 13544 11756
rect 13596 11744 13602 11756
rect 14645 11747 14703 11753
rect 13596 11716 13641 11744
rect 13596 11704 13602 11716
rect 14645 11713 14657 11747
rect 14691 11744 14703 11747
rect 15378 11744 15384 11756
rect 14691 11716 15384 11744
rect 14691 11713 14703 11716
rect 14645 11707 14703 11713
rect 15378 11704 15384 11716
rect 15436 11744 15442 11756
rect 15473 11747 15531 11753
rect 15473 11744 15485 11747
rect 15436 11716 15485 11744
rect 15436 11704 15442 11716
rect 15473 11713 15485 11716
rect 15519 11713 15531 11747
rect 15473 11707 15531 11713
rect 14734 11636 14740 11688
rect 14792 11676 14798 11688
rect 15197 11679 15255 11685
rect 15197 11676 15209 11679
rect 14792 11648 15209 11676
rect 14792 11636 14798 11648
rect 15197 11645 15209 11648
rect 15243 11676 15255 11679
rect 16500 11676 16528 11775
rect 16868 11753 16896 11852
rect 17497 11849 17509 11883
rect 17543 11880 17555 11883
rect 17586 11880 17592 11892
rect 17543 11852 17592 11880
rect 17543 11849 17555 11852
rect 17497 11843 17555 11849
rect 17586 11840 17592 11852
rect 17644 11880 17650 11892
rect 20625 11883 20683 11889
rect 17644 11852 18552 11880
rect 17644 11840 17650 11852
rect 18141 11815 18199 11821
rect 18141 11781 18153 11815
rect 18187 11781 18199 11815
rect 18141 11775 18199 11781
rect 16853 11747 16911 11753
rect 16853 11713 16865 11747
rect 16899 11713 16911 11747
rect 17034 11744 17040 11756
rect 16995 11716 17040 11744
rect 16853 11707 16911 11713
rect 17034 11704 17040 11716
rect 17092 11704 17098 11756
rect 18156 11676 18184 11775
rect 15243 11648 16528 11676
rect 16960 11648 18184 11676
rect 15243 11645 15255 11648
rect 15197 11639 15255 11645
rect 13170 11568 13176 11620
rect 13228 11608 13234 11620
rect 13722 11608 13728 11620
rect 13228 11580 13728 11608
rect 13228 11568 13234 11580
rect 13722 11568 13728 11580
rect 13780 11608 13786 11620
rect 13909 11611 13967 11617
rect 13909 11608 13921 11611
rect 13780 11580 13921 11608
rect 13780 11568 13786 11580
rect 13909 11577 13921 11580
rect 13955 11577 13967 11611
rect 13909 11571 13967 11577
rect 14918 11568 14924 11620
rect 14976 11608 14982 11620
rect 15381 11611 15439 11617
rect 15381 11608 15393 11611
rect 14976 11580 15393 11608
rect 14976 11568 14982 11580
rect 15381 11577 15393 11580
rect 15427 11608 15439 11611
rect 15562 11608 15568 11620
rect 15427 11580 15568 11608
rect 15427 11577 15439 11580
rect 15381 11571 15439 11577
rect 15562 11568 15568 11580
rect 15620 11568 15626 11620
rect 16022 11568 16028 11620
rect 16080 11608 16086 11620
rect 16960 11617 16988 11648
rect 16945 11611 17003 11617
rect 16945 11608 16957 11611
rect 16080 11580 16957 11608
rect 16080 11568 16086 11580
rect 16945 11577 16957 11580
rect 16991 11577 17003 11611
rect 18417 11611 18475 11617
rect 18417 11608 18429 11611
rect 16945 11571 17003 11577
rect 17788 11580 18429 11608
rect 17788 11552 17816 11580
rect 18417 11577 18429 11580
rect 18463 11577 18475 11611
rect 18524 11608 18552 11852
rect 20625 11849 20637 11883
rect 20671 11880 20683 11883
rect 20714 11880 20720 11892
rect 20671 11852 20720 11880
rect 20671 11849 20683 11852
rect 20625 11843 20683 11849
rect 20714 11840 20720 11852
rect 20772 11840 20778 11892
rect 20990 11880 20996 11892
rect 20951 11852 20996 11880
rect 20990 11840 20996 11852
rect 21048 11840 21054 11892
rect 22465 11883 22523 11889
rect 22465 11849 22477 11883
rect 22511 11880 22523 11883
rect 22738 11880 22744 11892
rect 22511 11852 22744 11880
rect 22511 11849 22523 11852
rect 22465 11843 22523 11849
rect 22738 11840 22744 11852
rect 22796 11840 22802 11892
rect 23477 11883 23535 11889
rect 23477 11849 23489 11883
rect 23523 11880 23535 11883
rect 23566 11880 23572 11892
rect 23523 11852 23572 11880
rect 23523 11849 23535 11852
rect 23477 11843 23535 11849
rect 23566 11840 23572 11852
rect 23624 11840 23630 11892
rect 24854 11840 24860 11892
rect 24912 11880 24918 11892
rect 25501 11883 25559 11889
rect 25501 11880 25513 11883
rect 24912 11852 25513 11880
rect 24912 11840 24918 11852
rect 25501 11849 25513 11852
rect 25547 11849 25559 11883
rect 25501 11843 25559 11849
rect 20073 11747 20131 11753
rect 20073 11713 20085 11747
rect 20119 11744 20131 11747
rect 20622 11744 20628 11756
rect 20119 11716 20628 11744
rect 20119 11713 20131 11716
rect 20073 11707 20131 11713
rect 20622 11704 20628 11716
rect 20680 11704 20686 11756
rect 23584 11744 23612 11840
rect 23584 11716 24256 11744
rect 20898 11636 20904 11688
rect 20956 11676 20962 11688
rect 21085 11679 21143 11685
rect 21085 11676 21097 11679
rect 20956 11648 21097 11676
rect 20956 11636 20962 11648
rect 21085 11645 21097 11648
rect 21131 11676 21143 11679
rect 21910 11676 21916 11688
rect 21131 11648 21916 11676
rect 21131 11645 21143 11648
rect 21085 11639 21143 11645
rect 21910 11636 21916 11648
rect 21968 11676 21974 11688
rect 23017 11679 23075 11685
rect 23017 11676 23029 11679
rect 21968 11648 23029 11676
rect 21968 11636 21974 11648
rect 23017 11645 23029 11648
rect 23063 11676 23075 11679
rect 23934 11676 23940 11688
rect 23063 11648 23940 11676
rect 23063 11645 23075 11648
rect 23017 11639 23075 11645
rect 23934 11636 23940 11648
rect 23992 11676 23998 11688
rect 24121 11679 24179 11685
rect 24121 11676 24133 11679
rect 23992 11648 24133 11676
rect 23992 11636 23998 11648
rect 24121 11645 24133 11648
rect 24167 11645 24179 11679
rect 24228 11676 24256 11716
rect 24377 11679 24435 11685
rect 24377 11676 24389 11679
rect 24228 11648 24389 11676
rect 24121 11639 24179 11645
rect 24377 11645 24389 11648
rect 24423 11645 24435 11679
rect 24377 11639 24435 11645
rect 18601 11611 18659 11617
rect 18601 11608 18613 11611
rect 18524 11580 18613 11608
rect 18417 11571 18475 11577
rect 18601 11577 18613 11580
rect 18647 11577 18659 11611
rect 18601 11571 18659 11577
rect 18693 11611 18751 11617
rect 18693 11577 18705 11611
rect 18739 11577 18751 11611
rect 18693 11571 18751 11577
rect 11425 11543 11483 11549
rect 11425 11509 11437 11543
rect 11471 11540 11483 11543
rect 11514 11540 11520 11552
rect 11471 11512 11520 11540
rect 11471 11509 11483 11512
rect 11425 11503 11483 11509
rect 11514 11500 11520 11512
rect 11572 11500 11578 11552
rect 13446 11540 13452 11552
rect 13407 11512 13452 11540
rect 13446 11500 13452 11512
rect 13504 11500 13510 11552
rect 15930 11540 15936 11552
rect 15891 11512 15936 11540
rect 15930 11500 15936 11512
rect 15988 11500 15994 11552
rect 17770 11540 17776 11552
rect 17731 11512 17776 11540
rect 17770 11500 17776 11512
rect 17828 11500 17834 11552
rect 18708 11540 18736 11571
rect 20346 11568 20352 11620
rect 20404 11608 20410 11620
rect 20622 11608 20628 11620
rect 20404 11580 20628 11608
rect 20404 11568 20410 11580
rect 20622 11568 20628 11580
rect 20680 11568 20686 11620
rect 21174 11568 21180 11620
rect 21232 11608 21238 11620
rect 21352 11611 21410 11617
rect 21352 11608 21364 11611
rect 21232 11580 21364 11608
rect 21232 11568 21238 11580
rect 21352 11577 21364 11580
rect 21398 11608 21410 11611
rect 22278 11608 22284 11620
rect 21398 11580 22284 11608
rect 21398 11577 21410 11580
rect 21352 11571 21410 11577
rect 22278 11568 22284 11580
rect 22336 11568 22342 11620
rect 19153 11543 19211 11549
rect 19153 11540 19165 11543
rect 18708 11512 19165 11540
rect 19153 11509 19165 11512
rect 19199 11540 19211 11543
rect 19426 11540 19432 11552
rect 19199 11512 19432 11540
rect 19199 11509 19211 11512
rect 19153 11503 19211 11509
rect 19426 11500 19432 11512
rect 19484 11500 19490 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 13446 11336 13452 11348
rect 12268 11308 13452 11336
rect 11330 11228 11336 11280
rect 11388 11268 11394 11280
rect 11425 11271 11483 11277
rect 11425 11268 11437 11271
rect 11388 11240 11437 11268
rect 11388 11228 11394 11240
rect 11425 11237 11437 11240
rect 11471 11268 11483 11271
rect 11790 11268 11796 11280
rect 11471 11240 11796 11268
rect 11471 11237 11483 11240
rect 11425 11231 11483 11237
rect 11790 11228 11796 11240
rect 11848 11228 11854 11280
rect 11146 11160 11152 11212
rect 11204 11200 11210 11212
rect 11241 11203 11299 11209
rect 11241 11200 11253 11203
rect 11204 11172 11253 11200
rect 11204 11160 11210 11172
rect 11241 11169 11253 11172
rect 11287 11169 11299 11203
rect 11241 11163 11299 11169
rect 11514 11132 11520 11144
rect 11475 11104 11520 11132
rect 11514 11092 11520 11104
rect 11572 11092 11578 11144
rect 12268 11073 12296 11308
rect 13446 11296 13452 11308
rect 13504 11296 13510 11348
rect 13538 11296 13544 11348
rect 13596 11336 13602 11348
rect 13817 11339 13875 11345
rect 13817 11336 13829 11339
rect 13596 11308 13829 11336
rect 13596 11296 13602 11308
rect 13817 11305 13829 11308
rect 13863 11305 13875 11339
rect 14918 11336 14924 11348
rect 14879 11308 14924 11336
rect 13817 11299 13875 11305
rect 14918 11296 14924 11308
rect 14976 11296 14982 11348
rect 16022 11336 16028 11348
rect 15983 11308 16028 11336
rect 16022 11296 16028 11308
rect 16080 11296 16086 11348
rect 16393 11339 16451 11345
rect 16393 11305 16405 11339
rect 16439 11336 16451 11339
rect 16942 11336 16948 11348
rect 16439 11308 16948 11336
rect 16439 11305 16451 11308
rect 16393 11299 16451 11305
rect 15565 11271 15623 11277
rect 15565 11237 15577 11271
rect 15611 11268 15623 11271
rect 16408 11268 16436 11299
rect 16942 11296 16948 11308
rect 17000 11296 17006 11348
rect 18601 11339 18659 11345
rect 18601 11305 18613 11339
rect 18647 11336 18659 11339
rect 18874 11336 18880 11348
rect 18647 11308 18880 11336
rect 18647 11305 18659 11308
rect 18601 11299 18659 11305
rect 18874 11296 18880 11308
rect 18932 11296 18938 11348
rect 22278 11336 22284 11348
rect 22239 11308 22284 11336
rect 22278 11296 22284 11308
rect 22336 11296 22342 11348
rect 22738 11296 22744 11348
rect 22796 11336 22802 11348
rect 22833 11339 22891 11345
rect 22833 11336 22845 11339
rect 22796 11308 22845 11336
rect 22796 11296 22802 11308
rect 22833 11305 22845 11308
rect 22879 11305 22891 11339
rect 22833 11299 22891 11305
rect 17037 11271 17095 11277
rect 17037 11268 17049 11271
rect 15611 11240 16436 11268
rect 16500 11240 17049 11268
rect 15611 11237 15623 11240
rect 15565 11231 15623 11237
rect 12342 11160 12348 11212
rect 12400 11200 12406 11212
rect 12693 11203 12751 11209
rect 12693 11200 12705 11203
rect 12400 11172 12705 11200
rect 12400 11160 12406 11172
rect 12693 11169 12705 11172
rect 12739 11169 12751 11203
rect 12693 11163 12751 11169
rect 12434 11132 12440 11144
rect 12395 11104 12440 11132
rect 12434 11092 12440 11104
rect 12492 11092 12498 11144
rect 10965 11067 11023 11073
rect 10965 11033 10977 11067
rect 11011 11064 11023 11067
rect 12253 11067 12311 11073
rect 12253 11064 12265 11067
rect 11011 11036 12265 11064
rect 11011 11033 11023 11036
rect 10965 11027 11023 11033
rect 12253 11033 12265 11036
rect 12299 11033 12311 11067
rect 12253 11027 12311 11033
rect 15562 10956 15568 11008
rect 15620 10996 15626 11008
rect 16500 10996 16528 11240
rect 17037 11237 17049 11240
rect 17083 11237 17095 11271
rect 17037 11231 17095 11237
rect 20717 11271 20775 11277
rect 20717 11237 20729 11271
rect 20763 11268 20775 11271
rect 20806 11268 20812 11280
rect 20763 11240 20812 11268
rect 20763 11237 20775 11240
rect 20717 11231 20775 11237
rect 20806 11228 20812 11240
rect 20864 11268 20870 11280
rect 21168 11271 21226 11277
rect 21168 11268 21180 11271
rect 20864 11240 21180 11268
rect 20864 11228 20870 11240
rect 21168 11237 21180 11240
rect 21214 11268 21226 11271
rect 21542 11268 21548 11280
rect 21214 11240 21548 11268
rect 21214 11237 21226 11240
rect 21168 11231 21226 11237
rect 21542 11228 21548 11240
rect 21600 11228 21606 11280
rect 16574 11160 16580 11212
rect 16632 11200 16638 11212
rect 16853 11203 16911 11209
rect 16853 11200 16865 11203
rect 16632 11172 16865 11200
rect 16632 11160 16638 11172
rect 16853 11169 16865 11172
rect 16899 11169 16911 11203
rect 16853 11163 16911 11169
rect 18417 11203 18475 11209
rect 18417 11169 18429 11203
rect 18463 11200 18475 11203
rect 18782 11200 18788 11212
rect 18463 11172 18788 11200
rect 18463 11169 18475 11172
rect 18417 11163 18475 11169
rect 16577 11067 16635 11073
rect 16577 11033 16589 11067
rect 16623 11064 16635 11067
rect 16758 11064 16764 11076
rect 16623 11036 16764 11064
rect 16623 11033 16635 11036
rect 16577 11027 16635 11033
rect 16758 11024 16764 11036
rect 16816 11024 16822 11076
rect 16868 11064 16896 11163
rect 18782 11160 18788 11172
rect 18840 11200 18846 11212
rect 19058 11200 19064 11212
rect 18840 11172 19064 11200
rect 18840 11160 18846 11172
rect 19058 11160 19064 11172
rect 19116 11160 19122 11212
rect 20898 11200 20904 11212
rect 20859 11172 20904 11200
rect 20898 11160 20904 11172
rect 20956 11160 20962 11212
rect 23934 11200 23940 11212
rect 23895 11172 23940 11200
rect 23934 11160 23940 11172
rect 23992 11160 23998 11212
rect 24193 11203 24251 11209
rect 24193 11200 24205 11203
rect 24044 11172 24205 11200
rect 17129 11135 17187 11141
rect 17129 11101 17141 11135
rect 17175 11132 17187 11135
rect 17310 11132 17316 11144
rect 17175 11104 17316 11132
rect 17175 11101 17187 11104
rect 17129 11095 17187 11101
rect 17310 11092 17316 11104
rect 17368 11092 17374 11144
rect 17954 11092 17960 11144
rect 18012 11132 18018 11144
rect 18693 11135 18751 11141
rect 18693 11132 18705 11135
rect 18012 11104 18705 11132
rect 18012 11092 18018 11104
rect 18693 11101 18705 11104
rect 18739 11101 18751 11135
rect 18693 11095 18751 11101
rect 19797 11135 19855 11141
rect 19797 11101 19809 11135
rect 19843 11132 19855 11135
rect 20714 11132 20720 11144
rect 19843 11104 20720 11132
rect 19843 11101 19855 11104
rect 19797 11095 19855 11101
rect 20714 11092 20720 11104
rect 20772 11092 20778 11144
rect 24044 11132 24072 11172
rect 24193 11169 24205 11172
rect 24239 11169 24251 11203
rect 24193 11163 24251 11169
rect 23676 11104 24072 11132
rect 18141 11067 18199 11073
rect 18141 11064 18153 11067
rect 16868 11036 18153 11064
rect 18141 11033 18153 11036
rect 18187 11033 18199 11067
rect 22738 11064 22744 11076
rect 18141 11027 18199 11033
rect 22112 11036 22744 11064
rect 17586 10996 17592 11008
rect 15620 10968 16528 10996
rect 17547 10968 17592 10996
rect 15620 10956 15626 10968
rect 17586 10956 17592 10968
rect 17644 10956 17650 11008
rect 17957 10999 18015 11005
rect 17957 10965 17969 10999
rect 18003 10996 18015 10999
rect 18046 10996 18052 11008
rect 18003 10968 18052 10996
rect 18003 10965 18015 10968
rect 17957 10959 18015 10965
rect 18046 10956 18052 10968
rect 18104 10996 18110 11008
rect 19061 10999 19119 11005
rect 19061 10996 19073 10999
rect 18104 10968 19073 10996
rect 18104 10956 18110 10968
rect 19061 10965 19073 10968
rect 19107 10965 19119 10999
rect 19061 10959 19119 10965
rect 21542 10956 21548 11008
rect 21600 10996 21606 11008
rect 22112 10996 22140 11036
rect 22738 11024 22744 11036
rect 22796 11024 22802 11076
rect 23676 11008 23704 11104
rect 24946 11024 24952 11076
rect 25004 11064 25010 11076
rect 25317 11067 25375 11073
rect 25317 11064 25329 11067
rect 25004 11036 25329 11064
rect 25004 11024 25010 11036
rect 25317 11033 25329 11036
rect 25363 11033 25375 11067
rect 25317 11027 25375 11033
rect 23658 10996 23664 11008
rect 21600 10968 22140 10996
rect 23619 10968 23664 10996
rect 21600 10956 21606 10968
rect 23658 10956 23664 10968
rect 23716 10956 23722 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 17865 10795 17923 10801
rect 17865 10761 17877 10795
rect 17911 10792 17923 10795
rect 17954 10792 17960 10804
rect 17911 10764 17960 10792
rect 17911 10761 17923 10764
rect 17865 10755 17923 10761
rect 17954 10752 17960 10764
rect 18012 10752 18018 10804
rect 18693 10795 18751 10801
rect 18693 10761 18705 10795
rect 18739 10792 18751 10795
rect 18782 10792 18788 10804
rect 18739 10764 18788 10792
rect 18739 10761 18751 10764
rect 18693 10755 18751 10761
rect 18782 10752 18788 10764
rect 18840 10752 18846 10804
rect 19886 10752 19892 10804
rect 19944 10792 19950 10804
rect 20162 10792 20168 10804
rect 19944 10764 20168 10792
rect 19944 10752 19950 10764
rect 20162 10752 20168 10764
rect 20220 10752 20226 10804
rect 20530 10752 20536 10804
rect 20588 10792 20594 10804
rect 21545 10795 21603 10801
rect 21545 10792 21557 10795
rect 20588 10764 21557 10792
rect 20588 10752 20594 10764
rect 21545 10761 21557 10764
rect 21591 10761 21603 10795
rect 21545 10755 21603 10761
rect 22094 10752 22100 10804
rect 22152 10792 22158 10804
rect 22465 10795 22523 10801
rect 22465 10792 22477 10795
rect 22152 10764 22477 10792
rect 22152 10752 22158 10764
rect 22465 10761 22477 10764
rect 22511 10761 22523 10795
rect 22465 10755 22523 10761
rect 23109 10795 23167 10801
rect 23109 10761 23121 10795
rect 23155 10792 23167 10795
rect 23658 10792 23664 10804
rect 23155 10764 23664 10792
rect 23155 10761 23167 10764
rect 23109 10755 23167 10761
rect 23658 10752 23664 10764
rect 23716 10752 23722 10804
rect 23934 10752 23940 10804
rect 23992 10792 23998 10804
rect 24765 10795 24823 10801
rect 24765 10792 24777 10795
rect 23992 10764 24777 10792
rect 23992 10752 23998 10764
rect 24765 10761 24777 10764
rect 24811 10761 24823 10795
rect 24765 10755 24823 10761
rect 16485 10727 16543 10733
rect 16485 10693 16497 10727
rect 16531 10724 16543 10727
rect 16574 10724 16580 10736
rect 16531 10696 16580 10724
rect 16531 10693 16543 10696
rect 16485 10687 16543 10693
rect 16574 10684 16580 10696
rect 16632 10684 16638 10736
rect 18325 10727 18383 10733
rect 18325 10693 18337 10727
rect 18371 10724 18383 10727
rect 18874 10724 18880 10736
rect 18371 10696 18880 10724
rect 18371 10693 18383 10696
rect 18325 10687 18383 10693
rect 18874 10684 18880 10696
rect 18932 10684 18938 10736
rect 20349 10727 20407 10733
rect 20349 10693 20361 10727
rect 20395 10724 20407 10727
rect 20806 10724 20812 10736
rect 20395 10696 20812 10724
rect 20395 10693 20407 10696
rect 20349 10687 20407 10693
rect 20806 10684 20812 10696
rect 20864 10684 20870 10736
rect 21266 10724 21272 10736
rect 21227 10696 21272 10724
rect 21266 10684 21272 10696
rect 21324 10724 21330 10736
rect 23753 10727 23811 10733
rect 21324 10696 21956 10724
rect 21324 10684 21330 10696
rect 12434 10616 12440 10668
rect 12492 10616 12498 10668
rect 15933 10659 15991 10665
rect 15933 10625 15945 10659
rect 15979 10656 15991 10659
rect 17037 10659 17095 10665
rect 17037 10656 17049 10659
rect 15979 10628 17049 10656
rect 15979 10625 15991 10628
rect 15933 10619 15991 10625
rect 17037 10625 17049 10628
rect 17083 10656 17095 10659
rect 17310 10656 17316 10668
rect 17083 10628 17316 10656
rect 17083 10625 17095 10628
rect 17037 10619 17095 10625
rect 17310 10616 17316 10628
rect 17368 10656 17374 10668
rect 17405 10659 17463 10665
rect 17405 10656 17417 10659
rect 17368 10628 17417 10656
rect 17368 10616 17374 10628
rect 17405 10625 17417 10628
rect 17451 10625 17463 10659
rect 17405 10619 17463 10625
rect 18046 10616 18052 10668
rect 18104 10656 18110 10668
rect 18969 10659 19027 10665
rect 18969 10656 18981 10659
rect 18104 10628 18981 10656
rect 18104 10616 18110 10628
rect 18969 10625 18981 10628
rect 19015 10625 19027 10659
rect 18969 10619 19027 10625
rect 19978 10616 19984 10668
rect 20036 10656 20042 10668
rect 21358 10656 21364 10668
rect 20036 10628 21364 10656
rect 20036 10616 20042 10628
rect 21358 10616 21364 10628
rect 21416 10616 21422 10668
rect 21928 10665 21956 10696
rect 23753 10693 23765 10727
rect 23799 10724 23811 10727
rect 24670 10724 24676 10736
rect 23799 10696 24676 10724
rect 23799 10693 23811 10696
rect 23753 10687 23811 10693
rect 24670 10684 24676 10696
rect 24728 10684 24734 10736
rect 21913 10659 21971 10665
rect 21913 10625 21925 10659
rect 21959 10656 21971 10659
rect 22002 10656 22008 10668
rect 21959 10628 22008 10656
rect 21959 10625 21971 10628
rect 21913 10619 21971 10625
rect 22002 10616 22008 10628
rect 22060 10616 22066 10668
rect 23477 10659 23535 10665
rect 23477 10625 23489 10659
rect 23523 10656 23535 10659
rect 24118 10656 24124 10668
rect 23523 10628 24124 10656
rect 23523 10625 23535 10628
rect 23477 10619 23535 10625
rect 24118 10616 24124 10628
rect 24176 10616 24182 10668
rect 10594 10588 10600 10600
rect 10555 10560 10600 10588
rect 10594 10548 10600 10560
rect 10652 10548 10658 10600
rect 12452 10588 12480 10616
rect 13538 10597 13544 10600
rect 12713 10591 12771 10597
rect 12713 10588 12725 10591
rect 12452 10560 12725 10588
rect 12713 10557 12725 10560
rect 12759 10588 12771 10591
rect 13173 10591 13231 10597
rect 13173 10588 13185 10591
rect 12759 10560 13185 10588
rect 12759 10557 12771 10560
rect 12713 10551 12771 10557
rect 13173 10557 13185 10560
rect 13219 10588 13231 10591
rect 13265 10591 13323 10597
rect 13265 10588 13277 10591
rect 13219 10560 13277 10588
rect 13219 10557 13231 10560
rect 13173 10551 13231 10557
rect 13265 10557 13277 10560
rect 13311 10557 13323 10591
rect 13532 10588 13544 10597
rect 13499 10560 13544 10588
rect 13265 10551 13323 10557
rect 13532 10551 13544 10560
rect 11333 10523 11391 10529
rect 11333 10489 11345 10523
rect 11379 10520 11391 10523
rect 12434 10520 12440 10532
rect 11379 10492 12440 10520
rect 11379 10489 11391 10492
rect 11333 10483 11391 10489
rect 12434 10480 12440 10492
rect 12492 10480 12498 10532
rect 13280 10520 13308 10551
rect 13538 10548 13544 10551
rect 13596 10548 13602 10600
rect 17586 10588 17592 10600
rect 16960 10560 17592 10588
rect 16022 10520 16028 10532
rect 13280 10492 16028 10520
rect 16022 10480 16028 10492
rect 16080 10480 16086 10532
rect 16301 10523 16359 10529
rect 16301 10489 16313 10523
rect 16347 10520 16359 10523
rect 16758 10520 16764 10532
rect 16347 10492 16764 10520
rect 16347 10489 16359 10492
rect 16301 10483 16359 10489
rect 16758 10480 16764 10492
rect 16816 10480 16822 10532
rect 16960 10529 16988 10560
rect 17586 10548 17592 10560
rect 17644 10548 17650 10600
rect 23658 10548 23664 10600
rect 23716 10588 23722 10600
rect 24305 10591 24363 10597
rect 24305 10588 24317 10591
rect 23716 10560 24317 10588
rect 23716 10548 23722 10560
rect 24305 10557 24317 10560
rect 24351 10557 24363 10591
rect 25222 10588 25228 10600
rect 25183 10560 25228 10588
rect 24305 10551 24363 10557
rect 25222 10548 25228 10560
rect 25280 10588 25286 10600
rect 25777 10591 25835 10597
rect 25777 10588 25789 10591
rect 25280 10560 25789 10588
rect 25280 10548 25286 10560
rect 25777 10557 25789 10560
rect 25823 10557 25835 10591
rect 25777 10551 25835 10557
rect 16945 10523 17003 10529
rect 16945 10489 16957 10523
rect 16991 10489 17003 10523
rect 16945 10483 17003 10489
rect 19150 10480 19156 10532
rect 19208 10529 19214 10532
rect 19208 10523 19272 10529
rect 19208 10489 19226 10523
rect 19260 10489 19272 10523
rect 20898 10520 20904 10532
rect 20859 10492 20904 10520
rect 19208 10483 19272 10489
rect 19208 10480 19214 10483
rect 20898 10480 20904 10492
rect 20956 10480 20962 10532
rect 22094 10480 22100 10532
rect 22152 10520 22158 10532
rect 22152 10492 22197 10520
rect 22152 10480 22158 10492
rect 10962 10452 10968 10464
rect 10923 10424 10968 10452
rect 10962 10412 10968 10424
rect 11020 10412 11026 10464
rect 12158 10452 12164 10464
rect 12119 10424 12164 10452
rect 12158 10412 12164 10424
rect 12216 10412 12222 10464
rect 14645 10455 14703 10461
rect 14645 10421 14657 10455
rect 14691 10452 14703 10455
rect 14734 10452 14740 10464
rect 14691 10424 14740 10452
rect 14691 10421 14703 10424
rect 14645 10415 14703 10421
rect 14734 10412 14740 10424
rect 14792 10412 14798 10464
rect 15562 10452 15568 10464
rect 15523 10424 15568 10452
rect 15562 10412 15568 10424
rect 15620 10412 15626 10464
rect 20916 10452 20944 10480
rect 22005 10455 22063 10461
rect 22005 10452 22017 10455
rect 20916 10424 22017 10452
rect 22005 10421 22017 10424
rect 22051 10421 22063 10455
rect 22005 10415 22063 10421
rect 23658 10412 23664 10464
rect 23716 10452 23722 10464
rect 24213 10455 24271 10461
rect 24213 10452 24225 10455
rect 23716 10424 24225 10452
rect 23716 10412 23722 10424
rect 24213 10421 24225 10424
rect 24259 10421 24271 10455
rect 24213 10415 24271 10421
rect 24762 10412 24768 10464
rect 24820 10452 24826 10464
rect 25409 10455 25467 10461
rect 25409 10452 25421 10455
rect 24820 10424 25421 10452
rect 24820 10412 24826 10424
rect 25409 10421 25421 10424
rect 25455 10421 25467 10455
rect 25409 10415 25467 10421
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 10965 10251 11023 10257
rect 10965 10217 10977 10251
rect 11011 10248 11023 10251
rect 11514 10248 11520 10260
rect 11011 10220 11520 10248
rect 11011 10217 11023 10220
rect 10965 10211 11023 10217
rect 11514 10208 11520 10220
rect 11572 10248 11578 10260
rect 12158 10248 12164 10260
rect 11572 10220 12164 10248
rect 11572 10208 11578 10220
rect 12158 10208 12164 10220
rect 12216 10208 12222 10260
rect 12986 10208 12992 10260
rect 13044 10248 13050 10260
rect 13541 10251 13599 10257
rect 13541 10248 13553 10251
rect 13044 10220 13553 10248
rect 13044 10208 13050 10220
rect 13541 10217 13553 10220
rect 13587 10248 13599 10251
rect 13814 10248 13820 10260
rect 13587 10220 13820 10248
rect 13587 10217 13599 10220
rect 13541 10211 13599 10217
rect 13814 10208 13820 10220
rect 13872 10208 13878 10260
rect 15841 10251 15899 10257
rect 15841 10217 15853 10251
rect 15887 10248 15899 10251
rect 16482 10248 16488 10260
rect 15887 10220 16488 10248
rect 15887 10217 15899 10220
rect 15841 10211 15899 10217
rect 16482 10208 16488 10220
rect 16540 10208 16546 10260
rect 17310 10248 17316 10260
rect 17271 10220 17316 10248
rect 17310 10208 17316 10220
rect 17368 10208 17374 10260
rect 18230 10208 18236 10260
rect 18288 10248 18294 10260
rect 18969 10251 19027 10257
rect 18969 10248 18981 10251
rect 18288 10220 18981 10248
rect 18288 10208 18294 10220
rect 18969 10217 18981 10220
rect 19015 10248 19027 10251
rect 19242 10248 19248 10260
rect 19015 10220 19248 10248
rect 19015 10217 19027 10220
rect 18969 10211 19027 10217
rect 19242 10208 19248 10220
rect 19300 10208 19306 10260
rect 20438 10208 20444 10260
rect 20496 10248 20502 10260
rect 21453 10251 21511 10257
rect 21453 10248 21465 10251
rect 20496 10220 21465 10248
rect 20496 10208 20502 10220
rect 21453 10217 21465 10220
rect 21499 10217 21511 10251
rect 22094 10248 22100 10260
rect 21453 10211 21511 10217
rect 21928 10220 22100 10248
rect 13630 10140 13636 10192
rect 13688 10180 13694 10192
rect 14001 10183 14059 10189
rect 14001 10180 14013 10183
rect 13688 10152 14013 10180
rect 13688 10140 13694 10152
rect 14001 10149 14013 10152
rect 14047 10149 14059 10183
rect 14001 10143 14059 10149
rect 17770 10140 17776 10192
rect 17828 10180 17834 10192
rect 18785 10183 18843 10189
rect 18785 10180 18797 10183
rect 17828 10152 18797 10180
rect 17828 10140 17834 10152
rect 18785 10149 18797 10152
rect 18831 10149 18843 10183
rect 18785 10143 18843 10149
rect 20717 10183 20775 10189
rect 20717 10149 20729 10183
rect 20763 10180 20775 10183
rect 20806 10180 20812 10192
rect 20763 10152 20812 10180
rect 20763 10149 20775 10152
rect 20717 10143 20775 10149
rect 20806 10140 20812 10152
rect 20864 10140 20870 10192
rect 21542 10180 21548 10192
rect 21503 10152 21548 10180
rect 21542 10140 21548 10152
rect 21600 10140 21606 10192
rect 16200 10115 16258 10121
rect 16200 10081 16212 10115
rect 16246 10112 16258 10115
rect 16942 10112 16948 10124
rect 16246 10084 16948 10112
rect 16246 10081 16258 10084
rect 16200 10075 16258 10081
rect 16942 10072 16948 10084
rect 17000 10112 17006 10124
rect 17954 10112 17960 10124
rect 17000 10084 17960 10112
rect 17000 10072 17006 10084
rect 17954 10072 17960 10084
rect 18012 10112 18018 10124
rect 18233 10115 18291 10121
rect 18233 10112 18245 10115
rect 18012 10084 18245 10112
rect 18012 10072 18018 10084
rect 18233 10081 18245 10084
rect 18279 10112 18291 10115
rect 19061 10115 19119 10121
rect 19061 10112 19073 10115
rect 18279 10084 19073 10112
rect 18279 10081 18291 10084
rect 18233 10075 18291 10081
rect 19061 10081 19073 10084
rect 19107 10081 19119 10115
rect 20824 10112 20852 10140
rect 21928 10121 21956 10220
rect 22094 10208 22100 10220
rect 22152 10208 22158 10260
rect 23017 10251 23075 10257
rect 23017 10217 23029 10251
rect 23063 10248 23075 10251
rect 23290 10248 23296 10260
rect 23063 10220 23296 10248
rect 23063 10217 23075 10220
rect 23017 10211 23075 10217
rect 23290 10208 23296 10220
rect 23348 10208 23354 10260
rect 23658 10180 23664 10192
rect 23619 10152 23664 10180
rect 23658 10140 23664 10152
rect 23716 10140 23722 10192
rect 23750 10140 23756 10192
rect 23808 10180 23814 10192
rect 24210 10180 24216 10192
rect 23808 10152 24216 10180
rect 23808 10140 23814 10152
rect 24210 10140 24216 10152
rect 24268 10180 24274 10192
rect 24397 10183 24455 10189
rect 24397 10180 24409 10183
rect 24268 10152 24409 10180
rect 24268 10140 24274 10152
rect 24397 10149 24409 10152
rect 24443 10149 24455 10183
rect 24397 10143 24455 10149
rect 24581 10183 24639 10189
rect 24581 10149 24593 10183
rect 24627 10180 24639 10183
rect 24670 10180 24676 10192
rect 24627 10152 24676 10180
rect 24627 10149 24639 10152
rect 24581 10143 24639 10149
rect 24670 10140 24676 10152
rect 24728 10140 24734 10192
rect 21913 10115 21971 10121
rect 21913 10112 21925 10115
rect 20824 10084 21925 10112
rect 19061 10075 19119 10081
rect 21913 10081 21925 10084
rect 21959 10081 21971 10115
rect 22830 10112 22836 10124
rect 22791 10084 22836 10112
rect 21913 10075 21971 10081
rect 22830 10072 22836 10084
rect 22888 10072 22894 10124
rect 13541 10047 13599 10053
rect 13541 10013 13553 10047
rect 13587 10013 13599 10047
rect 13541 10007 13599 10013
rect 13633 10047 13691 10053
rect 13633 10013 13645 10047
rect 13679 10044 13691 10047
rect 14734 10044 14740 10056
rect 13679 10016 14740 10044
rect 13679 10013 13691 10016
rect 13633 10007 13691 10013
rect 13556 9976 13584 10007
rect 14734 10004 14740 10016
rect 14792 10004 14798 10056
rect 15933 10047 15991 10053
rect 15933 10013 15945 10047
rect 15979 10013 15991 10047
rect 15933 10007 15991 10013
rect 13722 9976 13728 9988
rect 13556 9948 13728 9976
rect 13722 9936 13728 9948
rect 13780 9936 13786 9988
rect 13078 9908 13084 9920
rect 13039 9880 13084 9908
rect 13078 9868 13084 9880
rect 13136 9868 13142 9920
rect 15948 9908 15976 10007
rect 20990 10004 20996 10056
rect 21048 10044 21054 10056
rect 21453 10047 21511 10053
rect 21453 10044 21465 10047
rect 21048 10016 21465 10044
rect 21048 10004 21054 10016
rect 21453 10013 21465 10016
rect 21499 10044 21511 10047
rect 21726 10044 21732 10056
rect 21499 10016 21732 10044
rect 21499 10013 21511 10016
rect 21453 10007 21511 10013
rect 21726 10004 21732 10016
rect 21784 10004 21790 10056
rect 22373 10047 22431 10053
rect 22373 10013 22385 10047
rect 22419 10044 22431 10047
rect 23106 10044 23112 10056
rect 22419 10016 23112 10044
rect 22419 10013 22431 10016
rect 22373 10007 22431 10013
rect 23106 10004 23112 10016
rect 23164 10004 23170 10056
rect 23934 10004 23940 10056
rect 23992 10044 23998 10056
rect 24673 10047 24731 10053
rect 24673 10044 24685 10047
rect 23992 10016 24685 10044
rect 23992 10004 23998 10016
rect 24673 10013 24685 10016
rect 24719 10044 24731 10047
rect 24946 10044 24952 10056
rect 24719 10016 24952 10044
rect 24719 10013 24731 10016
rect 24673 10007 24731 10013
rect 24946 10004 24952 10016
rect 25004 10004 25010 10056
rect 17586 9936 17592 9988
rect 17644 9976 17650 9988
rect 18509 9979 18567 9985
rect 18509 9976 18521 9979
rect 17644 9948 18521 9976
rect 17644 9936 17650 9948
rect 18509 9945 18521 9948
rect 18555 9945 18567 9979
rect 18509 9939 18567 9945
rect 16114 9908 16120 9920
rect 15948 9880 16120 9908
rect 16114 9868 16120 9880
rect 16172 9908 16178 9920
rect 18046 9908 18052 9920
rect 16172 9880 18052 9908
rect 16172 9868 16178 9880
rect 18046 9868 18052 9880
rect 18104 9868 18110 9920
rect 19150 9868 19156 9920
rect 19208 9908 19214 9920
rect 19429 9911 19487 9917
rect 19429 9908 19441 9911
rect 19208 9880 19441 9908
rect 19208 9868 19214 9880
rect 19429 9877 19441 9880
rect 19475 9877 19487 9911
rect 19429 9871 19487 9877
rect 20806 9868 20812 9920
rect 20864 9908 20870 9920
rect 20993 9911 21051 9917
rect 20993 9908 21005 9911
rect 20864 9880 21005 9908
rect 20864 9868 20870 9880
rect 20993 9877 21005 9880
rect 21039 9877 21051 9911
rect 22554 9908 22560 9920
rect 22515 9880 22560 9908
rect 20993 9871 21051 9877
rect 22554 9868 22560 9880
rect 22612 9868 22618 9920
rect 24118 9908 24124 9920
rect 24079 9880 24124 9908
rect 24118 9868 24124 9880
rect 24176 9868 24182 9920
rect 25222 9908 25228 9920
rect 25183 9880 25228 9908
rect 25222 9868 25228 9880
rect 25280 9868 25286 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 15841 9707 15899 9713
rect 15841 9673 15853 9707
rect 15887 9704 15899 9707
rect 16853 9707 16911 9713
rect 16853 9704 16865 9707
rect 15887 9676 16865 9704
rect 15887 9673 15899 9676
rect 15841 9667 15899 9673
rect 16853 9673 16865 9676
rect 16899 9704 16911 9707
rect 16942 9704 16948 9716
rect 16899 9676 16948 9704
rect 16899 9673 16911 9676
rect 16853 9667 16911 9673
rect 16942 9664 16948 9676
rect 17000 9664 17006 9716
rect 17310 9664 17316 9716
rect 17368 9704 17374 9716
rect 17405 9707 17463 9713
rect 17405 9704 17417 9707
rect 17368 9676 17417 9704
rect 17368 9664 17374 9676
rect 17405 9673 17417 9676
rect 17451 9673 17463 9707
rect 17405 9667 17463 9673
rect 12434 9596 12440 9648
rect 12492 9636 12498 9648
rect 12713 9639 12771 9645
rect 12713 9636 12725 9639
rect 12492 9608 12725 9636
rect 12492 9596 12498 9608
rect 12713 9605 12725 9608
rect 12759 9605 12771 9639
rect 12713 9599 12771 9605
rect 12989 9639 13047 9645
rect 12989 9605 13001 9639
rect 13035 9636 13047 9639
rect 13722 9636 13728 9648
rect 13035 9608 13728 9636
rect 13035 9605 13047 9608
rect 12989 9599 13047 9605
rect 12728 9568 12756 9599
rect 13722 9596 13728 9608
rect 13780 9596 13786 9648
rect 13814 9596 13820 9648
rect 13872 9636 13878 9648
rect 13909 9639 13967 9645
rect 13909 9636 13921 9639
rect 13872 9608 13921 9636
rect 13872 9596 13878 9608
rect 13909 9605 13921 9608
rect 13955 9605 13967 9639
rect 13909 9599 13967 9605
rect 16022 9596 16028 9648
rect 16080 9636 16086 9648
rect 16393 9639 16451 9645
rect 16393 9636 16405 9639
rect 16080 9608 16405 9636
rect 16080 9596 16086 9608
rect 16393 9605 16405 9608
rect 16439 9605 16451 9639
rect 16393 9599 16451 9605
rect 13357 9571 13415 9577
rect 13357 9568 13369 9571
rect 12728 9540 13369 9568
rect 13357 9537 13369 9540
rect 13403 9537 13415 9571
rect 13357 9531 13415 9537
rect 13541 9571 13599 9577
rect 13541 9537 13553 9571
rect 13587 9568 13599 9571
rect 13630 9568 13636 9580
rect 13587 9540 13636 9568
rect 13587 9537 13599 9540
rect 13541 9531 13599 9537
rect 12253 9503 12311 9509
rect 12253 9469 12265 9503
rect 12299 9500 12311 9503
rect 13556 9500 13584 9531
rect 13630 9528 13636 9540
rect 13688 9528 13694 9580
rect 16758 9528 16764 9580
rect 16816 9568 16822 9580
rect 16945 9571 17003 9577
rect 16945 9568 16957 9571
rect 16816 9540 16957 9568
rect 16816 9528 16822 9540
rect 16945 9537 16957 9540
rect 16991 9537 17003 9571
rect 17420 9568 17448 9667
rect 17954 9664 17960 9716
rect 18012 9704 18018 9716
rect 19150 9704 19156 9716
rect 18012 9676 19156 9704
rect 18012 9664 18018 9676
rect 19150 9664 19156 9676
rect 19208 9704 19214 9716
rect 19429 9707 19487 9713
rect 19429 9704 19441 9707
rect 19208 9676 19441 9704
rect 19208 9664 19214 9676
rect 19429 9673 19441 9676
rect 19475 9673 19487 9707
rect 20990 9704 20996 9716
rect 19429 9667 19487 9673
rect 20640 9676 20996 9704
rect 17770 9636 17776 9648
rect 17731 9608 17776 9636
rect 17770 9596 17776 9608
rect 17828 9596 17834 9648
rect 19334 9596 19340 9648
rect 19392 9636 19398 9648
rect 19981 9639 20039 9645
rect 19981 9636 19993 9639
rect 19392 9608 19993 9636
rect 19392 9596 19398 9608
rect 19981 9605 19993 9608
rect 20027 9605 20039 9639
rect 19981 9599 20039 9605
rect 20533 9639 20591 9645
rect 20533 9605 20545 9639
rect 20579 9636 20591 9639
rect 20640 9636 20668 9676
rect 20990 9664 20996 9676
rect 21048 9664 21054 9716
rect 21542 9704 21548 9716
rect 21503 9676 21548 9704
rect 21542 9664 21548 9676
rect 21600 9664 21606 9716
rect 22830 9704 22836 9716
rect 21928 9676 22836 9704
rect 20579 9608 20668 9636
rect 20579 9605 20591 9608
rect 20533 9599 20591 9605
rect 20714 9596 20720 9648
rect 20772 9636 20778 9648
rect 21821 9639 21879 9645
rect 21821 9636 21833 9639
rect 20772 9608 21833 9636
rect 20772 9596 20778 9608
rect 21821 9605 21833 9608
rect 21867 9636 21879 9639
rect 21928 9636 21956 9676
rect 22830 9664 22836 9676
rect 22888 9664 22894 9716
rect 23109 9707 23167 9713
rect 23109 9673 23121 9707
rect 23155 9704 23167 9707
rect 23290 9704 23296 9716
rect 23155 9676 23296 9704
rect 23155 9673 23167 9676
rect 23109 9667 23167 9673
rect 23290 9664 23296 9676
rect 23348 9664 23354 9716
rect 24210 9664 24216 9716
rect 24268 9704 24274 9716
rect 24268 9676 24808 9704
rect 24268 9664 24274 9676
rect 21867 9608 21956 9636
rect 21867 9605 21879 9608
rect 21821 9599 21879 9605
rect 22094 9596 22100 9648
rect 22152 9636 22158 9648
rect 23753 9639 23811 9645
rect 22152 9608 22197 9636
rect 22152 9596 22158 9608
rect 23753 9605 23765 9639
rect 23799 9605 23811 9639
rect 24780 9636 24808 9676
rect 25777 9639 25835 9645
rect 25777 9636 25789 9639
rect 24780 9608 25789 9636
rect 23753 9599 23811 9605
rect 25777 9605 25789 9608
rect 25823 9605 25835 9639
rect 25777 9599 25835 9605
rect 17420 9540 18184 9568
rect 16945 9531 17003 9537
rect 14734 9509 14740 9512
rect 12299 9472 13584 9500
rect 14369 9503 14427 9509
rect 12299 9469 12311 9472
rect 12253 9463 12311 9469
rect 14369 9469 14381 9503
rect 14415 9500 14427 9503
rect 14461 9503 14519 9509
rect 14461 9500 14473 9503
rect 14415 9472 14473 9500
rect 14415 9469 14427 9472
rect 14369 9463 14427 9469
rect 14461 9469 14473 9472
rect 14507 9469 14519 9503
rect 14728 9500 14740 9509
rect 14695 9472 14740 9500
rect 14461 9463 14519 9469
rect 14728 9463 14740 9472
rect 13354 9392 13360 9444
rect 13412 9432 13418 9444
rect 13449 9435 13507 9441
rect 13449 9432 13461 9435
rect 13412 9404 13461 9432
rect 13412 9392 13418 9404
rect 13449 9401 13461 9404
rect 13495 9401 13507 9435
rect 14476 9432 14504 9463
rect 14734 9460 14740 9463
rect 14792 9460 14798 9512
rect 18046 9500 18052 9512
rect 18007 9472 18052 9500
rect 18046 9460 18052 9472
rect 18104 9460 18110 9512
rect 18156 9500 18184 9540
rect 20438 9528 20444 9580
rect 20496 9568 20502 9580
rect 20809 9571 20867 9577
rect 20809 9568 20821 9571
rect 20496 9540 20821 9568
rect 20496 9528 20502 9540
rect 20809 9537 20821 9540
rect 20855 9537 20867 9571
rect 22554 9568 22560 9580
rect 22515 9540 22560 9568
rect 20809 9531 20867 9537
rect 22554 9528 22560 9540
rect 22612 9528 22618 9580
rect 18305 9503 18363 9509
rect 18305 9500 18317 9503
rect 18156 9472 18317 9500
rect 18305 9469 18317 9472
rect 18351 9469 18363 9503
rect 23768 9500 23796 9599
rect 23934 9528 23940 9580
rect 23992 9568 23998 9580
rect 24673 9571 24731 9577
rect 24673 9568 24685 9571
rect 23992 9540 24685 9568
rect 23992 9528 23998 9540
rect 24673 9537 24685 9540
rect 24719 9537 24731 9571
rect 24673 9531 24731 9537
rect 24026 9500 24032 9512
rect 18305 9463 18363 9469
rect 22572 9472 23796 9500
rect 23987 9472 24032 9500
rect 16022 9432 16028 9444
rect 14476 9404 16028 9432
rect 13449 9395 13507 9401
rect 16022 9392 16028 9404
rect 16080 9392 16086 9444
rect 22572 9441 22600 9472
rect 24026 9460 24032 9472
rect 24084 9460 24090 9512
rect 25222 9500 25228 9512
rect 25183 9472 25228 9500
rect 25222 9460 25228 9472
rect 25280 9460 25286 9512
rect 22557 9435 22615 9441
rect 22557 9401 22569 9435
rect 22603 9401 22615 9435
rect 22557 9395 22615 9401
rect 20990 9364 20996 9376
rect 20951 9336 20996 9364
rect 20990 9324 20996 9336
rect 21048 9324 21054 9376
rect 21910 9324 21916 9376
rect 21968 9364 21974 9376
rect 22572 9364 22600 9395
rect 22646 9392 22652 9444
rect 22704 9432 22710 9444
rect 22704 9404 22749 9432
rect 22704 9392 22710 9404
rect 23106 9392 23112 9444
rect 23164 9432 23170 9444
rect 24305 9435 24363 9441
rect 24305 9432 24317 9435
rect 23164 9404 24317 9432
rect 23164 9392 23170 9404
rect 24305 9401 24317 9404
rect 24351 9432 24363 9435
rect 25041 9435 25099 9441
rect 25041 9432 25053 9435
rect 24351 9404 25053 9432
rect 24351 9401 24363 9404
rect 24305 9395 24363 9401
rect 25041 9401 25053 9404
rect 25087 9401 25099 9435
rect 25041 9395 25099 9401
rect 23474 9364 23480 9376
rect 21968 9336 22600 9364
rect 23435 9336 23480 9364
rect 21968 9324 21974 9336
rect 23474 9324 23480 9336
rect 23532 9364 23538 9376
rect 24213 9367 24271 9373
rect 24213 9364 24225 9367
rect 23532 9336 24225 9364
rect 23532 9324 23538 9336
rect 24213 9333 24225 9336
rect 24259 9333 24271 9367
rect 25406 9364 25412 9376
rect 25367 9336 25412 9364
rect 24213 9327 24271 9333
rect 25406 9324 25412 9336
rect 25464 9324 25470 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 13354 9160 13360 9172
rect 13315 9132 13360 9160
rect 13354 9120 13360 9132
rect 13412 9120 13418 9172
rect 13722 9160 13728 9172
rect 13683 9132 13728 9160
rect 13722 9120 13728 9132
rect 13780 9120 13786 9172
rect 14553 9163 14611 9169
rect 14553 9129 14565 9163
rect 14599 9160 14611 9163
rect 14734 9160 14740 9172
rect 14599 9132 14740 9160
rect 14599 9129 14611 9132
rect 14553 9123 14611 9129
rect 13081 9095 13139 9101
rect 13081 9061 13093 9095
rect 13127 9092 13139 9095
rect 14568 9092 14596 9123
rect 14734 9120 14740 9132
rect 14792 9120 14798 9172
rect 16850 9160 16856 9172
rect 16811 9132 16856 9160
rect 16850 9120 16856 9132
rect 16908 9120 16914 9172
rect 18046 9160 18052 9172
rect 18007 9132 18052 9160
rect 18046 9120 18052 9132
rect 18104 9120 18110 9172
rect 20346 9160 20352 9172
rect 20307 9132 20352 9160
rect 20346 9120 20352 9132
rect 20404 9120 20410 9172
rect 20717 9163 20775 9169
rect 20717 9129 20729 9163
rect 20763 9160 20775 9163
rect 21910 9160 21916 9172
rect 20763 9132 21916 9160
rect 20763 9129 20775 9132
rect 20717 9123 20775 9129
rect 21910 9120 21916 9132
rect 21968 9120 21974 9172
rect 22097 9163 22155 9169
rect 22097 9129 22109 9163
rect 22143 9160 22155 9163
rect 22646 9160 22652 9172
rect 22143 9132 22652 9160
rect 22143 9129 22155 9132
rect 22097 9123 22155 9129
rect 22646 9120 22652 9132
rect 22704 9160 22710 9172
rect 23750 9160 23756 9172
rect 22704 9132 23756 9160
rect 22704 9120 22710 9132
rect 23750 9120 23756 9132
rect 23808 9120 23814 9172
rect 24026 9120 24032 9172
rect 24084 9160 24090 9172
rect 24305 9163 24363 9169
rect 24305 9160 24317 9163
rect 24084 9132 24317 9160
rect 24084 9120 24090 9132
rect 24305 9129 24317 9132
rect 24351 9129 24363 9163
rect 24670 9160 24676 9172
rect 24631 9132 24676 9160
rect 24305 9123 24363 9129
rect 24670 9120 24676 9132
rect 24728 9120 24734 9172
rect 25409 9163 25467 9169
rect 25409 9129 25421 9163
rect 25455 9160 25467 9163
rect 25774 9160 25780 9172
rect 25455 9132 25780 9160
rect 25455 9129 25467 9132
rect 25409 9123 25467 9129
rect 25774 9120 25780 9132
rect 25832 9120 25838 9172
rect 13127 9064 14596 9092
rect 13127 9061 13139 9064
rect 13081 9055 13139 9061
rect 16574 9052 16580 9104
rect 16632 9092 16638 9104
rect 16669 9095 16727 9101
rect 16669 9092 16681 9095
rect 16632 9064 16681 9092
rect 16632 9052 16638 9064
rect 16669 9061 16681 9064
rect 16715 9061 16727 9095
rect 16942 9092 16948 9104
rect 16855 9064 16948 9092
rect 16669 9055 16727 9061
rect 16942 9052 16948 9064
rect 17000 9092 17006 9104
rect 17954 9092 17960 9104
rect 17000 9064 17960 9092
rect 17000 9052 17006 9064
rect 17954 9052 17960 9064
rect 18012 9052 18018 9104
rect 18322 9052 18328 9104
rect 18380 9092 18386 9104
rect 18570 9095 18628 9101
rect 18570 9092 18582 9095
rect 18380 9064 18582 9092
rect 18380 9052 18386 9064
rect 18570 9061 18582 9064
rect 18616 9061 18628 9095
rect 25222 9092 25228 9104
rect 25183 9064 25228 9092
rect 18570 9055 18628 9061
rect 25222 9052 25228 9064
rect 25280 9052 25286 9104
rect 21266 9024 21272 9036
rect 21227 8996 21272 9024
rect 21266 8984 21272 8996
rect 21324 8984 21330 9036
rect 21726 8984 21732 9036
rect 21784 9024 21790 9036
rect 22186 9024 22192 9036
rect 21784 8996 22192 9024
rect 21784 8984 21790 8996
rect 22186 8984 22192 8996
rect 22244 9024 22250 9036
rect 22373 9027 22431 9033
rect 22373 9024 22385 9027
rect 22244 8996 22385 9024
rect 22244 8984 22250 8996
rect 22373 8993 22385 8996
rect 22419 8993 22431 9027
rect 22373 8987 22431 8993
rect 22462 8984 22468 9036
rect 22520 9024 22526 9036
rect 22640 9027 22698 9033
rect 22640 9024 22652 9027
rect 22520 8996 22652 9024
rect 22520 8984 22526 8996
rect 22640 8993 22652 8996
rect 22686 9024 22698 9027
rect 23106 9024 23112 9036
rect 22686 8996 23112 9024
rect 22686 8993 22698 8996
rect 22640 8987 22698 8993
rect 23106 8984 23112 8996
rect 23164 8984 23170 9036
rect 18046 8916 18052 8968
rect 18104 8956 18110 8968
rect 18325 8959 18383 8965
rect 18325 8956 18337 8959
rect 18104 8928 18337 8956
rect 18104 8916 18110 8928
rect 18325 8925 18337 8928
rect 18371 8925 18383 8959
rect 25498 8956 25504 8968
rect 25459 8928 25504 8956
rect 18325 8919 18383 8925
rect 25498 8916 25504 8928
rect 25556 8916 25562 8968
rect 16390 8820 16396 8832
rect 16351 8792 16396 8820
rect 16390 8780 16396 8792
rect 16448 8780 16454 8832
rect 19705 8823 19763 8829
rect 19705 8789 19717 8823
rect 19751 8820 19763 8823
rect 19978 8820 19984 8832
rect 19751 8792 19984 8820
rect 19751 8789 19763 8792
rect 19705 8783 19763 8789
rect 19978 8780 19984 8792
rect 20036 8780 20042 8832
rect 20346 8780 20352 8832
rect 20404 8820 20410 8832
rect 20530 8820 20536 8832
rect 20404 8792 20536 8820
rect 20404 8780 20410 8792
rect 20530 8780 20536 8792
rect 20588 8780 20594 8832
rect 21174 8820 21180 8832
rect 21135 8792 21180 8820
rect 21174 8780 21180 8792
rect 21232 8780 21238 8832
rect 21450 8820 21456 8832
rect 21411 8792 21456 8820
rect 21450 8780 21456 8792
rect 21508 8780 21514 8832
rect 24854 8780 24860 8832
rect 24912 8820 24918 8832
rect 24949 8823 25007 8829
rect 24949 8820 24961 8823
rect 24912 8792 24961 8820
rect 24912 8780 24918 8792
rect 24949 8789 24961 8792
rect 24995 8789 25007 8823
rect 24949 8783 25007 8789
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 15562 8576 15568 8628
rect 15620 8616 15626 8628
rect 16485 8619 16543 8625
rect 16485 8616 16497 8619
rect 15620 8588 16497 8616
rect 15620 8576 15626 8588
rect 16485 8585 16497 8588
rect 16531 8585 16543 8619
rect 16485 8579 16543 8585
rect 16574 8576 16580 8628
rect 16632 8616 16638 8628
rect 17405 8619 17463 8625
rect 17405 8616 17417 8619
rect 16632 8588 17417 8616
rect 16632 8576 16638 8588
rect 17405 8585 17417 8588
rect 17451 8585 17463 8619
rect 17405 8579 17463 8585
rect 17865 8619 17923 8625
rect 17865 8585 17877 8619
rect 17911 8616 17923 8619
rect 18322 8616 18328 8628
rect 17911 8588 18328 8616
rect 17911 8585 17923 8588
rect 17865 8579 17923 8585
rect 18322 8576 18328 8588
rect 18380 8576 18386 8628
rect 19061 8619 19119 8625
rect 19061 8585 19073 8619
rect 19107 8616 19119 8619
rect 19518 8616 19524 8628
rect 19107 8588 19524 8616
rect 19107 8585 19119 8588
rect 19061 8579 19119 8585
rect 19518 8576 19524 8588
rect 19576 8576 19582 8628
rect 22462 8616 22468 8628
rect 22423 8588 22468 8616
rect 22462 8576 22468 8588
rect 22520 8576 22526 8628
rect 25222 8576 25228 8628
rect 25280 8616 25286 8628
rect 25961 8619 26019 8625
rect 25961 8616 25973 8619
rect 25280 8588 25973 8616
rect 25280 8576 25286 8588
rect 25961 8585 25973 8588
rect 26007 8585 26019 8619
rect 25961 8579 26019 8585
rect 15933 8551 15991 8557
rect 15933 8517 15945 8551
rect 15979 8548 15991 8551
rect 16942 8548 16948 8560
rect 15979 8520 16948 8548
rect 15979 8517 15991 8520
rect 15933 8511 15991 8517
rect 16942 8508 16948 8520
rect 17000 8508 17006 8560
rect 19334 8548 19340 8560
rect 19295 8520 19340 8548
rect 19334 8508 19340 8520
rect 19392 8508 19398 8560
rect 15565 8483 15623 8489
rect 15565 8449 15577 8483
rect 15611 8480 15623 8483
rect 16850 8480 16856 8492
rect 15611 8452 16856 8480
rect 15611 8449 15623 8452
rect 15565 8443 15623 8449
rect 16850 8440 16856 8452
rect 16908 8440 16914 8492
rect 17034 8480 17040 8492
rect 16995 8452 17040 8480
rect 17034 8440 17040 8452
rect 17092 8440 17098 8492
rect 18046 8440 18052 8492
rect 18104 8480 18110 8492
rect 18325 8483 18383 8489
rect 18325 8480 18337 8483
rect 18104 8452 18337 8480
rect 18104 8440 18110 8452
rect 18325 8449 18337 8452
rect 18371 8449 18383 8483
rect 19352 8480 19380 8508
rect 19536 8480 19564 8576
rect 19613 8551 19671 8557
rect 19613 8517 19625 8551
rect 19659 8548 19671 8551
rect 20530 8548 20536 8560
rect 19659 8520 20536 8548
rect 19659 8517 19671 8520
rect 19613 8511 19671 8517
rect 20530 8508 20536 8520
rect 20588 8508 20594 8560
rect 22186 8508 22192 8560
rect 22244 8548 22250 8560
rect 23017 8551 23075 8557
rect 23017 8548 23029 8551
rect 22244 8520 23029 8548
rect 22244 8508 22250 8520
rect 23017 8517 23029 8520
rect 23063 8548 23075 8551
rect 23385 8551 23443 8557
rect 23385 8548 23397 8551
rect 23063 8520 23397 8548
rect 23063 8517 23075 8520
rect 23017 8511 23075 8517
rect 23385 8517 23397 8520
rect 23431 8548 23443 8551
rect 25685 8551 25743 8557
rect 23431 8520 23704 8548
rect 23431 8517 23443 8520
rect 23385 8511 23443 8517
rect 23676 8492 23704 8520
rect 25685 8517 25697 8551
rect 25731 8548 25743 8551
rect 25774 8548 25780 8560
rect 25731 8520 25780 8548
rect 25731 8517 25743 8520
rect 25685 8511 25743 8517
rect 25774 8508 25780 8520
rect 25832 8508 25838 8560
rect 19981 8483 20039 8489
rect 19981 8480 19993 8483
rect 19352 8452 19472 8480
rect 19536 8452 19993 8480
rect 18325 8443 18383 8449
rect 16574 8372 16580 8424
rect 16632 8412 16638 8424
rect 17218 8412 17224 8424
rect 16632 8384 17224 8412
rect 16632 8372 16638 8384
rect 16298 8344 16304 8356
rect 16211 8316 16304 8344
rect 16298 8304 16304 8316
rect 16356 8344 16362 8356
rect 16758 8344 16764 8356
rect 16356 8316 16764 8344
rect 16356 8304 16362 8316
rect 16758 8304 16764 8316
rect 16816 8304 16822 8356
rect 16960 8353 16988 8384
rect 17218 8372 17224 8384
rect 17276 8372 17282 8424
rect 18509 8415 18567 8421
rect 18509 8381 18521 8415
rect 18555 8412 18567 8415
rect 19334 8412 19340 8424
rect 18555 8384 19340 8412
rect 18555 8381 18567 8384
rect 18509 8375 18567 8381
rect 19334 8372 19340 8384
rect 19392 8372 19398 8424
rect 16945 8347 17003 8353
rect 16945 8313 16957 8347
rect 16991 8313 17003 8347
rect 19444 8344 19472 8452
rect 19981 8449 19993 8452
rect 20027 8449 20039 8483
rect 23658 8480 23664 8492
rect 23571 8452 23664 8480
rect 19981 8443 20039 8449
rect 23658 8440 23664 8452
rect 23716 8440 23722 8492
rect 20990 8412 20996 8424
rect 20088 8384 20996 8412
rect 20088 8353 20116 8384
rect 20990 8372 20996 8384
rect 21048 8372 21054 8424
rect 21085 8415 21143 8421
rect 21085 8381 21097 8415
rect 21131 8412 21143 8415
rect 21726 8412 21732 8424
rect 21131 8384 21732 8412
rect 21131 8381 21143 8384
rect 21085 8375 21143 8381
rect 20073 8347 20131 8353
rect 20073 8344 20085 8347
rect 19444 8316 20085 8344
rect 16945 8307 17003 8313
rect 20073 8313 20085 8316
rect 20119 8313 20131 8347
rect 20073 8307 20131 8313
rect 20165 8347 20223 8353
rect 20165 8313 20177 8347
rect 20211 8313 20223 8347
rect 21100 8344 21128 8375
rect 21726 8372 21732 8384
rect 21784 8372 21790 8424
rect 23750 8372 23756 8424
rect 23808 8412 23814 8424
rect 23917 8415 23975 8421
rect 23917 8412 23929 8415
rect 23808 8384 23929 8412
rect 23808 8372 23814 8384
rect 23917 8381 23929 8384
rect 23963 8381 23975 8415
rect 23917 8375 23975 8381
rect 20165 8307 20223 8313
rect 20916 8316 21128 8344
rect 20180 8276 20208 8307
rect 20916 8288 20944 8316
rect 21174 8304 21180 8356
rect 21232 8344 21238 8356
rect 21330 8347 21388 8353
rect 21330 8344 21342 8347
rect 21232 8316 21342 8344
rect 21232 8304 21238 8316
rect 21330 8313 21342 8316
rect 21376 8313 21388 8347
rect 25498 8344 25504 8356
rect 21330 8307 21388 8313
rect 25148 8316 25504 8344
rect 25148 8288 25176 8316
rect 25498 8304 25504 8316
rect 25556 8344 25562 8356
rect 26329 8347 26387 8353
rect 26329 8344 26341 8347
rect 25556 8316 26341 8344
rect 25556 8304 25562 8316
rect 26329 8313 26341 8316
rect 26375 8313 26387 8347
rect 26329 8307 26387 8313
rect 20622 8276 20628 8288
rect 20180 8248 20628 8276
rect 20622 8236 20628 8248
rect 20680 8236 20686 8288
rect 20898 8276 20904 8288
rect 20859 8248 20904 8276
rect 20898 8236 20904 8248
rect 20956 8236 20962 8288
rect 25041 8279 25099 8285
rect 25041 8245 25053 8279
rect 25087 8276 25099 8279
rect 25130 8276 25136 8288
rect 25087 8248 25136 8276
rect 25087 8245 25099 8248
rect 25041 8239 25099 8245
rect 25130 8236 25136 8248
rect 25188 8236 25194 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 16482 8072 16488 8084
rect 16443 8044 16488 8072
rect 16482 8032 16488 8044
rect 16540 8032 16546 8084
rect 16853 8075 16911 8081
rect 16853 8041 16865 8075
rect 16899 8072 16911 8075
rect 17034 8072 17040 8084
rect 16899 8044 17040 8072
rect 16899 8041 16911 8044
rect 16853 8035 16911 8041
rect 17034 8032 17040 8044
rect 17092 8032 17098 8084
rect 22462 8032 22468 8084
rect 22520 8072 22526 8084
rect 22833 8075 22891 8081
rect 22833 8072 22845 8075
rect 22520 8044 22845 8072
rect 22520 8032 22526 8044
rect 22833 8041 22845 8044
rect 22879 8041 22891 8075
rect 23750 8072 23756 8084
rect 23711 8044 23756 8072
rect 22833 8035 22891 8041
rect 23750 8032 23756 8044
rect 23808 8032 23814 8084
rect 11054 7964 11060 8016
rect 11112 8004 11118 8016
rect 18506 8004 18512 8016
rect 11112 7976 18512 8004
rect 11112 7964 11118 7976
rect 18506 7964 18512 7976
rect 18564 7964 18570 8016
rect 19334 7964 19340 8016
rect 19392 8004 19398 8016
rect 19613 8007 19671 8013
rect 19613 8004 19625 8007
rect 19392 7976 19625 8004
rect 19392 7964 19398 7976
rect 19613 7973 19625 7976
rect 19659 7973 19671 8007
rect 19794 8004 19800 8016
rect 19755 7976 19800 8004
rect 19613 7967 19671 7973
rect 19794 7964 19800 7976
rect 19852 8004 19858 8016
rect 20714 8004 20720 8016
rect 19852 7976 20720 8004
rect 19852 7964 19858 7976
rect 20714 7964 20720 7976
rect 20772 7964 20778 8016
rect 23385 8007 23443 8013
rect 23385 7973 23397 8007
rect 23431 8004 23443 8007
rect 24762 8004 24768 8016
rect 23431 7976 24768 8004
rect 23431 7973 23443 7976
rect 23385 7967 23443 7973
rect 24762 7964 24768 7976
rect 24820 7964 24826 8016
rect 17957 7939 18015 7945
rect 17957 7905 17969 7939
rect 18003 7936 18015 7939
rect 18598 7936 18604 7948
rect 18003 7908 18604 7936
rect 18003 7905 18015 7908
rect 17957 7899 18015 7905
rect 18598 7896 18604 7908
rect 18656 7936 18662 7948
rect 18693 7939 18751 7945
rect 18693 7936 18705 7939
rect 18656 7908 18705 7936
rect 18656 7896 18662 7908
rect 18693 7905 18705 7908
rect 18739 7905 18751 7939
rect 18693 7899 18751 7905
rect 19889 7939 19947 7945
rect 19889 7905 19901 7939
rect 19935 7936 19947 7939
rect 19978 7936 19984 7948
rect 19935 7908 19984 7936
rect 19935 7905 19947 7908
rect 19889 7899 19947 7905
rect 19978 7896 19984 7908
rect 20036 7936 20042 7948
rect 20622 7936 20628 7948
rect 20036 7908 20628 7936
rect 20036 7896 20042 7908
rect 20622 7896 20628 7908
rect 20680 7936 20686 7948
rect 21168 7939 21226 7945
rect 21168 7936 21180 7939
rect 20680 7908 21180 7936
rect 20680 7896 20686 7908
rect 21168 7905 21180 7908
rect 21214 7936 21226 7939
rect 21910 7936 21916 7948
rect 21214 7908 21916 7936
rect 21214 7905 21226 7908
rect 21168 7899 21226 7905
rect 21910 7896 21916 7908
rect 21968 7896 21974 7948
rect 23658 7896 23664 7948
rect 23716 7936 23722 7948
rect 23937 7939 23995 7945
rect 23937 7936 23949 7939
rect 23716 7908 23949 7936
rect 23716 7896 23722 7908
rect 23937 7905 23949 7908
rect 23983 7905 23995 7939
rect 23937 7899 23995 7905
rect 24204 7939 24262 7945
rect 24204 7905 24216 7939
rect 24250 7936 24262 7939
rect 25130 7936 25136 7948
rect 24250 7908 25136 7936
rect 24250 7905 24262 7908
rect 24204 7899 24262 7905
rect 25130 7896 25136 7908
rect 25188 7896 25194 7948
rect 16945 7871 17003 7877
rect 16945 7837 16957 7871
rect 16991 7868 17003 7871
rect 18046 7868 18052 7880
rect 16991 7840 18052 7868
rect 16991 7837 17003 7840
rect 16945 7831 17003 7837
rect 18046 7828 18052 7840
rect 18104 7828 18110 7880
rect 18230 7868 18236 7880
rect 18191 7840 18236 7868
rect 18230 7828 18236 7840
rect 18288 7828 18294 7880
rect 20714 7828 20720 7880
rect 20772 7868 20778 7880
rect 20898 7868 20904 7880
rect 20772 7840 20904 7868
rect 20772 7828 20778 7840
rect 20898 7828 20904 7840
rect 20956 7828 20962 7880
rect 14645 7735 14703 7741
rect 14645 7701 14657 7735
rect 14691 7732 14703 7735
rect 15562 7732 15568 7744
rect 14691 7704 15568 7732
rect 14691 7701 14703 7704
rect 14645 7695 14703 7701
rect 15562 7692 15568 7704
rect 15620 7692 15626 7744
rect 19337 7735 19395 7741
rect 19337 7701 19349 7735
rect 19383 7732 19395 7735
rect 20533 7735 20591 7741
rect 20533 7732 20545 7735
rect 19383 7704 20545 7732
rect 19383 7701 19395 7704
rect 19337 7695 19395 7701
rect 20533 7701 20545 7704
rect 20579 7732 20591 7735
rect 20898 7732 20904 7744
rect 20579 7704 20904 7732
rect 20579 7701 20591 7704
rect 20533 7695 20591 7701
rect 20898 7692 20904 7704
rect 20956 7692 20962 7744
rect 21174 7692 21180 7744
rect 21232 7732 21238 7744
rect 22281 7735 22339 7741
rect 22281 7732 22293 7735
rect 21232 7704 22293 7732
rect 21232 7692 21238 7704
rect 22281 7701 22293 7704
rect 22327 7701 22339 7735
rect 25314 7732 25320 7744
rect 25275 7704 25320 7732
rect 22281 7695 22339 7701
rect 25314 7692 25320 7704
rect 25372 7692 25378 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 14366 7528 14372 7540
rect 14327 7500 14372 7528
rect 14366 7488 14372 7500
rect 14424 7488 14430 7540
rect 15746 7488 15752 7540
rect 15804 7528 15810 7540
rect 15841 7531 15899 7537
rect 15841 7528 15853 7531
rect 15804 7500 15853 7528
rect 15804 7488 15810 7500
rect 15841 7497 15853 7500
rect 15887 7497 15899 7531
rect 19426 7528 19432 7540
rect 19387 7500 19432 7528
rect 15841 7491 15899 7497
rect 14550 7420 14556 7472
rect 14608 7460 14614 7472
rect 14645 7463 14703 7469
rect 14645 7460 14657 7463
rect 14608 7432 14657 7460
rect 14608 7420 14614 7432
rect 14645 7429 14657 7432
rect 14691 7429 14703 7463
rect 14645 7423 14703 7429
rect 14642 7284 14648 7336
rect 14700 7324 14706 7336
rect 14921 7327 14979 7333
rect 14921 7324 14933 7327
rect 14700 7296 14933 7324
rect 14700 7284 14706 7296
rect 14921 7293 14933 7296
rect 14967 7293 14979 7327
rect 15856 7324 15884 7491
rect 19426 7488 19432 7500
rect 19484 7488 19490 7540
rect 20714 7488 20720 7540
rect 20772 7528 20778 7540
rect 21545 7531 21603 7537
rect 21545 7528 21557 7531
rect 20772 7500 21557 7528
rect 20772 7488 20778 7500
rect 21545 7497 21557 7500
rect 21591 7497 21603 7531
rect 21910 7528 21916 7540
rect 21871 7500 21916 7528
rect 21545 7491 21603 7497
rect 21910 7488 21916 7500
rect 21968 7488 21974 7540
rect 23477 7531 23535 7537
rect 23477 7497 23489 7531
rect 23523 7528 23535 7531
rect 23658 7528 23664 7540
rect 23523 7500 23664 7528
rect 23523 7497 23535 7500
rect 23477 7491 23535 7497
rect 23658 7488 23664 7500
rect 23716 7488 23722 7540
rect 16482 7460 16488 7472
rect 16443 7432 16488 7460
rect 16482 7420 16488 7432
rect 16540 7420 16546 7472
rect 20162 7420 20168 7472
rect 20220 7460 20226 7472
rect 20346 7460 20352 7472
rect 20220 7432 20352 7460
rect 20220 7420 20226 7432
rect 20346 7420 20352 7432
rect 20404 7420 20410 7472
rect 20622 7460 20628 7472
rect 20583 7432 20628 7460
rect 20622 7420 20628 7432
rect 20680 7420 20686 7472
rect 23198 7420 23204 7472
rect 23256 7460 23262 7472
rect 24029 7463 24087 7469
rect 24029 7460 24041 7463
rect 23256 7432 24041 7460
rect 23256 7420 23262 7432
rect 24029 7429 24041 7432
rect 24075 7429 24087 7463
rect 24029 7423 24087 7429
rect 20254 7352 20260 7404
rect 20312 7352 20318 7404
rect 20441 7395 20499 7401
rect 20441 7361 20453 7395
rect 20487 7392 20499 7395
rect 21174 7392 21180 7404
rect 20487 7364 21180 7392
rect 20487 7361 20499 7364
rect 20441 7355 20499 7361
rect 21174 7352 21180 7364
rect 21232 7352 21238 7404
rect 22557 7395 22615 7401
rect 22557 7361 22569 7395
rect 22603 7392 22615 7395
rect 23382 7392 23388 7404
rect 22603 7364 23388 7392
rect 22603 7361 22615 7364
rect 22557 7355 22615 7361
rect 23382 7352 23388 7364
rect 23440 7352 23446 7404
rect 24489 7395 24547 7401
rect 24489 7361 24501 7395
rect 24535 7392 24547 7395
rect 24762 7392 24768 7404
rect 24535 7364 24768 7392
rect 24535 7361 24547 7364
rect 24489 7355 24547 7361
rect 24762 7352 24768 7364
rect 24820 7352 24826 7404
rect 25041 7395 25099 7401
rect 25041 7361 25053 7395
rect 25087 7392 25099 7395
rect 25130 7392 25136 7404
rect 25087 7364 25136 7392
rect 25087 7361 25099 7364
rect 25041 7355 25099 7361
rect 25130 7352 25136 7364
rect 25188 7352 25194 7404
rect 17862 7324 17868 7336
rect 15856 7296 16988 7324
rect 17823 7296 17868 7324
rect 14921 7287 14979 7293
rect 14366 7216 14372 7268
rect 14424 7256 14430 7268
rect 15105 7259 15163 7265
rect 15105 7256 15117 7259
rect 14424 7228 15117 7256
rect 14424 7216 14430 7228
rect 15105 7225 15117 7228
rect 15151 7225 15163 7259
rect 15105 7219 15163 7225
rect 15197 7259 15255 7265
rect 15197 7225 15209 7259
rect 15243 7256 15255 7259
rect 15562 7256 15568 7268
rect 15243 7228 15568 7256
rect 15243 7225 15255 7228
rect 15197 7219 15255 7225
rect 15562 7216 15568 7228
rect 15620 7216 15626 7268
rect 16960 7265 16988 7296
rect 17862 7284 17868 7296
rect 17920 7324 17926 7336
rect 18049 7327 18107 7333
rect 18049 7324 18061 7327
rect 17920 7296 18061 7324
rect 17920 7284 17926 7296
rect 18049 7293 18061 7296
rect 18095 7293 18107 7327
rect 18049 7287 18107 7293
rect 16761 7259 16819 7265
rect 16761 7225 16773 7259
rect 16807 7225 16819 7259
rect 16761 7219 16819 7225
rect 16945 7259 17003 7265
rect 16945 7225 16957 7259
rect 16991 7225 17003 7259
rect 16945 7219 17003 7225
rect 17037 7259 17095 7265
rect 17037 7225 17049 7259
rect 17083 7225 17095 7259
rect 17037 7219 17095 7225
rect 16206 7188 16212 7200
rect 16167 7160 16212 7188
rect 16206 7148 16212 7160
rect 16264 7188 16270 7200
rect 16776 7188 16804 7219
rect 16264 7160 16804 7188
rect 17052 7188 17080 7219
rect 18138 7216 18144 7268
rect 18196 7256 18202 7268
rect 18294 7259 18352 7265
rect 18294 7256 18306 7259
rect 18196 7228 18306 7256
rect 18196 7216 18202 7228
rect 18294 7225 18306 7228
rect 18340 7225 18352 7259
rect 18294 7219 18352 7225
rect 19794 7216 19800 7268
rect 19852 7256 19858 7268
rect 19852 7228 20116 7256
rect 19852 7216 19858 7228
rect 20088 7200 20116 7228
rect 20272 7200 20300 7352
rect 20898 7324 20904 7336
rect 20859 7296 20904 7324
rect 20898 7284 20904 7296
rect 20956 7284 20962 7336
rect 22281 7327 22339 7333
rect 22281 7293 22293 7327
rect 22327 7324 22339 7327
rect 23198 7324 23204 7336
rect 22327 7296 23204 7324
rect 22327 7293 22339 7296
rect 22281 7287 22339 7293
rect 23198 7284 23204 7296
rect 23256 7284 23262 7336
rect 24578 7324 24584 7336
rect 24491 7296 24584 7324
rect 24578 7284 24584 7296
rect 24636 7324 24642 7336
rect 25314 7324 25320 7336
rect 24636 7296 25320 7324
rect 24636 7284 24642 7296
rect 25314 7284 25320 7296
rect 25372 7284 25378 7336
rect 25498 7324 25504 7336
rect 25459 7296 25504 7324
rect 25498 7284 25504 7296
rect 25556 7324 25562 7336
rect 26053 7327 26111 7333
rect 26053 7324 26065 7327
rect 25556 7296 26065 7324
rect 25556 7284 25562 7296
rect 26053 7293 26065 7296
rect 26099 7293 26111 7327
rect 26053 7287 26111 7293
rect 20530 7216 20536 7268
rect 20588 7256 20594 7268
rect 21085 7259 21143 7265
rect 21085 7256 21097 7259
rect 20588 7228 21097 7256
rect 20588 7216 20594 7228
rect 21085 7225 21097 7228
rect 21131 7225 21143 7259
rect 21085 7219 21143 7225
rect 23109 7259 23167 7265
rect 23109 7225 23121 7259
rect 23155 7256 23167 7259
rect 24596 7256 24624 7284
rect 23155 7228 24624 7256
rect 24872 7228 25084 7256
rect 23155 7225 23167 7228
rect 23109 7219 23167 7225
rect 17494 7188 17500 7200
rect 17052 7160 17500 7188
rect 16264 7148 16270 7160
rect 17494 7148 17500 7160
rect 17552 7148 17558 7200
rect 20070 7188 20076 7200
rect 20031 7160 20076 7188
rect 20070 7148 20076 7160
rect 20128 7148 20134 7200
rect 20254 7148 20260 7200
rect 20312 7148 20318 7200
rect 24489 7191 24547 7197
rect 24489 7157 24501 7191
rect 24535 7188 24547 7191
rect 24872 7188 24900 7228
rect 25056 7200 25084 7228
rect 24535 7160 24900 7188
rect 24535 7157 24547 7160
rect 24489 7151 24547 7157
rect 25038 7148 25044 7200
rect 25096 7188 25102 7200
rect 25317 7191 25375 7197
rect 25317 7188 25329 7191
rect 25096 7160 25329 7188
rect 25096 7148 25102 7160
rect 25317 7157 25329 7160
rect 25363 7157 25375 7191
rect 25682 7188 25688 7200
rect 25643 7160 25688 7188
rect 25317 7151 25375 7157
rect 25682 7148 25688 7160
rect 25740 7148 25746 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 14642 6984 14648 6996
rect 14603 6956 14648 6984
rect 14642 6944 14648 6956
rect 14700 6944 14706 6996
rect 18138 6984 18144 6996
rect 18099 6956 18144 6984
rect 18138 6944 18144 6956
rect 18196 6944 18202 6996
rect 19334 6944 19340 6996
rect 19392 6984 19398 6996
rect 19521 6987 19579 6993
rect 19521 6984 19533 6987
rect 19392 6956 19533 6984
rect 19392 6944 19398 6956
rect 19521 6953 19533 6956
rect 19567 6953 19579 6987
rect 19978 6984 19984 6996
rect 19939 6956 19984 6984
rect 19521 6947 19579 6953
rect 19978 6944 19984 6956
rect 20036 6944 20042 6996
rect 23198 6984 23204 6996
rect 23159 6956 23204 6984
rect 23198 6944 23204 6956
rect 23256 6944 23262 6996
rect 24578 6944 24584 6996
rect 24636 6984 24642 6996
rect 24673 6987 24731 6993
rect 24673 6984 24685 6987
rect 24636 6956 24685 6984
rect 24636 6944 24642 6956
rect 24673 6953 24685 6956
rect 24719 6953 24731 6987
rect 24673 6947 24731 6953
rect 16482 6876 16488 6928
rect 16540 6916 16546 6928
rect 19015 6919 19073 6925
rect 19015 6916 19027 6919
rect 16540 6888 19027 6916
rect 16540 6876 16546 6888
rect 19015 6885 19027 6888
rect 19061 6916 19073 6919
rect 19242 6916 19248 6928
rect 19061 6888 19248 6916
rect 19061 6885 19073 6888
rect 19015 6879 19073 6885
rect 19242 6876 19248 6888
rect 19300 6876 19306 6928
rect 23845 6919 23903 6925
rect 23845 6885 23857 6919
rect 23891 6885 23903 6919
rect 25409 6919 25467 6925
rect 25409 6916 25421 6919
rect 23845 6879 23903 6885
rect 25148 6888 25421 6916
rect 8021 6851 8079 6857
rect 8021 6817 8033 6851
rect 8067 6848 8079 6851
rect 8110 6848 8116 6860
rect 8067 6820 8116 6848
rect 8067 6817 8079 6820
rect 8021 6811 8079 6817
rect 8110 6808 8116 6820
rect 8168 6808 8174 6860
rect 16298 6857 16304 6860
rect 16292 6848 16304 6857
rect 16259 6820 16304 6848
rect 16292 6811 16304 6820
rect 16298 6808 16304 6811
rect 16356 6808 16362 6860
rect 18046 6808 18052 6860
rect 18104 6848 18110 6860
rect 18506 6848 18512 6860
rect 18104 6820 18512 6848
rect 18104 6808 18110 6820
rect 18506 6808 18512 6820
rect 18564 6848 18570 6860
rect 18877 6851 18935 6857
rect 18877 6848 18889 6851
rect 18564 6820 18889 6848
rect 18564 6808 18570 6820
rect 18877 6817 18889 6820
rect 18923 6817 18935 6851
rect 20530 6848 20536 6860
rect 20491 6820 20536 6848
rect 18877 6811 18935 6817
rect 20530 6808 20536 6820
rect 20588 6808 20594 6860
rect 20898 6848 20904 6860
rect 20859 6820 20904 6848
rect 20898 6808 20904 6820
rect 20956 6808 20962 6860
rect 21266 6808 21272 6860
rect 21324 6848 21330 6860
rect 21453 6851 21511 6857
rect 21453 6848 21465 6851
rect 21324 6820 21465 6848
rect 21324 6808 21330 6820
rect 21453 6817 21465 6820
rect 21499 6817 21511 6851
rect 21453 6811 21511 6817
rect 22005 6851 22063 6857
rect 22005 6817 22017 6851
rect 22051 6848 22063 6851
rect 22094 6848 22100 6860
rect 22051 6820 22100 6848
rect 22051 6817 22063 6820
rect 22005 6811 22063 6817
rect 22094 6808 22100 6820
rect 22152 6848 22158 6860
rect 22741 6851 22799 6857
rect 22741 6848 22753 6851
rect 22152 6820 22753 6848
rect 22152 6808 22158 6820
rect 22741 6817 22753 6820
rect 22787 6817 22799 6851
rect 22741 6811 22799 6817
rect 23290 6808 23296 6860
rect 23348 6848 23354 6860
rect 23860 6848 23888 6879
rect 23348 6820 23888 6848
rect 23348 6808 23354 6820
rect 24762 6808 24768 6860
rect 24820 6848 24826 6860
rect 25148 6848 25176 6888
rect 25409 6885 25421 6888
rect 25455 6885 25467 6919
rect 25409 6879 25467 6885
rect 24820 6820 25176 6848
rect 25225 6851 25283 6857
rect 24820 6808 24826 6820
rect 25225 6817 25237 6851
rect 25271 6848 25283 6851
rect 25314 6848 25320 6860
rect 25271 6820 25320 6848
rect 25271 6817 25283 6820
rect 25225 6811 25283 6817
rect 25314 6808 25320 6820
rect 25372 6848 25378 6860
rect 25866 6848 25872 6860
rect 25372 6820 25872 6848
rect 25372 6808 25378 6820
rect 25866 6808 25872 6820
rect 25924 6808 25930 6860
rect 16022 6780 16028 6792
rect 15983 6752 16028 6780
rect 16022 6740 16028 6752
rect 16080 6740 16086 6792
rect 18230 6740 18236 6792
rect 18288 6780 18294 6792
rect 19150 6780 19156 6792
rect 18288 6752 19156 6780
rect 18288 6740 18294 6752
rect 19150 6740 19156 6752
rect 19208 6740 19214 6792
rect 20916 6780 20944 6808
rect 22189 6783 22247 6789
rect 22189 6780 22201 6783
rect 20916 6752 22201 6780
rect 22189 6749 22201 6752
rect 22235 6749 22247 6783
rect 22189 6743 22247 6749
rect 22278 6740 22284 6792
rect 22336 6780 22342 6792
rect 23753 6783 23811 6789
rect 23753 6780 23765 6783
rect 22336 6752 23765 6780
rect 22336 6740 22342 6752
rect 23753 6749 23765 6752
rect 23799 6749 23811 6783
rect 23934 6780 23940 6792
rect 23895 6752 23940 6780
rect 23753 6743 23811 6749
rect 23934 6740 23940 6752
rect 23992 6740 23998 6792
rect 25130 6740 25136 6792
rect 25188 6780 25194 6792
rect 25498 6780 25504 6792
rect 25188 6752 25504 6780
rect 25188 6740 25194 6752
rect 25498 6740 25504 6752
rect 25556 6740 25562 6792
rect 8202 6712 8208 6724
rect 8163 6684 8208 6712
rect 8202 6672 8208 6684
rect 8260 6672 8266 6724
rect 17405 6715 17463 6721
rect 17405 6681 17417 6715
rect 17451 6712 17463 6715
rect 17494 6712 17500 6724
rect 17451 6684 17500 6712
rect 17451 6681 17463 6684
rect 17405 6675 17463 6681
rect 17494 6672 17500 6684
rect 17552 6712 17558 6724
rect 18138 6712 18144 6724
rect 17552 6684 18144 6712
rect 17552 6672 17558 6684
rect 18138 6672 18144 6684
rect 18196 6672 18202 6724
rect 18598 6712 18604 6724
rect 18559 6684 18604 6712
rect 18598 6672 18604 6684
rect 18656 6672 18662 6724
rect 24949 6715 25007 6721
rect 24949 6681 24961 6715
rect 24995 6712 25007 6715
rect 25038 6712 25044 6724
rect 24995 6684 25044 6712
rect 24995 6681 25007 6684
rect 24949 6675 25007 6681
rect 25038 6672 25044 6684
rect 25096 6672 25102 6724
rect 21082 6644 21088 6656
rect 21043 6616 21088 6644
rect 21082 6604 21088 6616
rect 21140 6604 21146 6656
rect 23385 6647 23443 6653
rect 23385 6613 23397 6647
rect 23431 6644 23443 6647
rect 23474 6644 23480 6656
rect 23431 6616 23480 6644
rect 23431 6613 23443 6616
rect 23385 6607 23443 6613
rect 23474 6604 23480 6616
rect 23532 6604 23538 6656
rect 24118 6604 24124 6656
rect 24176 6644 24182 6656
rect 24305 6647 24363 6653
rect 24305 6644 24317 6647
rect 24176 6616 24317 6644
rect 24176 6604 24182 6616
rect 24305 6613 24317 6616
rect 24351 6613 24363 6647
rect 24305 6607 24363 6613
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 14553 6443 14611 6449
rect 14553 6409 14565 6443
rect 14599 6440 14611 6443
rect 16022 6440 16028 6452
rect 14599 6412 16028 6440
rect 14599 6409 14611 6412
rect 14553 6403 14611 6409
rect 13630 6304 13636 6316
rect 13591 6276 13636 6304
rect 13630 6264 13636 6276
rect 13688 6264 13694 6316
rect 14660 6313 14688 6412
rect 16022 6400 16028 6412
rect 16080 6440 16086 6452
rect 16669 6443 16727 6449
rect 16669 6440 16681 6443
rect 16080 6412 16681 6440
rect 16080 6400 16086 6412
rect 16669 6409 16681 6412
rect 16715 6440 16727 6443
rect 17862 6440 17868 6452
rect 16715 6412 17868 6440
rect 16715 6409 16727 6412
rect 16669 6403 16727 6409
rect 17862 6400 17868 6412
rect 17920 6400 17926 6452
rect 19150 6400 19156 6452
rect 19208 6440 19214 6452
rect 19429 6443 19487 6449
rect 19429 6440 19441 6443
rect 19208 6412 19441 6440
rect 19208 6400 19214 6412
rect 19429 6409 19441 6412
rect 19475 6409 19487 6443
rect 19429 6403 19487 6409
rect 20073 6443 20131 6449
rect 20073 6409 20085 6443
rect 20119 6440 20131 6443
rect 20898 6440 20904 6452
rect 20119 6412 20904 6440
rect 20119 6409 20131 6412
rect 20073 6403 20131 6409
rect 20898 6400 20904 6412
rect 20956 6400 20962 6452
rect 21910 6440 21916 6452
rect 21871 6412 21916 6440
rect 21910 6400 21916 6412
rect 21968 6400 21974 6452
rect 22278 6400 22284 6452
rect 22336 6440 22342 6452
rect 22925 6443 22983 6449
rect 22925 6440 22937 6443
rect 22336 6412 22937 6440
rect 22336 6400 22342 6412
rect 22925 6409 22937 6412
rect 22971 6409 22983 6443
rect 23290 6440 23296 6452
rect 23251 6412 23296 6440
rect 22925 6403 22983 6409
rect 23290 6400 23296 6412
rect 23348 6440 23354 6452
rect 23750 6440 23756 6452
rect 23348 6412 23756 6440
rect 23348 6400 23354 6412
rect 23750 6400 23756 6412
rect 23808 6400 23814 6452
rect 24029 6443 24087 6449
rect 24029 6409 24041 6443
rect 24075 6440 24087 6443
rect 24762 6440 24768 6452
rect 24075 6412 24768 6440
rect 24075 6409 24087 6412
rect 24029 6403 24087 6409
rect 14645 6307 14703 6313
rect 14645 6273 14657 6307
rect 14691 6273 14703 6307
rect 17880 6304 17908 6400
rect 23566 6332 23572 6384
rect 23624 6372 23630 6384
rect 24044 6372 24072 6403
rect 24762 6400 24768 6412
rect 24820 6400 24826 6452
rect 25498 6400 25504 6452
rect 25556 6440 25562 6452
rect 26053 6443 26111 6449
rect 26053 6440 26065 6443
rect 25556 6412 26065 6440
rect 25556 6400 25562 6412
rect 26053 6409 26065 6412
rect 26099 6409 26111 6443
rect 26053 6403 26111 6409
rect 23624 6344 24072 6372
rect 23624 6332 23630 6344
rect 18049 6307 18107 6313
rect 18049 6304 18061 6307
rect 17880 6276 18061 6304
rect 14645 6267 14703 6273
rect 18049 6273 18061 6276
rect 18095 6273 18107 6307
rect 24118 6304 24124 6316
rect 24079 6276 24124 6304
rect 18049 6267 18107 6273
rect 13357 6239 13415 6245
rect 13357 6205 13369 6239
rect 13403 6205 13415 6239
rect 18064 6236 18092 6267
rect 24118 6264 24124 6276
rect 24176 6264 24182 6316
rect 20349 6239 20407 6245
rect 20349 6236 20361 6239
rect 18064 6208 20361 6236
rect 13357 6199 13415 6205
rect 20349 6205 20361 6208
rect 20395 6236 20407 6239
rect 20530 6236 20536 6248
rect 20395 6208 20536 6236
rect 20395 6205 20407 6208
rect 20349 6199 20407 6205
rect 8113 6103 8171 6109
rect 8113 6069 8125 6103
rect 8159 6100 8171 6103
rect 8202 6100 8208 6112
rect 8159 6072 8208 6100
rect 8159 6069 8171 6072
rect 8113 6063 8171 6069
rect 8202 6060 8208 6072
rect 8260 6060 8266 6112
rect 13372 6100 13400 6199
rect 20530 6196 20536 6208
rect 20588 6196 20594 6248
rect 22649 6239 22707 6245
rect 22649 6205 22661 6239
rect 22695 6236 22707 6239
rect 23934 6236 23940 6248
rect 22695 6208 23940 6236
rect 22695 6205 22707 6208
rect 22649 6199 22707 6205
rect 23934 6196 23940 6208
rect 23992 6196 23998 6248
rect 24388 6239 24446 6245
rect 24388 6205 24400 6239
rect 24434 6236 24446 6239
rect 24670 6236 24676 6248
rect 24434 6208 24676 6236
rect 24434 6205 24446 6208
rect 24388 6199 24446 6205
rect 24670 6196 24676 6208
rect 24728 6196 24734 6248
rect 14918 6177 14924 6180
rect 14912 6168 14924 6177
rect 14879 6140 14924 6168
rect 14912 6131 14924 6140
rect 14918 6128 14924 6131
rect 14976 6128 14982 6180
rect 16298 6168 16304 6180
rect 16040 6140 16304 6168
rect 14185 6103 14243 6109
rect 14185 6100 14197 6103
rect 13372 6072 14197 6100
rect 14185 6069 14197 6072
rect 14231 6100 14243 6103
rect 14274 6100 14280 6112
rect 14231 6072 14280 6100
rect 14231 6069 14243 6072
rect 14185 6063 14243 6069
rect 14274 6060 14280 6072
rect 14332 6060 14338 6112
rect 15470 6060 15476 6112
rect 15528 6100 15534 6112
rect 16040 6109 16068 6140
rect 16298 6128 16304 6140
rect 16356 6168 16362 6180
rect 16945 6171 17003 6177
rect 16945 6168 16957 6171
rect 16356 6140 16957 6168
rect 16356 6128 16362 6140
rect 16945 6137 16957 6140
rect 16991 6137 17003 6171
rect 16945 6131 17003 6137
rect 18138 6128 18144 6180
rect 18196 6168 18202 6180
rect 20806 6177 20812 6180
rect 18294 6171 18352 6177
rect 18294 6168 18306 6171
rect 18196 6140 18306 6168
rect 18196 6128 18202 6140
rect 18294 6137 18306 6140
rect 18340 6137 18352 6171
rect 20800 6168 20812 6177
rect 20767 6140 20812 6168
rect 18294 6131 18352 6137
rect 20800 6131 20812 6140
rect 20806 6128 20812 6131
rect 20864 6128 20870 6180
rect 16025 6103 16083 6109
rect 16025 6100 16037 6103
rect 15528 6072 16037 6100
rect 15528 6060 15534 6072
rect 16025 6069 16037 6072
rect 16071 6069 16083 6103
rect 16025 6063 16083 6069
rect 24670 6060 24676 6112
rect 24728 6100 24734 6112
rect 25501 6103 25559 6109
rect 25501 6100 25513 6103
rect 24728 6072 25513 6100
rect 24728 6060 24734 6072
rect 25501 6069 25513 6072
rect 25547 6069 25559 6103
rect 25501 6063 25559 6069
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 18138 5896 18144 5908
rect 18099 5868 18144 5896
rect 18138 5856 18144 5868
rect 18196 5856 18202 5908
rect 18506 5896 18512 5908
rect 18467 5868 18512 5896
rect 18506 5856 18512 5868
rect 18564 5856 18570 5908
rect 19242 5896 19248 5908
rect 19203 5868 19248 5896
rect 19242 5856 19248 5868
rect 19300 5856 19306 5908
rect 19889 5899 19947 5905
rect 19889 5865 19901 5899
rect 19935 5896 19947 5899
rect 19978 5896 19984 5908
rect 19935 5868 19984 5896
rect 19935 5865 19947 5868
rect 19889 5859 19947 5865
rect 19978 5856 19984 5868
rect 20036 5856 20042 5908
rect 20625 5899 20683 5905
rect 20625 5865 20637 5899
rect 20671 5896 20683 5899
rect 20806 5896 20812 5908
rect 20671 5868 20812 5896
rect 20671 5865 20683 5868
rect 20625 5859 20683 5865
rect 20806 5856 20812 5868
rect 20864 5896 20870 5908
rect 22094 5896 22100 5908
rect 20864 5868 22100 5896
rect 20864 5856 20870 5868
rect 22094 5856 22100 5868
rect 22152 5856 22158 5908
rect 22281 5899 22339 5905
rect 22281 5865 22293 5899
rect 22327 5896 22339 5899
rect 22370 5896 22376 5908
rect 22327 5868 22376 5896
rect 22327 5865 22339 5868
rect 22281 5859 22339 5865
rect 22370 5856 22376 5868
rect 22428 5856 22434 5908
rect 25314 5896 25320 5908
rect 25275 5868 25320 5896
rect 25314 5856 25320 5868
rect 25372 5856 25378 5908
rect 13998 5788 14004 5840
rect 14056 5828 14062 5840
rect 15562 5837 15568 5840
rect 14185 5831 14243 5837
rect 14185 5828 14197 5831
rect 14056 5800 14197 5828
rect 14056 5788 14062 5800
rect 14185 5797 14197 5800
rect 14231 5797 14243 5831
rect 15556 5828 15568 5837
rect 15523 5800 15568 5828
rect 14185 5791 14243 5797
rect 15556 5791 15568 5800
rect 15562 5788 15568 5791
rect 15620 5788 15626 5840
rect 18969 5831 19027 5837
rect 18969 5797 18981 5831
rect 19015 5828 19027 5831
rect 19150 5828 19156 5840
rect 19015 5800 19156 5828
rect 19015 5797 19027 5800
rect 18969 5791 19027 5797
rect 19150 5788 19156 5800
rect 19208 5788 19214 5840
rect 23566 5828 23572 5840
rect 20916 5800 23572 5828
rect 13906 5720 13912 5772
rect 13964 5760 13970 5772
rect 14277 5763 14335 5769
rect 14277 5760 14289 5763
rect 13964 5732 14289 5760
rect 13964 5720 13970 5732
rect 14277 5729 14289 5732
rect 14323 5760 14335 5763
rect 14645 5763 14703 5769
rect 14645 5760 14657 5763
rect 14323 5732 14657 5760
rect 14323 5729 14335 5732
rect 14277 5723 14335 5729
rect 14645 5729 14657 5732
rect 14691 5760 14703 5763
rect 14918 5760 14924 5772
rect 14691 5732 14924 5760
rect 14691 5729 14703 5732
rect 14645 5723 14703 5729
rect 14918 5720 14924 5732
rect 14976 5760 14982 5772
rect 15378 5760 15384 5772
rect 14976 5732 15384 5760
rect 14976 5720 14982 5732
rect 15378 5720 15384 5732
rect 15436 5720 15442 5772
rect 19705 5763 19763 5769
rect 19705 5729 19717 5763
rect 19751 5760 19763 5763
rect 19794 5760 19800 5772
rect 19751 5732 19800 5760
rect 19751 5729 19763 5732
rect 19705 5723 19763 5729
rect 19794 5720 19800 5732
rect 19852 5720 19858 5772
rect 20530 5720 20536 5772
rect 20588 5760 20594 5772
rect 20714 5760 20720 5772
rect 20588 5732 20720 5760
rect 20588 5720 20594 5732
rect 20714 5720 20720 5732
rect 20772 5760 20778 5772
rect 20916 5769 20944 5800
rect 20901 5763 20959 5769
rect 20901 5760 20913 5763
rect 20772 5732 20913 5760
rect 20772 5720 20778 5732
rect 20901 5729 20913 5732
rect 20947 5729 20959 5763
rect 20901 5723 20959 5729
rect 21168 5763 21226 5769
rect 21168 5729 21180 5763
rect 21214 5760 21226 5763
rect 21542 5760 21548 5772
rect 21214 5732 21548 5760
rect 21214 5729 21226 5732
rect 21168 5723 21226 5729
rect 21542 5720 21548 5732
rect 21600 5720 21606 5772
rect 23400 5769 23428 5800
rect 23566 5788 23572 5800
rect 23624 5828 23630 5840
rect 24118 5828 24124 5840
rect 23624 5800 24124 5828
rect 23624 5788 23630 5800
rect 24118 5788 24124 5800
rect 24176 5788 24182 5840
rect 23385 5763 23443 5769
rect 23385 5729 23397 5763
rect 23431 5729 23443 5763
rect 23385 5723 23443 5729
rect 23652 5763 23710 5769
rect 23652 5729 23664 5763
rect 23698 5760 23710 5763
rect 23934 5760 23940 5772
rect 23698 5732 23940 5760
rect 23698 5729 23710 5732
rect 23652 5723 23710 5729
rect 23934 5720 23940 5732
rect 23992 5760 23998 5772
rect 24670 5760 24676 5772
rect 23992 5732 24676 5760
rect 23992 5720 23998 5732
rect 24670 5720 24676 5732
rect 24728 5720 24734 5772
rect 14182 5692 14188 5704
rect 14143 5664 14188 5692
rect 14182 5652 14188 5664
rect 14240 5652 14246 5704
rect 15289 5695 15347 5701
rect 15289 5661 15301 5695
rect 15335 5661 15347 5695
rect 15289 5655 15347 5661
rect 13725 5627 13783 5633
rect 13725 5593 13737 5627
rect 13771 5624 13783 5627
rect 14826 5624 14832 5636
rect 13771 5596 14832 5624
rect 13771 5593 13783 5596
rect 13725 5587 13783 5593
rect 14826 5584 14832 5596
rect 14884 5624 14890 5636
rect 15013 5627 15071 5633
rect 15013 5624 15025 5627
rect 14884 5596 15025 5624
rect 14884 5584 14890 5596
rect 15013 5593 15025 5596
rect 15059 5593 15071 5627
rect 15013 5587 15071 5593
rect 15304 5556 15332 5655
rect 16022 5556 16028 5568
rect 15304 5528 16028 5556
rect 16022 5516 16028 5528
rect 16080 5516 16086 5568
rect 16574 5516 16580 5568
rect 16632 5556 16638 5568
rect 16669 5559 16727 5565
rect 16669 5556 16681 5559
rect 16632 5528 16681 5556
rect 16632 5516 16638 5528
rect 16669 5525 16681 5528
rect 16715 5525 16727 5559
rect 24762 5556 24768 5568
rect 24723 5528 24768 5556
rect 16669 5519 16727 5525
rect 24762 5516 24768 5528
rect 24820 5516 24826 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 13265 5355 13323 5361
rect 13265 5321 13277 5355
rect 13311 5352 13323 5355
rect 13906 5352 13912 5364
rect 13311 5324 13912 5352
rect 13311 5321 13323 5324
rect 13265 5315 13323 5321
rect 13906 5312 13912 5324
rect 13964 5312 13970 5364
rect 14182 5352 14188 5364
rect 14143 5324 14188 5352
rect 14182 5312 14188 5324
rect 14240 5312 14246 5364
rect 14274 5312 14280 5364
rect 14332 5352 14338 5364
rect 14461 5355 14519 5361
rect 14461 5352 14473 5355
rect 14332 5324 14473 5352
rect 14332 5312 14338 5324
rect 14461 5321 14473 5324
rect 14507 5321 14519 5355
rect 14461 5315 14519 5321
rect 15841 5355 15899 5361
rect 15841 5321 15853 5355
rect 15887 5352 15899 5355
rect 16482 5352 16488 5364
rect 15887 5324 16488 5352
rect 15887 5321 15899 5324
rect 15841 5315 15899 5321
rect 13357 5219 13415 5225
rect 13357 5185 13369 5219
rect 13403 5216 13415 5219
rect 14200 5216 14228 5312
rect 15194 5244 15200 5296
rect 15252 5284 15258 5296
rect 15856 5284 15884 5315
rect 16482 5312 16488 5324
rect 16540 5312 16546 5364
rect 20530 5352 20536 5364
rect 20491 5324 20536 5352
rect 20530 5312 20536 5324
rect 20588 5312 20594 5364
rect 22094 5312 22100 5364
rect 22152 5352 22158 5364
rect 23017 5355 23075 5361
rect 23017 5352 23029 5355
rect 22152 5324 23029 5352
rect 22152 5312 22158 5324
rect 23017 5321 23029 5324
rect 23063 5352 23075 5355
rect 24762 5352 24768 5364
rect 23063 5324 24768 5352
rect 23063 5321 23075 5324
rect 23017 5315 23075 5321
rect 24320 5296 24348 5324
rect 24762 5312 24768 5324
rect 24820 5312 24826 5364
rect 15252 5256 15884 5284
rect 16025 5287 16083 5293
rect 15252 5244 15258 5256
rect 16025 5253 16037 5287
rect 16071 5253 16083 5287
rect 19794 5284 19800 5296
rect 19755 5256 19800 5284
rect 16025 5247 16083 5253
rect 14826 5216 14832 5228
rect 13403 5188 14228 5216
rect 14787 5188 14832 5216
rect 13403 5185 13415 5188
rect 13357 5179 13415 5185
rect 14826 5176 14832 5188
rect 14884 5176 14890 5228
rect 15473 5219 15531 5225
rect 15473 5185 15485 5219
rect 15519 5216 15531 5219
rect 15565 5219 15623 5225
rect 15565 5216 15577 5219
rect 15519 5188 15577 5216
rect 15519 5185 15531 5188
rect 15473 5179 15531 5185
rect 15565 5185 15577 5188
rect 15611 5185 15623 5219
rect 15565 5179 15623 5185
rect 16040 5148 16068 5247
rect 19794 5244 19800 5256
rect 19852 5244 19858 5296
rect 23477 5287 23535 5293
rect 23477 5253 23489 5287
rect 23523 5284 23535 5287
rect 23566 5284 23572 5296
rect 23523 5256 23572 5284
rect 23523 5253 23535 5256
rect 23477 5247 23535 5253
rect 23566 5244 23572 5256
rect 23624 5244 23630 5296
rect 23753 5287 23811 5293
rect 23753 5253 23765 5287
rect 23799 5253 23811 5287
rect 23753 5247 23811 5253
rect 16482 5216 16488 5228
rect 16443 5188 16488 5216
rect 16482 5176 16488 5188
rect 16540 5176 16546 5228
rect 19337 5219 19395 5225
rect 19337 5216 19349 5219
rect 18616 5188 19349 5216
rect 14936 5120 16068 5148
rect 14826 5040 14832 5092
rect 14884 5080 14890 5092
rect 14936 5089 14964 5120
rect 18322 5108 18328 5160
rect 18380 5148 18386 5160
rect 18616 5157 18644 5188
rect 19337 5185 19349 5188
rect 19383 5185 19395 5219
rect 20990 5216 20996 5228
rect 20951 5188 20996 5216
rect 19337 5179 19395 5185
rect 20990 5176 20996 5188
rect 21048 5176 21054 5228
rect 18601 5151 18659 5157
rect 18601 5148 18613 5151
rect 18380 5120 18613 5148
rect 18380 5108 18386 5120
rect 18601 5117 18613 5120
rect 18647 5117 18659 5151
rect 18874 5148 18880 5160
rect 18835 5120 18880 5148
rect 18601 5111 18659 5117
rect 18874 5108 18880 5120
rect 18932 5108 18938 5160
rect 20257 5151 20315 5157
rect 20257 5117 20269 5151
rect 20303 5148 20315 5151
rect 20622 5148 20628 5160
rect 20303 5120 20628 5148
rect 20303 5117 20315 5120
rect 20257 5111 20315 5117
rect 20622 5108 20628 5120
rect 20680 5148 20686 5160
rect 20717 5151 20775 5157
rect 20717 5148 20729 5151
rect 20680 5120 20729 5148
rect 20680 5108 20686 5120
rect 20717 5117 20729 5120
rect 20763 5117 20775 5151
rect 22465 5151 22523 5157
rect 22465 5148 22477 5151
rect 20717 5111 20775 5117
rect 22296 5120 22477 5148
rect 22296 5092 22324 5120
rect 22465 5117 22477 5120
rect 22511 5117 22523 5151
rect 23768 5148 23796 5247
rect 24302 5244 24308 5296
rect 24360 5244 24366 5296
rect 24670 5284 24676 5296
rect 24631 5256 24676 5284
rect 24670 5244 24676 5256
rect 24728 5244 24734 5296
rect 23842 5176 23848 5228
rect 23900 5216 23906 5228
rect 24213 5219 24271 5225
rect 24213 5216 24225 5219
rect 23900 5188 24225 5216
rect 23900 5176 23906 5188
rect 24213 5185 24225 5188
rect 24259 5216 24271 5219
rect 25041 5219 25099 5225
rect 25041 5216 25053 5219
rect 24259 5188 25053 5216
rect 24259 5185 24271 5188
rect 24213 5179 24271 5185
rect 25041 5185 25053 5188
rect 25087 5185 25099 5219
rect 25406 5216 25412 5228
rect 25367 5188 25412 5216
rect 25041 5179 25099 5185
rect 25406 5176 25412 5188
rect 25464 5176 25470 5228
rect 25225 5151 25283 5157
rect 25225 5148 25237 5151
rect 23768 5120 25237 5148
rect 22465 5111 22523 5117
rect 25225 5117 25237 5120
rect 25271 5148 25283 5151
rect 25961 5151 26019 5157
rect 25961 5148 25973 5151
rect 25271 5120 25973 5148
rect 25271 5117 25283 5120
rect 25225 5111 25283 5117
rect 25961 5117 25973 5120
rect 26007 5117 26019 5151
rect 25961 5111 26019 5117
rect 14921 5083 14979 5089
rect 14921 5080 14933 5083
rect 14884 5052 14933 5080
rect 14884 5040 14890 5052
rect 14921 5049 14933 5052
rect 14967 5049 14979 5083
rect 14921 5043 14979 5049
rect 15010 5040 15016 5092
rect 15068 5080 15074 5092
rect 15470 5080 15476 5092
rect 15068 5052 15476 5080
rect 15068 5040 15074 5052
rect 15470 5040 15476 5052
rect 15528 5040 15534 5092
rect 15565 5083 15623 5089
rect 15565 5049 15577 5083
rect 15611 5080 15623 5083
rect 16022 5080 16028 5092
rect 15611 5052 16028 5080
rect 15611 5049 15623 5052
rect 15565 5043 15623 5049
rect 16022 5040 16028 5052
rect 16080 5040 16086 5092
rect 16574 5080 16580 5092
rect 16535 5052 16580 5080
rect 16574 5040 16580 5052
rect 16632 5040 16638 5092
rect 22278 5080 22284 5092
rect 22239 5052 22284 5080
rect 22278 5040 22284 5052
rect 22336 5040 22342 5092
rect 24302 5080 24308 5092
rect 24263 5052 24308 5080
rect 24302 5040 24308 5052
rect 24360 5040 24366 5092
rect 13906 5012 13912 5024
rect 13867 4984 13912 5012
rect 13906 4972 13912 4984
rect 13964 4972 13970 5024
rect 14550 4972 14556 5024
rect 14608 5012 14614 5024
rect 16485 5015 16543 5021
rect 16485 5012 16497 5015
rect 14608 4984 16497 5012
rect 14608 4972 14614 4984
rect 16485 4981 16497 4984
rect 16531 5012 16543 5015
rect 16945 5015 17003 5021
rect 16945 5012 16957 5015
rect 16531 4984 16957 5012
rect 16531 4981 16543 4984
rect 16485 4975 16543 4981
rect 16945 4981 16957 4984
rect 16991 4981 17003 5015
rect 21542 5012 21548 5024
rect 21503 4984 21548 5012
rect 16945 4975 17003 4981
rect 21542 4972 21548 4984
rect 21600 4972 21606 5024
rect 22646 5012 22652 5024
rect 22607 4984 22652 5012
rect 22646 4972 22652 4984
rect 22704 4972 22710 5024
rect 23474 4972 23480 5024
rect 23532 5012 23538 5024
rect 24210 5012 24216 5024
rect 23532 4984 24216 5012
rect 23532 4972 23538 4984
rect 24210 4972 24216 4984
rect 24268 4972 24274 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 14826 4808 14832 4820
rect 14787 4780 14832 4808
rect 14826 4768 14832 4780
rect 14884 4768 14890 4820
rect 15378 4768 15384 4820
rect 15436 4808 15442 4820
rect 16209 4811 16267 4817
rect 16209 4808 16221 4811
rect 15436 4780 16221 4808
rect 15436 4768 15442 4780
rect 16209 4777 16221 4780
rect 16255 4808 16267 4811
rect 16574 4808 16580 4820
rect 16255 4780 16580 4808
rect 16255 4777 16267 4780
rect 16209 4771 16267 4777
rect 16574 4768 16580 4780
rect 16632 4768 16638 4820
rect 23014 4768 23020 4820
rect 23072 4808 23078 4820
rect 23845 4811 23903 4817
rect 23845 4808 23857 4811
rect 23072 4780 23857 4808
rect 23072 4768 23078 4780
rect 23845 4777 23857 4780
rect 23891 4777 23903 4811
rect 23845 4771 23903 4777
rect 24210 4768 24216 4820
rect 24268 4808 24274 4820
rect 24305 4811 24363 4817
rect 24305 4808 24317 4811
rect 24268 4780 24317 4808
rect 24268 4768 24274 4780
rect 24305 4777 24317 4780
rect 24351 4777 24363 4811
rect 24305 4771 24363 4777
rect 14461 4743 14519 4749
rect 14461 4709 14473 4743
rect 14507 4740 14519 4743
rect 15010 4740 15016 4752
rect 14507 4712 15016 4740
rect 14507 4709 14519 4712
rect 14461 4703 14519 4709
rect 15010 4700 15016 4712
rect 15068 4700 15074 4752
rect 15562 4700 15568 4752
rect 15620 4740 15626 4752
rect 15841 4743 15899 4749
rect 15841 4740 15853 4743
rect 15620 4712 15853 4740
rect 15620 4700 15626 4712
rect 15841 4709 15853 4712
rect 15887 4709 15899 4743
rect 23934 4740 23940 4752
rect 23895 4712 23940 4740
rect 15841 4703 15899 4709
rect 23934 4700 23940 4712
rect 23992 4700 23998 4752
rect 13354 4672 13360 4684
rect 13315 4644 13360 4672
rect 13354 4632 13360 4644
rect 13412 4632 13418 4684
rect 15289 4675 15347 4681
rect 15289 4641 15301 4675
rect 15335 4672 15347 4675
rect 15654 4672 15660 4684
rect 15335 4644 15660 4672
rect 15335 4641 15347 4644
rect 15289 4635 15347 4641
rect 15654 4632 15660 4644
rect 15712 4632 15718 4684
rect 19794 4672 19800 4684
rect 19755 4644 19800 4672
rect 19794 4632 19800 4644
rect 19852 4632 19858 4684
rect 21818 4672 21824 4684
rect 21779 4644 21824 4672
rect 21818 4632 21824 4644
rect 21876 4632 21882 4684
rect 23658 4672 23664 4684
rect 23619 4644 23664 4672
rect 23658 4632 23664 4644
rect 23716 4632 23722 4684
rect 24857 4675 24915 4681
rect 24857 4641 24869 4675
rect 24903 4672 24915 4675
rect 25222 4672 25228 4684
rect 24903 4644 25228 4672
rect 24903 4641 24915 4644
rect 24857 4635 24915 4641
rect 25222 4632 25228 4644
rect 25280 4632 25286 4684
rect 23385 4539 23443 4545
rect 23385 4505 23397 4539
rect 23431 4536 23443 4539
rect 23842 4536 23848 4548
rect 23431 4508 23848 4536
rect 23431 4505 23443 4508
rect 23385 4499 23443 4505
rect 23842 4496 23848 4508
rect 23900 4496 23906 4548
rect 13538 4468 13544 4480
rect 13499 4440 13544 4468
rect 13538 4428 13544 4440
rect 13596 4428 13602 4480
rect 15473 4471 15531 4477
rect 15473 4437 15485 4471
rect 15519 4468 15531 4471
rect 15562 4468 15568 4480
rect 15519 4440 15568 4468
rect 15519 4437 15531 4440
rect 15473 4431 15531 4437
rect 15562 4428 15568 4440
rect 15620 4428 15626 4480
rect 22005 4471 22063 4477
rect 22005 4437 22017 4471
rect 22051 4468 22063 4471
rect 22094 4468 22100 4480
rect 22051 4440 22100 4468
rect 22051 4437 22063 4440
rect 22005 4431 22063 4437
rect 22094 4428 22100 4440
rect 22152 4428 22158 4480
rect 25038 4468 25044 4480
rect 24999 4440 25044 4468
rect 25038 4428 25044 4440
rect 25096 4428 25102 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 21818 4264 21824 4276
rect 21779 4236 21824 4264
rect 21818 4224 21824 4236
rect 21876 4224 21882 4276
rect 23658 4224 23664 4276
rect 23716 4264 23722 4276
rect 23845 4267 23903 4273
rect 23845 4264 23857 4267
rect 23716 4236 23857 4264
rect 23716 4224 23722 4236
rect 23845 4233 23857 4236
rect 23891 4233 23903 4267
rect 23845 4227 23903 4233
rect 4890 4088 4896 4140
rect 4948 4128 4954 4140
rect 5350 4128 5356 4140
rect 4948 4100 5356 4128
rect 4948 4088 4954 4100
rect 5350 4088 5356 4100
rect 5408 4088 5414 4140
rect 13265 4131 13323 4137
rect 13265 4097 13277 4131
rect 13311 4128 13323 4131
rect 13446 4128 13452 4140
rect 13311 4100 13452 4128
rect 13311 4097 13323 4100
rect 13265 4091 13323 4097
rect 4246 4020 4252 4072
rect 4304 4060 4310 4072
rect 5442 4060 5448 4072
rect 4304 4032 5448 4060
rect 4304 4020 4310 4032
rect 5442 4020 5448 4032
rect 5500 4020 5506 4072
rect 13372 4069 13400 4100
rect 13446 4088 13452 4100
rect 13504 4088 13510 4140
rect 15286 4128 15292 4140
rect 14752 4100 15292 4128
rect 14752 4069 14780 4100
rect 15286 4088 15292 4100
rect 15344 4088 15350 4140
rect 19337 4131 19395 4137
rect 19337 4128 19349 4131
rect 18708 4100 19349 4128
rect 13357 4063 13415 4069
rect 13357 4029 13369 4063
rect 13403 4060 13415 4063
rect 14737 4063 14795 4069
rect 13403 4032 13437 4060
rect 13403 4029 13415 4032
rect 13357 4023 13415 4029
rect 14737 4029 14749 4063
rect 14783 4029 14795 4063
rect 15838 4060 15844 4072
rect 15799 4032 15844 4060
rect 14737 4023 14795 4029
rect 15838 4020 15844 4032
rect 15896 4060 15902 4072
rect 18708 4069 18736 4100
rect 19337 4097 19349 4100
rect 19383 4128 19395 4131
rect 20162 4128 20168 4140
rect 19383 4100 20168 4128
rect 19383 4097 19395 4100
rect 19337 4091 19395 4097
rect 20162 4088 20168 4100
rect 20220 4088 20226 4140
rect 23014 4088 23020 4140
rect 23072 4128 23078 4140
rect 23198 4128 23204 4140
rect 23072 4100 23204 4128
rect 23072 4088 23078 4100
rect 23198 4088 23204 4100
rect 23256 4128 23262 4140
rect 23293 4131 23351 4137
rect 23293 4128 23305 4131
rect 23256 4100 23305 4128
rect 23256 4088 23262 4100
rect 23293 4097 23305 4100
rect 23339 4097 23351 4131
rect 25958 4128 25964 4140
rect 23293 4091 23351 4097
rect 25424 4100 25964 4128
rect 16577 4063 16635 4069
rect 16577 4060 16589 4063
rect 15896 4032 16589 4060
rect 15896 4020 15902 4032
rect 16577 4029 16589 4032
rect 16623 4029 16635 4063
rect 16577 4023 16635 4029
rect 18693 4063 18751 4069
rect 18693 4029 18705 4063
rect 18739 4029 18751 4063
rect 19794 4060 19800 4072
rect 19755 4032 19800 4060
rect 18693 4023 18751 4029
rect 19794 4020 19800 4032
rect 19852 4060 19858 4072
rect 20349 4063 20407 4069
rect 20349 4060 20361 4063
rect 19852 4032 20361 4060
rect 19852 4020 19858 4032
rect 20349 4029 20361 4032
rect 20395 4029 20407 4063
rect 20349 4023 20407 4029
rect 20438 4020 20444 4072
rect 20496 4060 20502 4072
rect 20901 4063 20959 4069
rect 20901 4060 20913 4063
rect 20496 4032 20913 4060
rect 20496 4020 20502 4032
rect 20901 4029 20913 4032
rect 20947 4060 20959 4063
rect 21453 4063 21511 4069
rect 21453 4060 21465 4063
rect 20947 4032 21465 4060
rect 20947 4029 20959 4032
rect 20901 4023 20959 4029
rect 21453 4029 21465 4032
rect 21499 4029 21511 4063
rect 21453 4023 21511 4029
rect 22373 4063 22431 4069
rect 22373 4029 22385 4063
rect 22419 4060 22431 4063
rect 22465 4063 22523 4069
rect 22465 4060 22477 4063
rect 22419 4032 22477 4060
rect 22419 4029 22431 4032
rect 22373 4023 22431 4029
rect 22465 4029 22477 4032
rect 22511 4060 22523 4063
rect 22554 4060 22560 4072
rect 22511 4032 22560 4060
rect 22511 4029 22523 4032
rect 22465 4023 22523 4029
rect 22554 4020 22560 4032
rect 22612 4020 22618 4072
rect 23750 4020 23756 4072
rect 23808 4060 23814 4072
rect 24305 4063 24363 4069
rect 24305 4060 24317 4063
rect 23808 4032 24317 4060
rect 23808 4020 23814 4032
rect 24305 4029 24317 4032
rect 24351 4060 24363 4063
rect 24857 4063 24915 4069
rect 24857 4060 24869 4063
rect 24351 4032 24869 4060
rect 24351 4029 24363 4032
rect 24305 4023 24363 4029
rect 24857 4029 24869 4032
rect 24903 4029 24915 4063
rect 25222 4060 25228 4072
rect 25183 4032 25228 4060
rect 24857 4023 24915 4029
rect 25222 4020 25228 4032
rect 25280 4020 25286 4072
rect 25424 4069 25452 4100
rect 25958 4088 25964 4100
rect 26016 4088 26022 4140
rect 25409 4063 25467 4069
rect 25409 4029 25421 4063
rect 25455 4029 25467 4063
rect 25409 4023 25467 4029
rect 13630 3992 13636 4004
rect 13591 3964 13636 3992
rect 13630 3952 13636 3964
rect 13688 3952 13694 4004
rect 16114 3992 16120 4004
rect 16075 3964 16120 3992
rect 16114 3952 16120 3964
rect 16172 3952 16178 4004
rect 26878 3992 26884 4004
rect 25608 3964 26884 3992
rect 13354 3884 13360 3936
rect 13412 3924 13418 3936
rect 14093 3927 14151 3933
rect 14093 3924 14105 3927
rect 13412 3896 14105 3924
rect 13412 3884 13418 3896
rect 14093 3893 14105 3896
rect 14139 3893 14151 3927
rect 14918 3924 14924 3936
rect 14879 3896 14924 3924
rect 14093 3887 14151 3893
rect 14918 3884 14924 3896
rect 14976 3884 14982 3936
rect 15654 3924 15660 3936
rect 15615 3896 15660 3924
rect 15654 3884 15660 3896
rect 15712 3884 15718 3936
rect 18874 3924 18880 3936
rect 18835 3896 18880 3924
rect 18874 3884 18880 3896
rect 18932 3884 18938 3936
rect 19978 3924 19984 3936
rect 19939 3896 19984 3924
rect 19978 3884 19984 3896
rect 20036 3884 20042 3936
rect 21082 3924 21088 3936
rect 21043 3896 21088 3924
rect 21082 3884 21088 3896
rect 21140 3884 21146 3936
rect 21818 3884 21824 3936
rect 21876 3924 21882 3936
rect 22186 3924 22192 3936
rect 21876 3896 22192 3924
rect 21876 3884 21882 3896
rect 22186 3884 22192 3896
rect 22244 3884 22250 3936
rect 22646 3924 22652 3936
rect 22607 3896 22652 3924
rect 22646 3884 22652 3896
rect 22704 3884 22710 3936
rect 24486 3924 24492 3936
rect 24447 3896 24492 3924
rect 24486 3884 24492 3896
rect 24544 3884 24550 3936
rect 25608 3933 25636 3964
rect 26878 3952 26884 3964
rect 26936 3952 26942 4004
rect 25593 3927 25651 3933
rect 25593 3893 25605 3927
rect 25639 3893 25651 3927
rect 25593 3887 25651 3893
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 18509 3723 18567 3729
rect 18509 3689 18521 3723
rect 18555 3720 18567 3723
rect 18690 3720 18696 3732
rect 18555 3692 18696 3720
rect 18555 3689 18567 3692
rect 18509 3683 18567 3689
rect 18690 3680 18696 3692
rect 18748 3680 18754 3732
rect 20438 3720 20444 3732
rect 20399 3692 20444 3720
rect 20438 3680 20444 3692
rect 20496 3680 20502 3732
rect 23934 3720 23940 3732
rect 23895 3692 23940 3720
rect 23934 3680 23940 3692
rect 23992 3680 23998 3732
rect 13630 3652 13636 3664
rect 13591 3624 13636 3652
rect 13630 3612 13636 3624
rect 13688 3612 13694 3664
rect 10226 3584 10232 3596
rect 10187 3556 10232 3584
rect 10226 3544 10232 3556
rect 10284 3544 10290 3596
rect 12253 3587 12311 3593
rect 12253 3553 12265 3587
rect 12299 3584 12311 3587
rect 12710 3584 12716 3596
rect 12299 3556 12716 3584
rect 12299 3553 12311 3556
rect 12253 3547 12311 3553
rect 12710 3544 12716 3556
rect 12768 3544 12774 3596
rect 13078 3544 13084 3596
rect 13136 3584 13142 3596
rect 13357 3587 13415 3593
rect 13357 3584 13369 3587
rect 13136 3556 13369 3584
rect 13136 3544 13142 3556
rect 13357 3553 13369 3556
rect 13403 3553 13415 3587
rect 13357 3547 13415 3553
rect 15933 3587 15991 3593
rect 15933 3553 15945 3587
rect 15979 3584 15991 3587
rect 16022 3584 16028 3596
rect 15979 3556 16028 3584
rect 15979 3553 15991 3556
rect 15933 3547 15991 3553
rect 16022 3544 16028 3556
rect 16080 3584 16086 3596
rect 16390 3584 16396 3596
rect 16080 3556 16396 3584
rect 16080 3544 16086 3556
rect 16390 3544 16396 3556
rect 16448 3544 16454 3596
rect 17218 3584 17224 3596
rect 17179 3556 17224 3584
rect 17218 3544 17224 3556
rect 17276 3544 17282 3596
rect 18322 3584 18328 3596
rect 18283 3556 18328 3584
rect 18322 3544 18328 3556
rect 18380 3544 18386 3596
rect 19429 3587 19487 3593
rect 19429 3553 19441 3587
rect 19475 3584 19487 3587
rect 20346 3584 20352 3596
rect 19475 3556 20352 3584
rect 19475 3553 19487 3556
rect 19429 3547 19487 3553
rect 20346 3544 20352 3556
rect 20404 3544 20410 3596
rect 20901 3587 20959 3593
rect 20901 3553 20913 3587
rect 20947 3584 20959 3587
rect 21174 3584 21180 3596
rect 20947 3556 21180 3584
rect 20947 3553 20959 3556
rect 20901 3547 20959 3553
rect 21174 3544 21180 3556
rect 21232 3544 21238 3596
rect 22002 3584 22008 3596
rect 21963 3556 22008 3584
rect 22002 3544 22008 3556
rect 22060 3544 22066 3596
rect 22922 3544 22928 3596
rect 22980 3584 22986 3596
rect 23109 3587 23167 3593
rect 23109 3584 23121 3587
rect 22980 3556 23121 3584
rect 22980 3544 22986 3556
rect 23109 3553 23121 3556
rect 23155 3584 23167 3587
rect 23290 3584 23296 3596
rect 23155 3556 23296 3584
rect 23155 3553 23167 3556
rect 23109 3547 23167 3553
rect 23290 3544 23296 3556
rect 23348 3544 23354 3596
rect 23385 3587 23443 3593
rect 23385 3553 23397 3587
rect 23431 3584 23443 3587
rect 24581 3587 24639 3593
rect 24581 3584 24593 3587
rect 23431 3556 24593 3584
rect 23431 3553 23443 3556
rect 23385 3547 23443 3553
rect 24581 3553 24593 3556
rect 24627 3584 24639 3587
rect 24762 3584 24768 3596
rect 24627 3556 24768 3584
rect 24627 3553 24639 3556
rect 24581 3547 24639 3553
rect 24762 3544 24768 3556
rect 24820 3544 24826 3596
rect 10505 3519 10563 3525
rect 10505 3485 10517 3519
rect 10551 3516 10563 3519
rect 11054 3516 11060 3528
rect 10551 3488 11060 3516
rect 10551 3485 10563 3488
rect 10505 3479 10563 3485
rect 11054 3476 11060 3488
rect 11112 3476 11118 3528
rect 15378 3476 15384 3528
rect 15436 3516 15442 3528
rect 16117 3519 16175 3525
rect 16117 3516 16129 3519
rect 15436 3488 16129 3516
rect 15436 3476 15442 3488
rect 16117 3485 16129 3488
rect 16163 3485 16175 3519
rect 19610 3516 19616 3528
rect 19571 3488 19616 3516
rect 16117 3479 16175 3485
rect 19610 3476 19616 3488
rect 19668 3476 19674 3528
rect 12437 3383 12495 3389
rect 12437 3349 12449 3383
rect 12483 3380 12495 3383
rect 14274 3380 14280 3392
rect 12483 3352 14280 3380
rect 12483 3349 12495 3352
rect 12437 3343 12495 3349
rect 14274 3340 14280 3352
rect 14332 3340 14338 3392
rect 17405 3383 17463 3389
rect 17405 3349 17417 3383
rect 17451 3380 17463 3383
rect 17586 3380 17592 3392
rect 17451 3352 17592 3380
rect 17451 3349 17463 3352
rect 17405 3343 17463 3349
rect 17586 3340 17592 3352
rect 17644 3340 17650 3392
rect 21082 3380 21088 3392
rect 21043 3352 21088 3380
rect 21082 3340 21088 3352
rect 21140 3340 21146 3392
rect 22189 3383 22247 3389
rect 22189 3349 22201 3383
rect 22235 3380 22247 3383
rect 23382 3380 23388 3392
rect 22235 3352 23388 3380
rect 22235 3349 22247 3352
rect 22189 3343 22247 3349
rect 23382 3340 23388 3352
rect 23440 3340 23446 3392
rect 24118 3340 24124 3392
rect 24176 3380 24182 3392
rect 24765 3383 24823 3389
rect 24765 3380 24777 3383
rect 24176 3352 24777 3380
rect 24176 3340 24182 3352
rect 24765 3349 24777 3352
rect 24811 3349 24823 3383
rect 24765 3343 24823 3349
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 10226 3176 10232 3188
rect 10187 3148 10232 3176
rect 10226 3136 10232 3148
rect 10284 3136 10290 3188
rect 13078 3136 13084 3188
rect 13136 3176 13142 3188
rect 14001 3179 14059 3185
rect 14001 3176 14013 3179
rect 13136 3148 14013 3176
rect 13136 3136 13142 3148
rect 14001 3145 14013 3148
rect 14047 3145 14059 3179
rect 16022 3176 16028 3188
rect 15983 3148 16028 3176
rect 14001 3139 14059 3145
rect 16022 3136 16028 3148
rect 16080 3136 16086 3188
rect 16666 3176 16672 3188
rect 16627 3148 16672 3176
rect 16666 3136 16672 3148
rect 16724 3136 16730 3188
rect 17218 3136 17224 3188
rect 17276 3176 17282 3188
rect 17405 3179 17463 3185
rect 17405 3176 17417 3179
rect 17276 3148 17417 3176
rect 17276 3136 17282 3148
rect 17405 3145 17417 3148
rect 17451 3145 17463 3179
rect 18322 3176 18328 3188
rect 18283 3148 18328 3176
rect 17405 3139 17463 3145
rect 18322 3136 18328 3148
rect 18380 3136 18386 3188
rect 18414 3136 18420 3188
rect 18472 3176 18478 3188
rect 18693 3179 18751 3185
rect 18693 3176 18705 3179
rect 18472 3148 18705 3176
rect 18472 3136 18478 3148
rect 18693 3145 18705 3148
rect 18739 3145 18751 3179
rect 19426 3176 19432 3188
rect 19387 3148 19432 3176
rect 18693 3139 18751 3145
rect 19426 3136 19432 3148
rect 19484 3136 19490 3188
rect 20257 3179 20315 3185
rect 20257 3145 20269 3179
rect 20303 3176 20315 3179
rect 20346 3176 20352 3188
rect 20303 3148 20352 3176
rect 20303 3145 20315 3148
rect 20257 3139 20315 3145
rect 20346 3136 20352 3148
rect 20404 3136 20410 3188
rect 21174 3176 21180 3188
rect 21135 3148 21180 3176
rect 21174 3136 21180 3148
rect 21232 3136 21238 3188
rect 23106 3176 23112 3188
rect 23067 3148 23112 3176
rect 23106 3136 23112 3148
rect 23164 3136 23170 3188
rect 23290 3136 23296 3188
rect 23348 3176 23354 3188
rect 23385 3179 23443 3185
rect 23385 3176 23397 3179
rect 23348 3148 23397 3176
rect 23348 3136 23354 3148
rect 23385 3145 23397 3148
rect 23431 3145 23443 3179
rect 23385 3139 23443 3145
rect 24026 3136 24032 3188
rect 24084 3176 24090 3188
rect 24397 3179 24455 3185
rect 24397 3176 24409 3179
rect 24084 3148 24409 3176
rect 24084 3136 24090 3148
rect 24397 3145 24409 3148
rect 24443 3145 24455 3179
rect 24762 3176 24768 3188
rect 24723 3148 24768 3176
rect 24397 3139 24455 3145
rect 24762 3136 24768 3148
rect 24820 3136 24826 3188
rect 13262 3108 13268 3120
rect 12912 3080 13268 3108
rect 7742 2932 7748 2984
rect 7800 2972 7806 2984
rect 8665 2975 8723 2981
rect 8665 2972 8677 2975
rect 7800 2944 8677 2972
rect 7800 2932 7806 2944
rect 8665 2941 8677 2944
rect 8711 2972 8723 2975
rect 9401 2975 9459 2981
rect 9401 2972 9413 2975
rect 8711 2944 9413 2972
rect 8711 2941 8723 2944
rect 8665 2935 8723 2941
rect 9401 2941 9413 2944
rect 9447 2941 9459 2975
rect 9401 2935 9459 2941
rect 10042 2932 10048 2984
rect 10100 2972 10106 2984
rect 12912 2981 12940 3080
rect 13262 3068 13268 3080
rect 13320 3108 13326 3120
rect 13633 3111 13691 3117
rect 13633 3108 13645 3111
rect 13320 3080 13645 3108
rect 13320 3068 13326 3080
rect 13633 3077 13645 3080
rect 13679 3077 13691 3111
rect 13633 3071 13691 3077
rect 13173 3043 13231 3049
rect 13173 3009 13185 3043
rect 13219 3040 13231 3043
rect 13354 3040 13360 3052
rect 13219 3012 13360 3040
rect 13219 3009 13231 3012
rect 13173 3003 13231 3009
rect 13354 3000 13360 3012
rect 13412 3000 13418 3052
rect 22097 3043 22155 3049
rect 22097 3009 22109 3043
rect 22143 3040 22155 3043
rect 23845 3043 23903 3049
rect 23845 3040 23857 3043
rect 22143 3012 23857 3040
rect 22143 3009 22155 3012
rect 22097 3003 22155 3009
rect 23845 3009 23857 3012
rect 23891 3009 23903 3043
rect 23845 3003 23903 3009
rect 10873 2975 10931 2981
rect 10873 2972 10885 2975
rect 10100 2944 10885 2972
rect 10100 2932 10106 2944
rect 10873 2941 10885 2944
rect 10919 2972 10931 2975
rect 11609 2975 11667 2981
rect 11609 2972 11621 2975
rect 10919 2944 11621 2972
rect 10919 2941 10931 2944
rect 10873 2935 10931 2941
rect 11609 2941 11621 2944
rect 11655 2941 11667 2975
rect 11609 2935 11667 2941
rect 12897 2975 12955 2981
rect 12897 2941 12909 2975
rect 12943 2941 12955 2975
rect 12897 2935 12955 2941
rect 14734 2932 14740 2984
rect 14792 2972 14798 2984
rect 14829 2975 14887 2981
rect 14829 2972 14841 2975
rect 14792 2944 14841 2972
rect 14792 2932 14798 2944
rect 14829 2941 14841 2944
rect 14875 2972 14887 2975
rect 15565 2975 15623 2981
rect 15565 2972 15577 2975
rect 14875 2944 15577 2972
rect 14875 2941 14887 2944
rect 14829 2935 14887 2941
rect 15565 2941 15577 2944
rect 15611 2941 15623 2975
rect 15565 2935 15623 2941
rect 16666 2932 16672 2984
rect 16724 2972 16730 2984
rect 16853 2975 16911 2981
rect 16853 2972 16865 2975
rect 16724 2944 16865 2972
rect 16724 2932 16730 2944
rect 16853 2941 16865 2944
rect 16899 2941 16911 2975
rect 16853 2935 16911 2941
rect 18141 2975 18199 2981
rect 18141 2941 18153 2975
rect 18187 2941 18199 2975
rect 19242 2972 19248 2984
rect 19203 2944 19248 2972
rect 18141 2935 18199 2941
rect 8941 2907 8999 2913
rect 8941 2873 8953 2907
rect 8987 2904 8999 2907
rect 9582 2904 9588 2916
rect 8987 2876 9588 2904
rect 8987 2873 8999 2876
rect 8941 2867 8999 2873
rect 9582 2864 9588 2876
rect 9640 2864 9646 2916
rect 11149 2907 11207 2913
rect 11149 2873 11161 2907
rect 11195 2904 11207 2907
rect 12434 2904 12440 2916
rect 11195 2876 12440 2904
rect 11195 2873 11207 2876
rect 11149 2867 11207 2873
rect 12434 2864 12440 2876
rect 12492 2864 12498 2916
rect 12710 2904 12716 2916
rect 12623 2876 12716 2904
rect 12710 2864 12716 2876
rect 12768 2904 12774 2916
rect 15105 2907 15163 2913
rect 15105 2904 15117 2907
rect 12768 2876 15117 2904
rect 12768 2864 12774 2876
rect 15105 2873 15117 2876
rect 15151 2873 15163 2907
rect 17770 2904 17776 2916
rect 17731 2876 17776 2904
rect 15105 2867 15163 2873
rect 17770 2864 17776 2876
rect 17828 2904 17834 2916
rect 18156 2904 18184 2935
rect 19242 2932 19248 2944
rect 19300 2972 19306 2984
rect 19797 2975 19855 2981
rect 19797 2972 19809 2975
rect 19300 2944 19809 2972
rect 19300 2932 19306 2944
rect 19797 2941 19809 2944
rect 19843 2941 19855 2975
rect 19797 2935 19855 2941
rect 20349 2975 20407 2981
rect 20349 2941 20361 2975
rect 20395 2972 20407 2975
rect 20438 2972 20444 2984
rect 20395 2944 20444 2972
rect 20395 2941 20407 2944
rect 20349 2935 20407 2941
rect 20438 2932 20444 2944
rect 20496 2932 20502 2984
rect 20622 2904 20628 2916
rect 17828 2876 18184 2904
rect 20583 2876 20628 2904
rect 17828 2864 17834 2876
rect 20622 2864 20628 2876
rect 20680 2864 20686 2916
rect 22002 2864 22008 2916
rect 22060 2904 22066 2916
rect 22112 2904 22140 3003
rect 22281 2975 22339 2981
rect 22281 2941 22293 2975
rect 22327 2972 22339 2975
rect 23106 2972 23112 2984
rect 22327 2944 23112 2972
rect 22327 2941 22339 2944
rect 22281 2935 22339 2941
rect 23106 2932 23112 2944
rect 23164 2932 23170 2984
rect 23661 2975 23719 2981
rect 23661 2941 23673 2975
rect 23707 2972 23719 2975
rect 24026 2972 24032 2984
rect 23707 2944 24032 2972
rect 23707 2941 23719 2944
rect 23661 2935 23719 2941
rect 24026 2932 24032 2944
rect 24084 2932 24090 2984
rect 24854 2932 24860 2984
rect 24912 2972 24918 2984
rect 24949 2975 25007 2981
rect 24949 2972 24961 2975
rect 24912 2944 24961 2972
rect 24912 2932 24918 2944
rect 24949 2941 24961 2944
rect 24995 2972 25007 2975
rect 25501 2975 25559 2981
rect 25501 2972 25513 2975
rect 24995 2944 25513 2972
rect 24995 2941 25007 2944
rect 24949 2935 25007 2941
rect 25501 2941 25513 2944
rect 25547 2941 25559 2975
rect 25501 2935 25559 2941
rect 22060 2876 22140 2904
rect 22060 2864 22066 2876
rect 22186 2864 22192 2916
rect 22244 2904 22250 2916
rect 22557 2907 22615 2913
rect 22557 2904 22569 2907
rect 22244 2876 22569 2904
rect 22244 2864 22250 2876
rect 22557 2873 22569 2876
rect 22603 2873 22615 2907
rect 22557 2867 22615 2873
rect 17034 2836 17040 2848
rect 16995 2808 17040 2836
rect 17034 2796 17040 2808
rect 17092 2796 17098 2848
rect 24854 2796 24860 2848
rect 24912 2836 24918 2848
rect 25133 2839 25191 2845
rect 25133 2836 25145 2839
rect 24912 2808 25145 2836
rect 24912 2796 24918 2808
rect 25133 2805 25145 2808
rect 25179 2805 25191 2839
rect 25133 2799 25191 2805
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 14921 2635 14979 2641
rect 14921 2601 14933 2635
rect 14967 2632 14979 2635
rect 15378 2632 15384 2644
rect 14967 2604 15384 2632
rect 14967 2601 14979 2604
rect 14921 2595 14979 2601
rect 11054 2456 11060 2508
rect 11112 2496 11118 2508
rect 11149 2499 11207 2505
rect 11149 2496 11161 2499
rect 11112 2468 11161 2496
rect 11112 2456 11118 2468
rect 11149 2465 11161 2468
rect 11195 2496 11207 2499
rect 11701 2499 11759 2505
rect 11701 2496 11713 2499
rect 11195 2468 11713 2496
rect 11195 2465 11207 2468
rect 11149 2459 11207 2465
rect 11701 2465 11713 2468
rect 11747 2465 11759 2499
rect 11701 2459 11759 2465
rect 12434 2456 12440 2508
rect 12492 2496 12498 2508
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12492 2468 12633 2496
rect 12492 2456 12498 2468
rect 12621 2465 12633 2468
rect 12667 2496 12679 2499
rect 13173 2499 13231 2505
rect 13173 2496 13185 2499
rect 12667 2468 13185 2496
rect 12667 2465 12679 2468
rect 12621 2459 12679 2465
rect 13173 2465 13185 2468
rect 13219 2465 13231 2499
rect 13173 2459 13231 2465
rect 14277 2499 14335 2505
rect 14277 2465 14289 2499
rect 14323 2496 14335 2499
rect 14936 2496 14964 2595
rect 15378 2592 15384 2604
rect 15436 2592 15442 2644
rect 16206 2632 16212 2644
rect 16167 2604 16212 2632
rect 16206 2592 16212 2604
rect 16264 2592 16270 2644
rect 17773 2635 17831 2641
rect 17773 2601 17785 2635
rect 17819 2632 17831 2635
rect 17862 2632 17868 2644
rect 17819 2604 17868 2632
rect 17819 2601 17831 2604
rect 17773 2595 17831 2601
rect 14323 2468 14964 2496
rect 14323 2465 14335 2468
rect 14277 2459 14335 2465
rect 15930 2456 15936 2508
rect 15988 2496 15994 2508
rect 16025 2499 16083 2505
rect 16025 2496 16037 2499
rect 15988 2468 16037 2496
rect 15988 2456 15994 2468
rect 16025 2465 16037 2468
rect 16071 2496 16083 2499
rect 16577 2499 16635 2505
rect 16577 2496 16589 2499
rect 16071 2468 16589 2496
rect 16071 2465 16083 2468
rect 16025 2459 16083 2465
rect 16577 2465 16589 2468
rect 16623 2465 16635 2499
rect 16577 2459 16635 2465
rect 17129 2499 17187 2505
rect 17129 2465 17141 2499
rect 17175 2496 17187 2499
rect 17788 2496 17816 2595
rect 17862 2592 17868 2604
rect 17920 2592 17926 2644
rect 18782 2632 18788 2644
rect 18743 2604 18788 2632
rect 18782 2592 18788 2604
rect 18840 2592 18846 2644
rect 20254 2632 20260 2644
rect 20215 2604 20260 2632
rect 20254 2592 20260 2604
rect 20312 2592 20318 2644
rect 22373 2635 22431 2641
rect 22373 2601 22385 2635
rect 22419 2632 22431 2635
rect 22554 2632 22560 2644
rect 22419 2604 22560 2632
rect 22419 2601 22431 2604
rect 22373 2595 22431 2601
rect 17175 2468 17816 2496
rect 18601 2499 18659 2505
rect 17175 2465 17187 2468
rect 17129 2459 17187 2465
rect 18601 2465 18613 2499
rect 18647 2496 18659 2499
rect 18690 2496 18696 2508
rect 18647 2468 18696 2496
rect 18647 2465 18659 2468
rect 18601 2459 18659 2465
rect 18690 2456 18696 2468
rect 18748 2496 18754 2508
rect 19153 2499 19211 2505
rect 19153 2496 19165 2499
rect 18748 2468 19165 2496
rect 18748 2456 18754 2468
rect 19153 2465 19165 2468
rect 19199 2465 19211 2499
rect 19153 2459 19211 2465
rect 19705 2499 19763 2505
rect 19705 2465 19717 2499
rect 19751 2496 19763 2499
rect 20272 2496 20300 2592
rect 19751 2468 20300 2496
rect 21729 2499 21787 2505
rect 19751 2465 19763 2468
rect 19705 2459 19763 2465
rect 21729 2465 21741 2499
rect 21775 2496 21787 2499
rect 22388 2496 22416 2595
rect 22554 2592 22560 2604
rect 22612 2592 22618 2644
rect 23014 2632 23020 2644
rect 22975 2604 23020 2632
rect 23014 2592 23020 2604
rect 23072 2592 23078 2644
rect 22830 2496 22836 2508
rect 21775 2468 22416 2496
rect 22791 2468 22836 2496
rect 21775 2465 21787 2468
rect 21729 2459 21787 2465
rect 22830 2456 22836 2468
rect 22888 2496 22894 2508
rect 23385 2499 23443 2505
rect 23385 2496 23397 2499
rect 22888 2468 23397 2496
rect 22888 2456 22894 2468
rect 23385 2465 23397 2468
rect 23431 2465 23443 2499
rect 24578 2496 24584 2508
rect 24539 2468 24584 2496
rect 23385 2459 23443 2465
rect 24578 2456 24584 2468
rect 24636 2496 24642 2508
rect 25133 2499 25191 2505
rect 25133 2496 25145 2499
rect 24636 2468 25145 2496
rect 24636 2456 24642 2468
rect 25133 2465 25145 2468
rect 25179 2465 25191 2499
rect 25133 2459 25191 2465
rect 12802 2360 12808 2372
rect 12763 2332 12808 2360
rect 12802 2320 12808 2332
rect 12860 2320 12866 2372
rect 14461 2363 14519 2369
rect 14461 2329 14473 2363
rect 14507 2360 14519 2363
rect 16850 2360 16856 2372
rect 14507 2332 16856 2360
rect 14507 2329 14519 2332
rect 14461 2323 14519 2329
rect 16850 2320 16856 2332
rect 16908 2320 16914 2372
rect 17313 2363 17371 2369
rect 17313 2329 17325 2363
rect 17359 2360 17371 2363
rect 19518 2360 19524 2372
rect 17359 2332 19524 2360
rect 17359 2329 17371 2332
rect 17313 2323 17371 2329
rect 19518 2320 19524 2332
rect 19576 2320 19582 2372
rect 19889 2363 19947 2369
rect 19889 2329 19901 2363
rect 19935 2360 19947 2363
rect 20898 2360 20904 2372
rect 19935 2332 20904 2360
rect 19935 2329 19947 2332
rect 19889 2323 19947 2329
rect 20898 2320 20904 2332
rect 20956 2320 20962 2372
rect 11330 2292 11336 2304
rect 11291 2264 11336 2292
rect 11330 2252 11336 2264
rect 11388 2252 11394 2304
rect 21910 2292 21916 2304
rect 21871 2264 21916 2292
rect 21910 2252 21916 2264
rect 21968 2252 21974 2304
rect 24762 2292 24768 2304
rect 24723 2264 24768 2292
rect 24762 2252 24768 2264
rect 24820 2252 24826 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 13538 552 13544 604
rect 13596 592 13602 604
rect 13906 592 13912 604
rect 13596 564 13912 592
rect 13596 552 13602 564
rect 13906 552 13912 564
rect 13964 552 13970 604
<< via1 >>
rect 12992 27412 13044 27464
rect 13176 27412 13228 27464
rect 22192 26256 22244 26308
rect 24584 26256 24636 26308
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 15936 25440 15988 25492
rect 20076 25440 20128 25492
rect 9956 25372 10008 25424
rect 10324 25347 10376 25356
rect 10324 25313 10333 25347
rect 10333 25313 10367 25347
rect 10367 25313 10376 25347
rect 10324 25304 10376 25313
rect 12716 25304 12768 25356
rect 19156 25347 19208 25356
rect 19156 25313 19165 25347
rect 19165 25313 19199 25347
rect 19199 25313 19208 25347
rect 19156 25304 19208 25313
rect 19984 25304 20036 25356
rect 24768 25304 24820 25356
rect 9864 25236 9916 25288
rect 11060 25236 11112 25288
rect 16212 25236 16264 25288
rect 10876 25168 10928 25220
rect 11244 25100 11296 25152
rect 12440 25100 12492 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 12716 24896 12768 24948
rect 9956 24871 10008 24880
rect 6000 24760 6052 24812
rect 9956 24837 9965 24871
rect 9965 24837 9999 24871
rect 9999 24837 10008 24871
rect 9956 24828 10008 24837
rect 10324 24871 10376 24880
rect 10324 24837 10333 24871
rect 10333 24837 10367 24871
rect 10367 24837 10376 24871
rect 10324 24828 10376 24837
rect 10784 24828 10836 24880
rect 8300 24760 8352 24812
rect 10876 24735 10928 24744
rect 7196 24667 7248 24676
rect 7196 24633 7205 24667
rect 7205 24633 7239 24667
rect 7239 24633 7248 24667
rect 7196 24624 7248 24633
rect 10876 24701 10885 24735
rect 10885 24701 10919 24735
rect 10919 24701 10928 24735
rect 10876 24692 10928 24701
rect 14004 24760 14056 24812
rect 19524 24760 19576 24812
rect 19984 24803 20036 24812
rect 19984 24769 19993 24803
rect 19993 24769 20027 24803
rect 20027 24769 20036 24803
rect 19984 24760 20036 24769
rect 21548 24760 21600 24812
rect 23572 24828 23624 24880
rect 22468 24760 22520 24812
rect 11060 24667 11112 24676
rect 11060 24633 11069 24667
rect 11069 24633 11103 24667
rect 11103 24633 11112 24667
rect 11060 24624 11112 24633
rect 11244 24624 11296 24676
rect 11980 24624 12032 24676
rect 13084 24624 13136 24676
rect 14096 24624 14148 24676
rect 7564 24556 7616 24608
rect 9864 24556 9916 24608
rect 10048 24556 10100 24608
rect 14556 24556 14608 24608
rect 16304 24692 16356 24744
rect 17776 24692 17828 24744
rect 18512 24692 18564 24744
rect 20904 24692 20956 24744
rect 22284 24692 22336 24744
rect 15476 24556 15528 24608
rect 16488 24624 16540 24676
rect 19156 24624 19208 24676
rect 16304 24599 16356 24608
rect 16304 24565 16313 24599
rect 16313 24565 16347 24599
rect 16347 24565 16356 24599
rect 16304 24556 16356 24565
rect 17868 24556 17920 24608
rect 18604 24599 18656 24608
rect 18604 24565 18613 24599
rect 18613 24565 18647 24599
rect 18647 24565 18656 24599
rect 18604 24556 18656 24565
rect 19432 24599 19484 24608
rect 19432 24565 19441 24599
rect 19441 24565 19475 24599
rect 19475 24565 19484 24599
rect 20076 24599 20128 24608
rect 19432 24556 19484 24565
rect 20076 24565 20085 24599
rect 20085 24565 20119 24599
rect 20119 24565 20128 24599
rect 20076 24556 20128 24565
rect 20352 24556 20404 24608
rect 21364 24556 21416 24608
rect 23388 24624 23440 24676
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 6368 24352 6420 24404
rect 7196 24352 7248 24404
rect 7564 24395 7616 24404
rect 7564 24361 7573 24395
rect 7573 24361 7607 24395
rect 7607 24361 7616 24395
rect 7564 24352 7616 24361
rect 8300 24395 8352 24404
rect 8300 24361 8309 24395
rect 8309 24361 8343 24395
rect 8343 24361 8352 24395
rect 8300 24352 8352 24361
rect 13084 24395 13136 24404
rect 13084 24361 13093 24395
rect 13093 24361 13127 24395
rect 13127 24361 13136 24395
rect 13084 24352 13136 24361
rect 17316 24352 17368 24404
rect 19248 24352 19300 24404
rect 21548 24395 21600 24404
rect 21548 24361 21557 24395
rect 21557 24361 21591 24395
rect 21591 24361 21600 24395
rect 21548 24352 21600 24361
rect 22744 24395 22796 24404
rect 22744 24361 22753 24395
rect 22753 24361 22787 24395
rect 22787 24361 22796 24395
rect 22744 24352 22796 24361
rect 24124 24352 24176 24404
rect 26884 24352 26936 24404
rect 9864 24284 9916 24336
rect 10876 24284 10928 24336
rect 14004 24284 14056 24336
rect 15844 24327 15896 24336
rect 15844 24293 15853 24327
rect 15853 24293 15887 24327
rect 15887 24293 15896 24327
rect 15844 24284 15896 24293
rect 19616 24327 19668 24336
rect 19616 24293 19625 24327
rect 19625 24293 19659 24327
rect 19659 24293 19668 24327
rect 19616 24284 19668 24293
rect 8024 24216 8076 24268
rect 12256 24216 12308 24268
rect 13544 24216 13596 24268
rect 16856 24259 16908 24268
rect 16856 24225 16865 24259
rect 16865 24225 16899 24259
rect 16899 24225 16908 24259
rect 16856 24216 16908 24225
rect 17592 24216 17644 24268
rect 19432 24216 19484 24268
rect 22560 24259 22612 24268
rect 22560 24225 22569 24259
rect 22569 24225 22603 24259
rect 22603 24225 22612 24259
rect 22560 24216 22612 24225
rect 24216 24216 24268 24268
rect 24860 24216 24912 24268
rect 8116 24148 8168 24200
rect 9680 24148 9732 24200
rect 10508 24191 10560 24200
rect 10508 24157 10517 24191
rect 10517 24157 10551 24191
rect 10551 24157 10560 24191
rect 10508 24148 10560 24157
rect 14464 24148 14516 24200
rect 15752 24191 15804 24200
rect 15752 24157 15761 24191
rect 15761 24157 15795 24191
rect 15795 24157 15804 24191
rect 15752 24148 15804 24157
rect 15936 24191 15988 24200
rect 15936 24157 15945 24191
rect 15945 24157 15979 24191
rect 15979 24157 15988 24191
rect 15936 24148 15988 24157
rect 19524 24191 19576 24200
rect 19524 24157 19533 24191
rect 19533 24157 19567 24191
rect 19567 24157 19576 24191
rect 19524 24148 19576 24157
rect 21456 24191 21508 24200
rect 21456 24157 21465 24191
rect 21465 24157 21499 24191
rect 21499 24157 21508 24191
rect 21456 24148 21508 24157
rect 21640 24191 21692 24200
rect 21640 24157 21649 24191
rect 21649 24157 21683 24191
rect 21683 24157 21692 24191
rect 21640 24148 21692 24157
rect 19064 24080 19116 24132
rect 21088 24123 21140 24132
rect 21088 24089 21097 24123
rect 21097 24089 21131 24123
rect 21131 24089 21140 24123
rect 21088 24080 21140 24089
rect 7840 24055 7892 24064
rect 7840 24021 7849 24055
rect 7849 24021 7883 24055
rect 7883 24021 7892 24055
rect 7840 24012 7892 24021
rect 10416 24055 10468 24064
rect 10416 24021 10425 24055
rect 10425 24021 10459 24055
rect 10459 24021 10468 24055
rect 10416 24012 10468 24021
rect 10784 24012 10836 24064
rect 11980 24012 12032 24064
rect 12440 24055 12492 24064
rect 12440 24021 12449 24055
rect 12449 24021 12483 24055
rect 12483 24021 12492 24055
rect 12440 24012 12492 24021
rect 13820 24012 13872 24064
rect 15384 24055 15436 24064
rect 15384 24021 15393 24055
rect 15393 24021 15427 24055
rect 15427 24021 15436 24055
rect 15384 24012 15436 24021
rect 16396 24055 16448 24064
rect 16396 24021 16405 24055
rect 16405 24021 16439 24055
rect 16439 24021 16448 24055
rect 16396 24012 16448 24021
rect 18880 24055 18932 24064
rect 18880 24021 18889 24055
rect 18889 24021 18923 24055
rect 18923 24021 18932 24055
rect 18880 24012 18932 24021
rect 19156 24055 19208 24064
rect 19156 24021 19165 24055
rect 19165 24021 19199 24055
rect 19199 24021 19208 24055
rect 19156 24012 19208 24021
rect 19340 24012 19392 24064
rect 19984 24012 20036 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 9864 23851 9916 23860
rect 9864 23817 9873 23851
rect 9873 23817 9907 23851
rect 9907 23817 9916 23851
rect 9864 23808 9916 23817
rect 10508 23808 10560 23860
rect 12256 23851 12308 23860
rect 10048 23740 10100 23792
rect 9864 23672 9916 23724
rect 10140 23672 10192 23724
rect 10968 23715 11020 23724
rect 7656 23604 7708 23656
rect 8300 23604 8352 23656
rect 10968 23681 10977 23715
rect 10977 23681 11011 23715
rect 11011 23681 11020 23715
rect 10968 23672 11020 23681
rect 12256 23817 12265 23851
rect 12265 23817 12299 23851
rect 12299 23817 12308 23851
rect 12256 23808 12308 23817
rect 12624 23851 12676 23860
rect 12624 23817 12633 23851
rect 12633 23817 12667 23851
rect 12667 23817 12676 23851
rect 12624 23808 12676 23817
rect 14464 23808 14516 23860
rect 15936 23808 15988 23860
rect 16488 23851 16540 23860
rect 16488 23817 16497 23851
rect 16497 23817 16531 23851
rect 16531 23817 16540 23851
rect 16488 23808 16540 23817
rect 21548 23808 21600 23860
rect 22100 23808 22152 23860
rect 24676 23808 24728 23860
rect 24952 23851 25004 23860
rect 24952 23817 24961 23851
rect 24961 23817 24995 23851
rect 24995 23817 25004 23851
rect 24952 23808 25004 23817
rect 18328 23783 18380 23792
rect 18328 23749 18337 23783
rect 18337 23749 18371 23783
rect 18371 23749 18380 23783
rect 18328 23740 18380 23749
rect 21456 23740 21508 23792
rect 23296 23740 23348 23792
rect 16396 23672 16448 23724
rect 18972 23672 19024 23724
rect 8116 23536 8168 23588
rect 10416 23536 10468 23588
rect 7012 23468 7064 23520
rect 8024 23468 8076 23520
rect 9588 23468 9640 23520
rect 10140 23511 10192 23520
rect 10140 23477 10149 23511
rect 10149 23477 10183 23511
rect 10183 23477 10192 23511
rect 10140 23468 10192 23477
rect 12440 23647 12492 23656
rect 12440 23613 12449 23647
rect 12449 23613 12483 23647
rect 12483 23613 12492 23647
rect 12440 23604 12492 23613
rect 13636 23604 13688 23656
rect 17868 23604 17920 23656
rect 20996 23604 21048 23656
rect 14096 23536 14148 23588
rect 16120 23536 16172 23588
rect 18880 23579 18932 23588
rect 12348 23468 12400 23520
rect 15108 23468 15160 23520
rect 15844 23468 15896 23520
rect 18880 23545 18889 23579
rect 18889 23545 18923 23579
rect 18923 23545 18932 23579
rect 18880 23536 18932 23545
rect 17592 23468 17644 23520
rect 19064 23468 19116 23520
rect 19432 23468 19484 23520
rect 21272 23511 21324 23520
rect 21272 23477 21281 23511
rect 21281 23477 21315 23511
rect 21315 23477 21324 23511
rect 21272 23468 21324 23477
rect 24216 23647 24268 23656
rect 24216 23613 24225 23647
rect 24225 23613 24259 23647
rect 24259 23613 24268 23647
rect 24216 23604 24268 23613
rect 23940 23536 23992 23588
rect 23112 23468 23164 23520
rect 23480 23511 23532 23520
rect 23480 23477 23489 23511
rect 23489 23477 23523 23511
rect 23523 23477 23532 23511
rect 23480 23468 23532 23477
rect 23848 23468 23900 23520
rect 24860 23468 24912 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 8300 23264 8352 23316
rect 11060 23264 11112 23316
rect 12624 23264 12676 23316
rect 13268 23264 13320 23316
rect 14004 23307 14056 23316
rect 14004 23273 14013 23307
rect 14013 23273 14047 23307
rect 14047 23273 14056 23307
rect 14004 23264 14056 23273
rect 15108 23307 15160 23316
rect 15108 23273 15117 23307
rect 15117 23273 15151 23307
rect 15151 23273 15160 23307
rect 15108 23264 15160 23273
rect 19524 23264 19576 23316
rect 22560 23264 22612 23316
rect 22836 23264 22888 23316
rect 24768 23307 24820 23316
rect 24768 23273 24777 23307
rect 24777 23273 24811 23307
rect 24811 23273 24820 23307
rect 24768 23264 24820 23273
rect 11980 23196 12032 23248
rect 14464 23196 14516 23248
rect 15936 23196 15988 23248
rect 21272 23239 21324 23248
rect 21272 23205 21306 23239
rect 21306 23205 21324 23239
rect 21272 23196 21324 23205
rect 6644 23128 6696 23180
rect 8208 23128 8260 23180
rect 12072 23128 12124 23180
rect 7012 23103 7064 23112
rect 7012 23069 7021 23103
rect 7021 23069 7055 23103
rect 7055 23069 7064 23103
rect 7012 23060 7064 23069
rect 9680 23060 9732 23112
rect 12440 23060 12492 23112
rect 13268 23103 13320 23112
rect 13268 23069 13277 23103
rect 13277 23069 13311 23103
rect 13311 23069 13320 23103
rect 13268 23060 13320 23069
rect 14188 23103 14240 23112
rect 14188 23069 14197 23103
rect 14197 23069 14231 23103
rect 14231 23069 14240 23103
rect 14188 23060 14240 23069
rect 15292 23103 15344 23112
rect 15292 23069 15301 23103
rect 15301 23069 15335 23103
rect 15335 23069 15344 23103
rect 15292 23060 15344 23069
rect 20996 23171 21048 23180
rect 20996 23137 21005 23171
rect 21005 23137 21039 23171
rect 21039 23137 21048 23171
rect 20996 23128 21048 23137
rect 24860 23128 24912 23180
rect 17684 23060 17736 23112
rect 9588 22924 9640 22976
rect 10876 22924 10928 22976
rect 12072 22967 12124 22976
rect 12072 22933 12081 22967
rect 12081 22933 12115 22967
rect 12115 22933 12124 22967
rect 12072 22924 12124 22933
rect 12808 22924 12860 22976
rect 16672 22967 16724 22976
rect 16672 22933 16681 22967
rect 16681 22933 16715 22967
rect 16715 22933 16724 22967
rect 16672 22924 16724 22933
rect 16856 22924 16908 22976
rect 18880 22924 18932 22976
rect 19432 22924 19484 22976
rect 20720 22967 20772 22976
rect 20720 22933 20729 22967
rect 20729 22933 20763 22967
rect 20763 22933 20772 22967
rect 20720 22924 20772 22933
rect 21640 22924 21692 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 6644 22763 6696 22772
rect 6644 22729 6653 22763
rect 6653 22729 6687 22763
rect 6687 22729 6696 22763
rect 6644 22720 6696 22729
rect 11980 22720 12032 22772
rect 13268 22720 13320 22772
rect 14464 22763 14516 22772
rect 14464 22729 14473 22763
rect 14473 22729 14507 22763
rect 14507 22729 14516 22763
rect 14464 22720 14516 22729
rect 16948 22763 17000 22772
rect 16948 22729 16957 22763
rect 16957 22729 16991 22763
rect 16991 22729 17000 22763
rect 16948 22720 17000 22729
rect 20996 22720 21048 22772
rect 24676 22720 24728 22772
rect 10324 22695 10376 22704
rect 10324 22661 10333 22695
rect 10333 22661 10367 22695
rect 10367 22661 10376 22695
rect 10324 22652 10376 22661
rect 11060 22652 11112 22704
rect 11796 22695 11848 22704
rect 11796 22661 11805 22695
rect 11805 22661 11839 22695
rect 11839 22661 11848 22695
rect 11796 22652 11848 22661
rect 12532 22695 12584 22704
rect 12532 22661 12541 22695
rect 12541 22661 12575 22695
rect 12575 22661 12584 22695
rect 12532 22652 12584 22661
rect 14556 22652 14608 22704
rect 21640 22652 21692 22704
rect 10876 22627 10928 22636
rect 10876 22593 10885 22627
rect 10885 22593 10919 22627
rect 10919 22593 10928 22627
rect 10876 22584 10928 22593
rect 13084 22627 13136 22636
rect 13084 22593 13093 22627
rect 13093 22593 13127 22627
rect 13127 22593 13136 22627
rect 13084 22584 13136 22593
rect 16672 22584 16724 22636
rect 21364 22584 21416 22636
rect 7012 22516 7064 22568
rect 8024 22559 8076 22568
rect 8024 22525 8058 22559
rect 8058 22525 8076 22559
rect 8024 22516 8076 22525
rect 10140 22516 10192 22568
rect 12808 22491 12860 22500
rect 12808 22457 12817 22491
rect 12817 22457 12851 22491
rect 12851 22457 12860 22491
rect 12808 22448 12860 22457
rect 15384 22559 15436 22568
rect 15384 22525 15393 22559
rect 15393 22525 15427 22559
rect 15427 22525 15436 22559
rect 15384 22516 15436 22525
rect 16764 22559 16816 22568
rect 16764 22525 16773 22559
rect 16773 22525 16807 22559
rect 16807 22525 16816 22559
rect 16764 22516 16816 22525
rect 13452 22448 13504 22500
rect 15292 22448 15344 22500
rect 17684 22448 17736 22500
rect 21272 22516 21324 22568
rect 18696 22448 18748 22500
rect 21364 22491 21416 22500
rect 21364 22457 21373 22491
rect 21373 22457 21407 22491
rect 21407 22457 21416 22491
rect 21364 22448 21416 22457
rect 21548 22491 21600 22500
rect 21548 22457 21557 22491
rect 21557 22457 21591 22491
rect 21591 22457 21600 22491
rect 21548 22448 21600 22457
rect 7656 22423 7708 22432
rect 7656 22389 7665 22423
rect 7665 22389 7699 22423
rect 7699 22389 7708 22423
rect 7656 22380 7708 22389
rect 8300 22380 8352 22432
rect 9680 22423 9732 22432
rect 9680 22389 9689 22423
rect 9689 22389 9723 22423
rect 9723 22389 9732 22423
rect 9680 22380 9732 22389
rect 10784 22423 10836 22432
rect 10784 22389 10793 22423
rect 10793 22389 10827 22423
rect 10827 22389 10836 22423
rect 10784 22380 10836 22389
rect 15108 22380 15160 22432
rect 19432 22380 19484 22432
rect 24216 22380 24268 22432
rect 24860 22380 24912 22432
rect 25780 22380 25832 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 6644 22219 6696 22228
rect 6644 22185 6653 22219
rect 6653 22185 6687 22219
rect 6687 22185 6696 22219
rect 6644 22176 6696 22185
rect 7840 22176 7892 22228
rect 10140 22176 10192 22228
rect 11888 22176 11940 22228
rect 12624 22176 12676 22228
rect 16304 22176 16356 22228
rect 16764 22176 16816 22228
rect 17224 22176 17276 22228
rect 17776 22219 17828 22228
rect 17776 22185 17785 22219
rect 17785 22185 17819 22219
rect 17819 22185 17828 22219
rect 17776 22176 17828 22185
rect 8024 22108 8076 22160
rect 8300 22151 8352 22160
rect 8300 22117 8309 22151
rect 8309 22117 8343 22151
rect 8343 22117 8352 22151
rect 11796 22151 11848 22160
rect 8300 22108 8352 22117
rect 11796 22117 11805 22151
rect 11805 22117 11839 22151
rect 11839 22117 11848 22151
rect 11796 22108 11848 22117
rect 14004 22151 14056 22160
rect 14004 22117 14013 22151
rect 14013 22117 14047 22151
rect 14047 22117 14056 22151
rect 14004 22108 14056 22117
rect 14648 22108 14700 22160
rect 17868 22151 17920 22160
rect 17868 22117 17877 22151
rect 17877 22117 17911 22151
rect 17911 22117 17920 22151
rect 17868 22108 17920 22117
rect 18696 22108 18748 22160
rect 19248 22176 19300 22228
rect 21272 22176 21324 22228
rect 19340 22151 19392 22160
rect 19340 22117 19349 22151
rect 19349 22117 19383 22151
rect 19383 22117 19392 22151
rect 19340 22108 19392 22117
rect 22192 22151 22244 22160
rect 22192 22117 22201 22151
rect 22201 22117 22235 22151
rect 22235 22117 22244 22151
rect 22192 22108 22244 22117
rect 11520 22083 11572 22092
rect 11520 22049 11529 22083
rect 11529 22049 11563 22083
rect 11563 22049 11572 22083
rect 11520 22040 11572 22049
rect 11704 22040 11756 22092
rect 13820 22040 13872 22092
rect 15108 22040 15160 22092
rect 19156 22040 19208 22092
rect 23020 22040 23072 22092
rect 7380 21972 7432 22024
rect 8208 21972 8260 22024
rect 14096 22015 14148 22024
rect 12072 21904 12124 21956
rect 13544 21947 13596 21956
rect 13544 21913 13553 21947
rect 13553 21913 13587 21947
rect 13587 21913 13596 21947
rect 13544 21904 13596 21913
rect 14096 21981 14105 22015
rect 14105 21981 14139 22015
rect 14139 21981 14148 22015
rect 14096 21972 14148 21981
rect 16212 22015 16264 22024
rect 16212 21981 16221 22015
rect 16221 21981 16255 22015
rect 16255 21981 16264 22015
rect 16212 21972 16264 21981
rect 16396 21972 16448 22024
rect 17776 22015 17828 22024
rect 17776 21981 17785 22015
rect 17785 21981 17819 22015
rect 17819 21981 17828 22015
rect 17776 21972 17828 21981
rect 14188 21904 14240 21956
rect 15752 21947 15804 21956
rect 15752 21913 15761 21947
rect 15761 21913 15795 21947
rect 15795 21913 15804 21947
rect 15752 21904 15804 21913
rect 19432 22015 19484 22024
rect 18880 21947 18932 21956
rect 18880 21913 18889 21947
rect 18889 21913 18923 21947
rect 18923 21913 18932 21947
rect 18880 21904 18932 21913
rect 19432 21981 19441 22015
rect 19441 21981 19475 22015
rect 19475 21981 19484 22015
rect 19432 21972 19484 21981
rect 22376 21972 22428 22024
rect 23204 22015 23256 22024
rect 23204 21981 23213 22015
rect 23213 21981 23247 22015
rect 23247 21981 23256 22015
rect 23204 21972 23256 21981
rect 7748 21879 7800 21888
rect 7748 21845 7757 21879
rect 7757 21845 7791 21879
rect 7791 21845 7800 21879
rect 7748 21836 7800 21845
rect 11336 21836 11388 21888
rect 13176 21879 13228 21888
rect 13176 21845 13185 21879
rect 13185 21845 13219 21879
rect 13219 21845 13228 21879
rect 13176 21836 13228 21845
rect 15568 21879 15620 21888
rect 15568 21845 15577 21879
rect 15577 21845 15611 21879
rect 15611 21845 15620 21879
rect 15568 21836 15620 21845
rect 16028 21836 16080 21888
rect 16488 21836 16540 21888
rect 16672 21879 16724 21888
rect 16672 21845 16681 21879
rect 16681 21845 16715 21879
rect 16715 21845 16724 21879
rect 16672 21836 16724 21845
rect 20168 21879 20220 21888
rect 20168 21845 20177 21879
rect 20177 21845 20211 21879
rect 20211 21845 20220 21879
rect 20168 21836 20220 21845
rect 21548 21836 21600 21888
rect 23480 21836 23532 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 14004 21632 14056 21684
rect 14740 21632 14792 21684
rect 16212 21632 16264 21684
rect 17224 21632 17276 21684
rect 17776 21675 17828 21684
rect 17776 21641 17785 21675
rect 17785 21641 17819 21675
rect 17819 21641 17828 21675
rect 17776 21632 17828 21641
rect 19340 21675 19392 21684
rect 19340 21641 19349 21675
rect 19349 21641 19383 21675
rect 19383 21641 19392 21675
rect 19340 21632 19392 21641
rect 20352 21675 20404 21684
rect 20352 21641 20361 21675
rect 20361 21641 20395 21675
rect 20395 21641 20404 21675
rect 20352 21632 20404 21641
rect 12808 21607 12860 21616
rect 7656 21496 7708 21548
rect 12808 21573 12817 21607
rect 12817 21573 12851 21607
rect 12851 21573 12860 21607
rect 12808 21564 12860 21573
rect 13912 21564 13964 21616
rect 11152 21539 11204 21548
rect 11152 21505 11161 21539
rect 11161 21505 11195 21539
rect 11195 21505 11204 21539
rect 11152 21496 11204 21505
rect 11336 21539 11388 21548
rect 11336 21505 11345 21539
rect 11345 21505 11379 21539
rect 11379 21505 11388 21539
rect 11336 21496 11388 21505
rect 17592 21564 17644 21616
rect 16856 21539 16908 21548
rect 16856 21505 16865 21539
rect 16865 21505 16899 21539
rect 16899 21505 16908 21539
rect 16856 21496 16908 21505
rect 21732 21564 21784 21616
rect 18972 21496 19024 21548
rect 19984 21496 20036 21548
rect 21180 21496 21232 21548
rect 22468 21496 22520 21548
rect 24216 21539 24268 21548
rect 24216 21505 24225 21539
rect 24225 21505 24259 21539
rect 24259 21505 24268 21539
rect 24216 21496 24268 21505
rect 14188 21471 14240 21480
rect 14188 21437 14197 21471
rect 14197 21437 14231 21471
rect 14231 21437 14240 21471
rect 14188 21428 14240 21437
rect 16488 21428 16540 21480
rect 16672 21471 16724 21480
rect 16672 21437 16681 21471
rect 16681 21437 16715 21471
rect 16715 21437 16724 21471
rect 16672 21428 16724 21437
rect 18696 21428 18748 21480
rect 20352 21428 20404 21480
rect 20720 21428 20772 21480
rect 8300 21360 8352 21412
rect 11060 21360 11112 21412
rect 11888 21360 11940 21412
rect 13176 21360 13228 21412
rect 13544 21360 13596 21412
rect 15568 21360 15620 21412
rect 16580 21360 16632 21412
rect 23756 21428 23808 21480
rect 24676 21471 24728 21480
rect 24676 21437 24685 21471
rect 24685 21437 24719 21471
rect 24719 21437 24728 21471
rect 24676 21428 24728 21437
rect 22560 21360 22612 21412
rect 22744 21360 22796 21412
rect 23204 21403 23256 21412
rect 23204 21369 23213 21403
rect 23213 21369 23247 21403
rect 23247 21369 23256 21403
rect 23204 21360 23256 21369
rect 9128 21292 9180 21344
rect 9772 21292 9824 21344
rect 11980 21292 12032 21344
rect 12256 21335 12308 21344
rect 12256 21301 12265 21335
rect 12265 21301 12299 21335
rect 12299 21301 12308 21335
rect 12256 21292 12308 21301
rect 14740 21292 14792 21344
rect 15660 21335 15712 21344
rect 15660 21301 15669 21335
rect 15669 21301 15703 21335
rect 15703 21301 15712 21335
rect 15660 21292 15712 21301
rect 16120 21335 16172 21344
rect 16120 21301 16129 21335
rect 16129 21301 16163 21335
rect 16163 21301 16172 21335
rect 16120 21292 16172 21301
rect 19064 21292 19116 21344
rect 20076 21292 20128 21344
rect 20812 21335 20864 21344
rect 20812 21301 20821 21335
rect 20821 21301 20855 21335
rect 20855 21301 20864 21335
rect 20812 21292 20864 21301
rect 21180 21335 21232 21344
rect 21180 21301 21189 21335
rect 21189 21301 21223 21335
rect 21223 21301 21232 21335
rect 21180 21292 21232 21301
rect 22008 21292 22060 21344
rect 23020 21292 23072 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 7380 21131 7432 21140
rect 7380 21097 7389 21131
rect 7389 21097 7423 21131
rect 7423 21097 7432 21131
rect 7380 21088 7432 21097
rect 7840 21088 7892 21140
rect 9128 21131 9180 21140
rect 8392 21063 8444 21072
rect 8392 21029 8401 21063
rect 8401 21029 8435 21063
rect 8435 21029 8444 21063
rect 8392 21020 8444 21029
rect 8484 21020 8536 21072
rect 9128 21097 9137 21131
rect 9137 21097 9171 21131
rect 9171 21097 9180 21131
rect 9128 21088 9180 21097
rect 11152 21088 11204 21140
rect 11520 21088 11572 21140
rect 11796 21088 11848 21140
rect 12256 21088 12308 21140
rect 13544 21088 13596 21140
rect 14096 21131 14148 21140
rect 14096 21097 14105 21131
rect 14105 21097 14139 21131
rect 14139 21097 14148 21131
rect 14096 21088 14148 21097
rect 16396 21088 16448 21140
rect 17592 21131 17644 21140
rect 17592 21097 17601 21131
rect 17601 21097 17635 21131
rect 17635 21097 17644 21131
rect 17592 21088 17644 21097
rect 19340 21088 19392 21140
rect 20812 21088 20864 21140
rect 22008 21131 22060 21140
rect 11336 21020 11388 21072
rect 12072 21020 12124 21072
rect 15476 21020 15528 21072
rect 16764 21020 16816 21072
rect 17776 21020 17828 21072
rect 17868 21020 17920 21072
rect 18144 21063 18196 21072
rect 18144 21029 18153 21063
rect 18153 21029 18187 21063
rect 18187 21029 18196 21063
rect 18144 21020 18196 21029
rect 19432 21020 19484 21072
rect 19524 21020 19576 21072
rect 22008 21097 22017 21131
rect 22017 21097 22051 21131
rect 22051 21097 22060 21131
rect 22008 21088 22060 21097
rect 22192 21088 22244 21140
rect 15844 20952 15896 21004
rect 20168 20952 20220 21004
rect 20812 20952 20864 21004
rect 22560 21088 22612 21140
rect 23020 21088 23072 21140
rect 22928 21020 22980 21072
rect 23848 21020 23900 21072
rect 22468 20952 22520 21004
rect 9864 20884 9916 20936
rect 11704 20927 11756 20936
rect 11704 20893 11713 20927
rect 11713 20893 11747 20927
rect 11747 20893 11756 20927
rect 11704 20884 11756 20893
rect 13820 20884 13872 20936
rect 15292 20927 15344 20936
rect 15292 20893 15301 20927
rect 15301 20893 15335 20927
rect 15335 20893 15344 20927
rect 15292 20884 15344 20893
rect 18328 20884 18380 20936
rect 20720 20884 20772 20936
rect 21916 20884 21968 20936
rect 22008 20816 22060 20868
rect 8116 20791 8168 20800
rect 8116 20757 8125 20791
rect 8125 20757 8159 20791
rect 8159 20757 8168 20791
rect 8116 20748 8168 20757
rect 13544 20748 13596 20800
rect 16580 20748 16632 20800
rect 17960 20748 18012 20800
rect 19984 20748 20036 20800
rect 21456 20748 21508 20800
rect 22192 20748 22244 20800
rect 24860 20884 24912 20936
rect 22744 20748 22796 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 8208 20544 8260 20596
rect 12072 20587 12124 20596
rect 12072 20553 12081 20587
rect 12081 20553 12115 20587
rect 12115 20553 12124 20587
rect 12072 20544 12124 20553
rect 17868 20544 17920 20596
rect 20628 20544 20680 20596
rect 15476 20519 15528 20528
rect 15476 20485 15485 20519
rect 15485 20485 15519 20519
rect 15519 20485 15528 20519
rect 15476 20476 15528 20485
rect 25504 20519 25556 20528
rect 25504 20485 25513 20519
rect 25513 20485 25547 20519
rect 25547 20485 25556 20519
rect 25504 20476 25556 20485
rect 8760 20451 8812 20460
rect 8760 20417 8769 20451
rect 8769 20417 8803 20451
rect 8803 20417 8812 20451
rect 8760 20408 8812 20417
rect 20812 20408 20864 20460
rect 11704 20340 11756 20392
rect 12992 20340 13044 20392
rect 9128 20272 9180 20324
rect 13544 20272 13596 20324
rect 8484 20247 8536 20256
rect 8484 20213 8493 20247
rect 8493 20213 8527 20247
rect 8527 20213 8536 20247
rect 8484 20204 8536 20213
rect 10140 20247 10192 20256
rect 10140 20213 10149 20247
rect 10149 20213 10183 20247
rect 10183 20213 10192 20247
rect 10140 20204 10192 20213
rect 10692 20204 10744 20256
rect 11704 20247 11756 20256
rect 11704 20213 11713 20247
rect 11713 20213 11747 20247
rect 11747 20213 11756 20247
rect 11704 20204 11756 20213
rect 15844 20340 15896 20392
rect 17500 20340 17552 20392
rect 19524 20340 19576 20392
rect 20996 20340 21048 20392
rect 22744 20340 22796 20392
rect 23940 20383 23992 20392
rect 23940 20349 23949 20383
rect 23949 20349 23983 20383
rect 23983 20349 23992 20383
rect 23940 20340 23992 20349
rect 15752 20315 15804 20324
rect 15752 20281 15761 20315
rect 15761 20281 15795 20315
rect 15795 20281 15804 20315
rect 15752 20272 15804 20281
rect 15936 20315 15988 20324
rect 15936 20281 15945 20315
rect 15945 20281 15979 20315
rect 15979 20281 15988 20315
rect 15936 20272 15988 20281
rect 18328 20315 18380 20324
rect 18328 20281 18362 20315
rect 18362 20281 18380 20315
rect 18328 20272 18380 20281
rect 21180 20272 21232 20324
rect 15292 20247 15344 20256
rect 15292 20213 15301 20247
rect 15301 20213 15335 20247
rect 15335 20213 15344 20247
rect 15292 20204 15344 20213
rect 16304 20204 16356 20256
rect 16948 20247 17000 20256
rect 16948 20213 16957 20247
rect 16957 20213 16991 20247
rect 16991 20213 17000 20247
rect 16948 20204 17000 20213
rect 19432 20247 19484 20256
rect 19432 20213 19441 20247
rect 19441 20213 19475 20247
rect 19475 20213 19484 20247
rect 19432 20204 19484 20213
rect 22468 20247 22520 20256
rect 22468 20213 22477 20247
rect 22477 20213 22511 20247
rect 22511 20213 22520 20247
rect 22468 20204 22520 20213
rect 23388 20247 23440 20256
rect 23388 20213 23397 20247
rect 23397 20213 23431 20247
rect 23431 20213 23440 20247
rect 23388 20204 23440 20213
rect 24124 20204 24176 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 8760 20043 8812 20052
rect 8760 20009 8769 20043
rect 8769 20009 8803 20043
rect 8803 20009 8812 20043
rect 8760 20000 8812 20009
rect 12072 20000 12124 20052
rect 13360 20000 13412 20052
rect 13728 20000 13780 20052
rect 15844 20043 15896 20052
rect 15844 20009 15853 20043
rect 15853 20009 15887 20043
rect 15887 20009 15896 20043
rect 15844 20000 15896 20009
rect 19340 20043 19392 20052
rect 19340 20009 19349 20043
rect 19349 20009 19383 20043
rect 19383 20009 19392 20043
rect 19340 20000 19392 20009
rect 21364 20000 21416 20052
rect 22100 20000 22152 20052
rect 22744 20000 22796 20052
rect 23480 20000 23532 20052
rect 15752 19932 15804 19984
rect 16948 19932 17000 19984
rect 19248 19932 19300 19984
rect 20536 19932 20588 19984
rect 8760 19864 8812 19916
rect 10600 19864 10652 19916
rect 10784 19907 10836 19916
rect 10784 19873 10818 19907
rect 10818 19873 10836 19907
rect 10784 19864 10836 19873
rect 12348 19864 12400 19916
rect 13728 19864 13780 19916
rect 16580 19907 16632 19916
rect 16580 19873 16614 19907
rect 16614 19873 16632 19907
rect 16580 19864 16632 19873
rect 21180 19864 21232 19916
rect 22560 19932 22612 19984
rect 22928 19932 22980 19984
rect 24860 19975 24912 19984
rect 24860 19941 24869 19975
rect 24869 19941 24903 19975
rect 24903 19941 24912 19975
rect 24860 19932 24912 19941
rect 22468 19864 22520 19916
rect 23388 19907 23440 19916
rect 23388 19873 23397 19907
rect 23397 19873 23431 19907
rect 23431 19873 23440 19907
rect 23388 19864 23440 19873
rect 24124 19864 24176 19916
rect 13544 19796 13596 19848
rect 15660 19796 15712 19848
rect 16304 19839 16356 19848
rect 16304 19805 16313 19839
rect 16313 19805 16347 19839
rect 16347 19805 16356 19839
rect 16304 19796 16356 19805
rect 18328 19839 18380 19848
rect 18328 19805 18337 19839
rect 18337 19805 18371 19839
rect 18371 19805 18380 19839
rect 18328 19796 18380 19805
rect 19064 19796 19116 19848
rect 23296 19839 23348 19848
rect 23296 19805 23305 19839
rect 23305 19805 23339 19839
rect 23339 19805 23348 19839
rect 23296 19796 23348 19805
rect 24768 19839 24820 19848
rect 24768 19805 24777 19839
rect 24777 19805 24811 19839
rect 24811 19805 24820 19839
rect 24768 19796 24820 19805
rect 13084 19771 13136 19780
rect 13084 19737 13093 19771
rect 13093 19737 13127 19771
rect 13127 19737 13136 19771
rect 13084 19728 13136 19737
rect 18880 19771 18932 19780
rect 18880 19737 18889 19771
rect 18889 19737 18923 19771
rect 18923 19737 18932 19771
rect 18880 19728 18932 19737
rect 22928 19728 22980 19780
rect 24676 19728 24728 19780
rect 8208 19660 8260 19712
rect 12532 19703 12584 19712
rect 12532 19669 12541 19703
rect 12541 19669 12575 19703
rect 12575 19669 12584 19703
rect 12532 19660 12584 19669
rect 14096 19703 14148 19712
rect 14096 19669 14105 19703
rect 14105 19669 14139 19703
rect 14139 19669 14148 19703
rect 14096 19660 14148 19669
rect 19800 19703 19852 19712
rect 19800 19669 19809 19703
rect 19809 19669 19843 19703
rect 19843 19669 19852 19703
rect 19800 19660 19852 19669
rect 21180 19660 21232 19712
rect 22376 19660 22428 19712
rect 23848 19703 23900 19712
rect 23848 19669 23857 19703
rect 23857 19669 23891 19703
rect 23891 19669 23900 19703
rect 23848 19660 23900 19669
rect 24124 19703 24176 19712
rect 24124 19669 24133 19703
rect 24133 19669 24167 19703
rect 24167 19669 24176 19703
rect 24124 19660 24176 19669
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 8760 19456 8812 19508
rect 12808 19456 12860 19508
rect 13360 19456 13412 19508
rect 19340 19456 19392 19508
rect 20260 19456 20312 19508
rect 21456 19499 21508 19508
rect 21456 19465 21465 19499
rect 21465 19465 21499 19499
rect 21499 19465 21508 19499
rect 21456 19456 21508 19465
rect 23296 19456 23348 19508
rect 24124 19456 24176 19508
rect 13176 19388 13228 19440
rect 23940 19431 23992 19440
rect 23940 19397 23949 19431
rect 23949 19397 23983 19431
rect 23983 19397 23992 19431
rect 23940 19388 23992 19397
rect 13268 19320 13320 19372
rect 18880 19320 18932 19372
rect 8392 19227 8444 19236
rect 8392 19193 8401 19227
rect 8401 19193 8435 19227
rect 8435 19193 8444 19227
rect 8392 19184 8444 19193
rect 9680 19252 9732 19304
rect 10140 19252 10192 19304
rect 12348 19252 12400 19304
rect 12532 19252 12584 19304
rect 12716 19295 12768 19304
rect 12716 19261 12725 19295
rect 12725 19261 12759 19295
rect 12759 19261 12768 19295
rect 12716 19252 12768 19261
rect 14096 19295 14148 19304
rect 14096 19261 14130 19295
rect 14130 19261 14148 19295
rect 14096 19252 14148 19261
rect 8116 19159 8168 19168
rect 8116 19125 8149 19159
rect 8149 19125 8168 19159
rect 8576 19159 8628 19168
rect 8116 19116 8168 19125
rect 8576 19125 8585 19159
rect 8585 19125 8619 19159
rect 8619 19125 8628 19159
rect 8576 19116 8628 19125
rect 9680 19116 9732 19168
rect 10784 19116 10836 19168
rect 12992 19116 13044 19168
rect 13360 19116 13412 19168
rect 15292 19184 15344 19236
rect 15752 19227 15804 19236
rect 15752 19193 15761 19227
rect 15761 19193 15795 19227
rect 15795 19193 15804 19227
rect 15752 19184 15804 19193
rect 14280 19116 14332 19168
rect 15844 19116 15896 19168
rect 16212 19116 16264 19168
rect 16672 19227 16724 19236
rect 16672 19193 16681 19227
rect 16681 19193 16715 19227
rect 16715 19193 16724 19227
rect 17960 19252 18012 19304
rect 19800 19320 19852 19372
rect 20536 19320 20588 19372
rect 20996 19320 21048 19372
rect 19340 19252 19392 19304
rect 20168 19252 20220 19304
rect 21732 19295 21784 19304
rect 21732 19261 21741 19295
rect 21741 19261 21775 19295
rect 21775 19261 21784 19295
rect 21732 19252 21784 19261
rect 16672 19184 16724 19193
rect 17776 19116 17828 19168
rect 17960 19116 18012 19168
rect 18880 19184 18932 19236
rect 19984 19227 20036 19236
rect 19984 19193 19993 19227
rect 19993 19193 20027 19227
rect 20027 19193 20036 19227
rect 19984 19184 20036 19193
rect 20352 19184 20404 19236
rect 22008 19227 22060 19236
rect 22008 19193 22017 19227
rect 22017 19193 22051 19227
rect 22051 19193 22060 19227
rect 22008 19184 22060 19193
rect 22468 19184 22520 19236
rect 23848 19184 23900 19236
rect 24492 19184 24544 19236
rect 24860 19184 24912 19236
rect 19432 19116 19484 19168
rect 20168 19159 20220 19168
rect 20168 19125 20177 19159
rect 20177 19125 20211 19159
rect 20211 19125 20220 19159
rect 20168 19116 20220 19125
rect 21364 19116 21416 19168
rect 21916 19159 21968 19168
rect 21916 19125 21925 19159
rect 21925 19125 21959 19159
rect 21959 19125 21968 19159
rect 21916 19116 21968 19125
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 8300 18912 8352 18964
rect 10692 18955 10744 18964
rect 10692 18921 10701 18955
rect 10701 18921 10735 18955
rect 10735 18921 10744 18955
rect 10692 18912 10744 18921
rect 13544 18955 13596 18964
rect 13544 18921 13553 18955
rect 13553 18921 13587 18955
rect 13587 18921 13596 18955
rect 13544 18912 13596 18921
rect 14464 18912 14516 18964
rect 16212 18912 16264 18964
rect 16580 18912 16632 18964
rect 19064 18955 19116 18964
rect 19064 18921 19073 18955
rect 19073 18921 19107 18955
rect 19107 18921 19116 18955
rect 19064 18912 19116 18921
rect 21180 18955 21232 18964
rect 21180 18921 21189 18955
rect 21189 18921 21223 18955
rect 21223 18921 21232 18955
rect 21180 18912 21232 18921
rect 22008 18912 22060 18964
rect 22928 18955 22980 18964
rect 22928 18921 22937 18955
rect 22937 18921 22971 18955
rect 22971 18921 22980 18955
rect 22928 18912 22980 18921
rect 23480 18912 23532 18964
rect 10140 18844 10192 18896
rect 12164 18844 12216 18896
rect 14096 18844 14148 18896
rect 10600 18708 10652 18760
rect 8576 18640 8628 18692
rect 10784 18572 10836 18624
rect 12624 18751 12676 18760
rect 12624 18717 12633 18751
rect 12633 18717 12667 18751
rect 12667 18717 12676 18751
rect 12624 18708 12676 18717
rect 14280 18751 14332 18760
rect 14280 18717 14289 18751
rect 14289 18717 14323 18751
rect 14323 18717 14332 18751
rect 14280 18708 14332 18717
rect 12440 18572 12492 18624
rect 13360 18572 13412 18624
rect 13728 18615 13780 18624
rect 13728 18581 13737 18615
rect 13737 18581 13771 18615
rect 13771 18581 13780 18615
rect 13728 18572 13780 18581
rect 14832 18572 14884 18624
rect 21732 18844 21784 18896
rect 22376 18887 22428 18896
rect 22376 18853 22385 18887
rect 22385 18853 22419 18887
rect 22419 18853 22428 18887
rect 22376 18844 22428 18853
rect 24492 18887 24544 18896
rect 24492 18853 24501 18887
rect 24501 18853 24535 18887
rect 24535 18853 24544 18887
rect 24492 18844 24544 18853
rect 24952 18844 25004 18896
rect 15660 18819 15712 18828
rect 15660 18785 15669 18819
rect 15669 18785 15703 18819
rect 15703 18785 15712 18819
rect 15660 18776 15712 18785
rect 16764 18776 16816 18828
rect 22192 18819 22244 18828
rect 22192 18785 22201 18819
rect 22201 18785 22235 18819
rect 22235 18785 22244 18819
rect 22192 18776 22244 18785
rect 24216 18819 24268 18828
rect 24216 18785 24225 18819
rect 24225 18785 24259 18819
rect 24259 18785 24268 18819
rect 24216 18776 24268 18785
rect 15936 18751 15988 18760
rect 15936 18717 15945 18751
rect 15945 18717 15979 18751
rect 15979 18717 15988 18751
rect 15936 18708 15988 18717
rect 16304 18708 16356 18760
rect 17132 18751 17184 18760
rect 17132 18717 17141 18751
rect 17141 18717 17175 18751
rect 17175 18717 17184 18751
rect 17132 18708 17184 18717
rect 20628 18708 20680 18760
rect 22468 18751 22520 18760
rect 22468 18717 22477 18751
rect 22477 18717 22511 18751
rect 22511 18717 22520 18751
rect 22468 18708 22520 18717
rect 24584 18708 24636 18760
rect 25044 18708 25096 18760
rect 19340 18640 19392 18692
rect 20168 18640 20220 18692
rect 22100 18640 22152 18692
rect 24768 18640 24820 18692
rect 15384 18615 15436 18624
rect 15384 18581 15393 18615
rect 15393 18581 15427 18615
rect 15427 18581 15436 18615
rect 15384 18572 15436 18581
rect 18512 18615 18564 18624
rect 18512 18581 18521 18615
rect 18521 18581 18555 18615
rect 18555 18581 18564 18615
rect 18512 18572 18564 18581
rect 20352 18572 20404 18624
rect 21180 18572 21232 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 8392 18368 8444 18420
rect 10600 18411 10652 18420
rect 10600 18377 10609 18411
rect 10609 18377 10643 18411
rect 10643 18377 10652 18411
rect 10600 18368 10652 18377
rect 12716 18368 12768 18420
rect 14096 18368 14148 18420
rect 15660 18368 15712 18420
rect 19984 18368 20036 18420
rect 24216 18368 24268 18420
rect 24860 18368 24912 18420
rect 19524 18343 19576 18352
rect 19524 18309 19533 18343
rect 19533 18309 19567 18343
rect 19567 18309 19576 18343
rect 23480 18343 23532 18352
rect 19524 18300 19576 18309
rect 9496 18232 9548 18284
rect 10140 18275 10192 18284
rect 10140 18241 10149 18275
rect 10149 18241 10183 18275
rect 10183 18241 10192 18275
rect 10140 18232 10192 18241
rect 11520 18232 11572 18284
rect 12440 18275 12492 18284
rect 12440 18241 12449 18275
rect 12449 18241 12483 18275
rect 12483 18241 12492 18275
rect 12440 18232 12492 18241
rect 23480 18309 23489 18343
rect 23489 18309 23523 18343
rect 23523 18309 23532 18343
rect 23480 18300 23532 18309
rect 22836 18232 22888 18284
rect 24952 18275 25004 18284
rect 24952 18241 24961 18275
rect 24961 18241 24995 18275
rect 24995 18241 25004 18275
rect 25320 18275 25372 18284
rect 24952 18232 25004 18241
rect 25320 18241 25329 18275
rect 25329 18241 25363 18275
rect 25363 18241 25372 18275
rect 25320 18232 25372 18241
rect 9864 18207 9916 18216
rect 9864 18173 9873 18207
rect 9873 18173 9907 18207
rect 9907 18173 9916 18207
rect 9864 18164 9916 18173
rect 12164 18207 12216 18216
rect 12164 18173 12173 18207
rect 12173 18173 12207 18207
rect 12207 18173 12216 18207
rect 12164 18164 12216 18173
rect 16304 18164 16356 18216
rect 22100 18207 22152 18216
rect 22100 18173 22109 18207
rect 22109 18173 22143 18207
rect 22143 18173 22152 18207
rect 22100 18164 22152 18173
rect 24032 18164 24084 18216
rect 24676 18207 24728 18216
rect 24676 18173 24685 18207
rect 24685 18173 24719 18207
rect 24719 18173 24728 18207
rect 24676 18164 24728 18173
rect 12716 18139 12768 18148
rect 12716 18105 12750 18139
rect 12750 18105 12768 18139
rect 12716 18096 12768 18105
rect 9312 18071 9364 18080
rect 9312 18037 9321 18071
rect 9321 18037 9355 18071
rect 9355 18037 9364 18071
rect 9312 18028 9364 18037
rect 10692 18028 10744 18080
rect 11336 18071 11388 18080
rect 11336 18037 11345 18071
rect 11345 18037 11379 18071
rect 11379 18037 11388 18071
rect 11336 18028 11388 18037
rect 14280 18028 14332 18080
rect 15936 18096 15988 18148
rect 18144 18096 18196 18148
rect 18604 18139 18656 18148
rect 18604 18105 18613 18139
rect 18613 18105 18647 18139
rect 18647 18105 18656 18139
rect 18604 18096 18656 18105
rect 19524 18096 19576 18148
rect 23480 18096 23532 18148
rect 24768 18096 24820 18148
rect 16764 18028 16816 18080
rect 17132 18028 17184 18080
rect 17500 18071 17552 18080
rect 17500 18037 17509 18071
rect 17509 18037 17543 18071
rect 17543 18037 17552 18071
rect 17500 18028 17552 18037
rect 18328 18028 18380 18080
rect 21180 18028 21232 18080
rect 22468 18028 22520 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 9496 17867 9548 17876
rect 9496 17833 9505 17867
rect 9505 17833 9539 17867
rect 9539 17833 9548 17867
rect 9496 17824 9548 17833
rect 9772 17756 9824 17808
rect 11060 17756 11112 17808
rect 11520 17824 11572 17876
rect 14280 17824 14332 17876
rect 14464 17867 14516 17876
rect 14464 17833 14473 17867
rect 14473 17833 14507 17867
rect 14507 17833 14516 17867
rect 14464 17824 14516 17833
rect 15844 17867 15896 17876
rect 15844 17833 15853 17867
rect 15853 17833 15887 17867
rect 15887 17833 15896 17867
rect 15844 17824 15896 17833
rect 18144 17867 18196 17876
rect 18144 17833 18153 17867
rect 18153 17833 18187 17867
rect 18187 17833 18196 17867
rect 18144 17824 18196 17833
rect 19524 17824 19576 17876
rect 22376 17824 22428 17876
rect 23572 17824 23624 17876
rect 23848 17824 23900 17876
rect 25320 17867 25372 17876
rect 25320 17833 25329 17867
rect 25329 17833 25363 17867
rect 25363 17833 25372 17867
rect 25320 17824 25372 17833
rect 18512 17756 18564 17808
rect 10324 17663 10376 17672
rect 10324 17629 10333 17663
rect 10333 17629 10367 17663
rect 10367 17629 10376 17663
rect 10324 17620 10376 17629
rect 10416 17663 10468 17672
rect 10416 17629 10425 17663
rect 10425 17629 10459 17663
rect 10459 17629 10468 17663
rect 10416 17620 10468 17629
rect 10784 17620 10836 17672
rect 11152 17620 11204 17672
rect 14740 17688 14792 17740
rect 15384 17688 15436 17740
rect 21180 17731 21232 17740
rect 21180 17697 21214 17731
rect 21214 17697 21232 17731
rect 21180 17688 21232 17697
rect 24216 17731 24268 17740
rect 24216 17697 24250 17731
rect 24250 17697 24268 17731
rect 24216 17688 24268 17697
rect 15568 17620 15620 17672
rect 16764 17620 16816 17672
rect 18328 17663 18380 17672
rect 18328 17629 18337 17663
rect 18337 17629 18371 17663
rect 18371 17629 18380 17663
rect 18328 17620 18380 17629
rect 20904 17663 20956 17672
rect 20904 17629 20913 17663
rect 20913 17629 20947 17663
rect 20947 17629 20956 17663
rect 20904 17620 20956 17629
rect 23664 17620 23716 17672
rect 10968 17552 11020 17604
rect 16488 17552 16540 17604
rect 11704 17484 11756 17536
rect 12256 17484 12308 17536
rect 12716 17527 12768 17536
rect 12716 17493 12725 17527
rect 12725 17493 12759 17527
rect 12759 17493 12768 17527
rect 12716 17484 12768 17493
rect 13084 17484 13136 17536
rect 14832 17484 14884 17536
rect 17040 17484 17092 17536
rect 22284 17527 22336 17536
rect 22284 17493 22293 17527
rect 22293 17493 22327 17527
rect 22327 17493 22336 17527
rect 22284 17484 22336 17493
rect 22468 17484 22520 17536
rect 23756 17527 23808 17536
rect 23756 17493 23765 17527
rect 23765 17493 23799 17527
rect 23799 17493 23808 17527
rect 23756 17484 23808 17493
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 10416 17280 10468 17332
rect 11796 17280 11848 17332
rect 12256 17323 12308 17332
rect 12256 17289 12265 17323
rect 12265 17289 12299 17323
rect 12299 17289 12308 17323
rect 12256 17280 12308 17289
rect 12532 17323 12584 17332
rect 12532 17289 12541 17323
rect 12541 17289 12575 17323
rect 12575 17289 12584 17323
rect 12532 17280 12584 17289
rect 15568 17280 15620 17332
rect 15844 17280 15896 17332
rect 18512 17280 18564 17332
rect 19340 17280 19392 17332
rect 21732 17323 21784 17332
rect 14096 17255 14148 17264
rect 14096 17221 14105 17255
rect 14105 17221 14139 17255
rect 14139 17221 14148 17255
rect 14096 17212 14148 17221
rect 16488 17255 16540 17264
rect 16488 17221 16497 17255
rect 16497 17221 16531 17255
rect 16531 17221 16540 17255
rect 16488 17212 16540 17221
rect 18328 17255 18380 17264
rect 18328 17221 18337 17255
rect 18337 17221 18371 17255
rect 18371 17221 18380 17255
rect 18328 17212 18380 17221
rect 11336 17187 11388 17196
rect 11336 17153 11345 17187
rect 11345 17153 11379 17187
rect 11379 17153 11388 17187
rect 11336 17144 11388 17153
rect 13084 17187 13136 17196
rect 13084 17153 13093 17187
rect 13093 17153 13127 17187
rect 13127 17153 13136 17187
rect 13084 17144 13136 17153
rect 14464 17144 14516 17196
rect 14832 17144 14884 17196
rect 17040 17187 17092 17196
rect 17040 17153 17049 17187
rect 17049 17153 17083 17187
rect 17083 17153 17092 17187
rect 17040 17144 17092 17153
rect 19064 17187 19116 17196
rect 19064 17153 19073 17187
rect 19073 17153 19107 17187
rect 19107 17153 19116 17187
rect 19064 17144 19116 17153
rect 19524 17144 19576 17196
rect 11152 17076 11204 17128
rect 16764 17119 16816 17128
rect 10324 17008 10376 17060
rect 11244 17008 11296 17060
rect 11796 17008 11848 17060
rect 13820 17008 13872 17060
rect 14372 17008 14424 17060
rect 16764 17085 16773 17119
rect 16773 17085 16807 17119
rect 16807 17085 16816 17119
rect 16764 17076 16816 17085
rect 20628 17187 20680 17196
rect 20628 17153 20637 17187
rect 20637 17153 20671 17187
rect 20671 17153 20680 17187
rect 20628 17144 20680 17153
rect 21732 17289 21741 17323
rect 21741 17289 21775 17323
rect 21775 17289 21784 17323
rect 21732 17280 21784 17289
rect 22376 17280 22428 17332
rect 14832 17008 14884 17060
rect 19156 17008 19208 17060
rect 23664 17119 23716 17128
rect 23664 17085 23673 17119
rect 23673 17085 23707 17119
rect 23707 17085 23716 17119
rect 23664 17076 23716 17085
rect 22468 17051 22520 17060
rect 22468 17017 22477 17051
rect 22477 17017 22511 17051
rect 22511 17017 22520 17051
rect 22468 17008 22520 17017
rect 9772 16940 9824 16992
rect 10968 16940 11020 16992
rect 11520 16940 11572 16992
rect 12992 16983 13044 16992
rect 12992 16949 13001 16983
rect 13001 16949 13035 16983
rect 13035 16949 13044 16983
rect 12992 16940 13044 16949
rect 16948 16983 17000 16992
rect 16948 16949 16957 16983
rect 16957 16949 16991 16983
rect 16991 16949 17000 16983
rect 16948 16940 17000 16949
rect 20628 16983 20680 16992
rect 20628 16949 20637 16983
rect 20637 16949 20671 16983
rect 20671 16949 20680 16983
rect 20628 16940 20680 16949
rect 20904 16940 20956 16992
rect 21916 16940 21968 16992
rect 23756 17008 23808 17060
rect 23112 16940 23164 16992
rect 23296 16940 23348 16992
rect 23664 16940 23716 16992
rect 24676 16940 24728 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 10784 16736 10836 16788
rect 10968 16779 11020 16788
rect 10968 16745 10977 16779
rect 10977 16745 11011 16779
rect 11011 16745 11020 16779
rect 10968 16736 11020 16745
rect 10140 16668 10192 16720
rect 10508 16668 10560 16720
rect 11152 16668 11204 16720
rect 11612 16668 11664 16720
rect 11520 16600 11572 16652
rect 16488 16736 16540 16788
rect 16948 16736 17000 16788
rect 19064 16736 19116 16788
rect 21180 16779 21232 16788
rect 21180 16745 21189 16779
rect 21189 16745 21223 16779
rect 21223 16745 21232 16779
rect 21180 16736 21232 16745
rect 23664 16736 23716 16788
rect 24216 16736 24268 16788
rect 14004 16668 14056 16720
rect 14740 16711 14792 16720
rect 14740 16677 14749 16711
rect 14749 16677 14783 16711
rect 14783 16677 14792 16711
rect 14740 16668 14792 16677
rect 15844 16711 15896 16720
rect 15844 16677 15853 16711
rect 15853 16677 15887 16711
rect 15887 16677 15896 16711
rect 15844 16668 15896 16677
rect 16856 16668 16908 16720
rect 18512 16668 18564 16720
rect 19248 16668 19300 16720
rect 19524 16668 19576 16720
rect 22284 16668 22336 16720
rect 9588 16532 9640 16584
rect 10508 16575 10560 16584
rect 10508 16541 10517 16575
rect 10517 16541 10551 16575
rect 10551 16541 10560 16575
rect 10508 16532 10560 16541
rect 11060 16532 11112 16584
rect 13176 16532 13228 16584
rect 15384 16600 15436 16652
rect 16764 16600 16816 16652
rect 17040 16643 17092 16652
rect 17040 16609 17049 16643
rect 17049 16609 17083 16643
rect 17083 16609 17092 16643
rect 17040 16600 17092 16609
rect 21916 16600 21968 16652
rect 24768 16736 24820 16788
rect 24860 16668 24912 16720
rect 25412 16600 25464 16652
rect 15936 16575 15988 16584
rect 15936 16541 15945 16575
rect 15945 16541 15979 16575
rect 15979 16541 15988 16575
rect 15936 16532 15988 16541
rect 18604 16532 18656 16584
rect 19984 16532 20036 16584
rect 20444 16532 20496 16584
rect 25320 16532 25372 16584
rect 20628 16464 20680 16516
rect 13912 16396 13964 16448
rect 18972 16396 19024 16448
rect 20444 16439 20496 16448
rect 20444 16405 20453 16439
rect 20453 16405 20487 16439
rect 20487 16405 20496 16439
rect 20444 16396 20496 16405
rect 21272 16396 21324 16448
rect 23112 16396 23164 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 9588 16235 9640 16244
rect 9588 16201 9597 16235
rect 9597 16201 9631 16235
rect 9631 16201 9640 16235
rect 9588 16192 9640 16201
rect 10508 16192 10560 16244
rect 10968 16192 11020 16244
rect 12992 16192 13044 16244
rect 13176 16235 13228 16244
rect 13176 16201 13185 16235
rect 13185 16201 13219 16235
rect 13219 16201 13228 16235
rect 13176 16192 13228 16201
rect 11612 16056 11664 16108
rect 12440 16056 12492 16108
rect 14832 16192 14884 16244
rect 17500 16235 17552 16244
rect 17500 16201 17509 16235
rect 17509 16201 17543 16235
rect 17543 16201 17552 16235
rect 17500 16192 17552 16201
rect 18420 16235 18472 16244
rect 18420 16201 18429 16235
rect 18429 16201 18463 16235
rect 18463 16201 18472 16235
rect 18420 16192 18472 16201
rect 18604 16192 18656 16244
rect 22100 16192 22152 16244
rect 23296 16192 23348 16244
rect 23480 16235 23532 16244
rect 23480 16201 23489 16235
rect 23489 16201 23523 16235
rect 23523 16201 23532 16235
rect 23480 16192 23532 16201
rect 25412 16235 25464 16244
rect 25412 16201 25421 16235
rect 25421 16201 25455 16235
rect 25455 16201 25464 16235
rect 25412 16192 25464 16201
rect 15108 16124 15160 16176
rect 15844 16124 15896 16176
rect 19340 16124 19392 16176
rect 21548 16167 21600 16176
rect 21548 16133 21557 16167
rect 21557 16133 21591 16167
rect 21591 16133 21600 16167
rect 21548 16124 21600 16133
rect 21180 16056 21232 16108
rect 13912 16031 13964 16040
rect 13912 15997 13946 16031
rect 13946 15997 13964 16031
rect 11152 15963 11204 15972
rect 11152 15929 11161 15963
rect 11161 15929 11195 15963
rect 11195 15929 11204 15963
rect 11152 15920 11204 15929
rect 10692 15895 10744 15904
rect 10692 15861 10701 15895
rect 10701 15861 10735 15895
rect 10735 15861 10744 15895
rect 10692 15852 10744 15861
rect 11428 15852 11480 15904
rect 11520 15852 11572 15904
rect 13912 15988 13964 15997
rect 15936 15988 15988 16040
rect 18972 16031 19024 16040
rect 18972 15997 18981 16031
rect 18981 15997 19015 16031
rect 19015 15997 19024 16031
rect 18972 15988 19024 15997
rect 21272 15988 21324 16040
rect 16580 15920 16632 15972
rect 16948 15963 17000 15972
rect 16948 15929 16957 15963
rect 16957 15929 16991 15963
rect 16991 15929 17000 15963
rect 16948 15920 17000 15929
rect 14832 15852 14884 15904
rect 17684 15920 17736 15972
rect 18696 15963 18748 15972
rect 18696 15929 18705 15963
rect 18705 15929 18739 15963
rect 18739 15929 18748 15963
rect 18696 15920 18748 15929
rect 20352 15920 20404 15972
rect 20536 15963 20588 15972
rect 20536 15929 20545 15963
rect 20545 15929 20579 15963
rect 20579 15929 20588 15963
rect 20536 15920 20588 15929
rect 21824 15963 21876 15972
rect 21824 15929 21833 15963
rect 21833 15929 21867 15963
rect 21867 15929 21876 15963
rect 21824 15920 21876 15929
rect 23296 15988 23348 16040
rect 24032 16031 24084 16040
rect 24032 15997 24041 16031
rect 24041 15997 24075 16031
rect 24075 15997 24084 16031
rect 24032 15988 24084 15997
rect 24676 15988 24728 16040
rect 19432 15895 19484 15904
rect 19432 15861 19441 15895
rect 19441 15861 19475 15895
rect 19475 15861 19484 15895
rect 19432 15852 19484 15861
rect 20444 15895 20496 15904
rect 20444 15861 20453 15895
rect 20453 15861 20487 15895
rect 20487 15861 20496 15895
rect 20444 15852 20496 15861
rect 24676 15852 24728 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 10140 15648 10192 15700
rect 13820 15648 13872 15700
rect 15108 15691 15160 15700
rect 15108 15657 15117 15691
rect 15117 15657 15151 15691
rect 15151 15657 15160 15691
rect 15108 15648 15160 15657
rect 16580 15648 16632 15700
rect 17684 15648 17736 15700
rect 23388 15648 23440 15700
rect 24032 15691 24084 15700
rect 24032 15657 24041 15691
rect 24041 15657 24075 15691
rect 24075 15657 24084 15691
rect 24032 15648 24084 15657
rect 25412 15691 25464 15700
rect 12072 15580 12124 15632
rect 14188 15580 14240 15632
rect 14740 15580 14792 15632
rect 18144 15580 18196 15632
rect 18328 15580 18380 15632
rect 18880 15580 18932 15632
rect 20812 15580 20864 15632
rect 21548 15580 21600 15632
rect 21732 15580 21784 15632
rect 22836 15623 22888 15632
rect 22836 15589 22845 15623
rect 22845 15589 22879 15623
rect 22879 15589 22888 15623
rect 22836 15580 22888 15589
rect 25412 15657 25421 15691
rect 25421 15657 25455 15691
rect 25455 15657 25464 15691
rect 25412 15648 25464 15657
rect 24768 15580 24820 15632
rect 12164 15555 12216 15564
rect 12164 15521 12173 15555
rect 12173 15521 12207 15555
rect 12207 15521 12216 15555
rect 12164 15512 12216 15521
rect 12440 15555 12492 15564
rect 12440 15521 12449 15555
rect 12449 15521 12483 15555
rect 12483 15521 12492 15555
rect 15568 15555 15620 15564
rect 12440 15512 12492 15521
rect 15568 15521 15602 15555
rect 15602 15521 15620 15555
rect 15568 15512 15620 15521
rect 11428 15444 11480 15496
rect 13820 15487 13872 15496
rect 13820 15453 13829 15487
rect 13829 15453 13863 15487
rect 13863 15453 13872 15487
rect 13820 15444 13872 15453
rect 14188 15444 14240 15496
rect 14832 15444 14884 15496
rect 17776 15487 17828 15496
rect 17776 15453 17785 15487
rect 17785 15453 17819 15487
rect 17819 15453 17828 15487
rect 17776 15444 17828 15453
rect 20536 15444 20588 15496
rect 22008 15444 22060 15496
rect 23112 15487 23164 15496
rect 23112 15453 23121 15487
rect 23121 15453 23155 15487
rect 23155 15453 23164 15487
rect 23112 15444 23164 15453
rect 24860 15444 24912 15496
rect 10784 15419 10836 15428
rect 10784 15385 10793 15419
rect 10793 15385 10827 15419
rect 10827 15385 10836 15419
rect 10784 15376 10836 15385
rect 11060 15376 11112 15428
rect 13636 15376 13688 15428
rect 22192 15376 22244 15428
rect 13452 15351 13504 15360
rect 13452 15317 13461 15351
rect 13461 15317 13495 15351
rect 13495 15317 13504 15351
rect 13452 15308 13504 15317
rect 14096 15308 14148 15360
rect 15936 15308 15988 15360
rect 17040 15308 17092 15360
rect 18052 15308 18104 15360
rect 20352 15308 20404 15360
rect 20720 15308 20772 15360
rect 23940 15308 23992 15360
rect 24216 15308 24268 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 11612 15104 11664 15156
rect 12164 15104 12216 15156
rect 12808 15104 12860 15156
rect 13728 15104 13780 15156
rect 15384 15147 15436 15156
rect 15384 15113 15393 15147
rect 15393 15113 15427 15147
rect 15427 15113 15436 15147
rect 15384 15104 15436 15113
rect 15568 15104 15620 15156
rect 12716 15036 12768 15088
rect 12072 14968 12124 15020
rect 17684 15104 17736 15156
rect 18052 15104 18104 15156
rect 22836 15147 22888 15156
rect 22836 15113 22845 15147
rect 22845 15113 22879 15147
rect 22879 15113 22888 15147
rect 22836 15104 22888 15113
rect 24032 15104 24084 15156
rect 24768 15104 24820 15156
rect 25412 15104 25464 15156
rect 17132 15036 17184 15088
rect 18144 15036 18196 15088
rect 22560 15079 22612 15088
rect 22560 15045 22569 15079
rect 22569 15045 22603 15079
rect 22603 15045 22612 15079
rect 22560 15036 22612 15045
rect 23388 15036 23440 15088
rect 23756 15079 23808 15088
rect 23756 15045 23765 15079
rect 23765 15045 23799 15079
rect 23799 15045 23808 15079
rect 23756 15036 23808 15045
rect 19248 15011 19300 15020
rect 19248 14977 19257 15011
rect 19257 14977 19291 15011
rect 19291 14977 19300 15011
rect 19248 14968 19300 14977
rect 24216 15011 24268 15020
rect 12440 14900 12492 14952
rect 13360 14900 13412 14952
rect 13820 14900 13872 14952
rect 20260 14943 20312 14952
rect 14096 14875 14148 14884
rect 14096 14841 14105 14875
rect 14105 14841 14139 14875
rect 14139 14841 14148 14875
rect 14096 14832 14148 14841
rect 14188 14875 14240 14884
rect 14188 14841 14197 14875
rect 14197 14841 14231 14875
rect 14231 14841 14240 14875
rect 14188 14832 14240 14841
rect 15936 14832 15988 14884
rect 20260 14909 20269 14943
rect 20269 14909 20303 14943
rect 20303 14909 20312 14943
rect 20260 14900 20312 14909
rect 24216 14977 24225 15011
rect 24225 14977 24259 15011
rect 24259 14977 24268 15011
rect 24216 14968 24268 14977
rect 20536 14943 20588 14952
rect 20536 14909 20570 14943
rect 20570 14909 20588 14943
rect 20536 14900 20588 14909
rect 23940 14900 23992 14952
rect 18604 14875 18656 14884
rect 18604 14841 18613 14875
rect 18613 14841 18647 14875
rect 18647 14841 18656 14875
rect 18604 14832 18656 14841
rect 13268 14764 13320 14816
rect 14832 14807 14884 14816
rect 14832 14773 14841 14807
rect 14841 14773 14875 14807
rect 14875 14773 14884 14807
rect 14832 14764 14884 14773
rect 17776 14807 17828 14816
rect 17776 14773 17785 14807
rect 17785 14773 17819 14807
rect 17819 14773 17828 14807
rect 17776 14764 17828 14773
rect 19248 14807 19300 14816
rect 19248 14773 19257 14807
rect 19257 14773 19291 14807
rect 19291 14773 19300 14807
rect 19248 14764 19300 14773
rect 20260 14764 20312 14816
rect 20904 14764 20956 14816
rect 23480 14764 23532 14816
rect 24676 14807 24728 14816
rect 24676 14773 24685 14807
rect 24685 14773 24719 14807
rect 24719 14773 24728 14807
rect 24676 14764 24728 14773
rect 25228 14807 25280 14816
rect 25228 14773 25237 14807
rect 25237 14773 25271 14807
rect 25271 14773 25280 14807
rect 25228 14764 25280 14773
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 12716 14560 12768 14612
rect 13360 14560 13412 14612
rect 14280 14560 14332 14612
rect 15568 14560 15620 14612
rect 17132 14560 17184 14612
rect 19156 14560 19208 14612
rect 19248 14560 19300 14612
rect 20628 14560 20680 14612
rect 22100 14560 22152 14612
rect 23112 14560 23164 14612
rect 24216 14560 24268 14612
rect 14004 14535 14056 14544
rect 14004 14501 14013 14535
rect 14013 14501 14047 14535
rect 14047 14501 14056 14535
rect 14004 14492 14056 14501
rect 12164 14424 12216 14476
rect 13360 14424 13412 14476
rect 14372 14492 14424 14544
rect 15844 14535 15896 14544
rect 15844 14501 15853 14535
rect 15853 14501 15887 14535
rect 15887 14501 15896 14535
rect 15844 14492 15896 14501
rect 17500 14492 17552 14544
rect 18604 14492 18656 14544
rect 21180 14535 21232 14544
rect 21180 14501 21214 14535
rect 21214 14501 21232 14535
rect 21180 14492 21232 14501
rect 24032 14535 24084 14544
rect 24032 14501 24066 14535
rect 24066 14501 24084 14535
rect 24032 14492 24084 14501
rect 18972 14424 19024 14476
rect 20628 14424 20680 14476
rect 23848 14424 23900 14476
rect 11796 14356 11848 14408
rect 13452 14356 13504 14408
rect 14280 14399 14332 14408
rect 14280 14365 14289 14399
rect 14289 14365 14323 14399
rect 14323 14365 14332 14399
rect 14280 14356 14332 14365
rect 15752 14399 15804 14408
rect 15752 14365 15761 14399
rect 15761 14365 15795 14399
rect 15795 14365 15804 14399
rect 15752 14356 15804 14365
rect 17776 14399 17828 14408
rect 17776 14365 17785 14399
rect 17785 14365 17819 14399
rect 17819 14365 17828 14399
rect 17776 14356 17828 14365
rect 20904 14399 20956 14408
rect 20904 14365 20913 14399
rect 20913 14365 20947 14399
rect 20947 14365 20956 14399
rect 20904 14356 20956 14365
rect 13820 14288 13872 14340
rect 13268 14220 13320 14272
rect 14096 14220 14148 14272
rect 18144 14220 18196 14272
rect 23480 14220 23532 14272
rect 23940 14220 23992 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 11796 14059 11848 14068
rect 11796 14025 11805 14059
rect 11805 14025 11839 14059
rect 11839 14025 11848 14059
rect 11796 14016 11848 14025
rect 12164 14059 12216 14068
rect 12164 14025 12173 14059
rect 12173 14025 12207 14059
rect 12207 14025 12216 14059
rect 12164 14016 12216 14025
rect 12716 14059 12768 14068
rect 12716 14025 12725 14059
rect 12725 14025 12759 14059
rect 12759 14025 12768 14059
rect 12716 14016 12768 14025
rect 13360 14059 13412 14068
rect 13360 14025 13369 14059
rect 13369 14025 13403 14059
rect 13403 14025 13412 14059
rect 13360 14016 13412 14025
rect 14004 14016 14056 14068
rect 14188 14016 14240 14068
rect 15752 14059 15804 14068
rect 15752 14025 15761 14059
rect 15761 14025 15795 14059
rect 15795 14025 15804 14059
rect 15752 14016 15804 14025
rect 16488 14059 16540 14068
rect 16488 14025 16497 14059
rect 16497 14025 16531 14059
rect 16531 14025 16540 14059
rect 16488 14016 16540 14025
rect 17500 14059 17552 14068
rect 17500 14025 17509 14059
rect 17509 14025 17543 14059
rect 17543 14025 17552 14059
rect 17500 14016 17552 14025
rect 18420 14059 18472 14068
rect 18420 14025 18429 14059
rect 18429 14025 18463 14059
rect 18463 14025 18472 14059
rect 18420 14016 18472 14025
rect 18972 14059 19024 14068
rect 18972 14025 18981 14059
rect 18981 14025 19015 14059
rect 19015 14025 19024 14059
rect 18972 14016 19024 14025
rect 20168 14016 20220 14068
rect 20444 14016 20496 14068
rect 20904 14016 20956 14068
rect 21916 14016 21968 14068
rect 23112 14059 23164 14068
rect 23112 14025 23121 14059
rect 23121 14025 23155 14059
rect 23155 14025 23164 14059
rect 23112 14016 23164 14025
rect 24032 14016 24084 14068
rect 12808 13923 12860 13932
rect 12808 13889 12817 13923
rect 12817 13889 12851 13923
rect 12851 13889 12860 13923
rect 12808 13880 12860 13889
rect 16580 13880 16632 13932
rect 17224 13948 17276 14000
rect 19248 13948 19300 14000
rect 23204 13948 23256 14000
rect 17132 13880 17184 13932
rect 19432 13880 19484 13932
rect 21180 13880 21232 13932
rect 23572 13948 23624 14000
rect 23848 13880 23900 13932
rect 23940 13880 23992 13932
rect 13820 13855 13872 13864
rect 13820 13821 13829 13855
rect 13829 13821 13863 13855
rect 13863 13821 13872 13855
rect 13820 13812 13872 13821
rect 14280 13744 14332 13796
rect 20536 13812 20588 13864
rect 22284 13812 22336 13864
rect 18236 13744 18288 13796
rect 19340 13744 19392 13796
rect 20168 13744 20220 13796
rect 20996 13787 21048 13796
rect 20996 13753 21005 13787
rect 21005 13753 21039 13787
rect 21039 13753 21048 13787
rect 20996 13744 21048 13753
rect 22468 13744 22520 13796
rect 23756 13812 23808 13864
rect 24400 13855 24452 13864
rect 24400 13821 24423 13855
rect 24423 13821 24452 13855
rect 24400 13812 24452 13821
rect 17132 13676 17184 13728
rect 17776 13719 17828 13728
rect 17776 13685 17785 13719
rect 17785 13685 17819 13719
rect 17819 13685 17828 13719
rect 17776 13676 17828 13685
rect 22100 13676 22152 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 12164 13472 12216 13524
rect 12440 13472 12492 13524
rect 13820 13472 13872 13524
rect 14832 13472 14884 13524
rect 15844 13472 15896 13524
rect 16212 13472 16264 13524
rect 16488 13515 16540 13524
rect 16488 13481 16497 13515
rect 16497 13481 16531 13515
rect 16531 13481 16540 13515
rect 16488 13472 16540 13481
rect 17408 13472 17460 13524
rect 17684 13472 17736 13524
rect 17868 13472 17920 13524
rect 18420 13472 18472 13524
rect 19432 13515 19484 13524
rect 19432 13481 19441 13515
rect 19441 13481 19475 13515
rect 19475 13481 19484 13515
rect 19432 13472 19484 13481
rect 11152 13404 11204 13456
rect 12348 13404 12400 13456
rect 17316 13447 17368 13456
rect 17316 13413 17325 13447
rect 17325 13413 17359 13447
rect 17359 13413 17368 13447
rect 17316 13404 17368 13413
rect 18052 13404 18104 13456
rect 20444 13472 20496 13524
rect 20996 13472 21048 13524
rect 21180 13472 21232 13524
rect 21824 13472 21876 13524
rect 22100 13515 22152 13524
rect 22100 13481 22109 13515
rect 22109 13481 22143 13515
rect 22143 13481 22152 13515
rect 23112 13515 23164 13524
rect 22100 13472 22152 13481
rect 23112 13481 23121 13515
rect 23121 13481 23155 13515
rect 23155 13481 23164 13515
rect 23112 13472 23164 13481
rect 24400 13472 24452 13524
rect 19616 13404 19668 13456
rect 20076 13404 20128 13456
rect 22652 13404 22704 13456
rect 23848 13447 23900 13456
rect 23848 13413 23857 13447
rect 23857 13413 23891 13447
rect 23891 13413 23900 13447
rect 23848 13404 23900 13413
rect 25228 13404 25280 13456
rect 18696 13336 18748 13388
rect 23112 13336 23164 13388
rect 24124 13336 24176 13388
rect 24860 13336 24912 13388
rect 25688 13404 25740 13456
rect 11428 13311 11480 13320
rect 11428 13277 11437 13311
rect 11437 13277 11471 13311
rect 11471 13277 11480 13311
rect 11428 13268 11480 13277
rect 15752 13311 15804 13320
rect 15752 13277 15761 13311
rect 15761 13277 15795 13311
rect 15795 13277 15804 13311
rect 15752 13268 15804 13277
rect 17408 13311 17460 13320
rect 17408 13277 17417 13311
rect 17417 13277 17451 13311
rect 17451 13277 17460 13311
rect 17408 13268 17460 13277
rect 19064 13268 19116 13320
rect 21364 13311 21416 13320
rect 21364 13277 21373 13311
rect 21373 13277 21407 13311
rect 21407 13277 21416 13311
rect 21364 13268 21416 13277
rect 22284 13268 22336 13320
rect 22468 13311 22520 13320
rect 22468 13277 22477 13311
rect 22477 13277 22511 13311
rect 22511 13277 22520 13311
rect 22468 13268 22520 13277
rect 17776 13200 17828 13252
rect 23480 13200 23532 13252
rect 14280 13175 14332 13184
rect 14280 13141 14289 13175
rect 14289 13141 14323 13175
rect 14323 13141 14332 13175
rect 14280 13132 14332 13141
rect 15292 13132 15344 13184
rect 15568 13132 15620 13184
rect 19984 13132 20036 13184
rect 20168 13175 20220 13184
rect 20168 13141 20177 13175
rect 20177 13141 20211 13175
rect 20211 13141 20220 13175
rect 20168 13132 20220 13141
rect 21732 13132 21784 13184
rect 24216 13175 24268 13184
rect 24216 13141 24225 13175
rect 24225 13141 24259 13175
rect 24259 13141 24268 13175
rect 24216 13132 24268 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 11152 12971 11204 12980
rect 11152 12937 11161 12971
rect 11161 12937 11195 12971
rect 11195 12937 11204 12971
rect 11152 12928 11204 12937
rect 15292 12928 15344 12980
rect 17040 12971 17092 12980
rect 17040 12937 17049 12971
rect 17049 12937 17083 12971
rect 17083 12937 17092 12971
rect 17040 12928 17092 12937
rect 17408 12928 17460 12980
rect 17868 12928 17920 12980
rect 19064 12971 19116 12980
rect 19064 12937 19073 12971
rect 19073 12937 19107 12971
rect 19107 12937 19116 12971
rect 19064 12928 19116 12937
rect 20352 12928 20404 12980
rect 22652 12971 22704 12980
rect 12440 12860 12492 12912
rect 17684 12860 17736 12912
rect 18052 12860 18104 12912
rect 17408 12792 17460 12844
rect 20444 12860 20496 12912
rect 21180 12903 21232 12912
rect 21180 12869 21189 12903
rect 21189 12869 21223 12903
rect 21223 12869 21232 12903
rect 21180 12860 21232 12869
rect 20720 12792 20772 12844
rect 21364 12792 21416 12844
rect 22652 12937 22661 12971
rect 22661 12937 22695 12971
rect 22695 12937 22704 12971
rect 22652 12928 22704 12937
rect 24860 12971 24912 12980
rect 24860 12937 24869 12971
rect 24869 12937 24903 12971
rect 24903 12937 24912 12971
rect 24860 12928 24912 12937
rect 25688 12971 25740 12980
rect 25688 12937 25697 12971
rect 25697 12937 25731 12971
rect 25731 12937 25740 12971
rect 25688 12928 25740 12937
rect 23756 12903 23808 12912
rect 23756 12869 23765 12903
rect 23765 12869 23799 12903
rect 23799 12869 23808 12903
rect 23756 12860 23808 12869
rect 24216 12835 24268 12844
rect 24216 12801 24225 12835
rect 24225 12801 24259 12835
rect 24259 12801 24268 12835
rect 24216 12792 24268 12801
rect 11428 12724 11480 12776
rect 12440 12767 12492 12776
rect 12440 12733 12449 12767
rect 12449 12733 12483 12767
rect 12483 12733 12492 12767
rect 12440 12724 12492 12733
rect 12532 12656 12584 12708
rect 18420 12767 18472 12776
rect 18420 12733 18429 12767
rect 18429 12733 18463 12767
rect 18463 12733 18472 12767
rect 18420 12724 18472 12733
rect 18604 12724 18656 12776
rect 19984 12724 20036 12776
rect 20812 12724 20864 12776
rect 15384 12656 15436 12708
rect 18696 12699 18748 12708
rect 18696 12665 18705 12699
rect 18705 12665 18739 12699
rect 18739 12665 18748 12699
rect 18696 12656 18748 12665
rect 19340 12656 19392 12708
rect 20720 12699 20772 12708
rect 20720 12665 20729 12699
rect 20729 12665 20763 12699
rect 20763 12665 20772 12699
rect 20720 12656 20772 12665
rect 21088 12656 21140 12708
rect 21364 12656 21416 12708
rect 24308 12699 24360 12708
rect 24308 12665 24317 12699
rect 24317 12665 24351 12699
rect 24351 12665 24360 12699
rect 24308 12656 24360 12665
rect 12348 12588 12400 12640
rect 13912 12588 13964 12640
rect 14924 12631 14976 12640
rect 14924 12597 14933 12631
rect 14933 12597 14967 12631
rect 14967 12597 14976 12631
rect 14924 12588 14976 12597
rect 17684 12588 17736 12640
rect 20168 12588 20220 12640
rect 20536 12588 20588 12640
rect 22284 12588 22336 12640
rect 23112 12631 23164 12640
rect 23112 12597 23121 12631
rect 23121 12597 23155 12631
rect 23155 12597 23164 12631
rect 23112 12588 23164 12597
rect 25044 12588 25096 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 17408 12427 17460 12436
rect 17408 12393 17417 12427
rect 17417 12393 17451 12427
rect 17451 12393 17460 12427
rect 17408 12384 17460 12393
rect 17776 12427 17828 12436
rect 17776 12393 17785 12427
rect 17785 12393 17819 12427
rect 17819 12393 17828 12427
rect 17776 12384 17828 12393
rect 17868 12384 17920 12436
rect 20720 12384 20772 12436
rect 21180 12384 21232 12436
rect 23848 12427 23900 12436
rect 23848 12393 23857 12427
rect 23857 12393 23891 12427
rect 23891 12393 23900 12427
rect 23848 12384 23900 12393
rect 25228 12384 25280 12436
rect 12256 12359 12308 12368
rect 12256 12325 12265 12359
rect 12265 12325 12299 12359
rect 12299 12325 12308 12359
rect 12256 12316 12308 12325
rect 12348 12359 12400 12368
rect 12348 12325 12357 12359
rect 12357 12325 12391 12359
rect 12391 12325 12400 12359
rect 13820 12359 13872 12368
rect 12348 12316 12400 12325
rect 13820 12325 13829 12359
rect 13829 12325 13863 12359
rect 13863 12325 13872 12359
rect 13820 12316 13872 12325
rect 14188 12316 14240 12368
rect 14924 12316 14976 12368
rect 13912 12291 13964 12300
rect 13912 12257 13921 12291
rect 13921 12257 13955 12291
rect 13955 12257 13964 12291
rect 15936 12316 15988 12368
rect 18696 12316 18748 12368
rect 19432 12316 19484 12368
rect 20076 12316 20128 12368
rect 20996 12316 21048 12368
rect 21548 12316 21600 12368
rect 13912 12248 13964 12257
rect 17040 12248 17092 12300
rect 17132 12248 17184 12300
rect 17960 12248 18012 12300
rect 20720 12248 20772 12300
rect 21272 12291 21324 12300
rect 21272 12257 21281 12291
rect 21281 12257 21315 12291
rect 21315 12257 21324 12291
rect 21272 12248 21324 12257
rect 22744 12291 22796 12300
rect 22744 12257 22778 12291
rect 22778 12257 22796 12291
rect 22744 12248 22796 12257
rect 12164 12223 12216 12232
rect 12164 12189 12173 12223
rect 12173 12189 12207 12223
rect 12207 12189 12216 12223
rect 12164 12180 12216 12189
rect 13728 12223 13780 12232
rect 13728 12189 13737 12223
rect 13737 12189 13771 12223
rect 13771 12189 13780 12223
rect 13728 12180 13780 12189
rect 20260 12180 20312 12232
rect 20904 12180 20956 12232
rect 21548 12223 21600 12232
rect 21548 12189 21557 12223
rect 21557 12189 21591 12223
rect 21591 12189 21600 12223
rect 21548 12180 21600 12189
rect 13544 12112 13596 12164
rect 20812 12112 20864 12164
rect 11796 12087 11848 12096
rect 11796 12053 11805 12087
rect 11805 12053 11839 12087
rect 11839 12053 11848 12087
rect 11796 12044 11848 12053
rect 13360 12087 13412 12096
rect 13360 12053 13369 12087
rect 13369 12053 13403 12087
rect 13403 12053 13412 12087
rect 13360 12044 13412 12053
rect 13452 12044 13504 12096
rect 14740 12087 14792 12096
rect 14740 12053 14749 12087
rect 14749 12053 14783 12087
rect 14783 12053 14792 12087
rect 14740 12044 14792 12053
rect 15384 12044 15436 12096
rect 21180 12044 21232 12096
rect 21916 12044 21968 12096
rect 24308 12112 24360 12164
rect 23664 12044 23716 12096
rect 24860 12044 24912 12096
rect 25136 12087 25188 12096
rect 25136 12053 25145 12087
rect 25145 12053 25179 12087
rect 25179 12053 25188 12087
rect 25136 12044 25188 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 12072 11840 12124 11892
rect 12256 11840 12308 11892
rect 13820 11840 13872 11892
rect 13912 11840 13964 11892
rect 15752 11840 15804 11892
rect 12992 11815 13044 11824
rect 12992 11781 13001 11815
rect 13001 11781 13035 11815
rect 13035 11781 13044 11815
rect 12992 11772 13044 11781
rect 14832 11772 14884 11824
rect 11796 11704 11848 11756
rect 13452 11704 13504 11756
rect 13544 11747 13596 11756
rect 13544 11713 13553 11747
rect 13553 11713 13587 11747
rect 13587 11713 13596 11747
rect 13544 11704 13596 11713
rect 15384 11704 15436 11756
rect 14740 11636 14792 11688
rect 17592 11840 17644 11892
rect 17040 11747 17092 11756
rect 17040 11713 17049 11747
rect 17049 11713 17083 11747
rect 17083 11713 17092 11747
rect 17040 11704 17092 11713
rect 13176 11568 13228 11620
rect 13728 11568 13780 11620
rect 14924 11568 14976 11620
rect 15568 11568 15620 11620
rect 16028 11568 16080 11620
rect 20720 11840 20772 11892
rect 20996 11883 21048 11892
rect 20996 11849 21005 11883
rect 21005 11849 21039 11883
rect 21039 11849 21048 11883
rect 20996 11840 21048 11849
rect 22744 11840 22796 11892
rect 23572 11840 23624 11892
rect 24860 11840 24912 11892
rect 20628 11704 20680 11756
rect 20904 11636 20956 11688
rect 21916 11636 21968 11688
rect 23940 11679 23992 11688
rect 23940 11645 23949 11679
rect 23949 11645 23983 11679
rect 23983 11645 23992 11679
rect 23940 11636 23992 11645
rect 11520 11500 11572 11552
rect 13452 11543 13504 11552
rect 13452 11509 13461 11543
rect 13461 11509 13495 11543
rect 13495 11509 13504 11543
rect 13452 11500 13504 11509
rect 15936 11543 15988 11552
rect 15936 11509 15945 11543
rect 15945 11509 15979 11543
rect 15979 11509 15988 11543
rect 15936 11500 15988 11509
rect 17776 11543 17828 11552
rect 17776 11509 17785 11543
rect 17785 11509 17819 11543
rect 17819 11509 17828 11543
rect 17776 11500 17828 11509
rect 20352 11568 20404 11620
rect 20628 11568 20680 11620
rect 21180 11568 21232 11620
rect 22284 11568 22336 11620
rect 19432 11543 19484 11552
rect 19432 11509 19441 11543
rect 19441 11509 19475 11543
rect 19475 11509 19484 11543
rect 19432 11500 19484 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 11336 11228 11388 11280
rect 11796 11228 11848 11280
rect 11152 11160 11204 11212
rect 11520 11135 11572 11144
rect 11520 11101 11529 11135
rect 11529 11101 11563 11135
rect 11563 11101 11572 11135
rect 11520 11092 11572 11101
rect 13452 11296 13504 11348
rect 13544 11296 13596 11348
rect 14924 11339 14976 11348
rect 14924 11305 14933 11339
rect 14933 11305 14967 11339
rect 14967 11305 14976 11339
rect 14924 11296 14976 11305
rect 16028 11339 16080 11348
rect 16028 11305 16037 11339
rect 16037 11305 16071 11339
rect 16071 11305 16080 11339
rect 16028 11296 16080 11305
rect 16948 11296 17000 11348
rect 18880 11296 18932 11348
rect 22284 11339 22336 11348
rect 22284 11305 22293 11339
rect 22293 11305 22327 11339
rect 22327 11305 22336 11339
rect 22284 11296 22336 11305
rect 22744 11296 22796 11348
rect 12348 11160 12400 11212
rect 12440 11135 12492 11144
rect 12440 11101 12449 11135
rect 12449 11101 12483 11135
rect 12483 11101 12492 11135
rect 12440 11092 12492 11101
rect 15568 10956 15620 11008
rect 20812 11228 20864 11280
rect 21548 11228 21600 11280
rect 16580 11160 16632 11212
rect 16764 11024 16816 11076
rect 18788 11160 18840 11212
rect 19064 11160 19116 11212
rect 20904 11203 20956 11212
rect 20904 11169 20913 11203
rect 20913 11169 20947 11203
rect 20947 11169 20956 11203
rect 20904 11160 20956 11169
rect 23940 11203 23992 11212
rect 23940 11169 23949 11203
rect 23949 11169 23983 11203
rect 23983 11169 23992 11203
rect 23940 11160 23992 11169
rect 17316 11092 17368 11144
rect 17960 11092 18012 11144
rect 20720 11092 20772 11144
rect 17592 10999 17644 11008
rect 17592 10965 17601 10999
rect 17601 10965 17635 10999
rect 17635 10965 17644 10999
rect 17592 10956 17644 10965
rect 18052 10956 18104 11008
rect 21548 10956 21600 11008
rect 22744 11024 22796 11076
rect 24952 11024 25004 11076
rect 23664 10999 23716 11008
rect 23664 10965 23673 10999
rect 23673 10965 23707 10999
rect 23707 10965 23716 10999
rect 23664 10956 23716 10965
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 17960 10752 18012 10804
rect 18788 10752 18840 10804
rect 19892 10752 19944 10804
rect 20168 10752 20220 10804
rect 20536 10752 20588 10804
rect 22100 10752 22152 10804
rect 23664 10752 23716 10804
rect 23940 10752 23992 10804
rect 16580 10684 16632 10736
rect 18880 10684 18932 10736
rect 20812 10684 20864 10736
rect 21272 10727 21324 10736
rect 21272 10693 21281 10727
rect 21281 10693 21315 10727
rect 21315 10693 21324 10727
rect 21272 10684 21324 10693
rect 12440 10616 12492 10668
rect 17316 10616 17368 10668
rect 18052 10616 18104 10668
rect 19984 10616 20036 10668
rect 21364 10616 21416 10668
rect 24676 10684 24728 10736
rect 22008 10616 22060 10668
rect 24124 10659 24176 10668
rect 24124 10625 24133 10659
rect 24133 10625 24167 10659
rect 24167 10625 24176 10659
rect 24124 10616 24176 10625
rect 10600 10591 10652 10600
rect 10600 10557 10609 10591
rect 10609 10557 10643 10591
rect 10643 10557 10652 10591
rect 10600 10548 10652 10557
rect 13544 10591 13596 10600
rect 13544 10557 13578 10591
rect 13578 10557 13596 10591
rect 12440 10480 12492 10532
rect 13544 10548 13596 10557
rect 16028 10480 16080 10532
rect 16764 10523 16816 10532
rect 16764 10489 16773 10523
rect 16773 10489 16807 10523
rect 16807 10489 16816 10523
rect 16764 10480 16816 10489
rect 17592 10548 17644 10600
rect 23664 10548 23716 10600
rect 25228 10591 25280 10600
rect 25228 10557 25237 10591
rect 25237 10557 25271 10591
rect 25271 10557 25280 10591
rect 25228 10548 25280 10557
rect 19156 10480 19208 10532
rect 20904 10523 20956 10532
rect 20904 10489 20913 10523
rect 20913 10489 20947 10523
rect 20947 10489 20956 10523
rect 20904 10480 20956 10489
rect 22100 10523 22152 10532
rect 22100 10489 22109 10523
rect 22109 10489 22143 10523
rect 22143 10489 22152 10523
rect 22100 10480 22152 10489
rect 10968 10455 11020 10464
rect 10968 10421 10977 10455
rect 10977 10421 11011 10455
rect 11011 10421 11020 10455
rect 10968 10412 11020 10421
rect 12164 10455 12216 10464
rect 12164 10421 12173 10455
rect 12173 10421 12207 10455
rect 12207 10421 12216 10455
rect 12164 10412 12216 10421
rect 14740 10412 14792 10464
rect 15568 10455 15620 10464
rect 15568 10421 15577 10455
rect 15577 10421 15611 10455
rect 15611 10421 15620 10455
rect 15568 10412 15620 10421
rect 23664 10412 23716 10464
rect 24768 10412 24820 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 11520 10208 11572 10260
rect 12164 10208 12216 10260
rect 12992 10208 13044 10260
rect 13820 10208 13872 10260
rect 16488 10208 16540 10260
rect 17316 10251 17368 10260
rect 17316 10217 17325 10251
rect 17325 10217 17359 10251
rect 17359 10217 17368 10251
rect 17316 10208 17368 10217
rect 18236 10208 18288 10260
rect 19248 10208 19300 10260
rect 20444 10208 20496 10260
rect 13636 10140 13688 10192
rect 17776 10140 17828 10192
rect 20812 10140 20864 10192
rect 21548 10183 21600 10192
rect 21548 10149 21557 10183
rect 21557 10149 21591 10183
rect 21591 10149 21600 10183
rect 21548 10140 21600 10149
rect 16948 10072 17000 10124
rect 17960 10072 18012 10124
rect 22100 10208 22152 10260
rect 23296 10208 23348 10260
rect 23664 10183 23716 10192
rect 23664 10149 23673 10183
rect 23673 10149 23707 10183
rect 23707 10149 23716 10183
rect 23664 10140 23716 10149
rect 23756 10140 23808 10192
rect 24216 10140 24268 10192
rect 24676 10140 24728 10192
rect 22836 10115 22888 10124
rect 22836 10081 22845 10115
rect 22845 10081 22879 10115
rect 22879 10081 22888 10115
rect 22836 10072 22888 10081
rect 14740 10004 14792 10056
rect 13728 9936 13780 9988
rect 13084 9911 13136 9920
rect 13084 9877 13093 9911
rect 13093 9877 13127 9911
rect 13127 9877 13136 9911
rect 13084 9868 13136 9877
rect 20996 10004 21048 10056
rect 21732 10004 21784 10056
rect 23112 10047 23164 10056
rect 23112 10013 23121 10047
rect 23121 10013 23155 10047
rect 23155 10013 23164 10047
rect 23112 10004 23164 10013
rect 23940 10004 23992 10056
rect 24952 10004 25004 10056
rect 17592 9936 17644 9988
rect 16120 9868 16172 9920
rect 18052 9868 18104 9920
rect 19156 9868 19208 9920
rect 20812 9868 20864 9920
rect 22560 9911 22612 9920
rect 22560 9877 22569 9911
rect 22569 9877 22603 9911
rect 22603 9877 22612 9911
rect 22560 9868 22612 9877
rect 24124 9911 24176 9920
rect 24124 9877 24133 9911
rect 24133 9877 24167 9911
rect 24167 9877 24176 9911
rect 24124 9868 24176 9877
rect 25228 9911 25280 9920
rect 25228 9877 25237 9911
rect 25237 9877 25271 9911
rect 25271 9877 25280 9911
rect 25228 9868 25280 9877
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 16948 9664 17000 9716
rect 17316 9664 17368 9716
rect 12440 9596 12492 9648
rect 13728 9596 13780 9648
rect 13820 9596 13872 9648
rect 16028 9596 16080 9648
rect 13636 9528 13688 9580
rect 16764 9528 16816 9580
rect 17960 9664 18012 9716
rect 19156 9664 19208 9716
rect 17776 9639 17828 9648
rect 17776 9605 17785 9639
rect 17785 9605 17819 9639
rect 17819 9605 17828 9639
rect 17776 9596 17828 9605
rect 19340 9596 19392 9648
rect 20996 9664 21048 9716
rect 21548 9707 21600 9716
rect 21548 9673 21557 9707
rect 21557 9673 21591 9707
rect 21591 9673 21600 9707
rect 21548 9664 21600 9673
rect 20720 9596 20772 9648
rect 22836 9664 22888 9716
rect 23296 9664 23348 9716
rect 24216 9664 24268 9716
rect 22100 9639 22152 9648
rect 22100 9605 22109 9639
rect 22109 9605 22143 9639
rect 22143 9605 22152 9639
rect 22100 9596 22152 9605
rect 14740 9503 14792 9512
rect 14740 9469 14774 9503
rect 14774 9469 14792 9503
rect 13360 9392 13412 9444
rect 14740 9460 14792 9469
rect 18052 9503 18104 9512
rect 18052 9469 18061 9503
rect 18061 9469 18095 9503
rect 18095 9469 18104 9503
rect 18052 9460 18104 9469
rect 20444 9528 20496 9580
rect 22560 9571 22612 9580
rect 22560 9537 22569 9571
rect 22569 9537 22603 9571
rect 22603 9537 22612 9571
rect 22560 9528 22612 9537
rect 23940 9528 23992 9580
rect 24032 9503 24084 9512
rect 16028 9392 16080 9444
rect 24032 9469 24041 9503
rect 24041 9469 24075 9503
rect 24075 9469 24084 9503
rect 24032 9460 24084 9469
rect 25228 9503 25280 9512
rect 25228 9469 25237 9503
rect 25237 9469 25271 9503
rect 25271 9469 25280 9503
rect 25228 9460 25280 9469
rect 20996 9367 21048 9376
rect 20996 9333 21005 9367
rect 21005 9333 21039 9367
rect 21039 9333 21048 9367
rect 20996 9324 21048 9333
rect 21916 9324 21968 9376
rect 22652 9435 22704 9444
rect 22652 9401 22661 9435
rect 22661 9401 22695 9435
rect 22695 9401 22704 9435
rect 22652 9392 22704 9401
rect 23112 9392 23164 9444
rect 23480 9367 23532 9376
rect 23480 9333 23489 9367
rect 23489 9333 23523 9367
rect 23523 9333 23532 9367
rect 23480 9324 23532 9333
rect 25412 9367 25464 9376
rect 25412 9333 25421 9367
rect 25421 9333 25455 9367
rect 25455 9333 25464 9367
rect 25412 9324 25464 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 13360 9163 13412 9172
rect 13360 9129 13369 9163
rect 13369 9129 13403 9163
rect 13403 9129 13412 9163
rect 13360 9120 13412 9129
rect 13728 9163 13780 9172
rect 13728 9129 13737 9163
rect 13737 9129 13771 9163
rect 13771 9129 13780 9163
rect 13728 9120 13780 9129
rect 14740 9120 14792 9172
rect 16856 9163 16908 9172
rect 16856 9129 16865 9163
rect 16865 9129 16899 9163
rect 16899 9129 16908 9163
rect 16856 9120 16908 9129
rect 18052 9163 18104 9172
rect 18052 9129 18061 9163
rect 18061 9129 18095 9163
rect 18095 9129 18104 9163
rect 18052 9120 18104 9129
rect 20352 9163 20404 9172
rect 20352 9129 20361 9163
rect 20361 9129 20395 9163
rect 20395 9129 20404 9163
rect 20352 9120 20404 9129
rect 21916 9120 21968 9172
rect 22652 9120 22704 9172
rect 23756 9163 23808 9172
rect 23756 9129 23765 9163
rect 23765 9129 23799 9163
rect 23799 9129 23808 9163
rect 23756 9120 23808 9129
rect 24032 9120 24084 9172
rect 24676 9163 24728 9172
rect 24676 9129 24685 9163
rect 24685 9129 24719 9163
rect 24719 9129 24728 9163
rect 24676 9120 24728 9129
rect 25780 9120 25832 9172
rect 16580 9052 16632 9104
rect 16948 9095 17000 9104
rect 16948 9061 16957 9095
rect 16957 9061 16991 9095
rect 16991 9061 17000 9095
rect 16948 9052 17000 9061
rect 17960 9052 18012 9104
rect 18328 9052 18380 9104
rect 25228 9095 25280 9104
rect 25228 9061 25237 9095
rect 25237 9061 25271 9095
rect 25271 9061 25280 9095
rect 25228 9052 25280 9061
rect 21272 9027 21324 9036
rect 21272 8993 21281 9027
rect 21281 8993 21315 9027
rect 21315 8993 21324 9027
rect 21272 8984 21324 8993
rect 21732 8984 21784 9036
rect 22192 8984 22244 9036
rect 22468 8984 22520 9036
rect 23112 8984 23164 9036
rect 18052 8916 18104 8968
rect 25504 8959 25556 8968
rect 25504 8925 25513 8959
rect 25513 8925 25547 8959
rect 25547 8925 25556 8959
rect 25504 8916 25556 8925
rect 16396 8823 16448 8832
rect 16396 8789 16405 8823
rect 16405 8789 16439 8823
rect 16439 8789 16448 8823
rect 16396 8780 16448 8789
rect 19984 8780 20036 8832
rect 20352 8780 20404 8832
rect 20536 8780 20588 8832
rect 21180 8823 21232 8832
rect 21180 8789 21189 8823
rect 21189 8789 21223 8823
rect 21223 8789 21232 8823
rect 21180 8780 21232 8789
rect 21456 8823 21508 8832
rect 21456 8789 21465 8823
rect 21465 8789 21499 8823
rect 21499 8789 21508 8823
rect 21456 8780 21508 8789
rect 24860 8780 24912 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 15568 8576 15620 8628
rect 16580 8576 16632 8628
rect 18328 8576 18380 8628
rect 19524 8576 19576 8628
rect 22468 8619 22520 8628
rect 22468 8585 22477 8619
rect 22477 8585 22511 8619
rect 22511 8585 22520 8619
rect 22468 8576 22520 8585
rect 25228 8576 25280 8628
rect 16948 8508 17000 8560
rect 19340 8551 19392 8560
rect 19340 8517 19349 8551
rect 19349 8517 19383 8551
rect 19383 8517 19392 8551
rect 19340 8508 19392 8517
rect 16856 8440 16908 8492
rect 17040 8483 17092 8492
rect 17040 8449 17049 8483
rect 17049 8449 17083 8483
rect 17083 8449 17092 8483
rect 17040 8440 17092 8449
rect 18052 8440 18104 8492
rect 20536 8508 20588 8560
rect 22192 8508 22244 8560
rect 25780 8508 25832 8560
rect 16580 8372 16632 8424
rect 16304 8347 16356 8356
rect 16304 8313 16313 8347
rect 16313 8313 16347 8347
rect 16347 8313 16356 8347
rect 16764 8347 16816 8356
rect 16304 8304 16356 8313
rect 16764 8313 16773 8347
rect 16773 8313 16807 8347
rect 16807 8313 16816 8347
rect 16764 8304 16816 8313
rect 17224 8372 17276 8424
rect 19340 8372 19392 8424
rect 23664 8483 23716 8492
rect 23664 8449 23673 8483
rect 23673 8449 23707 8483
rect 23707 8449 23716 8483
rect 23664 8440 23716 8449
rect 20996 8372 21048 8424
rect 21732 8372 21784 8424
rect 23756 8372 23808 8424
rect 21180 8304 21232 8356
rect 25504 8304 25556 8356
rect 20628 8279 20680 8288
rect 20628 8245 20637 8279
rect 20637 8245 20671 8279
rect 20671 8245 20680 8279
rect 20628 8236 20680 8245
rect 20904 8279 20956 8288
rect 20904 8245 20913 8279
rect 20913 8245 20947 8279
rect 20947 8245 20956 8279
rect 20904 8236 20956 8245
rect 25136 8236 25188 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 16488 8075 16540 8084
rect 16488 8041 16497 8075
rect 16497 8041 16531 8075
rect 16531 8041 16540 8075
rect 16488 8032 16540 8041
rect 17040 8032 17092 8084
rect 22468 8032 22520 8084
rect 23756 8075 23808 8084
rect 23756 8041 23765 8075
rect 23765 8041 23799 8075
rect 23799 8041 23808 8075
rect 23756 8032 23808 8041
rect 11060 7964 11112 8016
rect 18512 7964 18564 8016
rect 19340 7964 19392 8016
rect 19800 8007 19852 8016
rect 19800 7973 19809 8007
rect 19809 7973 19843 8007
rect 19843 7973 19852 8007
rect 19800 7964 19852 7973
rect 20720 7964 20772 8016
rect 24768 7964 24820 8016
rect 18604 7896 18656 7948
rect 19984 7896 20036 7948
rect 20628 7896 20680 7948
rect 21916 7896 21968 7948
rect 23664 7896 23716 7948
rect 25136 7896 25188 7948
rect 18052 7828 18104 7880
rect 18236 7871 18288 7880
rect 18236 7837 18245 7871
rect 18245 7837 18279 7871
rect 18279 7837 18288 7871
rect 18236 7828 18288 7837
rect 20720 7828 20772 7880
rect 20904 7871 20956 7880
rect 20904 7837 20913 7871
rect 20913 7837 20947 7871
rect 20947 7837 20956 7871
rect 20904 7828 20956 7837
rect 15568 7692 15620 7744
rect 20904 7692 20956 7744
rect 21180 7692 21232 7744
rect 25320 7735 25372 7744
rect 25320 7701 25329 7735
rect 25329 7701 25363 7735
rect 25363 7701 25372 7735
rect 25320 7692 25372 7701
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 14372 7531 14424 7540
rect 14372 7497 14381 7531
rect 14381 7497 14415 7531
rect 14415 7497 14424 7531
rect 14372 7488 14424 7497
rect 15752 7488 15804 7540
rect 19432 7531 19484 7540
rect 14556 7420 14608 7472
rect 14648 7284 14700 7336
rect 19432 7497 19441 7531
rect 19441 7497 19475 7531
rect 19475 7497 19484 7531
rect 19432 7488 19484 7497
rect 20720 7488 20772 7540
rect 21916 7531 21968 7540
rect 21916 7497 21925 7531
rect 21925 7497 21959 7531
rect 21959 7497 21968 7531
rect 21916 7488 21968 7497
rect 23664 7488 23716 7540
rect 16488 7463 16540 7472
rect 16488 7429 16497 7463
rect 16497 7429 16531 7463
rect 16531 7429 16540 7463
rect 16488 7420 16540 7429
rect 20168 7420 20220 7472
rect 20352 7420 20404 7472
rect 20628 7463 20680 7472
rect 20628 7429 20637 7463
rect 20637 7429 20671 7463
rect 20671 7429 20680 7463
rect 20628 7420 20680 7429
rect 23204 7420 23256 7472
rect 20260 7352 20312 7404
rect 21180 7395 21232 7404
rect 21180 7361 21189 7395
rect 21189 7361 21223 7395
rect 21223 7361 21232 7395
rect 21180 7352 21232 7361
rect 23388 7352 23440 7404
rect 24768 7352 24820 7404
rect 25136 7352 25188 7404
rect 17868 7327 17920 7336
rect 14372 7216 14424 7268
rect 15568 7216 15620 7268
rect 17868 7293 17877 7327
rect 17877 7293 17911 7327
rect 17911 7293 17920 7327
rect 17868 7284 17920 7293
rect 16212 7191 16264 7200
rect 16212 7157 16221 7191
rect 16221 7157 16255 7191
rect 16255 7157 16264 7191
rect 18144 7216 18196 7268
rect 19800 7216 19852 7268
rect 20904 7327 20956 7336
rect 20904 7293 20913 7327
rect 20913 7293 20947 7327
rect 20947 7293 20956 7327
rect 20904 7284 20956 7293
rect 23204 7284 23256 7336
rect 24584 7327 24636 7336
rect 24584 7293 24593 7327
rect 24593 7293 24627 7327
rect 24627 7293 24636 7327
rect 24584 7284 24636 7293
rect 25320 7284 25372 7336
rect 25504 7327 25556 7336
rect 25504 7293 25513 7327
rect 25513 7293 25547 7327
rect 25547 7293 25556 7327
rect 25504 7284 25556 7293
rect 20536 7216 20588 7268
rect 17500 7191 17552 7200
rect 16212 7148 16264 7157
rect 17500 7157 17509 7191
rect 17509 7157 17543 7191
rect 17543 7157 17552 7191
rect 17500 7148 17552 7157
rect 20076 7191 20128 7200
rect 20076 7157 20085 7191
rect 20085 7157 20119 7191
rect 20119 7157 20128 7191
rect 20076 7148 20128 7157
rect 20260 7148 20312 7200
rect 25044 7148 25096 7200
rect 25688 7191 25740 7200
rect 25688 7157 25697 7191
rect 25697 7157 25731 7191
rect 25731 7157 25740 7191
rect 25688 7148 25740 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 14648 6987 14700 6996
rect 14648 6953 14657 6987
rect 14657 6953 14691 6987
rect 14691 6953 14700 6987
rect 14648 6944 14700 6953
rect 18144 6987 18196 6996
rect 18144 6953 18153 6987
rect 18153 6953 18187 6987
rect 18187 6953 18196 6987
rect 18144 6944 18196 6953
rect 19340 6944 19392 6996
rect 19984 6987 20036 6996
rect 19984 6953 19993 6987
rect 19993 6953 20027 6987
rect 20027 6953 20036 6987
rect 19984 6944 20036 6953
rect 23204 6987 23256 6996
rect 23204 6953 23213 6987
rect 23213 6953 23247 6987
rect 23247 6953 23256 6987
rect 23204 6944 23256 6953
rect 24584 6944 24636 6996
rect 16488 6876 16540 6928
rect 19248 6876 19300 6928
rect 8116 6808 8168 6860
rect 16304 6851 16356 6860
rect 16304 6817 16338 6851
rect 16338 6817 16356 6851
rect 16304 6808 16356 6817
rect 18052 6808 18104 6860
rect 18512 6808 18564 6860
rect 20536 6851 20588 6860
rect 20536 6817 20545 6851
rect 20545 6817 20579 6851
rect 20579 6817 20588 6851
rect 20536 6808 20588 6817
rect 20904 6851 20956 6860
rect 20904 6817 20913 6851
rect 20913 6817 20947 6851
rect 20947 6817 20956 6851
rect 20904 6808 20956 6817
rect 21272 6808 21324 6860
rect 22100 6808 22152 6860
rect 23296 6808 23348 6860
rect 24768 6808 24820 6860
rect 25320 6808 25372 6860
rect 25872 6808 25924 6860
rect 16028 6783 16080 6792
rect 16028 6749 16037 6783
rect 16037 6749 16071 6783
rect 16071 6749 16080 6783
rect 16028 6740 16080 6749
rect 18236 6740 18288 6792
rect 19156 6783 19208 6792
rect 19156 6749 19165 6783
rect 19165 6749 19199 6783
rect 19199 6749 19208 6783
rect 19156 6740 19208 6749
rect 22284 6740 22336 6792
rect 23940 6783 23992 6792
rect 23940 6749 23949 6783
rect 23949 6749 23983 6783
rect 23983 6749 23992 6783
rect 23940 6740 23992 6749
rect 25136 6740 25188 6792
rect 25504 6783 25556 6792
rect 25504 6749 25513 6783
rect 25513 6749 25547 6783
rect 25547 6749 25556 6783
rect 25504 6740 25556 6749
rect 8208 6715 8260 6724
rect 8208 6681 8217 6715
rect 8217 6681 8251 6715
rect 8251 6681 8260 6715
rect 8208 6672 8260 6681
rect 17500 6672 17552 6724
rect 18144 6672 18196 6724
rect 18604 6715 18656 6724
rect 18604 6681 18613 6715
rect 18613 6681 18647 6715
rect 18647 6681 18656 6715
rect 18604 6672 18656 6681
rect 25044 6672 25096 6724
rect 21088 6647 21140 6656
rect 21088 6613 21097 6647
rect 21097 6613 21131 6647
rect 21131 6613 21140 6647
rect 21088 6604 21140 6613
rect 23480 6604 23532 6656
rect 24124 6604 24176 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 13636 6307 13688 6316
rect 13636 6273 13645 6307
rect 13645 6273 13679 6307
rect 13679 6273 13688 6307
rect 13636 6264 13688 6273
rect 16028 6400 16080 6452
rect 17868 6443 17920 6452
rect 17868 6409 17877 6443
rect 17877 6409 17911 6443
rect 17911 6409 17920 6443
rect 17868 6400 17920 6409
rect 19156 6400 19208 6452
rect 20904 6400 20956 6452
rect 21916 6443 21968 6452
rect 21916 6409 21925 6443
rect 21925 6409 21959 6443
rect 21959 6409 21968 6443
rect 21916 6400 21968 6409
rect 22284 6400 22336 6452
rect 23296 6443 23348 6452
rect 23296 6409 23305 6443
rect 23305 6409 23339 6443
rect 23339 6409 23348 6443
rect 23296 6400 23348 6409
rect 23756 6400 23808 6452
rect 23572 6332 23624 6384
rect 24768 6400 24820 6452
rect 25504 6400 25556 6452
rect 24124 6307 24176 6316
rect 24124 6273 24133 6307
rect 24133 6273 24167 6307
rect 24167 6273 24176 6307
rect 24124 6264 24176 6273
rect 20536 6239 20588 6248
rect 8208 6060 8260 6112
rect 20536 6205 20545 6239
rect 20545 6205 20579 6239
rect 20579 6205 20588 6239
rect 20536 6196 20588 6205
rect 23940 6196 23992 6248
rect 24676 6196 24728 6248
rect 14924 6171 14976 6180
rect 14924 6137 14958 6171
rect 14958 6137 14976 6171
rect 14924 6128 14976 6137
rect 14280 6060 14332 6112
rect 15476 6060 15528 6112
rect 16304 6128 16356 6180
rect 18144 6128 18196 6180
rect 20812 6171 20864 6180
rect 20812 6137 20846 6171
rect 20846 6137 20864 6171
rect 20812 6128 20864 6137
rect 24676 6060 24728 6112
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 18144 5899 18196 5908
rect 18144 5865 18153 5899
rect 18153 5865 18187 5899
rect 18187 5865 18196 5899
rect 18144 5856 18196 5865
rect 18512 5899 18564 5908
rect 18512 5865 18521 5899
rect 18521 5865 18555 5899
rect 18555 5865 18564 5899
rect 18512 5856 18564 5865
rect 19248 5899 19300 5908
rect 19248 5865 19257 5899
rect 19257 5865 19291 5899
rect 19291 5865 19300 5899
rect 19248 5856 19300 5865
rect 19984 5856 20036 5908
rect 20812 5856 20864 5908
rect 22100 5856 22152 5908
rect 22376 5856 22428 5908
rect 25320 5899 25372 5908
rect 25320 5865 25329 5899
rect 25329 5865 25363 5899
rect 25363 5865 25372 5899
rect 25320 5856 25372 5865
rect 14004 5788 14056 5840
rect 15568 5831 15620 5840
rect 15568 5797 15602 5831
rect 15602 5797 15620 5831
rect 15568 5788 15620 5797
rect 19156 5788 19208 5840
rect 13912 5720 13964 5772
rect 14924 5720 14976 5772
rect 15384 5720 15436 5772
rect 19800 5720 19852 5772
rect 20536 5720 20588 5772
rect 20720 5720 20772 5772
rect 21548 5720 21600 5772
rect 23572 5788 23624 5840
rect 24124 5788 24176 5840
rect 23940 5720 23992 5772
rect 24676 5720 24728 5772
rect 14188 5695 14240 5704
rect 14188 5661 14197 5695
rect 14197 5661 14231 5695
rect 14231 5661 14240 5695
rect 14188 5652 14240 5661
rect 14832 5584 14884 5636
rect 16028 5516 16080 5568
rect 16580 5516 16632 5568
rect 24768 5559 24820 5568
rect 24768 5525 24777 5559
rect 24777 5525 24811 5559
rect 24811 5525 24820 5559
rect 24768 5516 24820 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 13912 5312 13964 5364
rect 14188 5355 14240 5364
rect 14188 5321 14197 5355
rect 14197 5321 14231 5355
rect 14231 5321 14240 5355
rect 14188 5312 14240 5321
rect 14280 5312 14332 5364
rect 15200 5244 15252 5296
rect 16488 5312 16540 5364
rect 20536 5355 20588 5364
rect 20536 5321 20545 5355
rect 20545 5321 20579 5355
rect 20579 5321 20588 5355
rect 20536 5312 20588 5321
rect 22100 5312 22152 5364
rect 24768 5312 24820 5364
rect 19800 5287 19852 5296
rect 14832 5219 14884 5228
rect 14832 5185 14841 5219
rect 14841 5185 14875 5219
rect 14875 5185 14884 5219
rect 14832 5176 14884 5185
rect 19800 5253 19809 5287
rect 19809 5253 19843 5287
rect 19843 5253 19852 5287
rect 19800 5244 19852 5253
rect 23572 5244 23624 5296
rect 16488 5219 16540 5228
rect 16488 5185 16497 5219
rect 16497 5185 16531 5219
rect 16531 5185 16540 5219
rect 16488 5176 16540 5185
rect 14832 5040 14884 5092
rect 18328 5108 18380 5160
rect 20996 5219 21048 5228
rect 20996 5185 21005 5219
rect 21005 5185 21039 5219
rect 21039 5185 21048 5219
rect 20996 5176 21048 5185
rect 18880 5151 18932 5160
rect 18880 5117 18889 5151
rect 18889 5117 18923 5151
rect 18923 5117 18932 5151
rect 18880 5108 18932 5117
rect 20628 5108 20680 5160
rect 24308 5244 24360 5296
rect 24676 5287 24728 5296
rect 24676 5253 24685 5287
rect 24685 5253 24719 5287
rect 24719 5253 24728 5287
rect 24676 5244 24728 5253
rect 23848 5176 23900 5228
rect 25412 5219 25464 5228
rect 25412 5185 25421 5219
rect 25421 5185 25455 5219
rect 25455 5185 25464 5219
rect 25412 5176 25464 5185
rect 15016 5083 15068 5092
rect 15016 5049 15025 5083
rect 15025 5049 15059 5083
rect 15059 5049 15068 5083
rect 15016 5040 15068 5049
rect 15476 5040 15528 5092
rect 16028 5040 16080 5092
rect 16580 5083 16632 5092
rect 16580 5049 16589 5083
rect 16589 5049 16623 5083
rect 16623 5049 16632 5083
rect 16580 5040 16632 5049
rect 22284 5083 22336 5092
rect 22284 5049 22293 5083
rect 22293 5049 22327 5083
rect 22327 5049 22336 5083
rect 22284 5040 22336 5049
rect 24308 5083 24360 5092
rect 24308 5049 24317 5083
rect 24317 5049 24351 5083
rect 24351 5049 24360 5083
rect 24308 5040 24360 5049
rect 13912 5015 13964 5024
rect 13912 4981 13921 5015
rect 13921 4981 13955 5015
rect 13955 4981 13964 5015
rect 13912 4972 13964 4981
rect 14556 4972 14608 5024
rect 21548 5015 21600 5024
rect 21548 4981 21557 5015
rect 21557 4981 21591 5015
rect 21591 4981 21600 5015
rect 21548 4972 21600 4981
rect 22652 5015 22704 5024
rect 22652 4981 22661 5015
rect 22661 4981 22695 5015
rect 22695 4981 22704 5015
rect 22652 4972 22704 4981
rect 23480 4972 23532 5024
rect 24216 5015 24268 5024
rect 24216 4981 24225 5015
rect 24225 4981 24259 5015
rect 24259 4981 24268 5015
rect 24216 4972 24268 4981
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 14832 4811 14884 4820
rect 14832 4777 14841 4811
rect 14841 4777 14875 4811
rect 14875 4777 14884 4811
rect 14832 4768 14884 4777
rect 15384 4768 15436 4820
rect 16580 4768 16632 4820
rect 23020 4768 23072 4820
rect 24216 4768 24268 4820
rect 15016 4700 15068 4752
rect 15568 4700 15620 4752
rect 23940 4743 23992 4752
rect 23940 4709 23949 4743
rect 23949 4709 23983 4743
rect 23983 4709 23992 4743
rect 23940 4700 23992 4709
rect 13360 4675 13412 4684
rect 13360 4641 13369 4675
rect 13369 4641 13403 4675
rect 13403 4641 13412 4675
rect 13360 4632 13412 4641
rect 15660 4632 15712 4684
rect 19800 4675 19852 4684
rect 19800 4641 19809 4675
rect 19809 4641 19843 4675
rect 19843 4641 19852 4675
rect 19800 4632 19852 4641
rect 21824 4675 21876 4684
rect 21824 4641 21833 4675
rect 21833 4641 21867 4675
rect 21867 4641 21876 4675
rect 21824 4632 21876 4641
rect 23664 4675 23716 4684
rect 23664 4641 23673 4675
rect 23673 4641 23707 4675
rect 23707 4641 23716 4675
rect 23664 4632 23716 4641
rect 25228 4632 25280 4684
rect 23848 4496 23900 4548
rect 13544 4471 13596 4480
rect 13544 4437 13553 4471
rect 13553 4437 13587 4471
rect 13587 4437 13596 4471
rect 13544 4428 13596 4437
rect 15568 4428 15620 4480
rect 22100 4428 22152 4480
rect 25044 4471 25096 4480
rect 25044 4437 25053 4471
rect 25053 4437 25087 4471
rect 25087 4437 25096 4471
rect 25044 4428 25096 4437
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 21824 4267 21876 4276
rect 21824 4233 21833 4267
rect 21833 4233 21867 4267
rect 21867 4233 21876 4267
rect 21824 4224 21876 4233
rect 23664 4224 23716 4276
rect 4896 4088 4948 4140
rect 5356 4088 5408 4140
rect 4252 4020 4304 4072
rect 5448 4020 5500 4072
rect 13452 4088 13504 4140
rect 15292 4131 15344 4140
rect 15292 4097 15301 4131
rect 15301 4097 15335 4131
rect 15335 4097 15344 4131
rect 15292 4088 15344 4097
rect 15844 4063 15896 4072
rect 15844 4029 15853 4063
rect 15853 4029 15887 4063
rect 15887 4029 15896 4063
rect 20168 4088 20220 4140
rect 23020 4088 23072 4140
rect 23204 4088 23256 4140
rect 25964 4131 26016 4140
rect 15844 4020 15896 4029
rect 19800 4063 19852 4072
rect 19800 4029 19809 4063
rect 19809 4029 19843 4063
rect 19843 4029 19852 4063
rect 19800 4020 19852 4029
rect 20444 4020 20496 4072
rect 22560 4020 22612 4072
rect 23756 4020 23808 4072
rect 25228 4063 25280 4072
rect 25228 4029 25237 4063
rect 25237 4029 25271 4063
rect 25271 4029 25280 4063
rect 25228 4020 25280 4029
rect 25964 4097 25973 4131
rect 25973 4097 26007 4131
rect 26007 4097 26016 4131
rect 25964 4088 26016 4097
rect 13636 3995 13688 4004
rect 13636 3961 13645 3995
rect 13645 3961 13679 3995
rect 13679 3961 13688 3995
rect 13636 3952 13688 3961
rect 16120 3995 16172 4004
rect 16120 3961 16129 3995
rect 16129 3961 16163 3995
rect 16163 3961 16172 3995
rect 16120 3952 16172 3961
rect 13360 3884 13412 3936
rect 14924 3927 14976 3936
rect 14924 3893 14933 3927
rect 14933 3893 14967 3927
rect 14967 3893 14976 3927
rect 14924 3884 14976 3893
rect 15660 3927 15712 3936
rect 15660 3893 15669 3927
rect 15669 3893 15703 3927
rect 15703 3893 15712 3927
rect 15660 3884 15712 3893
rect 18880 3927 18932 3936
rect 18880 3893 18889 3927
rect 18889 3893 18923 3927
rect 18923 3893 18932 3927
rect 18880 3884 18932 3893
rect 19984 3927 20036 3936
rect 19984 3893 19993 3927
rect 19993 3893 20027 3927
rect 20027 3893 20036 3927
rect 19984 3884 20036 3893
rect 21088 3927 21140 3936
rect 21088 3893 21097 3927
rect 21097 3893 21131 3927
rect 21131 3893 21140 3927
rect 21088 3884 21140 3893
rect 21824 3884 21876 3936
rect 22192 3884 22244 3936
rect 22652 3927 22704 3936
rect 22652 3893 22661 3927
rect 22661 3893 22695 3927
rect 22695 3893 22704 3927
rect 22652 3884 22704 3893
rect 24492 3927 24544 3936
rect 24492 3893 24501 3927
rect 24501 3893 24535 3927
rect 24535 3893 24544 3927
rect 24492 3884 24544 3893
rect 26884 3952 26936 4004
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 18696 3680 18748 3732
rect 20444 3723 20496 3732
rect 20444 3689 20453 3723
rect 20453 3689 20487 3723
rect 20487 3689 20496 3723
rect 20444 3680 20496 3689
rect 23940 3723 23992 3732
rect 23940 3689 23949 3723
rect 23949 3689 23983 3723
rect 23983 3689 23992 3723
rect 23940 3680 23992 3689
rect 13636 3655 13688 3664
rect 13636 3621 13645 3655
rect 13645 3621 13679 3655
rect 13679 3621 13688 3655
rect 13636 3612 13688 3621
rect 10232 3587 10284 3596
rect 10232 3553 10241 3587
rect 10241 3553 10275 3587
rect 10275 3553 10284 3587
rect 10232 3544 10284 3553
rect 12716 3544 12768 3596
rect 13084 3544 13136 3596
rect 16028 3544 16080 3596
rect 16396 3544 16448 3596
rect 17224 3587 17276 3596
rect 17224 3553 17233 3587
rect 17233 3553 17267 3587
rect 17267 3553 17276 3587
rect 17224 3544 17276 3553
rect 18328 3587 18380 3596
rect 18328 3553 18337 3587
rect 18337 3553 18371 3587
rect 18371 3553 18380 3587
rect 18328 3544 18380 3553
rect 20352 3544 20404 3596
rect 21180 3544 21232 3596
rect 22008 3587 22060 3596
rect 22008 3553 22017 3587
rect 22017 3553 22051 3587
rect 22051 3553 22060 3587
rect 22008 3544 22060 3553
rect 22928 3544 22980 3596
rect 23296 3544 23348 3596
rect 24768 3544 24820 3596
rect 11060 3476 11112 3528
rect 15384 3476 15436 3528
rect 19616 3519 19668 3528
rect 19616 3485 19625 3519
rect 19625 3485 19659 3519
rect 19659 3485 19668 3519
rect 19616 3476 19668 3485
rect 14280 3340 14332 3392
rect 17592 3340 17644 3392
rect 21088 3383 21140 3392
rect 21088 3349 21097 3383
rect 21097 3349 21131 3383
rect 21131 3349 21140 3383
rect 21088 3340 21140 3349
rect 23388 3340 23440 3392
rect 24124 3340 24176 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 10232 3179 10284 3188
rect 10232 3145 10241 3179
rect 10241 3145 10275 3179
rect 10275 3145 10284 3179
rect 10232 3136 10284 3145
rect 13084 3136 13136 3188
rect 16028 3179 16080 3188
rect 16028 3145 16037 3179
rect 16037 3145 16071 3179
rect 16071 3145 16080 3179
rect 16028 3136 16080 3145
rect 16672 3179 16724 3188
rect 16672 3145 16681 3179
rect 16681 3145 16715 3179
rect 16715 3145 16724 3179
rect 16672 3136 16724 3145
rect 17224 3136 17276 3188
rect 18328 3179 18380 3188
rect 18328 3145 18337 3179
rect 18337 3145 18371 3179
rect 18371 3145 18380 3179
rect 18328 3136 18380 3145
rect 18420 3136 18472 3188
rect 19432 3179 19484 3188
rect 19432 3145 19441 3179
rect 19441 3145 19475 3179
rect 19475 3145 19484 3179
rect 19432 3136 19484 3145
rect 20352 3136 20404 3188
rect 21180 3179 21232 3188
rect 21180 3145 21189 3179
rect 21189 3145 21223 3179
rect 21223 3145 21232 3179
rect 21180 3136 21232 3145
rect 23112 3179 23164 3188
rect 23112 3145 23121 3179
rect 23121 3145 23155 3179
rect 23155 3145 23164 3179
rect 23112 3136 23164 3145
rect 23296 3136 23348 3188
rect 24032 3136 24084 3188
rect 24768 3179 24820 3188
rect 24768 3145 24777 3179
rect 24777 3145 24811 3179
rect 24811 3145 24820 3179
rect 24768 3136 24820 3145
rect 7748 2932 7800 2984
rect 10048 2932 10100 2984
rect 13268 3068 13320 3120
rect 13360 3000 13412 3052
rect 14740 2932 14792 2984
rect 16672 2932 16724 2984
rect 19248 2975 19300 2984
rect 9588 2864 9640 2916
rect 12440 2864 12492 2916
rect 12716 2907 12768 2916
rect 12716 2873 12725 2907
rect 12725 2873 12759 2907
rect 12759 2873 12768 2907
rect 12716 2864 12768 2873
rect 17776 2907 17828 2916
rect 17776 2873 17785 2907
rect 17785 2873 17819 2907
rect 17819 2873 17828 2907
rect 19248 2941 19257 2975
rect 19257 2941 19291 2975
rect 19291 2941 19300 2975
rect 19248 2932 19300 2941
rect 20444 2932 20496 2984
rect 20628 2907 20680 2916
rect 17776 2864 17828 2873
rect 20628 2873 20637 2907
rect 20637 2873 20671 2907
rect 20671 2873 20680 2907
rect 20628 2864 20680 2873
rect 22008 2864 22060 2916
rect 23112 2932 23164 2984
rect 24032 2932 24084 2984
rect 24860 2932 24912 2984
rect 22192 2864 22244 2916
rect 17040 2839 17092 2848
rect 17040 2805 17049 2839
rect 17049 2805 17083 2839
rect 17083 2805 17092 2839
rect 17040 2796 17092 2805
rect 24860 2796 24912 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 11060 2456 11112 2508
rect 12440 2456 12492 2508
rect 15384 2592 15436 2644
rect 16212 2635 16264 2644
rect 16212 2601 16221 2635
rect 16221 2601 16255 2635
rect 16255 2601 16264 2635
rect 16212 2592 16264 2601
rect 15936 2456 15988 2508
rect 17868 2592 17920 2644
rect 18788 2635 18840 2644
rect 18788 2601 18797 2635
rect 18797 2601 18831 2635
rect 18831 2601 18840 2635
rect 18788 2592 18840 2601
rect 20260 2635 20312 2644
rect 20260 2601 20269 2635
rect 20269 2601 20303 2635
rect 20303 2601 20312 2635
rect 20260 2592 20312 2601
rect 18696 2456 18748 2508
rect 22560 2592 22612 2644
rect 23020 2635 23072 2644
rect 23020 2601 23029 2635
rect 23029 2601 23063 2635
rect 23063 2601 23072 2635
rect 23020 2592 23072 2601
rect 22836 2499 22888 2508
rect 22836 2465 22845 2499
rect 22845 2465 22879 2499
rect 22879 2465 22888 2499
rect 22836 2456 22888 2465
rect 24584 2499 24636 2508
rect 24584 2465 24593 2499
rect 24593 2465 24627 2499
rect 24627 2465 24636 2499
rect 24584 2456 24636 2465
rect 12808 2363 12860 2372
rect 12808 2329 12817 2363
rect 12817 2329 12851 2363
rect 12851 2329 12860 2363
rect 12808 2320 12860 2329
rect 16856 2320 16908 2372
rect 19524 2320 19576 2372
rect 20904 2320 20956 2372
rect 11336 2295 11388 2304
rect 11336 2261 11345 2295
rect 11345 2261 11379 2295
rect 11379 2261 11388 2295
rect 11336 2252 11388 2261
rect 21916 2295 21968 2304
rect 21916 2261 21925 2295
rect 21925 2261 21959 2295
rect 21959 2261 21968 2295
rect 21916 2252 21968 2261
rect 24768 2295 24820 2304
rect 24768 2261 24777 2295
rect 24777 2261 24811 2295
rect 24811 2261 24820 2295
rect 24768 2252 24820 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 13544 552 13596 604
rect 13912 552 13964 604
<< metal2 >>
rect 294 27520 350 28000
rect 938 27520 994 28000
rect 1582 27520 1638 28000
rect 2318 27520 2374 28000
rect 2962 27520 3018 28000
rect 3698 27520 3754 28000
rect 4342 27520 4398 28000
rect 4986 27520 5042 28000
rect 5722 27520 5778 28000
rect 6366 27520 6422 28000
rect 7102 27520 7158 28000
rect 7746 27520 7802 28000
rect 8390 27520 8446 28000
rect 9126 27520 9182 28000
rect 9770 27520 9826 28000
rect 10506 27520 10562 28000
rect 11150 27520 11206 28000
rect 11886 27520 11942 28000
rect 12530 27520 12586 28000
rect 13174 27520 13230 28000
rect 13910 27520 13966 28000
rect 14554 27520 14610 28000
rect 15290 27520 15346 28000
rect 15934 27520 15990 28000
rect 16578 27520 16634 28000
rect 17314 27520 17370 28000
rect 17958 27520 18014 28000
rect 18694 27520 18750 28000
rect 19338 27520 19394 28000
rect 20074 27520 20130 28000
rect 20718 27520 20774 28000
rect 21362 27520 21418 28000
rect 22098 27520 22154 28000
rect 22742 27520 22798 28000
rect 23478 27520 23534 28000
rect 24122 27520 24178 28000
rect 24582 27704 24638 27713
rect 24582 27639 24638 27648
rect 308 19281 336 27520
rect 952 23633 980 27520
rect 1596 24449 1624 27520
rect 1582 24440 1638 24449
rect 1582 24375 1638 24384
rect 938 23624 994 23633
rect 938 23559 994 23568
rect 2332 20505 2360 27520
rect 2976 24857 3004 27520
rect 2962 24848 3018 24857
rect 2962 24783 3018 24792
rect 3712 23769 3740 27520
rect 4356 24177 4384 27520
rect 5000 24721 5028 27520
rect 5736 25242 5764 27520
rect 5736 25214 6040 25242
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 6012 24818 6040 25214
rect 6000 24812 6052 24818
rect 6000 24754 6052 24760
rect 4986 24712 5042 24721
rect 4986 24647 5042 24656
rect 6380 24410 6408 27520
rect 7116 24834 7144 27520
rect 7116 24806 7328 24834
rect 7196 24676 7248 24682
rect 7196 24618 7248 24624
rect 7208 24410 7236 24618
rect 6368 24404 6420 24410
rect 6368 24346 6420 24352
rect 7196 24404 7248 24410
rect 7196 24346 7248 24352
rect 4342 24168 4398 24177
rect 4342 24103 4398 24112
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 3698 23760 3754 23769
rect 3698 23695 3754 23704
rect 7012 23520 7064 23526
rect 7012 23462 7064 23468
rect 6644 23180 6696 23186
rect 6644 23122 6696 23128
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 6656 22778 6684 23122
rect 7024 23118 7052 23462
rect 7012 23112 7064 23118
rect 7012 23054 7064 23060
rect 6644 22772 6696 22778
rect 6644 22714 6696 22720
rect 7024 22574 7052 23054
rect 7012 22568 7064 22574
rect 7012 22510 7064 22516
rect 6642 22264 6698 22273
rect 6642 22199 6644 22208
rect 6696 22199 6698 22208
rect 6644 22170 6696 22176
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 2318 20496 2374 20505
rect 2318 20431 2374 20440
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 294 19272 350 19281
rect 294 19207 350 19216
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5446 15464 5502 15473
rect 5446 15399 5502 15408
rect 5354 15056 5410 15065
rect 5354 14991 5410 15000
rect 3606 8936 3662 8945
rect 3606 8871 3662 8880
rect 2226 7984 2282 7993
rect 2226 7919 2282 7928
rect 294 5264 350 5273
rect 294 5199 350 5208
rect 308 480 336 5199
rect 1674 4720 1730 4729
rect 1674 4655 1730 4664
rect 1582 4040 1638 4049
rect 1582 3975 1638 3984
rect 938 3768 994 3777
rect 938 3703 994 3712
rect 952 480 980 3703
rect 1596 480 1624 3975
rect 1688 3777 1716 4655
rect 1674 3768 1730 3777
rect 1674 3703 1730 3712
rect 2240 480 2268 7919
rect 2870 2952 2926 2961
rect 2870 2887 2926 2896
rect 2884 480 2912 2887
rect 3620 480 3648 8871
rect 4066 7984 4122 7993
rect 4066 7919 4122 7928
rect 4080 7041 4108 7919
rect 4066 7032 4122 7041
rect 4066 6967 4122 6976
rect 5368 4146 5396 14991
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 4252 4072 4304 4078
rect 4252 4014 4304 4020
rect 4264 480 4292 4014
rect 4908 480 4936 4082
rect 5460 4078 5488 15399
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 7208 13433 7236 24346
rect 7300 21185 7328 24806
rect 7564 24608 7616 24614
rect 7564 24550 7616 24556
rect 7576 24410 7604 24550
rect 7564 24404 7616 24410
rect 7564 24346 7616 24352
rect 7576 23644 7604 24346
rect 7656 23656 7708 23662
rect 7576 23616 7656 23644
rect 7656 23598 7708 23604
rect 7656 22432 7708 22438
rect 7656 22374 7708 22380
rect 7380 22024 7432 22030
rect 7380 21966 7432 21972
rect 7286 21176 7342 21185
rect 7392 21146 7420 21966
rect 7668 21554 7696 22374
rect 7760 22001 7788 27520
rect 8300 24812 8352 24818
rect 8300 24754 8352 24760
rect 8312 24410 8340 24754
rect 8300 24404 8352 24410
rect 8300 24346 8352 24352
rect 8024 24268 8076 24274
rect 8024 24210 8076 24216
rect 7840 24064 7892 24070
rect 7840 24006 7892 24012
rect 7852 22234 7880 24006
rect 8036 23526 8064 24210
rect 8116 24200 8168 24206
rect 8116 24142 8168 24148
rect 8128 23594 8156 24142
rect 8300 23656 8352 23662
rect 8300 23598 8352 23604
rect 8116 23588 8168 23594
rect 8116 23530 8168 23536
rect 8024 23520 8076 23526
rect 8024 23462 8076 23468
rect 8036 22574 8064 23462
rect 8128 22817 8156 23530
rect 8206 23352 8262 23361
rect 8312 23322 8340 23598
rect 8206 23287 8262 23296
rect 8300 23316 8352 23322
rect 8220 23186 8248 23287
rect 8300 23258 8352 23264
rect 8208 23180 8260 23186
rect 8208 23122 8260 23128
rect 8114 22808 8170 22817
rect 8114 22743 8170 22752
rect 8024 22568 8076 22574
rect 8024 22510 8076 22516
rect 8206 22536 8262 22545
rect 7840 22228 7892 22234
rect 7840 22170 7892 22176
rect 7746 21992 7802 22001
rect 7746 21927 7802 21936
rect 7748 21888 7800 21894
rect 7748 21830 7800 21836
rect 7656 21548 7708 21554
rect 7656 21490 7708 21496
rect 7286 21111 7342 21120
rect 7380 21140 7432 21146
rect 7380 21082 7432 21088
rect 7668 21049 7696 21490
rect 7654 21040 7710 21049
rect 7654 20975 7710 20984
rect 7194 13424 7250 13433
rect 7194 13359 7250 13368
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 6274 6352 6330 6361
rect 6274 6287 6330 6296
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5538 3088 5594 3097
rect 5538 3023 5594 3032
rect 5552 480 5580 3023
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 6288 480 6316 6287
rect 7562 5672 7618 5681
rect 7562 5607 7618 5616
rect 6918 4040 6974 4049
rect 6918 3975 6974 3984
rect 6932 480 6960 3975
rect 7576 480 7604 5607
rect 7760 2990 7788 21830
rect 7852 21146 7880 22170
rect 8036 22166 8064 22510
rect 8206 22471 8262 22480
rect 8024 22160 8076 22166
rect 8024 22102 8076 22108
rect 8220 22030 8248 22471
rect 8300 22432 8352 22438
rect 8300 22374 8352 22380
rect 8312 22166 8340 22374
rect 8300 22160 8352 22166
rect 8300 22102 8352 22108
rect 8208 22024 8260 22030
rect 8208 21966 8260 21972
rect 8312 21418 8340 22102
rect 8300 21412 8352 21418
rect 8300 21354 8352 21360
rect 7840 21140 7892 21146
rect 7840 21082 7892 21088
rect 8404 21078 8432 27520
rect 9140 21729 9168 27520
rect 9784 27418 9812 27520
rect 9784 27390 10180 27418
rect 9956 25424 10008 25430
rect 9956 25366 10008 25372
rect 9864 25288 9916 25294
rect 9864 25230 9916 25236
rect 9876 24614 9904 25230
rect 9968 24886 9996 25366
rect 9956 24880 10008 24886
rect 9954 24848 9956 24857
rect 10008 24848 10010 24857
rect 9954 24783 10010 24792
rect 9954 24712 10010 24721
rect 9954 24647 10010 24656
rect 9864 24608 9916 24614
rect 9864 24550 9916 24556
rect 9876 24342 9904 24550
rect 9864 24336 9916 24342
rect 9864 24278 9916 24284
rect 9680 24200 9732 24206
rect 9680 24142 9732 24148
rect 9588 23520 9640 23526
rect 9588 23462 9640 23468
rect 9600 22982 9628 23462
rect 9692 23118 9720 24142
rect 9876 23866 9904 24278
rect 9864 23860 9916 23866
rect 9864 23802 9916 23808
rect 9864 23724 9916 23730
rect 9864 23666 9916 23672
rect 9680 23112 9732 23118
rect 9680 23054 9732 23060
rect 9588 22976 9640 22982
rect 9588 22918 9640 22924
rect 9692 22438 9720 23054
rect 9680 22432 9732 22438
rect 9680 22374 9732 22380
rect 9126 21720 9182 21729
rect 9126 21655 9182 21664
rect 9128 21344 9180 21350
rect 9128 21286 9180 21292
rect 8482 21176 8538 21185
rect 9140 21146 9168 21286
rect 8482 21111 8538 21120
rect 9128 21140 9180 21146
rect 8496 21078 8524 21111
rect 9128 21082 9180 21088
rect 8392 21072 8444 21078
rect 8392 21014 8444 21020
rect 8484 21072 8536 21078
rect 8484 21014 8536 21020
rect 8758 21040 8814 21049
rect 8116 20800 8168 20806
rect 8404 20754 8432 21014
rect 8116 20742 8168 20748
rect 8128 19292 8156 20742
rect 8220 20726 8432 20754
rect 8220 20602 8248 20726
rect 8208 20596 8260 20602
rect 8208 20538 8260 20544
rect 8496 20262 8524 21014
rect 8758 20975 8814 20984
rect 8772 20466 8800 20975
rect 8760 20460 8812 20466
rect 8760 20402 8812 20408
rect 8484 20256 8536 20262
rect 8484 20198 8536 20204
rect 8496 19825 8524 20198
rect 8772 20058 8800 20402
rect 9140 20330 9168 21082
rect 9692 21049 9720 22374
rect 9770 21992 9826 22001
rect 9770 21927 9826 21936
rect 9784 21350 9812 21927
rect 9772 21344 9824 21350
rect 9772 21286 9824 21292
rect 9678 21040 9734 21049
rect 9876 21026 9904 23666
rect 9968 22001 9996 24647
rect 10048 24608 10100 24614
rect 10048 24550 10100 24556
rect 10060 24449 10088 24550
rect 10046 24440 10102 24449
rect 10046 24375 10102 24384
rect 10048 23792 10100 23798
rect 10048 23734 10100 23740
rect 9954 21992 10010 22001
rect 9954 21927 10010 21936
rect 9876 20998 9996 21026
rect 9678 20975 9734 20984
rect 9864 20936 9916 20942
rect 9864 20878 9916 20884
rect 9128 20324 9180 20330
rect 9128 20266 9180 20272
rect 8760 20052 8812 20058
rect 8760 19994 8812 20000
rect 8772 19922 8800 19994
rect 8760 19916 8812 19922
rect 8760 19858 8812 19864
rect 8482 19816 8538 19825
rect 8482 19751 8538 19760
rect 8208 19712 8260 19718
rect 8260 19660 8432 19666
rect 8208 19654 8432 19660
rect 8220 19638 8432 19654
rect 8128 19264 8340 19292
rect 8116 19168 8168 19174
rect 8116 19110 8168 19116
rect 8128 15994 8156 19110
rect 8312 18970 8340 19264
rect 8404 19242 8432 19638
rect 8772 19514 8800 19858
rect 8760 19508 8812 19514
rect 8760 19450 8812 19456
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 8392 19236 8444 19242
rect 8392 19178 8444 19184
rect 8300 18964 8352 18970
rect 8300 18906 8352 18912
rect 8404 18426 8432 19178
rect 9692 19174 9720 19246
rect 8576 19168 8628 19174
rect 8576 19110 8628 19116
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 8588 18698 8616 19110
rect 8576 18692 8628 18698
rect 8576 18634 8628 18640
rect 8392 18420 8444 18426
rect 8392 18362 8444 18368
rect 9496 18284 9548 18290
rect 9496 18226 9548 18232
rect 9312 18080 9364 18086
rect 9312 18022 9364 18028
rect 8036 15966 8156 15994
rect 8036 3641 8064 15966
rect 8942 7576 8998 7585
rect 8942 7511 8998 7520
rect 8116 6860 8168 6866
rect 8116 6802 8168 6808
rect 8128 6610 8156 6802
rect 8206 6760 8262 6769
rect 8206 6695 8208 6704
rect 8260 6695 8262 6704
rect 8208 6666 8260 6672
rect 8128 6582 8248 6610
rect 8220 6118 8248 6582
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 8022 3632 8078 3641
rect 8022 3567 8078 3576
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 8220 480 8248 6054
rect 8956 480 8984 7511
rect 9324 4049 9352 18022
rect 9508 17882 9536 18226
rect 9876 18222 9904 20878
rect 9864 18216 9916 18222
rect 9864 18158 9916 18164
rect 9496 17876 9548 17882
rect 9496 17818 9548 17824
rect 9772 17808 9824 17814
rect 9772 17750 9824 17756
rect 9784 16998 9812 17750
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9588 16584 9640 16590
rect 9588 16526 9640 16532
rect 9600 16250 9628 16526
rect 9588 16244 9640 16250
rect 9588 16186 9640 16192
rect 9784 15065 9812 16934
rect 9770 15056 9826 15065
rect 9770 14991 9826 15000
rect 9968 14929 9996 20998
rect 9954 14920 10010 14929
rect 9954 14855 10010 14864
rect 9494 5808 9550 5817
rect 9494 5743 9550 5752
rect 9310 4040 9366 4049
rect 9310 3975 9366 3984
rect 9508 1034 9536 5743
rect 10060 2990 10088 23734
rect 10152 23730 10180 27390
rect 10520 25786 10548 27520
rect 10520 25758 10732 25786
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10324 25356 10376 25362
rect 10324 25298 10376 25304
rect 10336 24886 10364 25298
rect 10324 24880 10376 24886
rect 10324 24822 10376 24828
rect 10336 24721 10364 24822
rect 10322 24712 10378 24721
rect 10322 24647 10378 24656
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10508 24200 10560 24206
rect 10508 24142 10560 24148
rect 10416 24064 10468 24070
rect 10416 24006 10468 24012
rect 10140 23724 10192 23730
rect 10140 23666 10192 23672
rect 10428 23594 10456 24006
rect 10520 23866 10548 24142
rect 10508 23860 10560 23866
rect 10508 23802 10560 23808
rect 10416 23588 10468 23594
rect 10416 23530 10468 23536
rect 10140 23520 10192 23526
rect 10140 23462 10192 23468
rect 10152 23361 10180 23462
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10138 23352 10194 23361
rect 10289 23344 10585 23364
rect 10138 23287 10194 23296
rect 10324 22704 10376 22710
rect 10324 22646 10376 22652
rect 10140 22568 10192 22574
rect 10336 22545 10364 22646
rect 10140 22510 10192 22516
rect 10322 22536 10378 22545
rect 10152 22273 10180 22510
rect 10322 22471 10378 22480
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10138 22264 10194 22273
rect 10289 22256 10585 22276
rect 10138 22199 10140 22208
rect 10192 22199 10194 22208
rect 10140 22170 10192 22176
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10704 20346 10732 25758
rect 11060 25288 11112 25294
rect 11060 25230 11112 25236
rect 10876 25220 10928 25226
rect 10876 25162 10928 25168
rect 10784 24880 10836 24886
rect 10784 24822 10836 24828
rect 10796 24070 10824 24822
rect 10888 24750 10916 25162
rect 10876 24744 10928 24750
rect 10876 24686 10928 24692
rect 11072 24682 11100 25230
rect 11060 24676 11112 24682
rect 11060 24618 11112 24624
rect 10876 24336 10928 24342
rect 10876 24278 10928 24284
rect 10784 24064 10836 24070
rect 10784 24006 10836 24012
rect 10888 23066 10916 24278
rect 10968 23724 11020 23730
rect 10968 23666 11020 23672
rect 10980 23304 11008 23666
rect 11060 23316 11112 23322
rect 10980 23276 11060 23304
rect 11060 23258 11112 23264
rect 10888 23038 11100 23066
rect 10876 22976 10928 22982
rect 10876 22918 10928 22924
rect 10888 22642 10916 22918
rect 11072 22710 11100 23038
rect 11060 22704 11112 22710
rect 11060 22646 11112 22652
rect 10876 22636 10928 22642
rect 10876 22578 10928 22584
rect 10784 22432 10836 22438
rect 10782 22400 10784 22409
rect 10836 22400 10838 22409
rect 10782 22335 10838 22344
rect 11164 21554 11192 27520
rect 11244 25152 11296 25158
rect 11244 25094 11296 25100
rect 11256 24682 11284 25094
rect 11900 24834 11928 27520
rect 12544 25514 12572 27520
rect 13188 27470 13216 27520
rect 12992 27464 13044 27470
rect 12992 27406 13044 27412
rect 13176 27464 13228 27470
rect 13176 27406 13228 27412
rect 12544 25486 12940 25514
rect 12716 25356 12768 25362
rect 12716 25298 12768 25304
rect 12440 25152 12492 25158
rect 12440 25094 12492 25100
rect 11624 24806 11928 24834
rect 11244 24676 11296 24682
rect 11244 24618 11296 24624
rect 11426 24032 11482 24041
rect 11426 23967 11482 23976
rect 11336 21888 11388 21894
rect 11336 21830 11388 21836
rect 11348 21554 11376 21830
rect 11152 21548 11204 21554
rect 11152 21490 11204 21496
rect 11336 21548 11388 21554
rect 11336 21490 11388 21496
rect 11060 21412 11112 21418
rect 11060 21354 11112 21360
rect 10704 20318 10916 20346
rect 10140 20256 10192 20262
rect 10140 20198 10192 20204
rect 10692 20256 10744 20262
rect 10692 20198 10744 20204
rect 10152 19310 10180 20198
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10600 19916 10652 19922
rect 10600 19858 10652 19864
rect 10612 19802 10640 19858
rect 10704 19802 10732 20198
rect 10784 19916 10836 19922
rect 10784 19858 10836 19864
rect 10612 19774 10732 19802
rect 10140 19304 10192 19310
rect 10140 19246 10192 19252
rect 10152 18902 10180 19246
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10704 18970 10732 19774
rect 10796 19174 10824 19858
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 10692 18964 10744 18970
rect 10692 18906 10744 18912
rect 10140 18896 10192 18902
rect 10140 18838 10192 18844
rect 10152 18290 10180 18838
rect 10600 18760 10652 18766
rect 10600 18702 10652 18708
rect 10690 18728 10746 18737
rect 10612 18465 10640 18702
rect 10690 18663 10746 18672
rect 10598 18456 10654 18465
rect 10598 18391 10600 18400
rect 10652 18391 10654 18400
rect 10600 18362 10652 18368
rect 10140 18284 10192 18290
rect 10140 18226 10192 18232
rect 10704 18086 10732 18663
rect 10784 18624 10836 18630
rect 10784 18566 10836 18572
rect 10692 18080 10744 18086
rect 10692 18022 10744 18028
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10796 17678 10824 18566
rect 10324 17672 10376 17678
rect 10324 17614 10376 17620
rect 10416 17672 10468 17678
rect 10416 17614 10468 17620
rect 10784 17672 10836 17678
rect 10784 17614 10836 17620
rect 10138 17096 10194 17105
rect 10336 17066 10364 17614
rect 10428 17338 10456 17614
rect 10416 17332 10468 17338
rect 10416 17274 10468 17280
rect 10138 17031 10194 17040
rect 10324 17060 10376 17066
rect 10152 16726 10180 17031
rect 10324 17002 10376 17008
rect 10782 16960 10838 16969
rect 10289 16892 10585 16912
rect 10782 16895 10838 16904
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10796 16794 10824 16895
rect 10784 16788 10836 16794
rect 10784 16730 10836 16736
rect 10140 16720 10192 16726
rect 10140 16662 10192 16668
rect 10508 16720 10560 16726
rect 10508 16662 10560 16668
rect 10152 15706 10180 16662
rect 10520 16590 10548 16662
rect 10508 16584 10560 16590
rect 10508 16526 10560 16532
rect 10520 16250 10548 16526
rect 10508 16244 10560 16250
rect 10508 16186 10560 16192
rect 10888 16130 10916 20318
rect 10966 18320 11022 18329
rect 10966 18255 11022 18264
rect 10980 17610 11008 18255
rect 11072 17814 11100 21354
rect 11164 21146 11192 21490
rect 11152 21140 11204 21146
rect 11152 21082 11204 21088
rect 11348 21078 11376 21490
rect 11336 21072 11388 21078
rect 11336 21014 11388 21020
rect 11336 18080 11388 18086
rect 11336 18022 11388 18028
rect 11060 17808 11112 17814
rect 11060 17750 11112 17756
rect 11152 17672 11204 17678
rect 11152 17614 11204 17620
rect 10968 17604 11020 17610
rect 10968 17546 11020 17552
rect 11164 17134 11192 17614
rect 11348 17202 11376 18022
rect 11336 17196 11388 17202
rect 11336 17138 11388 17144
rect 11152 17128 11204 17134
rect 11440 17082 11468 23967
rect 11520 22092 11572 22098
rect 11520 22034 11572 22040
rect 11532 21146 11560 22034
rect 11520 21140 11572 21146
rect 11520 21082 11572 21088
rect 11520 18284 11572 18290
rect 11520 18226 11572 18232
rect 11532 17882 11560 18226
rect 11520 17876 11572 17882
rect 11520 17818 11572 17824
rect 11152 17070 11204 17076
rect 10968 16992 11020 16998
rect 10968 16934 11020 16940
rect 10980 16794 11008 16934
rect 10968 16788 11020 16794
rect 10968 16730 11020 16736
rect 10980 16250 11008 16730
rect 11164 16726 11192 17070
rect 11244 17060 11296 17066
rect 11244 17002 11296 17008
rect 11348 17054 11468 17082
rect 11152 16720 11204 16726
rect 11152 16662 11204 16668
rect 11060 16584 11112 16590
rect 11060 16526 11112 16532
rect 10968 16244 11020 16250
rect 10968 16186 11020 16192
rect 10888 16102 11008 16130
rect 10692 15904 10744 15910
rect 10692 15846 10744 15852
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10600 10600 10652 10606
rect 10598 10568 10600 10577
rect 10652 10568 10654 10577
rect 10598 10503 10654 10512
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10230 3632 10286 3641
rect 10230 3567 10232 3576
rect 10284 3567 10286 3576
rect 10232 3538 10284 3544
rect 10244 3194 10272 3538
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 10048 2984 10100 2990
rect 10048 2926 10100 2932
rect 9588 2916 9640 2922
rect 9588 2858 9640 2864
rect 9600 1737 9628 2858
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 9586 1728 9642 1737
rect 9586 1663 9642 1672
rect 10704 1442 10732 15846
rect 10782 15464 10838 15473
rect 10782 15399 10784 15408
rect 10836 15399 10838 15408
rect 10784 15370 10836 15376
rect 10980 11098 11008 16102
rect 11072 15434 11100 16526
rect 11150 16144 11206 16153
rect 11150 16079 11206 16088
rect 11164 15978 11192 16079
rect 11152 15972 11204 15978
rect 11152 15914 11204 15920
rect 11060 15428 11112 15434
rect 11060 15370 11112 15376
rect 11152 13456 11204 13462
rect 11152 13398 11204 13404
rect 11164 12986 11192 13398
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 11256 12209 11284 17002
rect 11242 12200 11298 12209
rect 11242 12135 11298 12144
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 11164 11098 11192 11154
rect 10980 11070 11192 11098
rect 10980 10470 11008 11070
rect 11256 10792 11284 12135
rect 11348 11286 11376 17054
rect 11532 16998 11560 17818
rect 11624 17218 11652 24806
rect 12452 24698 12480 25094
rect 12728 24954 12756 25298
rect 12716 24948 12768 24954
rect 12716 24890 12768 24896
rect 11980 24676 12032 24682
rect 12452 24670 12572 24698
rect 11980 24618 12032 24624
rect 11992 24070 12020 24618
rect 12256 24268 12308 24274
rect 12256 24210 12308 24216
rect 11980 24064 12032 24070
rect 11980 24006 12032 24012
rect 11992 23254 12020 24006
rect 12268 23866 12296 24210
rect 12440 24064 12492 24070
rect 12440 24006 12492 24012
rect 12256 23860 12308 23866
rect 12256 23802 12308 23808
rect 12452 23662 12480 24006
rect 12440 23656 12492 23662
rect 12440 23598 12492 23604
rect 12348 23520 12400 23526
rect 12400 23468 12480 23474
rect 12348 23462 12480 23468
rect 12360 23446 12480 23462
rect 11980 23248 12032 23254
rect 11980 23190 12032 23196
rect 11886 23080 11942 23089
rect 11886 23015 11942 23024
rect 11796 22704 11848 22710
rect 11796 22646 11848 22652
rect 11808 22166 11836 22646
rect 11900 22234 11928 23015
rect 11992 22778 12020 23190
rect 12072 23180 12124 23186
rect 12072 23122 12124 23128
rect 12084 22982 12112 23122
rect 12452 23118 12480 23446
rect 12440 23112 12492 23118
rect 12440 23054 12492 23060
rect 12072 22976 12124 22982
rect 12072 22918 12124 22924
rect 11980 22772 12032 22778
rect 11980 22714 12032 22720
rect 11888 22228 11940 22234
rect 11888 22170 11940 22176
rect 11796 22160 11848 22166
rect 11702 22128 11758 22137
rect 11796 22102 11848 22108
rect 11702 22063 11704 22072
rect 11756 22063 11758 22072
rect 11704 22034 11756 22040
rect 11808 21146 11836 22102
rect 11900 21418 11928 22170
rect 12084 21962 12112 22918
rect 12544 22710 12572 24670
rect 12622 24168 12678 24177
rect 12622 24103 12678 24112
rect 12636 23866 12664 24103
rect 12624 23860 12676 23866
rect 12624 23802 12676 23808
rect 12624 23316 12676 23322
rect 12624 23258 12676 23264
rect 12532 22704 12584 22710
rect 12532 22646 12584 22652
rect 12636 22234 12664 23258
rect 12624 22228 12676 22234
rect 12624 22170 12676 22176
rect 12072 21956 12124 21962
rect 12072 21898 12124 21904
rect 11888 21412 11940 21418
rect 11888 21354 11940 21360
rect 11980 21344 12032 21350
rect 11980 21286 12032 21292
rect 12256 21344 12308 21350
rect 12256 21286 12308 21292
rect 11796 21140 11848 21146
rect 11796 21082 11848 21088
rect 11704 20936 11756 20942
rect 11704 20878 11756 20884
rect 11716 20398 11744 20878
rect 11704 20392 11756 20398
rect 11704 20334 11756 20340
rect 11716 20262 11744 20334
rect 11704 20256 11756 20262
rect 11704 20198 11756 20204
rect 11704 17536 11756 17542
rect 11756 17496 11836 17524
rect 11704 17478 11756 17484
rect 11808 17338 11836 17496
rect 11796 17332 11848 17338
rect 11796 17274 11848 17280
rect 11624 17190 11744 17218
rect 11520 16992 11572 16998
rect 11520 16934 11572 16940
rect 11532 16658 11560 16934
rect 11612 16720 11664 16726
rect 11612 16662 11664 16668
rect 11520 16652 11572 16658
rect 11520 16594 11572 16600
rect 11426 16008 11482 16017
rect 11426 15943 11482 15952
rect 11440 15910 11468 15943
rect 11532 15910 11560 16594
rect 11624 16114 11652 16662
rect 11612 16108 11664 16114
rect 11612 16050 11664 16056
rect 11428 15904 11480 15910
rect 11428 15846 11480 15852
rect 11520 15904 11572 15910
rect 11520 15846 11572 15852
rect 11440 15502 11468 15846
rect 11428 15496 11480 15502
rect 11428 15438 11480 15444
rect 11624 15162 11652 16050
rect 11612 15156 11664 15162
rect 11612 15098 11664 15104
rect 11610 13424 11666 13433
rect 11610 13359 11666 13368
rect 11428 13320 11480 13326
rect 11428 13262 11480 13268
rect 11440 12782 11468 13262
rect 11428 12776 11480 12782
rect 11428 12718 11480 12724
rect 11520 11552 11572 11558
rect 11520 11494 11572 11500
rect 11336 11280 11388 11286
rect 11336 11222 11388 11228
rect 11532 11150 11560 11494
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11256 10764 11468 10792
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 10980 9761 11008 10406
rect 10966 9752 11022 9761
rect 10966 9687 11022 9696
rect 11440 9058 11468 10764
rect 11532 10266 11560 11086
rect 11624 10441 11652 13359
rect 11610 10432 11666 10441
rect 11610 10367 11666 10376
rect 11520 10260 11572 10266
rect 11520 10202 11572 10208
rect 11716 9217 11744 17190
rect 11808 17066 11836 17274
rect 11796 17060 11848 17066
rect 11796 17002 11848 17008
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 11808 14074 11836 14350
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11992 13433 12020 21286
rect 12268 21146 12296 21286
rect 12256 21140 12308 21146
rect 12256 21082 12308 21088
rect 12072 21072 12124 21078
rect 12072 21014 12124 21020
rect 12084 20602 12112 21014
rect 12072 20596 12124 20602
rect 12072 20538 12124 20544
rect 12084 20058 12112 20538
rect 12072 20052 12124 20058
rect 12072 19994 12124 20000
rect 12348 19916 12400 19922
rect 12348 19858 12400 19864
rect 12360 19310 12388 19858
rect 12532 19712 12584 19718
rect 12532 19654 12584 19660
rect 12544 19310 12572 19654
rect 12728 19310 12756 24890
rect 12808 22976 12860 22982
rect 12808 22918 12860 22924
rect 12820 22506 12848 22918
rect 12808 22500 12860 22506
rect 12808 22442 12860 22448
rect 12820 22273 12848 22442
rect 12806 22264 12862 22273
rect 12806 22199 12862 22208
rect 12808 21616 12860 21622
rect 12808 21558 12860 21564
rect 12820 20913 12848 21558
rect 12806 20904 12862 20913
rect 12806 20839 12862 20848
rect 12808 19508 12860 19514
rect 12808 19450 12860 19456
rect 12348 19304 12400 19310
rect 12070 19272 12126 19281
rect 12348 19246 12400 19252
rect 12532 19304 12584 19310
rect 12532 19246 12584 19252
rect 12716 19304 12768 19310
rect 12716 19246 12768 19252
rect 12070 19207 12126 19216
rect 12084 15638 12112 19207
rect 12164 18896 12216 18902
rect 12164 18838 12216 18844
rect 12176 18222 12204 18838
rect 12440 18624 12492 18630
rect 12440 18566 12492 18572
rect 12452 18290 12480 18566
rect 12440 18284 12492 18290
rect 12440 18226 12492 18232
rect 12164 18216 12216 18222
rect 12162 18184 12164 18193
rect 12216 18184 12218 18193
rect 12162 18119 12218 18128
rect 12256 17536 12308 17542
rect 12256 17478 12308 17484
rect 12268 17338 12296 17478
rect 12544 17338 12572 19246
rect 12622 19000 12678 19009
rect 12622 18935 12678 18944
rect 12636 18766 12664 18935
rect 12624 18760 12676 18766
rect 12676 18720 12756 18748
rect 12624 18702 12676 18708
rect 12622 18456 12678 18465
rect 12728 18426 12756 18720
rect 12622 18391 12678 18400
rect 12716 18420 12768 18426
rect 12256 17332 12308 17338
rect 12256 17274 12308 17280
rect 12532 17332 12584 17338
rect 12532 17274 12584 17280
rect 12440 16108 12492 16114
rect 12440 16050 12492 16056
rect 12072 15632 12124 15638
rect 12072 15574 12124 15580
rect 12084 15026 12112 15574
rect 12452 15570 12480 16050
rect 12164 15564 12216 15570
rect 12164 15506 12216 15512
rect 12440 15564 12492 15570
rect 12440 15506 12492 15512
rect 12176 15162 12204 15506
rect 12164 15156 12216 15162
rect 12164 15098 12216 15104
rect 12072 15020 12124 15026
rect 12072 14962 12124 14968
rect 12176 14600 12204 15098
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12452 14770 12480 14894
rect 12360 14742 12480 14770
rect 12176 14572 12296 14600
rect 12164 14476 12216 14482
rect 12164 14418 12216 14424
rect 12176 14074 12204 14418
rect 12164 14068 12216 14074
rect 12164 14010 12216 14016
rect 12176 13530 12204 14010
rect 12164 13524 12216 13530
rect 12164 13466 12216 13472
rect 11978 13424 12034 13433
rect 11978 13359 12034 13368
rect 12268 13297 12296 14572
rect 12360 13462 12388 14742
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12348 13456 12400 13462
rect 12348 13398 12400 13404
rect 12254 13288 12310 13297
rect 12254 13223 12310 13232
rect 12268 12374 12296 13223
rect 12452 12918 12480 13466
rect 12440 12912 12492 12918
rect 12492 12860 12572 12866
rect 12440 12854 12572 12860
rect 12452 12838 12572 12854
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12348 12640 12400 12646
rect 12348 12582 12400 12588
rect 12360 12374 12388 12582
rect 12256 12368 12308 12374
rect 12162 12336 12218 12345
rect 12256 12310 12308 12316
rect 12348 12368 12400 12374
rect 12348 12310 12400 12316
rect 12162 12271 12218 12280
rect 12176 12238 12204 12271
rect 12164 12232 12216 12238
rect 12164 12174 12216 12180
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11808 11762 11836 12038
rect 12176 11914 12204 12174
rect 12084 11898 12204 11914
rect 12268 11898 12296 12310
rect 12072 11892 12204 11898
rect 12124 11886 12204 11892
rect 12256 11892 12308 11898
rect 12072 11834 12124 11840
rect 12256 11834 12308 11840
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 11796 11280 11848 11286
rect 11796 11222 11848 11228
rect 11808 10577 11836 11222
rect 12360 11218 12388 12310
rect 12348 11212 12400 11218
rect 12348 11154 12400 11160
rect 11794 10568 11850 10577
rect 11794 10503 11850 10512
rect 12164 10464 12216 10470
rect 12360 10452 12388 11154
rect 12452 11150 12480 12718
rect 12544 12714 12572 12838
rect 12532 12708 12584 12714
rect 12532 12650 12584 12656
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 12452 10674 12480 11086
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 12440 10532 12492 10538
rect 12440 10474 12492 10480
rect 12216 10424 12388 10452
rect 12164 10406 12216 10412
rect 12176 10266 12204 10406
rect 12164 10260 12216 10266
rect 12164 10202 12216 10208
rect 12452 9654 12480 10474
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 11702 9208 11758 9217
rect 11702 9143 11758 9152
rect 11440 9030 11744 9058
rect 11060 8016 11112 8022
rect 11060 7958 11112 7964
rect 10874 7168 10930 7177
rect 10874 7103 10930 7112
rect 10244 1414 10732 1442
rect 9508 1006 9628 1034
rect 9600 480 9628 1006
rect 10244 480 10272 1414
rect 10888 480 10916 7103
rect 11072 6361 11100 7958
rect 11058 6352 11114 6361
rect 11058 6287 11114 6296
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 11072 2514 11100 3470
rect 11060 2508 11112 2514
rect 11060 2450 11112 2456
rect 11336 2304 11388 2310
rect 11336 2246 11388 2252
rect 11348 1601 11376 2246
rect 11334 1592 11390 1601
rect 11334 1527 11390 1536
rect 11716 626 11744 9030
rect 12636 7857 12664 18391
rect 12716 18362 12768 18368
rect 12716 18148 12768 18154
rect 12716 18090 12768 18096
rect 12728 17542 12756 18090
rect 12716 17536 12768 17542
rect 12716 17478 12768 17484
rect 12820 16436 12848 19450
rect 12912 16561 12940 25486
rect 13004 20482 13032 27406
rect 13450 24712 13506 24721
rect 13084 24676 13136 24682
rect 13450 24647 13506 24656
rect 13084 24618 13136 24624
rect 13096 24410 13124 24618
rect 13084 24404 13136 24410
rect 13084 24346 13136 24352
rect 13096 24041 13124 24346
rect 13082 24032 13138 24041
rect 13082 23967 13138 23976
rect 13266 23352 13322 23361
rect 13266 23287 13268 23296
rect 13320 23287 13322 23296
rect 13268 23258 13320 23264
rect 13268 23112 13320 23118
rect 13268 23054 13320 23060
rect 13280 22778 13308 23054
rect 13268 22772 13320 22778
rect 13268 22714 13320 22720
rect 13082 22672 13138 22681
rect 13082 22607 13084 22616
rect 13136 22607 13138 22616
rect 13084 22578 13136 22584
rect 13464 22506 13492 24647
rect 13544 24268 13596 24274
rect 13544 24210 13596 24216
rect 13452 22500 13504 22506
rect 13452 22442 13504 22448
rect 13176 21888 13228 21894
rect 13176 21830 13228 21836
rect 13188 21418 13216 21830
rect 13176 21412 13228 21418
rect 13176 21354 13228 21360
rect 13004 20454 13216 20482
rect 12992 20392 13044 20398
rect 12992 20334 13044 20340
rect 13004 19174 13032 20334
rect 13082 20224 13138 20233
rect 13082 20159 13138 20168
rect 13096 19786 13124 20159
rect 13084 19780 13136 19786
rect 13084 19722 13136 19728
rect 13188 19446 13216 20454
rect 13360 20052 13412 20058
rect 13360 19994 13412 20000
rect 13372 19514 13400 19994
rect 13360 19508 13412 19514
rect 13360 19450 13412 19456
rect 13176 19440 13228 19446
rect 13176 19382 13228 19388
rect 13268 19372 13320 19378
rect 13268 19314 13320 19320
rect 12992 19168 13044 19174
rect 12992 19110 13044 19116
rect 13084 17536 13136 17542
rect 13084 17478 13136 17484
rect 13096 17202 13124 17478
rect 13084 17196 13136 17202
rect 13084 17138 13136 17144
rect 12992 16992 13044 16998
rect 12990 16960 12992 16969
rect 13044 16960 13046 16969
rect 12990 16895 13046 16904
rect 12898 16552 12954 16561
rect 12898 16487 12954 16496
rect 12820 16408 12940 16436
rect 12808 15156 12860 15162
rect 12808 15098 12860 15104
rect 12716 15088 12768 15094
rect 12716 15030 12768 15036
rect 12728 14618 12756 15030
rect 12716 14612 12768 14618
rect 12716 14554 12768 14560
rect 12728 14074 12756 14554
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 12820 13938 12848 15098
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 12622 7848 12678 7857
rect 12622 7783 12678 7792
rect 12912 5681 12940 16408
rect 13004 16250 13032 16895
rect 13176 16584 13228 16590
rect 13176 16526 13228 16532
rect 13188 16250 13216 16526
rect 12992 16244 13044 16250
rect 12992 16186 13044 16192
rect 13176 16244 13228 16250
rect 13176 16186 13228 16192
rect 13280 15688 13308 19314
rect 13360 19168 13412 19174
rect 13360 19110 13412 19116
rect 13372 18630 13400 19110
rect 13360 18624 13412 18630
rect 13360 18566 13412 18572
rect 13464 18465 13492 22442
rect 13556 21962 13584 24210
rect 13820 24064 13872 24070
rect 13820 24006 13872 24012
rect 13636 23656 13688 23662
rect 13636 23598 13688 23604
rect 13544 21956 13596 21962
rect 13544 21898 13596 21904
rect 13544 21412 13596 21418
rect 13544 21354 13596 21360
rect 13556 21146 13584 21354
rect 13544 21140 13596 21146
rect 13544 21082 13596 21088
rect 13556 20806 13584 21082
rect 13544 20800 13596 20806
rect 13544 20742 13596 20748
rect 13556 20330 13584 20742
rect 13544 20324 13596 20330
rect 13544 20266 13596 20272
rect 13556 19854 13584 20266
rect 13544 19848 13596 19854
rect 13544 19790 13596 19796
rect 13556 18970 13584 19790
rect 13648 19258 13676 23598
rect 13832 22098 13860 24006
rect 13820 22092 13872 22098
rect 13820 22034 13872 22040
rect 13924 21622 13952 27520
rect 14004 24812 14056 24818
rect 14004 24754 14056 24760
rect 14016 24342 14044 24754
rect 14096 24676 14148 24682
rect 14096 24618 14148 24624
rect 14004 24336 14056 24342
rect 14004 24278 14056 24284
rect 14016 23322 14044 24278
rect 14108 23594 14136 24618
rect 14568 24614 14596 27520
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14556 24608 14608 24614
rect 14556 24550 14608 24556
rect 14464 24200 14516 24206
rect 15304 24177 15332 27520
rect 15948 25498 15976 27520
rect 15936 25492 15988 25498
rect 15936 25434 15988 25440
rect 16212 25288 16264 25294
rect 16212 25230 16264 25236
rect 15476 24608 15528 24614
rect 15476 24550 15528 24556
rect 14464 24142 14516 24148
rect 15290 24168 15346 24177
rect 14476 23866 14504 24142
rect 15290 24103 15346 24112
rect 15384 24064 15436 24070
rect 15384 24006 15436 24012
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 14464 23860 14516 23866
rect 14464 23802 14516 23808
rect 14096 23588 14148 23594
rect 14096 23530 14148 23536
rect 14004 23316 14056 23322
rect 14004 23258 14056 23264
rect 14002 22808 14058 22817
rect 14002 22743 14058 22752
rect 14016 22166 14044 22743
rect 14004 22160 14056 22166
rect 14004 22102 14056 22108
rect 14016 21690 14044 22102
rect 14108 22030 14136 23530
rect 14476 23254 14504 23802
rect 15108 23520 15160 23526
rect 15108 23462 15160 23468
rect 15120 23322 15148 23462
rect 15108 23316 15160 23322
rect 15108 23258 15160 23264
rect 14464 23248 14516 23254
rect 14464 23190 14516 23196
rect 14188 23112 14240 23118
rect 14188 23054 14240 23060
rect 14200 22137 14228 23054
rect 14476 22778 14504 23190
rect 15292 23112 15344 23118
rect 15292 23054 15344 23060
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 14464 22772 14516 22778
rect 14464 22714 14516 22720
rect 14556 22704 14608 22710
rect 14556 22646 14608 22652
rect 14186 22128 14242 22137
rect 14186 22063 14242 22072
rect 14096 22024 14148 22030
rect 14096 21966 14148 21972
rect 14004 21684 14056 21690
rect 14004 21626 14056 21632
rect 13912 21616 13964 21622
rect 13912 21558 13964 21564
rect 14108 21146 14136 21966
rect 14188 21956 14240 21962
rect 14188 21898 14240 21904
rect 14200 21486 14228 21898
rect 14188 21480 14240 21486
rect 14186 21448 14188 21457
rect 14240 21448 14242 21457
rect 14186 21383 14242 21392
rect 14096 21140 14148 21146
rect 14096 21082 14148 21088
rect 13820 20936 13872 20942
rect 13820 20878 13872 20884
rect 13726 20088 13782 20097
rect 13726 20023 13728 20032
rect 13780 20023 13782 20032
rect 13728 19994 13780 20000
rect 13728 19916 13780 19922
rect 13832 19904 13860 20878
rect 13780 19876 13860 19904
rect 13728 19858 13780 19864
rect 14186 19816 14242 19825
rect 14186 19751 14242 19760
rect 14096 19712 14148 19718
rect 14096 19654 14148 19660
rect 14108 19310 14136 19654
rect 14096 19304 14148 19310
rect 13648 19230 14044 19258
rect 14096 19246 14148 19252
rect 13634 19000 13690 19009
rect 13544 18964 13596 18970
rect 13634 18935 13690 18944
rect 13544 18906 13596 18912
rect 13450 18456 13506 18465
rect 13450 18391 13506 18400
rect 13188 15660 13308 15688
rect 13648 15688 13676 18935
rect 13728 18624 13780 18630
rect 13728 18566 13780 18572
rect 13740 18057 13768 18566
rect 13726 18048 13782 18057
rect 13726 17983 13782 17992
rect 13820 17060 13872 17066
rect 13820 17002 13872 17008
rect 13832 15858 13860 17002
rect 14016 16726 14044 19230
rect 14108 18902 14136 19246
rect 14096 18896 14148 18902
rect 14096 18838 14148 18844
rect 14108 18426 14136 18838
rect 14096 18420 14148 18426
rect 14096 18362 14148 18368
rect 14096 17264 14148 17270
rect 14096 17206 14148 17212
rect 14108 17105 14136 17206
rect 14094 17096 14150 17105
rect 14094 17031 14150 17040
rect 14004 16720 14056 16726
rect 14004 16662 14056 16668
rect 13912 16448 13964 16454
rect 13912 16390 13964 16396
rect 13924 16046 13952 16390
rect 13912 16040 13964 16046
rect 13912 15982 13964 15988
rect 13832 15830 13952 15858
rect 13820 15700 13872 15706
rect 13648 15660 13820 15688
rect 13188 12889 13216 15660
rect 13648 15609 13676 15660
rect 13820 15642 13872 15648
rect 13266 15600 13322 15609
rect 13266 15535 13322 15544
rect 13634 15600 13690 15609
rect 13634 15535 13690 15544
rect 13280 14822 13308 15535
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 13636 15428 13688 15434
rect 13636 15370 13688 15376
rect 13452 15360 13504 15366
rect 13452 15302 13504 15308
rect 13360 14952 13412 14958
rect 13360 14894 13412 14900
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13372 14618 13400 14894
rect 13360 14612 13412 14618
rect 13360 14554 13412 14560
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 13268 14272 13320 14278
rect 13268 14214 13320 14220
rect 13174 12880 13230 12889
rect 13174 12815 13230 12824
rect 12992 11824 13044 11830
rect 12992 11766 13044 11772
rect 13004 10266 13032 11766
rect 13176 11620 13228 11626
rect 13176 11562 13228 11568
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 12898 5672 12954 5681
rect 12898 5607 12954 5616
rect 12898 4992 12954 5001
rect 12898 4927 12954 4936
rect 12716 3596 12768 3602
rect 12716 3538 12768 3544
rect 12728 2922 12756 3538
rect 12440 2916 12492 2922
rect 12440 2858 12492 2864
rect 12716 2916 12768 2922
rect 12716 2858 12768 2864
rect 12452 2514 12480 2858
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 12806 2408 12862 2417
rect 12806 2343 12808 2352
rect 12860 2343 12862 2352
rect 12808 2314 12860 2320
rect 12254 1864 12310 1873
rect 12254 1799 12310 1808
rect 11624 598 11744 626
rect 11624 480 11652 598
rect 12268 480 12296 1799
rect 12912 480 12940 4927
rect 13096 3602 13124 9862
rect 13188 5273 13216 11562
rect 13174 5264 13230 5273
rect 13174 5199 13230 5208
rect 13084 3596 13136 3602
rect 13084 3538 13136 3544
rect 13096 3194 13124 3538
rect 13084 3188 13136 3194
rect 13084 3130 13136 3136
rect 13280 3126 13308 14214
rect 13372 14074 13400 14418
rect 13464 14414 13492 15302
rect 13648 15042 13676 15370
rect 13728 15156 13780 15162
rect 13832 15144 13860 15438
rect 13780 15116 13860 15144
rect 13728 15098 13780 15104
rect 13648 15014 13860 15042
rect 13832 14958 13860 15014
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 13452 14408 13504 14414
rect 13452 14350 13504 14356
rect 13832 14346 13860 14894
rect 13820 14340 13872 14346
rect 13820 14282 13872 14288
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13832 13530 13860 13806
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13924 12730 13952 15830
rect 14200 15638 14228 19751
rect 14280 19168 14332 19174
rect 14280 19110 14332 19116
rect 14292 18766 14320 19110
rect 14464 18964 14516 18970
rect 14464 18906 14516 18912
rect 14280 18760 14332 18766
rect 14280 18702 14332 18708
rect 14292 18086 14320 18702
rect 14280 18080 14332 18086
rect 14280 18022 14332 18028
rect 14292 17882 14320 18022
rect 14476 17882 14504 18906
rect 14280 17876 14332 17882
rect 14280 17818 14332 17824
rect 14464 17876 14516 17882
rect 14464 17818 14516 17824
rect 14370 17776 14426 17785
rect 14370 17711 14426 17720
rect 14384 17066 14412 17711
rect 14464 17196 14516 17202
rect 14464 17138 14516 17144
rect 14372 17060 14424 17066
rect 14372 17002 14424 17008
rect 14188 15632 14240 15638
rect 14188 15574 14240 15580
rect 14188 15496 14240 15502
rect 14188 15438 14240 15444
rect 14096 15360 14148 15366
rect 14096 15302 14148 15308
rect 14002 14920 14058 14929
rect 14108 14890 14136 15302
rect 14200 14890 14228 15438
rect 14002 14855 14058 14864
rect 14096 14884 14148 14890
rect 14016 14550 14044 14855
rect 14096 14826 14148 14832
rect 14188 14884 14240 14890
rect 14188 14826 14240 14832
rect 14004 14544 14056 14550
rect 14004 14486 14056 14492
rect 14016 14074 14044 14486
rect 14108 14278 14136 14826
rect 14200 14600 14228 14826
rect 14370 14648 14426 14657
rect 14280 14612 14332 14618
rect 14200 14572 14280 14600
rect 14096 14272 14148 14278
rect 14096 14214 14148 14220
rect 14200 14074 14228 14572
rect 14370 14583 14426 14592
rect 14280 14554 14332 14560
rect 14384 14550 14412 14583
rect 14372 14544 14424 14550
rect 14372 14486 14424 14492
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14004 14068 14056 14074
rect 14004 14010 14056 14016
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 13832 12702 13952 12730
rect 13832 12481 13860 12702
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 13818 12472 13874 12481
rect 13818 12407 13874 12416
rect 13820 12368 13872 12374
rect 13820 12310 13872 12316
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13544 12164 13596 12170
rect 13544 12106 13596 12112
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 13372 9450 13400 12038
rect 13464 11762 13492 12038
rect 13556 11762 13584 12106
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13544 11756 13596 11762
rect 13544 11698 13596 11704
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13464 11354 13492 11494
rect 13556 11354 13584 11698
rect 13740 11665 13768 12174
rect 13832 11898 13860 12310
rect 13924 12306 13952 12582
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 13924 11898 13952 12242
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 13726 11656 13782 11665
rect 13726 11591 13728 11600
rect 13780 11591 13782 11600
rect 13728 11562 13780 11568
rect 13740 11531 13768 11562
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13556 10606 13584 11290
rect 13544 10600 13596 10606
rect 13544 10542 13596 10548
rect 13556 10282 13584 10542
rect 13556 10254 13676 10282
rect 13648 10198 13676 10254
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13636 10192 13688 10198
rect 13636 10134 13688 10140
rect 13542 9752 13598 9761
rect 13542 9687 13598 9696
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 13372 9178 13400 9386
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 13556 9081 13584 9687
rect 13648 9586 13676 10134
rect 13728 9988 13780 9994
rect 13728 9930 13780 9936
rect 13740 9654 13768 9930
rect 13832 9654 13860 10202
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13636 9580 13688 9586
rect 13636 9522 13688 9528
rect 13740 9178 13768 9590
rect 14016 9353 14044 14010
rect 14292 13802 14320 14350
rect 14280 13796 14332 13802
rect 14280 13738 14332 13744
rect 14292 13190 14320 13738
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 14476 13002 14504 17138
rect 14200 12974 14504 13002
rect 14200 12374 14228 12974
rect 14370 12880 14426 12889
rect 14370 12815 14426 12824
rect 14384 12481 14412 12815
rect 14370 12472 14426 12481
rect 14370 12407 14426 12416
rect 14188 12368 14240 12374
rect 14188 12310 14240 12316
rect 14002 9344 14058 9353
rect 14002 9279 14058 9288
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13542 9072 13598 9081
rect 13542 9007 13598 9016
rect 13450 8392 13506 8401
rect 13450 8327 13506 8336
rect 13360 4684 13412 4690
rect 13360 4626 13412 4632
rect 13372 3942 13400 4626
rect 13464 4146 13492 8327
rect 14384 7546 14412 12407
rect 14568 10033 14596 22646
rect 14646 22536 14702 22545
rect 15304 22506 15332 23054
rect 15396 22574 15424 24006
rect 15384 22568 15436 22574
rect 15384 22510 15436 22516
rect 14646 22471 14702 22480
rect 15292 22500 15344 22506
rect 14660 22166 14688 22471
rect 15292 22442 15344 22448
rect 15108 22432 15160 22438
rect 15108 22374 15160 22380
rect 14648 22160 14700 22166
rect 14648 22102 14700 22108
rect 14554 10024 14610 10033
rect 14554 9959 14610 9968
rect 14372 7540 14424 7546
rect 14372 7482 14424 7488
rect 14384 7274 14412 7482
rect 14556 7472 14608 7478
rect 14556 7414 14608 7420
rect 14372 7268 14424 7274
rect 14372 7210 14424 7216
rect 13634 6352 13690 6361
rect 13634 6287 13636 6296
rect 13688 6287 13690 6296
rect 13636 6258 13688 6264
rect 14280 6112 14332 6118
rect 14280 6054 14332 6060
rect 14004 5840 14056 5846
rect 14004 5782 14056 5788
rect 13912 5772 13964 5778
rect 13912 5714 13964 5720
rect 13924 5370 13952 5714
rect 13912 5364 13964 5370
rect 13912 5306 13964 5312
rect 13912 5024 13964 5030
rect 14016 5012 14044 5782
rect 14188 5704 14240 5710
rect 14188 5646 14240 5652
rect 14200 5370 14228 5646
rect 14292 5370 14320 6054
rect 14188 5364 14240 5370
rect 14188 5306 14240 5312
rect 14280 5364 14332 5370
rect 14280 5306 14332 5312
rect 14568 5030 14596 7414
rect 14660 7342 14688 22102
rect 15120 22098 15148 22374
rect 15108 22092 15160 22098
rect 15108 22034 15160 22040
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14738 21720 14794 21729
rect 14956 21712 15252 21732
rect 14738 21655 14740 21664
rect 14792 21655 14794 21664
rect 14740 21626 14792 21632
rect 14752 21350 14780 21626
rect 14740 21344 14792 21350
rect 14740 21286 14792 21292
rect 15304 20942 15332 22442
rect 15488 21078 15516 24550
rect 15844 24336 15896 24342
rect 15844 24278 15896 24284
rect 15752 24200 15804 24206
rect 15856 24177 15884 24278
rect 15936 24200 15988 24206
rect 15752 24142 15804 24148
rect 15842 24168 15898 24177
rect 15764 21962 15792 24142
rect 15936 24142 15988 24148
rect 15842 24103 15898 24112
rect 15856 23526 15884 24103
rect 15948 23866 15976 24142
rect 15936 23860 15988 23866
rect 15936 23802 15988 23808
rect 15844 23520 15896 23526
rect 15844 23462 15896 23468
rect 15948 23254 15976 23802
rect 16118 23624 16174 23633
rect 16118 23559 16120 23568
rect 16172 23559 16174 23568
rect 16120 23530 16172 23536
rect 15936 23248 15988 23254
rect 15936 23190 15988 23196
rect 16224 22030 16252 25230
rect 16304 24744 16356 24750
rect 16592 24698 16620 27520
rect 16304 24686 16356 24692
rect 16316 24614 16344 24686
rect 16500 24682 16620 24698
rect 16488 24676 16620 24682
rect 16540 24670 16620 24676
rect 16488 24618 16540 24624
rect 16304 24608 16356 24614
rect 16302 24576 16304 24585
rect 16356 24576 16358 24585
rect 16302 24511 16358 24520
rect 17328 24410 17356 27520
rect 17776 24744 17828 24750
rect 17972 24698 18000 27520
rect 18602 24848 18658 24857
rect 18602 24783 18658 24792
rect 17776 24686 17828 24692
rect 17316 24404 17368 24410
rect 17316 24346 17368 24352
rect 16486 24304 16542 24313
rect 16486 24239 16542 24248
rect 16856 24268 16908 24274
rect 16396 24064 16448 24070
rect 16396 24006 16448 24012
rect 16408 23769 16436 24006
rect 16500 23866 16528 24239
rect 16856 24210 16908 24216
rect 17592 24268 17644 24274
rect 17592 24210 17644 24216
rect 16488 23860 16540 23866
rect 16488 23802 16540 23808
rect 16394 23760 16450 23769
rect 16394 23695 16396 23704
rect 16448 23695 16450 23704
rect 16396 23666 16448 23672
rect 16408 23338 16436 23666
rect 16408 23310 16528 23338
rect 16394 22944 16450 22953
rect 16394 22879 16450 22888
rect 16304 22228 16356 22234
rect 16304 22170 16356 22176
rect 16212 22024 16264 22030
rect 16212 21966 16264 21972
rect 15752 21956 15804 21962
rect 15752 21898 15804 21904
rect 15568 21888 15620 21894
rect 15568 21830 15620 21836
rect 16028 21888 16080 21894
rect 16028 21830 16080 21836
rect 15580 21418 15608 21830
rect 15568 21412 15620 21418
rect 15568 21354 15620 21360
rect 15660 21344 15712 21350
rect 15660 21286 15712 21292
rect 15476 21072 15528 21078
rect 15476 21014 15528 21020
rect 15292 20936 15344 20942
rect 15292 20878 15344 20884
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15304 20262 15332 20878
rect 15672 20777 15700 21286
rect 15844 21004 15896 21010
rect 15844 20946 15896 20952
rect 15658 20768 15714 20777
rect 15658 20703 15714 20712
rect 15476 20528 15528 20534
rect 15476 20470 15528 20476
rect 15292 20256 15344 20262
rect 15292 20198 15344 20204
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15304 19242 15332 20198
rect 15292 19236 15344 19242
rect 15292 19178 15344 19184
rect 14832 18624 14884 18630
rect 14832 18566 14884 18572
rect 15384 18624 15436 18630
rect 15384 18566 15436 18572
rect 14844 18329 14872 18566
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14830 18320 14886 18329
rect 14830 18255 14886 18264
rect 15396 17746 15424 18566
rect 14740 17740 14792 17746
rect 14740 17682 14792 17688
rect 15384 17740 15436 17746
rect 15384 17682 15436 17688
rect 14752 16726 14780 17682
rect 14832 17536 14884 17542
rect 14832 17478 14884 17484
rect 14844 17241 14872 17478
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14830 17232 14886 17241
rect 14830 17167 14832 17176
rect 14884 17167 14886 17176
rect 14832 17138 14884 17144
rect 14832 17060 14884 17066
rect 14832 17002 14884 17008
rect 14740 16720 14792 16726
rect 14740 16662 14792 16668
rect 14844 16250 14872 17002
rect 15384 16652 15436 16658
rect 15384 16594 15436 16600
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 14832 16244 14884 16250
rect 14832 16186 14884 16192
rect 15108 16176 15160 16182
rect 15108 16118 15160 16124
rect 14832 15904 14884 15910
rect 14832 15846 14884 15852
rect 14740 15632 14792 15638
rect 14740 15574 14792 15580
rect 14752 13569 14780 15574
rect 14844 15502 14872 15846
rect 15120 15706 15148 16118
rect 15108 15700 15160 15706
rect 15108 15642 15160 15648
rect 14832 15496 14884 15502
rect 14832 15438 14884 15444
rect 14844 14822 14872 15438
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15396 15162 15424 16594
rect 15384 15156 15436 15162
rect 15384 15098 15436 15104
rect 14832 14816 14884 14822
rect 14832 14758 14884 14764
rect 14738 13560 14794 13569
rect 14844 13530 14872 14758
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14738 13495 14794 13504
rect 14832 13524 14884 13530
rect 14832 13466 14884 13472
rect 14844 12628 14872 13466
rect 15292 13184 15344 13190
rect 15292 13126 15344 13132
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15304 12986 15332 13126
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15384 12708 15436 12714
rect 15384 12650 15436 12656
rect 14924 12640 14976 12646
rect 14844 12600 14924 12628
rect 14924 12582 14976 12588
rect 15290 12608 15346 12617
rect 14936 12374 14964 12582
rect 15290 12543 15346 12552
rect 14924 12368 14976 12374
rect 14924 12310 14976 12316
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14752 11694 14780 12038
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14832 11824 14884 11830
rect 14832 11766 14884 11772
rect 14740 11688 14792 11694
rect 14740 11630 14792 11636
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14752 10062 14780 10406
rect 14740 10056 14792 10062
rect 14740 9998 14792 10004
rect 14752 9518 14780 9998
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 14752 9178 14780 9454
rect 14740 9172 14792 9178
rect 14740 9114 14792 9120
rect 14648 7336 14700 7342
rect 14648 7278 14700 7284
rect 14660 7002 14688 7278
rect 14648 6996 14700 7002
rect 14648 6938 14700 6944
rect 14844 5794 14872 11766
rect 14924 11620 14976 11626
rect 14924 11562 14976 11568
rect 14936 11354 14964 11562
rect 14924 11348 14976 11354
rect 14924 11290 14976 11296
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14924 6180 14976 6186
rect 14924 6122 14976 6128
rect 14752 5766 14872 5794
rect 14936 5778 14964 6122
rect 14924 5772 14976 5778
rect 13964 4984 14044 5012
rect 14556 5024 14608 5030
rect 13912 4966 13964 4972
rect 14556 4966 14608 4972
rect 13544 4480 13596 4486
rect 13544 4422 13596 4428
rect 13556 4185 13584 4422
rect 13542 4176 13598 4185
rect 13452 4140 13504 4146
rect 13542 4111 13598 4120
rect 13452 4082 13504 4088
rect 13634 4040 13690 4049
rect 13634 3975 13636 3984
rect 13688 3975 13690 3984
rect 13636 3946 13688 3952
rect 13360 3936 13412 3942
rect 13360 3878 13412 3884
rect 13634 3904 13690 3913
rect 13268 3120 13320 3126
rect 13268 3062 13320 3068
rect 13372 3058 13400 3878
rect 13634 3839 13690 3848
rect 13648 3670 13676 3839
rect 13636 3664 13688 3670
rect 13636 3606 13688 3612
rect 13360 3052 13412 3058
rect 13360 2994 13412 3000
rect 13924 610 13952 4966
rect 14280 3392 14332 3398
rect 14280 3334 14332 3340
rect 13544 604 13596 610
rect 13544 546 13596 552
rect 13912 604 13964 610
rect 13912 546 13964 552
rect 13556 480 13584 546
rect 14292 480 14320 3334
rect 14752 2990 14780 5766
rect 14924 5714 14976 5720
rect 14832 5636 14884 5642
rect 14832 5578 14884 5584
rect 14844 5234 14872 5578
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15200 5296 15252 5302
rect 15200 5238 15252 5244
rect 14832 5228 14884 5234
rect 14832 5170 14884 5176
rect 14832 5092 14884 5098
rect 14832 5034 14884 5040
rect 15016 5092 15068 5098
rect 15016 5034 15068 5040
rect 14844 4826 14872 5034
rect 14832 4820 14884 4826
rect 14832 4762 14884 4768
rect 15028 4758 15056 5034
rect 15212 5001 15240 5238
rect 15198 4992 15254 5001
rect 15198 4927 15254 4936
rect 15016 4752 15068 4758
rect 15016 4694 15068 4700
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14830 4176 14886 4185
rect 15304 4146 15332 12543
rect 15396 12102 15424 12650
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 15396 11762 15424 12038
rect 15384 11756 15436 11762
rect 15384 11698 15436 11704
rect 15488 8401 15516 20470
rect 15856 20398 15884 20946
rect 15934 20904 15990 20913
rect 15934 20839 15990 20848
rect 15844 20392 15896 20398
rect 15844 20334 15896 20340
rect 15752 20324 15804 20330
rect 15752 20266 15804 20272
rect 15764 20233 15792 20266
rect 15750 20224 15806 20233
rect 15750 20159 15806 20168
rect 15764 19990 15792 20159
rect 15856 20058 15884 20334
rect 15948 20330 15976 20839
rect 15936 20324 15988 20330
rect 15936 20266 15988 20272
rect 15844 20052 15896 20058
rect 15844 19994 15896 20000
rect 15752 19984 15804 19990
rect 15752 19926 15804 19932
rect 15660 19848 15712 19854
rect 15660 19790 15712 19796
rect 15672 18834 15700 19790
rect 15750 19272 15806 19281
rect 15750 19207 15752 19216
rect 15804 19207 15806 19216
rect 15752 19178 15804 19184
rect 15844 19168 15896 19174
rect 15842 19136 15844 19145
rect 15896 19136 15898 19145
rect 15764 19094 15842 19122
rect 15660 18828 15712 18834
rect 15660 18770 15712 18776
rect 15672 18426 15700 18770
rect 15660 18420 15712 18426
rect 15660 18362 15712 18368
rect 15658 18184 15714 18193
rect 15658 18119 15714 18128
rect 15568 17672 15620 17678
rect 15568 17614 15620 17620
rect 15580 17338 15608 17614
rect 15568 17332 15620 17338
rect 15568 17274 15620 17280
rect 15672 15858 15700 18119
rect 15764 15994 15792 19094
rect 15842 19071 15898 19080
rect 15856 19011 15884 19071
rect 15936 18760 15988 18766
rect 15936 18702 15988 18708
rect 15948 18154 15976 18702
rect 15936 18148 15988 18154
rect 15936 18090 15988 18096
rect 15842 18048 15898 18057
rect 15842 17983 15898 17992
rect 15856 17882 15884 17983
rect 15844 17876 15896 17882
rect 15844 17818 15896 17824
rect 15856 17338 15884 17818
rect 15844 17332 15896 17338
rect 15844 17274 15896 17280
rect 15844 16720 15896 16726
rect 15844 16662 15896 16668
rect 15856 16182 15884 16662
rect 15936 16584 15988 16590
rect 15936 16526 15988 16532
rect 15844 16176 15896 16182
rect 15844 16118 15896 16124
rect 15948 16046 15976 16526
rect 15936 16040 15988 16046
rect 15764 15966 15884 15994
rect 15936 15982 15988 15988
rect 15672 15830 15792 15858
rect 15568 15564 15620 15570
rect 15568 15506 15620 15512
rect 15580 15162 15608 15506
rect 15568 15156 15620 15162
rect 15568 15098 15620 15104
rect 15580 14618 15608 15098
rect 15658 14648 15714 14657
rect 15568 14612 15620 14618
rect 15658 14583 15714 14592
rect 15568 14554 15620 14560
rect 15568 13184 15620 13190
rect 15568 13126 15620 13132
rect 15580 11626 15608 13126
rect 15568 11620 15620 11626
rect 15568 11562 15620 11568
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 15580 10470 15608 10950
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 15580 8634 15608 10406
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15474 8392 15530 8401
rect 15474 8327 15530 8336
rect 15568 7744 15620 7750
rect 15568 7686 15620 7692
rect 15580 7313 15608 7686
rect 15566 7304 15622 7313
rect 15566 7239 15568 7248
rect 15620 7239 15622 7248
rect 15568 7210 15620 7216
rect 15476 6112 15528 6118
rect 15476 6054 15528 6060
rect 15384 5772 15436 5778
rect 15384 5714 15436 5720
rect 15396 4826 15424 5714
rect 15488 5098 15516 6054
rect 15580 5846 15608 7210
rect 15568 5840 15620 5846
rect 15568 5782 15620 5788
rect 15476 5092 15528 5098
rect 15476 5034 15528 5040
rect 15384 4820 15436 4826
rect 15384 4762 15436 4768
rect 15580 4758 15608 5782
rect 15672 4842 15700 14583
rect 15764 14414 15792 15830
rect 15856 14550 15884 15966
rect 15948 15366 15976 15982
rect 15936 15360 15988 15366
rect 15936 15302 15988 15308
rect 15934 14920 15990 14929
rect 15934 14855 15936 14864
rect 15988 14855 15990 14864
rect 15936 14826 15988 14832
rect 16040 14657 16068 21830
rect 16224 21690 16252 21966
rect 16212 21684 16264 21690
rect 16212 21626 16264 21632
rect 16120 21344 16172 21350
rect 16316 21332 16344 22170
rect 16408 22030 16436 22879
rect 16396 22024 16448 22030
rect 16396 21966 16448 21972
rect 16172 21304 16344 21332
rect 16120 21286 16172 21292
rect 16132 16017 16160 21286
rect 16408 21146 16436 21966
rect 16500 21894 16528 23310
rect 16868 22982 16896 24210
rect 17604 23526 17632 24210
rect 17592 23520 17644 23526
rect 16946 23488 17002 23497
rect 17592 23462 17644 23468
rect 16946 23423 17002 23432
rect 16672 22976 16724 22982
rect 16672 22918 16724 22924
rect 16856 22976 16908 22982
rect 16856 22918 16908 22924
rect 16684 22642 16712 22918
rect 16672 22636 16724 22642
rect 16672 22578 16724 22584
rect 16764 22568 16816 22574
rect 16764 22510 16816 22516
rect 16776 22234 16804 22510
rect 16764 22228 16816 22234
rect 16764 22170 16816 22176
rect 16488 21888 16540 21894
rect 16488 21830 16540 21836
rect 16672 21888 16724 21894
rect 16672 21830 16724 21836
rect 16684 21486 16712 21830
rect 16868 21554 16896 22918
rect 16960 22778 16988 23423
rect 17604 23089 17632 23462
rect 17684 23112 17736 23118
rect 17590 23080 17646 23089
rect 17684 23054 17736 23060
rect 17590 23015 17646 23024
rect 16948 22772 17000 22778
rect 16948 22714 17000 22720
rect 17696 22506 17724 23054
rect 17684 22500 17736 22506
rect 17684 22442 17736 22448
rect 17788 22234 17816 24686
rect 17880 24670 18000 24698
rect 18512 24744 18564 24750
rect 18512 24686 18564 24692
rect 17880 24614 17908 24670
rect 17868 24608 17920 24614
rect 17868 24550 17920 24556
rect 17958 24576 18014 24585
rect 17958 24511 18014 24520
rect 17868 23656 17920 23662
rect 17868 23598 17920 23604
rect 17224 22228 17276 22234
rect 17224 22170 17276 22176
rect 17776 22228 17828 22234
rect 17776 22170 17828 22176
rect 17236 21690 17264 22170
rect 17880 22166 17908 23598
rect 17972 22817 18000 24511
rect 18328 23792 18380 23798
rect 18328 23734 18380 23740
rect 18340 23361 18368 23734
rect 18326 23352 18382 23361
rect 18326 23287 18382 23296
rect 17958 22808 18014 22817
rect 17958 22743 18014 22752
rect 18524 22386 18552 24686
rect 18616 24614 18644 24783
rect 18604 24608 18656 24614
rect 18604 24550 18656 24556
rect 18708 23497 18736 27520
rect 19156 25356 19208 25362
rect 19156 25298 19208 25304
rect 19168 24682 19196 25298
rect 19156 24676 19208 24682
rect 19156 24618 19208 24624
rect 19168 24154 19196 24618
rect 19352 24426 19380 27520
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 20088 25498 20116 27520
rect 20076 25492 20128 25498
rect 20076 25434 20128 25440
rect 19984 25356 20036 25362
rect 19984 25298 20036 25304
rect 19996 24818 20024 25298
rect 20732 24857 20760 27520
rect 20718 24848 20774 24857
rect 19524 24812 19576 24818
rect 19524 24754 19576 24760
rect 19984 24812 20036 24818
rect 20718 24783 20774 24792
rect 19984 24754 20036 24760
rect 19430 24712 19486 24721
rect 19430 24647 19486 24656
rect 19444 24614 19472 24647
rect 19432 24608 19484 24614
rect 19432 24550 19484 24556
rect 19260 24410 19380 24426
rect 19248 24404 19380 24410
rect 19300 24398 19380 24404
rect 19248 24346 19300 24352
rect 19432 24268 19484 24274
rect 19432 24210 19484 24216
rect 19064 24132 19116 24138
rect 19168 24126 19288 24154
rect 19064 24074 19116 24080
rect 18880 24064 18932 24070
rect 18880 24006 18932 24012
rect 18892 23594 18920 24006
rect 18972 23724 19024 23730
rect 18972 23666 19024 23672
rect 18880 23588 18932 23594
rect 18880 23530 18932 23536
rect 18694 23488 18750 23497
rect 18694 23423 18750 23432
rect 18892 22982 18920 23530
rect 18880 22976 18932 22982
rect 18880 22918 18932 22924
rect 18892 22681 18920 22918
rect 18878 22672 18934 22681
rect 18878 22607 18934 22616
rect 18696 22500 18748 22506
rect 18696 22442 18748 22448
rect 18602 22400 18658 22409
rect 18524 22358 18602 22386
rect 18602 22335 18658 22344
rect 18142 22264 18198 22273
rect 18142 22199 18198 22208
rect 17868 22160 17920 22166
rect 17868 22102 17920 22108
rect 17776 22024 17828 22030
rect 17314 21992 17370 22001
rect 17776 21966 17828 21972
rect 17314 21927 17370 21936
rect 17224 21684 17276 21690
rect 17224 21626 17276 21632
rect 16856 21548 16908 21554
rect 16856 21490 16908 21496
rect 16488 21480 16540 21486
rect 16488 21422 16540 21428
rect 16672 21480 16724 21486
rect 16672 21422 16724 21428
rect 16396 21140 16448 21146
rect 16396 21082 16448 21088
rect 16304 20256 16356 20262
rect 16304 20198 16356 20204
rect 16316 19854 16344 20198
rect 16304 19848 16356 19854
rect 16304 19790 16356 19796
rect 16212 19168 16264 19174
rect 16212 19110 16264 19116
rect 16224 18970 16252 19110
rect 16212 18964 16264 18970
rect 16212 18906 16264 18912
rect 16316 18766 16344 19790
rect 16304 18760 16356 18766
rect 16304 18702 16356 18708
rect 16316 18222 16344 18702
rect 16304 18216 16356 18222
rect 16304 18158 16356 18164
rect 16500 17610 16528 21422
rect 16580 21412 16632 21418
rect 16580 21354 16632 21360
rect 16592 20806 16620 21354
rect 16764 21072 16816 21078
rect 16764 21014 16816 21020
rect 16580 20800 16632 20806
rect 16580 20742 16632 20748
rect 16592 19922 16620 20742
rect 16580 19916 16632 19922
rect 16580 19858 16632 19864
rect 16592 18970 16620 19858
rect 16776 19292 16804 21014
rect 16948 20256 17000 20262
rect 16948 20198 17000 20204
rect 16960 19990 16988 20198
rect 16948 19984 17000 19990
rect 16948 19926 17000 19932
rect 16776 19264 16896 19292
rect 16672 19236 16724 19242
rect 16672 19178 16724 19184
rect 16684 19145 16712 19178
rect 16670 19136 16726 19145
rect 16670 19071 16726 19080
rect 16580 18964 16632 18970
rect 16580 18906 16632 18912
rect 16764 18828 16816 18834
rect 16764 18770 16816 18776
rect 16776 18086 16804 18770
rect 16764 18080 16816 18086
rect 16764 18022 16816 18028
rect 16776 17678 16804 18022
rect 16764 17672 16816 17678
rect 16764 17614 16816 17620
rect 16488 17604 16540 17610
rect 16488 17546 16540 17552
rect 16488 17264 16540 17270
rect 16488 17206 16540 17212
rect 16762 17232 16818 17241
rect 16500 16794 16528 17206
rect 16762 17167 16818 17176
rect 16776 17134 16804 17167
rect 16764 17128 16816 17134
rect 16764 17070 16816 17076
rect 16488 16788 16540 16794
rect 16488 16730 16540 16736
rect 16776 16658 16804 17070
rect 16868 16726 16896 19264
rect 17132 18760 17184 18766
rect 17132 18702 17184 18708
rect 17144 18086 17172 18702
rect 17132 18080 17184 18086
rect 17132 18022 17184 18028
rect 17040 17536 17092 17542
rect 17040 17478 17092 17484
rect 17052 17202 17080 17478
rect 17040 17196 17092 17202
rect 17040 17138 17092 17144
rect 16948 16992 17000 16998
rect 16946 16960 16948 16969
rect 17000 16960 17002 16969
rect 16946 16895 17002 16904
rect 17052 16810 17080 17138
rect 16948 16788 17000 16794
rect 17052 16782 17172 16810
rect 16948 16730 17000 16736
rect 16856 16720 16908 16726
rect 16856 16662 16908 16668
rect 16764 16652 16816 16658
rect 16764 16594 16816 16600
rect 16854 16552 16910 16561
rect 16854 16487 16910 16496
rect 16118 16008 16174 16017
rect 16118 15943 16174 15952
rect 16580 15972 16632 15978
rect 16580 15914 16632 15920
rect 16592 15858 16620 15914
rect 16500 15830 16620 15858
rect 16026 14648 16082 14657
rect 16026 14583 16082 14592
rect 15844 14544 15896 14550
rect 15844 14486 15896 14492
rect 15752 14408 15804 14414
rect 15856 14385 15884 14486
rect 15752 14350 15804 14356
rect 15842 14376 15898 14385
rect 15764 14074 15792 14350
rect 15842 14311 15898 14320
rect 15752 14068 15804 14074
rect 15752 14010 15804 14016
rect 15856 13530 15884 14311
rect 16500 14074 16528 15830
rect 16592 15706 16620 15830
rect 16580 15700 16632 15706
rect 16580 15642 16632 15648
rect 16488 14068 16540 14074
rect 16488 14010 16540 14016
rect 16580 13932 16632 13938
rect 16580 13874 16632 13880
rect 15844 13524 15896 13530
rect 15844 13466 15896 13472
rect 16212 13524 16264 13530
rect 16212 13466 16264 13472
rect 16488 13524 16540 13530
rect 16592 13512 16620 13874
rect 16540 13484 16620 13512
rect 16488 13466 16540 13472
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 15764 11898 15792 13262
rect 15936 12368 15988 12374
rect 15936 12310 15988 12316
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 15948 11558 15976 12310
rect 16028 11620 16080 11626
rect 16028 11562 16080 11568
rect 15936 11552 15988 11558
rect 15936 11494 15988 11500
rect 15948 11234 15976 11494
rect 16040 11354 16068 11562
rect 16028 11348 16080 11354
rect 16028 11290 16080 11296
rect 15948 11206 16068 11234
rect 15934 10568 15990 10577
rect 16040 10538 16068 11206
rect 15934 10503 15990 10512
rect 16028 10532 16080 10538
rect 15842 10024 15898 10033
rect 15842 9959 15898 9968
rect 15750 7848 15806 7857
rect 15750 7783 15806 7792
rect 15764 7546 15792 7783
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15672 4814 15792 4842
rect 15568 4752 15620 4758
rect 15568 4694 15620 4700
rect 15660 4684 15712 4690
rect 15660 4626 15712 4632
rect 15568 4480 15620 4486
rect 15568 4422 15620 4428
rect 14830 4111 14886 4120
rect 15292 4140 15344 4146
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 14844 1986 14872 4111
rect 15292 4082 15344 4088
rect 14924 3936 14976 3942
rect 14924 3878 14976 3884
rect 14936 3505 14964 3878
rect 15384 3528 15436 3534
rect 14922 3496 14978 3505
rect 15384 3470 15436 3476
rect 14922 3431 14978 3440
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 15396 2650 15424 3470
rect 15384 2644 15436 2650
rect 15384 2586 15436 2592
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14844 1958 14964 1986
rect 14936 480 14964 1958
rect 15580 480 15608 4422
rect 15672 3942 15700 4626
rect 15660 3936 15712 3942
rect 15658 3904 15660 3913
rect 15712 3904 15714 3913
rect 15658 3839 15714 3848
rect 15764 3777 15792 4814
rect 15856 4078 15884 9959
rect 15844 4072 15896 4078
rect 15844 4014 15896 4020
rect 15750 3768 15806 3777
rect 15750 3703 15806 3712
rect 15948 2514 15976 10503
rect 16028 10474 16080 10480
rect 16040 9908 16068 10474
rect 16120 9920 16172 9926
rect 16040 9880 16120 9908
rect 16040 9654 16068 9880
rect 16120 9862 16172 9868
rect 16028 9648 16080 9654
rect 16028 9590 16080 9596
rect 16040 9450 16068 9590
rect 16028 9444 16080 9450
rect 16028 9386 16080 9392
rect 16224 8945 16252 13466
rect 16580 11212 16632 11218
rect 16500 11172 16580 11200
rect 16500 10266 16528 11172
rect 16580 11154 16632 11160
rect 16764 11076 16816 11082
rect 16764 11018 16816 11024
rect 16580 10736 16632 10742
rect 16580 10678 16632 10684
rect 16776 10690 16804 11018
rect 16868 10849 16896 16487
rect 16960 15978 16988 16730
rect 17040 16652 17092 16658
rect 17040 16594 17092 16600
rect 16948 15972 17000 15978
rect 16948 15914 17000 15920
rect 17052 15366 17080 16594
rect 17040 15360 17092 15366
rect 17040 15302 17092 15308
rect 17144 15094 17172 16782
rect 17132 15088 17184 15094
rect 17132 15030 17184 15036
rect 17144 14618 17172 15030
rect 17132 14612 17184 14618
rect 17132 14554 17184 14560
rect 17144 13938 17172 14554
rect 17236 14006 17264 21626
rect 17224 14000 17276 14006
rect 17224 13942 17276 13948
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 17328 13818 17356 21927
rect 17788 21690 17816 21966
rect 17776 21684 17828 21690
rect 17776 21626 17828 21632
rect 17592 21616 17644 21622
rect 17592 21558 17644 21564
rect 17604 21146 17632 21558
rect 17880 21162 17908 22102
rect 17592 21140 17644 21146
rect 17592 21082 17644 21088
rect 17788 21134 17908 21162
rect 17788 21078 17816 21134
rect 18156 21078 18184 22199
rect 17776 21072 17828 21078
rect 17776 21014 17828 21020
rect 17868 21072 17920 21078
rect 17868 21014 17920 21020
rect 18144 21072 18196 21078
rect 18144 21014 18196 21020
rect 17774 20768 17830 20777
rect 17774 20703 17830 20712
rect 17406 20496 17462 20505
rect 17406 20431 17462 20440
rect 17236 13790 17356 13818
rect 17132 13728 17184 13734
rect 17132 13670 17184 13676
rect 17040 12980 17092 12986
rect 17040 12922 17092 12928
rect 17052 12306 17080 12922
rect 17144 12306 17172 13670
rect 17040 12300 17092 12306
rect 17040 12242 17092 12248
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 17052 11762 17080 12242
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 16948 11348 17000 11354
rect 17052 11336 17080 11698
rect 17000 11308 17080 11336
rect 16948 11290 17000 11296
rect 16854 10840 16910 10849
rect 16854 10775 16910 10784
rect 16488 10260 16540 10266
rect 16488 10202 16540 10208
rect 16302 9208 16358 9217
rect 16302 9143 16358 9152
rect 16210 8936 16266 8945
rect 16210 8871 16266 8880
rect 16316 8362 16344 9143
rect 16592 9110 16620 10678
rect 16776 10662 16896 10690
rect 16764 10532 16816 10538
rect 16764 10474 16816 10480
rect 16776 9586 16804 10474
rect 16764 9580 16816 9586
rect 16764 9522 16816 9528
rect 16868 9178 16896 10662
rect 16948 10124 17000 10130
rect 16948 10066 17000 10072
rect 16960 9722 16988 10066
rect 16948 9716 17000 9722
rect 16948 9658 17000 9664
rect 16960 9602 16988 9658
rect 16960 9574 17080 9602
rect 16856 9172 16908 9178
rect 16856 9114 16908 9120
rect 16580 9104 16632 9110
rect 16580 9046 16632 9052
rect 16396 8832 16448 8838
rect 16396 8774 16448 8780
rect 16304 8356 16356 8362
rect 16304 8298 16356 8304
rect 16212 7200 16264 7206
rect 16210 7168 16212 7177
rect 16264 7168 16266 7177
rect 16210 7103 16266 7112
rect 16304 6860 16356 6866
rect 16304 6802 16356 6808
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 16040 6458 16068 6734
rect 16028 6452 16080 6458
rect 16028 6394 16080 6400
rect 16040 5574 16068 6394
rect 16316 6186 16344 6802
rect 16304 6180 16356 6186
rect 16304 6122 16356 6128
rect 16028 5568 16080 5574
rect 16028 5510 16080 5516
rect 16040 5098 16068 5510
rect 16028 5092 16080 5098
rect 16028 5034 16080 5040
rect 16120 4004 16172 4010
rect 16120 3946 16172 3952
rect 16132 3641 16160 3946
rect 16118 3632 16174 3641
rect 16028 3596 16080 3602
rect 16408 3602 16436 8774
rect 16592 8634 16620 9046
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 16868 8498 16896 9114
rect 16948 9104 17000 9110
rect 16948 9046 17000 9052
rect 16960 8566 16988 9046
rect 16948 8560 17000 8566
rect 16948 8502 17000 8508
rect 17052 8498 17080 9574
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 17040 8492 17092 8498
rect 17040 8434 17092 8440
rect 16580 8424 16632 8430
rect 16580 8366 16632 8372
rect 16592 8106 16620 8366
rect 16764 8356 16816 8362
rect 16764 8298 16816 8304
rect 16500 8090 16712 8106
rect 16488 8084 16712 8090
rect 16540 8078 16712 8084
rect 16488 8026 16540 8032
rect 16488 7472 16540 7478
rect 16488 7414 16540 7420
rect 16500 6934 16528 7414
rect 16488 6928 16540 6934
rect 16488 6870 16540 6876
rect 16580 5568 16632 5574
rect 16580 5510 16632 5516
rect 16486 5400 16542 5409
rect 16486 5335 16488 5344
rect 16540 5335 16542 5344
rect 16488 5306 16540 5312
rect 16500 5234 16528 5306
rect 16488 5228 16540 5234
rect 16488 5170 16540 5176
rect 16592 5098 16620 5510
rect 16580 5092 16632 5098
rect 16580 5034 16632 5040
rect 16592 4826 16620 5034
rect 16580 4820 16632 4826
rect 16580 4762 16632 4768
rect 16118 3567 16174 3576
rect 16396 3596 16448 3602
rect 16028 3538 16080 3544
rect 16396 3538 16448 3544
rect 16040 3194 16068 3538
rect 16118 3496 16174 3505
rect 16118 3431 16174 3440
rect 16028 3188 16080 3194
rect 16028 3130 16080 3136
rect 15936 2508 15988 2514
rect 15936 2450 15988 2456
rect 16132 1986 16160 3431
rect 16684 3194 16712 8078
rect 16776 6225 16804 8298
rect 17052 8090 17080 8434
rect 17236 8430 17264 13790
rect 17420 13530 17448 20431
rect 17500 20392 17552 20398
rect 17500 20334 17552 20340
rect 17512 18086 17540 20334
rect 17788 19258 17816 20703
rect 17880 20602 17908 21014
rect 18328 20936 18380 20942
rect 18328 20878 18380 20884
rect 17960 20800 18012 20806
rect 17960 20742 18012 20748
rect 17868 20596 17920 20602
rect 17868 20538 17920 20544
rect 17972 19310 18000 20742
rect 18340 20330 18368 20878
rect 18328 20324 18380 20330
rect 18328 20266 18380 20272
rect 18340 19854 18368 20266
rect 18328 19848 18380 19854
rect 18328 19790 18380 19796
rect 17960 19304 18012 19310
rect 17788 19230 17908 19258
rect 17960 19246 18012 19252
rect 17776 19168 17828 19174
rect 17776 19110 17828 19116
rect 17500 18080 17552 18086
rect 17788 18057 17816 19110
rect 17500 18022 17552 18028
rect 17774 18048 17830 18057
rect 17774 17983 17830 17992
rect 17498 16688 17554 16697
rect 17498 16623 17554 16632
rect 17512 16250 17540 16623
rect 17500 16244 17552 16250
rect 17552 16204 17632 16232
rect 17500 16186 17552 16192
rect 17500 14544 17552 14550
rect 17500 14486 17552 14492
rect 17512 14074 17540 14486
rect 17500 14068 17552 14074
rect 17500 14010 17552 14016
rect 17408 13524 17460 13530
rect 17408 13466 17460 13472
rect 17316 13456 17368 13462
rect 17316 13398 17368 13404
rect 17498 13424 17554 13433
rect 17328 12866 17356 13398
rect 17498 13359 17554 13368
rect 17408 13320 17460 13326
rect 17408 13262 17460 13268
rect 17420 12986 17448 13262
rect 17408 12980 17460 12986
rect 17408 12922 17460 12928
rect 17328 12850 17448 12866
rect 17328 12844 17460 12850
rect 17328 12838 17408 12844
rect 17408 12786 17460 12792
rect 17420 12442 17448 12786
rect 17408 12436 17460 12442
rect 17408 12378 17460 12384
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 17328 10674 17356 11086
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 17328 10266 17356 10610
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 17328 9722 17356 10202
rect 17512 9761 17540 13359
rect 17604 11898 17632 16204
rect 17684 15972 17736 15978
rect 17684 15914 17736 15920
rect 17696 15706 17724 15914
rect 17684 15700 17736 15706
rect 17684 15642 17736 15648
rect 17696 15162 17724 15642
rect 17776 15496 17828 15502
rect 17776 15438 17828 15444
rect 17684 15156 17736 15162
rect 17684 15098 17736 15104
rect 17788 14822 17816 15438
rect 17776 14816 17828 14822
rect 17776 14758 17828 14764
rect 17788 14414 17816 14758
rect 17776 14408 17828 14414
rect 17776 14350 17828 14356
rect 17788 13734 17816 14350
rect 17776 13728 17828 13734
rect 17776 13670 17828 13676
rect 17880 13530 17908 19230
rect 17960 19168 18012 19174
rect 17960 19110 18012 19116
rect 17684 13524 17736 13530
rect 17684 13466 17736 13472
rect 17868 13524 17920 13530
rect 17868 13466 17920 13472
rect 17696 12918 17724 13466
rect 17776 13252 17828 13258
rect 17776 13194 17828 13200
rect 17684 12912 17736 12918
rect 17684 12854 17736 12860
rect 17696 12646 17724 12854
rect 17684 12640 17736 12646
rect 17682 12608 17684 12617
rect 17736 12608 17738 12617
rect 17682 12543 17738 12552
rect 17788 12442 17816 13194
rect 17868 12980 17920 12986
rect 17868 12922 17920 12928
rect 17880 12442 17908 12922
rect 17972 12594 18000 19110
rect 18512 18624 18564 18630
rect 18512 18566 18564 18572
rect 18616 18578 18644 22335
rect 18708 22166 18736 22442
rect 18696 22160 18748 22166
rect 18696 22102 18748 22108
rect 18878 22128 18934 22137
rect 18708 21486 18736 22102
rect 18878 22063 18934 22072
rect 18892 21962 18920 22063
rect 18880 21956 18932 21962
rect 18880 21898 18932 21904
rect 18984 21554 19012 23666
rect 19076 23526 19104 24074
rect 19156 24064 19208 24070
rect 19156 24006 19208 24012
rect 19064 23520 19116 23526
rect 19064 23462 19116 23468
rect 18972 21548 19024 21554
rect 18972 21490 19024 21496
rect 18696 21480 18748 21486
rect 18696 21422 18748 21428
rect 19076 21350 19104 23462
rect 19168 22545 19196 24006
rect 19260 23225 19288 24126
rect 19340 24064 19392 24070
rect 19340 24006 19392 24012
rect 19246 23216 19302 23225
rect 19246 23151 19302 23160
rect 19246 23080 19302 23089
rect 19246 23015 19302 23024
rect 19154 22536 19210 22545
rect 19154 22471 19210 22480
rect 19260 22234 19288 23015
rect 19352 22273 19380 24006
rect 19444 23526 19472 24210
rect 19536 24206 19564 24754
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19616 24336 19668 24342
rect 19614 24304 19616 24313
rect 19668 24304 19670 24313
rect 19614 24239 19670 24248
rect 19524 24200 19576 24206
rect 19524 24142 19576 24148
rect 19432 23520 19484 23526
rect 19432 23462 19484 23468
rect 19444 22982 19472 23462
rect 19536 23322 19564 24142
rect 19996 24070 20024 24754
rect 20904 24744 20956 24750
rect 20904 24686 20956 24692
rect 20076 24608 20128 24614
rect 20076 24550 20128 24556
rect 20352 24608 20404 24614
rect 20352 24550 20404 24556
rect 20088 24313 20116 24550
rect 20074 24304 20130 24313
rect 20074 24239 20130 24248
rect 19984 24064 20036 24070
rect 19984 24006 20036 24012
rect 20258 23624 20314 23633
rect 20258 23559 20314 23568
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19524 23316 19576 23322
rect 19524 23258 19576 23264
rect 19522 23216 19578 23225
rect 19522 23151 19578 23160
rect 19432 22976 19484 22982
rect 19432 22918 19484 22924
rect 19444 22438 19472 22918
rect 19432 22432 19484 22438
rect 19432 22374 19484 22380
rect 19338 22264 19394 22273
rect 19248 22228 19300 22234
rect 19338 22199 19394 22208
rect 19248 22170 19300 22176
rect 19340 22160 19392 22166
rect 19340 22102 19392 22108
rect 19156 22092 19208 22098
rect 19156 22034 19208 22040
rect 19064 21344 19116 21350
rect 19064 21286 19116 21292
rect 19064 19848 19116 19854
rect 19064 19790 19116 19796
rect 18880 19780 18932 19786
rect 18880 19722 18932 19728
rect 18892 19378 18920 19722
rect 18880 19372 18932 19378
rect 18880 19314 18932 19320
rect 18880 19236 18932 19242
rect 18880 19178 18932 19184
rect 18144 18148 18196 18154
rect 18144 18090 18196 18096
rect 18156 17882 18184 18090
rect 18328 18080 18380 18086
rect 18234 18048 18290 18057
rect 18328 18022 18380 18028
rect 18234 17983 18290 17992
rect 18144 17876 18196 17882
rect 18144 17818 18196 17824
rect 18248 15994 18276 17983
rect 18340 17678 18368 18022
rect 18524 17814 18552 18566
rect 18616 18550 18736 18578
rect 18602 18456 18658 18465
rect 18602 18391 18658 18400
rect 18616 18154 18644 18391
rect 18604 18148 18656 18154
rect 18604 18090 18656 18096
rect 18708 18034 18736 18550
rect 18616 18006 18736 18034
rect 18512 17808 18564 17814
rect 18512 17750 18564 17756
rect 18328 17672 18380 17678
rect 18328 17614 18380 17620
rect 18340 17270 18368 17614
rect 18524 17338 18552 17750
rect 18512 17332 18564 17338
rect 18512 17274 18564 17280
rect 18328 17264 18380 17270
rect 18328 17206 18380 17212
rect 18418 17096 18474 17105
rect 18418 17031 18474 17040
rect 18432 16250 18460 17031
rect 18524 16726 18552 17274
rect 18512 16720 18564 16726
rect 18512 16662 18564 16668
rect 18616 16590 18644 18006
rect 18786 16960 18842 16969
rect 18786 16895 18842 16904
rect 18604 16584 18656 16590
rect 18604 16526 18656 16532
rect 18616 16250 18644 16526
rect 18420 16244 18472 16250
rect 18420 16186 18472 16192
rect 18604 16244 18656 16250
rect 18604 16186 18656 16192
rect 18248 15966 18460 15994
rect 18144 15632 18196 15638
rect 18144 15574 18196 15580
rect 18328 15632 18380 15638
rect 18328 15574 18380 15580
rect 18052 15360 18104 15366
rect 18052 15302 18104 15308
rect 18064 15162 18092 15302
rect 18052 15156 18104 15162
rect 18052 15098 18104 15104
rect 18156 15094 18184 15574
rect 18234 15192 18290 15201
rect 18234 15127 18290 15136
rect 18144 15088 18196 15094
rect 18144 15030 18196 15036
rect 18156 14278 18184 15030
rect 18144 14272 18196 14278
rect 18144 14214 18196 14220
rect 18248 13802 18276 15127
rect 18236 13796 18288 13802
rect 18236 13738 18288 13744
rect 18052 13456 18104 13462
rect 18052 13398 18104 13404
rect 18064 12918 18092 13398
rect 18052 12912 18104 12918
rect 18052 12854 18104 12860
rect 17972 12566 18092 12594
rect 17776 12436 17828 12442
rect 17776 12378 17828 12384
rect 17868 12436 17920 12442
rect 17868 12378 17920 12384
rect 18064 12356 18092 12566
rect 18064 12328 18184 12356
rect 17960 12300 18012 12306
rect 18012 12260 18092 12288
rect 17960 12242 18012 12248
rect 17592 11892 17644 11898
rect 17592 11834 17644 11840
rect 17774 11656 17830 11665
rect 17774 11591 17830 11600
rect 17788 11558 17816 11591
rect 17776 11552 17828 11558
rect 17776 11494 17828 11500
rect 17592 11008 17644 11014
rect 17592 10950 17644 10956
rect 17604 10606 17632 10950
rect 17592 10600 17644 10606
rect 17592 10542 17644 10548
rect 17604 9994 17632 10542
rect 17788 10198 17816 11494
rect 17960 11144 18012 11150
rect 17960 11086 18012 11092
rect 17972 10810 18000 11086
rect 18064 11014 18092 12260
rect 18052 11008 18104 11014
rect 18052 10950 18104 10956
rect 17960 10804 18012 10810
rect 17960 10746 18012 10752
rect 17776 10192 17828 10198
rect 17776 10134 17828 10140
rect 17592 9988 17644 9994
rect 17592 9930 17644 9936
rect 17498 9752 17554 9761
rect 17316 9716 17368 9722
rect 17498 9687 17554 9696
rect 17316 9658 17368 9664
rect 17788 9654 17816 10134
rect 17972 10130 18000 10746
rect 18064 10674 18092 10950
rect 18052 10668 18104 10674
rect 18052 10610 18104 10616
rect 17960 10124 18012 10130
rect 17960 10066 18012 10072
rect 18064 9926 18092 10610
rect 18052 9920 18104 9926
rect 18052 9862 18104 9868
rect 17960 9716 18012 9722
rect 17960 9658 18012 9664
rect 17776 9648 17828 9654
rect 17776 9590 17828 9596
rect 17972 9110 18000 9658
rect 18064 9518 18092 9862
rect 18156 9602 18184 12328
rect 18248 10266 18276 13738
rect 18236 10260 18288 10266
rect 18236 10202 18288 10208
rect 18156 9574 18276 9602
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 18064 9178 18092 9454
rect 18052 9172 18104 9178
rect 18052 9114 18104 9120
rect 17960 9104 18012 9110
rect 17960 9046 18012 9052
rect 18064 8974 18092 9114
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 18064 8498 18092 8910
rect 18052 8492 18104 8498
rect 17880 8452 18052 8480
rect 17224 8424 17276 8430
rect 17224 8366 17276 8372
rect 17040 8084 17092 8090
rect 17040 8026 17092 8032
rect 17880 7342 17908 8452
rect 18052 8434 18104 8440
rect 18248 8004 18276 9574
rect 18340 9110 18368 15574
rect 18432 14074 18460 15966
rect 18616 15858 18644 16186
rect 18694 16008 18750 16017
rect 18694 15943 18696 15952
rect 18748 15943 18750 15952
rect 18696 15914 18748 15920
rect 18616 15830 18736 15858
rect 18604 14884 18656 14890
rect 18604 14826 18656 14832
rect 18616 14550 18644 14826
rect 18604 14544 18656 14550
rect 18604 14486 18656 14492
rect 18708 14396 18736 15830
rect 18616 14368 18736 14396
rect 18420 14068 18472 14074
rect 18420 14010 18472 14016
rect 18420 13524 18472 13530
rect 18420 13466 18472 13472
rect 18432 12782 18460 13466
rect 18616 12889 18644 14368
rect 18696 13388 18748 13394
rect 18696 13330 18748 13336
rect 18602 12880 18658 12889
rect 18602 12815 18658 12824
rect 18420 12776 18472 12782
rect 18420 12718 18472 12724
rect 18604 12776 18656 12782
rect 18604 12718 18656 12724
rect 18418 12608 18474 12617
rect 18418 12543 18474 12552
rect 18432 9602 18460 12543
rect 18616 11121 18644 12718
rect 18708 12714 18736 13330
rect 18800 12730 18828 16895
rect 18892 15638 18920 19178
rect 19076 18970 19104 19790
rect 19064 18964 19116 18970
rect 19064 18906 19116 18912
rect 18970 17232 19026 17241
rect 19168 17218 19196 22034
rect 19352 21690 19380 22102
rect 19444 22030 19472 22374
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19340 21684 19392 21690
rect 19340 21626 19392 21632
rect 19352 21146 19380 21626
rect 19340 21140 19392 21146
rect 19340 21082 19392 21088
rect 19444 21078 19472 21966
rect 19536 21078 19564 23151
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 20168 21888 20220 21894
rect 20168 21830 20220 21836
rect 19984 21548 20036 21554
rect 19984 21490 20036 21496
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19432 21072 19484 21078
rect 19432 21014 19484 21020
rect 19524 21072 19576 21078
rect 19524 21014 19576 21020
rect 19996 20913 20024 21490
rect 20076 21344 20128 21350
rect 20076 21286 20128 21292
rect 20088 21185 20116 21286
rect 20074 21176 20130 21185
rect 20074 21111 20130 21120
rect 20074 21040 20130 21049
rect 20180 21010 20208 21830
rect 20074 20975 20130 20984
rect 20168 21004 20220 21010
rect 19982 20904 20038 20913
rect 19982 20839 20038 20848
rect 19984 20800 20036 20806
rect 19984 20742 20036 20748
rect 19524 20392 19576 20398
rect 19338 20360 19394 20369
rect 19524 20334 19576 20340
rect 19338 20295 19394 20304
rect 19352 20058 19380 20295
rect 19432 20256 19484 20262
rect 19432 20198 19484 20204
rect 19340 20052 19392 20058
rect 19340 19994 19392 20000
rect 19248 19984 19300 19990
rect 19248 19926 19300 19932
rect 19260 19394 19288 19926
rect 19352 19514 19380 19994
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 19260 19366 19380 19394
rect 19352 19310 19380 19366
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 19444 19174 19472 20198
rect 19432 19168 19484 19174
rect 19432 19110 19484 19116
rect 19340 18692 19392 18698
rect 19340 18634 19392 18640
rect 19352 17338 19380 18634
rect 19536 18358 19564 20334
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19800 19712 19852 19718
rect 19800 19654 19852 19660
rect 19812 19378 19840 19654
rect 19800 19372 19852 19378
rect 19800 19314 19852 19320
rect 19996 19242 20024 20742
rect 19984 19236 20036 19242
rect 19984 19178 20036 19184
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19996 18426 20024 19178
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 19524 18352 19576 18358
rect 19524 18294 19576 18300
rect 19524 18148 19576 18154
rect 19524 18090 19576 18096
rect 19536 17882 19564 18090
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19524 17876 19576 17882
rect 19524 17818 19576 17824
rect 19340 17332 19392 17338
rect 19340 17274 19392 17280
rect 18970 17167 19026 17176
rect 19064 17196 19116 17202
rect 18984 16538 19012 17167
rect 19168 17190 19288 17218
rect 19536 17202 19564 17818
rect 19064 17138 19116 17144
rect 19076 16794 19104 17138
rect 19156 17060 19208 17066
rect 19156 17002 19208 17008
rect 19064 16788 19116 16794
rect 19064 16730 19116 16736
rect 18984 16510 19104 16538
rect 18972 16448 19024 16454
rect 18972 16390 19024 16396
rect 18984 16046 19012 16390
rect 18972 16040 19024 16046
rect 18972 15982 19024 15988
rect 18880 15632 18932 15638
rect 18984 15609 19012 15982
rect 18880 15574 18932 15580
rect 18970 15600 19026 15609
rect 18970 15535 19026 15544
rect 19076 15144 19104 16510
rect 18892 15116 19104 15144
rect 18892 12866 18920 15116
rect 19168 15042 19196 17002
rect 19260 16726 19288 17190
rect 19524 17196 19576 17202
rect 19524 17138 19576 17144
rect 19536 16726 19564 17138
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19248 16720 19300 16726
rect 19246 16688 19248 16697
rect 19524 16720 19576 16726
rect 19300 16688 19302 16697
rect 19524 16662 19576 16668
rect 19246 16623 19302 16632
rect 19984 16584 20036 16590
rect 19984 16526 20036 16532
rect 19340 16176 19392 16182
rect 19340 16118 19392 16124
rect 19352 15144 19380 16118
rect 19432 15904 19484 15910
rect 19432 15846 19484 15852
rect 19444 15473 19472 15846
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19430 15464 19486 15473
rect 19430 15399 19486 15408
rect 19076 15014 19196 15042
rect 19260 15116 19380 15144
rect 19260 15026 19288 15116
rect 19248 15020 19300 15026
rect 18972 14476 19024 14482
rect 18972 14418 19024 14424
rect 18984 14074 19012 14418
rect 18972 14068 19024 14074
rect 18972 14010 19024 14016
rect 19076 13326 19104 15014
rect 19248 14962 19300 14968
rect 19260 14906 19288 14962
rect 19996 14929 20024 16526
rect 19168 14878 19288 14906
rect 19982 14920 20038 14929
rect 19168 14618 19196 14878
rect 19982 14855 20038 14864
rect 19248 14816 19300 14822
rect 19248 14758 19300 14764
rect 19260 14618 19288 14758
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19156 14612 19208 14618
rect 19156 14554 19208 14560
rect 19248 14612 19300 14618
rect 19248 14554 19300 14560
rect 19248 14000 19300 14006
rect 19248 13942 19300 13948
rect 19260 13784 19288 13942
rect 19432 13932 19484 13938
rect 19432 13874 19484 13880
rect 19340 13796 19392 13802
rect 19260 13756 19340 13784
rect 19340 13738 19392 13744
rect 19444 13530 19472 13874
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19432 13524 19484 13530
rect 19432 13466 19484 13472
rect 20088 13462 20116 20975
rect 20168 20946 20220 20952
rect 20180 19310 20208 20946
rect 20272 19666 20300 23559
rect 20364 21729 20392 24550
rect 20720 22976 20772 22982
rect 20718 22944 20720 22953
rect 20772 22944 20774 22953
rect 20718 22879 20774 22888
rect 20534 22808 20590 22817
rect 20534 22743 20590 22752
rect 20350 21720 20406 21729
rect 20350 21655 20352 21664
rect 20404 21655 20406 21664
rect 20352 21626 20404 21632
rect 20364 21486 20392 21626
rect 20352 21480 20404 21486
rect 20352 21422 20404 21428
rect 20548 19990 20576 22743
rect 20720 21480 20772 21486
rect 20718 21448 20720 21457
rect 20772 21448 20774 21457
rect 20718 21383 20774 21392
rect 20812 21344 20864 21350
rect 20812 21286 20864 21292
rect 20824 21146 20852 21286
rect 20812 21140 20864 21146
rect 20812 21082 20864 21088
rect 20812 21004 20864 21010
rect 20812 20946 20864 20952
rect 20720 20936 20772 20942
rect 20720 20878 20772 20884
rect 20628 20596 20680 20602
rect 20732 20584 20760 20878
rect 20680 20556 20760 20584
rect 20628 20538 20680 20544
rect 20824 20505 20852 20946
rect 20810 20496 20866 20505
rect 20810 20431 20812 20440
rect 20864 20431 20866 20440
rect 20812 20402 20864 20408
rect 20536 19984 20588 19990
rect 20536 19926 20588 19932
rect 20272 19638 20484 19666
rect 20260 19508 20312 19514
rect 20260 19450 20312 19456
rect 20168 19304 20220 19310
rect 20168 19246 20220 19252
rect 20168 19168 20220 19174
rect 20168 19110 20220 19116
rect 20180 18698 20208 19110
rect 20168 18692 20220 18698
rect 20168 18634 20220 18640
rect 20272 15042 20300 19450
rect 20352 19236 20404 19242
rect 20352 19178 20404 19184
rect 20364 18630 20392 19178
rect 20352 18624 20404 18630
rect 20352 18566 20404 18572
rect 20456 16590 20484 19638
rect 20548 19378 20576 19926
rect 20536 19372 20588 19378
rect 20536 19314 20588 19320
rect 20628 18760 20680 18766
rect 20916 18737 20944 24686
rect 21376 24614 21404 27520
rect 21548 24812 21600 24818
rect 21548 24754 21600 24760
rect 21364 24608 21416 24614
rect 21364 24550 21416 24556
rect 21560 24410 21588 24754
rect 21548 24404 21600 24410
rect 21548 24346 21600 24352
rect 21456 24200 21508 24206
rect 21086 24168 21142 24177
rect 21456 24142 21508 24148
rect 21086 24103 21088 24112
rect 21140 24103 21142 24112
rect 21088 24074 21140 24080
rect 21468 23798 21496 24142
rect 21560 23866 21588 24346
rect 21640 24200 21692 24206
rect 21640 24142 21692 24148
rect 21548 23860 21600 23866
rect 21548 23802 21600 23808
rect 21456 23792 21508 23798
rect 21456 23734 21508 23740
rect 20996 23656 21048 23662
rect 20996 23598 21048 23604
rect 21008 23186 21036 23598
rect 21272 23520 21324 23526
rect 21272 23462 21324 23468
rect 21284 23254 21312 23462
rect 21272 23248 21324 23254
rect 21272 23190 21324 23196
rect 20996 23180 21048 23186
rect 20996 23122 21048 23128
rect 21008 22778 21036 23122
rect 20996 22772 21048 22778
rect 20996 22714 21048 22720
rect 21008 20398 21036 22714
rect 21284 22574 21312 23190
rect 21364 22636 21416 22642
rect 21364 22578 21416 22584
rect 21272 22568 21324 22574
rect 21272 22510 21324 22516
rect 21284 22234 21312 22510
rect 21376 22506 21404 22578
rect 21364 22500 21416 22506
rect 21364 22442 21416 22448
rect 21272 22228 21324 22234
rect 21272 22170 21324 22176
rect 21376 22137 21404 22442
rect 21362 22128 21418 22137
rect 21362 22063 21418 22072
rect 21180 21548 21232 21554
rect 21180 21490 21232 21496
rect 21192 21350 21220 21490
rect 21180 21344 21232 21350
rect 21180 21286 21232 21292
rect 21192 21049 21220 21286
rect 21178 21040 21234 21049
rect 21178 20975 21234 20984
rect 21468 20890 21496 23734
rect 21652 22982 21680 24142
rect 22112 23866 22140 27520
rect 22192 26308 22244 26314
rect 22192 26250 22244 26256
rect 22100 23860 22152 23866
rect 22100 23802 22152 23808
rect 22204 23746 22232 26250
rect 22468 24812 22520 24818
rect 22468 24754 22520 24760
rect 22284 24744 22336 24750
rect 22284 24686 22336 24692
rect 22112 23718 22232 23746
rect 21914 23352 21970 23361
rect 21914 23287 21970 23296
rect 21640 22976 21692 22982
rect 21640 22918 21692 22924
rect 21640 22704 21692 22710
rect 21928 22681 21956 23287
rect 21640 22646 21692 22652
rect 21914 22672 21970 22681
rect 21546 22536 21602 22545
rect 21546 22471 21548 22480
rect 21600 22471 21602 22480
rect 21548 22442 21600 22448
rect 21548 21888 21600 21894
rect 21548 21830 21600 21836
rect 21376 20862 21496 20890
rect 20996 20392 21048 20398
rect 20996 20334 21048 20340
rect 21180 20324 21232 20330
rect 21180 20266 21232 20272
rect 21192 19922 21220 20266
rect 21376 20058 21404 20862
rect 21456 20800 21508 20806
rect 21456 20742 21508 20748
rect 21364 20052 21416 20058
rect 21364 19994 21416 20000
rect 21180 19916 21232 19922
rect 21180 19858 21232 19864
rect 21192 19718 21220 19858
rect 21180 19712 21232 19718
rect 21180 19654 21232 19660
rect 20996 19372 21048 19378
rect 20996 19314 21048 19320
rect 20628 18702 20680 18708
rect 20902 18728 20958 18737
rect 20640 17649 20668 18702
rect 20902 18663 20958 18672
rect 20904 17672 20956 17678
rect 20626 17640 20682 17649
rect 20904 17614 20956 17620
rect 20626 17575 20682 17584
rect 20626 17368 20682 17377
rect 20626 17303 20682 17312
rect 20640 17202 20668 17303
rect 20628 17196 20680 17202
rect 20628 17138 20680 17144
rect 20916 16998 20944 17614
rect 20628 16992 20680 16998
rect 20628 16934 20680 16940
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 20444 16584 20496 16590
rect 20444 16526 20496 16532
rect 20640 16522 20668 16934
rect 20628 16516 20680 16522
rect 20628 16458 20680 16464
rect 20444 16448 20496 16454
rect 20444 16390 20496 16396
rect 20352 15972 20404 15978
rect 20352 15914 20404 15920
rect 20364 15366 20392 15914
rect 20456 15910 20484 16390
rect 20536 15972 20588 15978
rect 20536 15914 20588 15920
rect 20444 15904 20496 15910
rect 20444 15846 20496 15852
rect 20352 15360 20404 15366
rect 20352 15302 20404 15308
rect 20180 15014 20300 15042
rect 20180 14074 20208 15014
rect 20260 14952 20312 14958
rect 20260 14894 20312 14900
rect 20272 14822 20300 14894
rect 20260 14816 20312 14822
rect 20260 14758 20312 14764
rect 20258 14648 20314 14657
rect 20258 14583 20314 14592
rect 20168 14068 20220 14074
rect 20168 14010 20220 14016
rect 20180 13802 20208 14010
rect 20168 13796 20220 13802
rect 20168 13738 20220 13744
rect 19616 13456 19668 13462
rect 19616 13398 19668 13404
rect 20076 13456 20128 13462
rect 20076 13398 20128 13404
rect 19064 13320 19116 13326
rect 19628 13308 19656 13398
rect 19064 13262 19116 13268
rect 19536 13280 19656 13308
rect 19076 12986 19104 13262
rect 19064 12980 19116 12986
rect 19064 12922 19116 12928
rect 18892 12838 19104 12866
rect 18878 12744 18934 12753
rect 18696 12708 18748 12714
rect 18800 12702 18878 12730
rect 18878 12679 18934 12688
rect 18696 12650 18748 12656
rect 18708 12374 18736 12650
rect 18696 12368 18748 12374
rect 18696 12310 18748 12316
rect 18892 11354 18920 12679
rect 18880 11348 18932 11354
rect 18880 11290 18932 11296
rect 18788 11212 18840 11218
rect 18788 11154 18840 11160
rect 18602 11112 18658 11121
rect 18602 11047 18658 11056
rect 18800 10810 18828 11154
rect 18788 10804 18840 10810
rect 18788 10746 18840 10752
rect 18892 10742 18920 11290
rect 19076 11218 19104 12838
rect 19340 12708 19392 12714
rect 19340 12650 19392 12656
rect 19352 11506 19380 12650
rect 19430 12472 19486 12481
rect 19430 12407 19486 12416
rect 19444 12374 19472 12407
rect 19432 12368 19484 12374
rect 19432 12310 19484 12316
rect 19432 11552 19484 11558
rect 19352 11500 19432 11506
rect 19352 11494 19484 11500
rect 19352 11478 19472 11494
rect 19064 11212 19116 11218
rect 19064 11154 19116 11160
rect 18880 10736 18932 10742
rect 18880 10678 18932 10684
rect 19156 10532 19208 10538
rect 19156 10474 19208 10480
rect 18786 10160 18842 10169
rect 18786 10095 18842 10104
rect 18800 9761 18828 10095
rect 19168 9926 19196 10474
rect 19248 10260 19300 10266
rect 19248 10202 19300 10208
rect 19156 9920 19208 9926
rect 19156 9862 19208 9868
rect 18786 9752 18842 9761
rect 19168 9722 19196 9862
rect 18786 9687 18842 9696
rect 19156 9716 19208 9722
rect 18432 9574 18552 9602
rect 18328 9104 18380 9110
rect 18328 9046 18380 9052
rect 18340 8634 18368 9046
rect 18328 8628 18380 8634
rect 18328 8570 18380 8576
rect 18524 8022 18552 9574
rect 18512 8016 18564 8022
rect 18248 7976 18368 8004
rect 18052 7880 18104 7886
rect 18236 7880 18288 7886
rect 18052 7822 18104 7828
rect 18234 7848 18236 7857
rect 18288 7848 18290 7857
rect 17958 7712 18014 7721
rect 17958 7647 18014 7656
rect 17868 7336 17920 7342
rect 17868 7278 17920 7284
rect 17500 7200 17552 7206
rect 17500 7142 17552 7148
rect 17512 6730 17540 7142
rect 17500 6724 17552 6730
rect 17500 6666 17552 6672
rect 17880 6458 17908 7278
rect 17972 6769 18000 7647
rect 18064 6866 18092 7822
rect 18234 7783 18290 7792
rect 18144 7268 18196 7274
rect 18144 7210 18196 7216
rect 18156 7002 18184 7210
rect 18144 6996 18196 7002
rect 18196 6956 18276 6984
rect 18144 6938 18196 6944
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 18248 6798 18276 6956
rect 18236 6792 18288 6798
rect 17958 6760 18014 6769
rect 18236 6734 18288 6740
rect 17958 6695 18014 6704
rect 18144 6724 18196 6730
rect 18144 6666 18196 6672
rect 17868 6452 17920 6458
rect 17868 6394 17920 6400
rect 16762 6216 16818 6225
rect 18156 6186 18184 6666
rect 16762 6151 16818 6160
rect 18144 6180 18196 6186
rect 18144 6122 18196 6128
rect 18156 5914 18184 6122
rect 18144 5908 18196 5914
rect 18144 5850 18196 5856
rect 18340 5166 18368 7976
rect 18512 7958 18564 7964
rect 18604 7948 18656 7954
rect 18604 7890 18656 7896
rect 18512 6860 18564 6866
rect 18512 6802 18564 6808
rect 18524 5914 18552 6802
rect 18616 6730 18644 7890
rect 18694 7440 18750 7449
rect 18694 7375 18750 7384
rect 18604 6724 18656 6730
rect 18604 6666 18656 6672
rect 18512 5908 18564 5914
rect 18512 5850 18564 5856
rect 18328 5160 18380 5166
rect 18328 5102 18380 5108
rect 18326 4720 18382 4729
rect 18326 4655 18382 4664
rect 17222 3768 17278 3777
rect 17222 3703 17278 3712
rect 17236 3602 17264 3703
rect 18340 3618 18368 4655
rect 18708 3738 18736 7375
rect 18696 3732 18748 3738
rect 18696 3674 18748 3680
rect 18800 3618 18828 9687
rect 19156 9658 19208 9664
rect 19260 9636 19288 10202
rect 19340 9648 19392 9654
rect 19260 9608 19340 9636
rect 19340 9590 19392 9596
rect 19338 9344 19394 9353
rect 19338 9279 19394 9288
rect 19352 8566 19380 9279
rect 19340 8560 19392 8566
rect 19340 8502 19392 8508
rect 19340 8424 19392 8430
rect 19340 8366 19392 8372
rect 19352 8022 19380 8366
rect 19340 8016 19392 8022
rect 19340 7958 19392 7964
rect 19352 7002 19380 7958
rect 19444 7546 19472 11478
rect 19536 8634 19564 13280
rect 20180 13274 20208 13738
rect 20088 13246 20208 13274
rect 19984 13184 20036 13190
rect 19984 13126 20036 13132
rect 19996 12782 20024 13126
rect 19984 12776 20036 12782
rect 19984 12718 20036 12724
rect 20088 12594 20116 13246
rect 20168 13184 20220 13190
rect 20168 13126 20220 13132
rect 20180 12646 20208 13126
rect 20272 12866 20300 14583
rect 20364 12986 20392 15302
rect 20456 14074 20484 15846
rect 20548 15502 20576 15914
rect 20536 15496 20588 15502
rect 20536 15438 20588 15444
rect 20548 14958 20576 15438
rect 20536 14952 20588 14958
rect 20640 14929 20668 16458
rect 20812 15632 20864 15638
rect 20812 15574 20864 15580
rect 20720 15360 20772 15366
rect 20720 15302 20772 15308
rect 20536 14894 20588 14900
rect 20626 14920 20682 14929
rect 20626 14855 20682 14864
rect 20640 14770 20668 14855
rect 20548 14742 20668 14770
rect 20444 14068 20496 14074
rect 20444 14010 20496 14016
rect 20548 13954 20576 14742
rect 20628 14612 20680 14618
rect 20732 14600 20760 15302
rect 20680 14572 20760 14600
rect 20628 14554 20680 14560
rect 20824 14498 20852 15574
rect 20904 14816 20956 14822
rect 20904 14758 20956 14764
rect 20640 14482 20852 14498
rect 20628 14476 20852 14482
rect 20680 14470 20852 14476
rect 20628 14418 20680 14424
rect 20916 14414 20944 14758
rect 20904 14408 20956 14414
rect 20904 14350 20956 14356
rect 20916 14074 20944 14350
rect 20904 14068 20956 14074
rect 20904 14010 20956 14016
rect 20456 13926 20576 13954
rect 20456 13530 20484 13926
rect 20536 13864 20588 13870
rect 20536 13806 20588 13812
rect 20444 13524 20496 13530
rect 20444 13466 20496 13472
rect 20548 13161 20576 13806
rect 21008 13802 21036 19314
rect 21192 18970 21220 19654
rect 21376 19174 21404 19994
rect 21468 19514 21496 20742
rect 21456 19508 21508 19514
rect 21456 19450 21508 19456
rect 21364 19168 21416 19174
rect 21364 19110 21416 19116
rect 21180 18964 21232 18970
rect 21180 18906 21232 18912
rect 21180 18624 21232 18630
rect 21180 18566 21232 18572
rect 21192 18086 21220 18566
rect 21180 18080 21232 18086
rect 21180 18022 21232 18028
rect 21192 17746 21220 18022
rect 21180 17740 21232 17746
rect 21180 17682 21232 17688
rect 21192 16794 21220 17682
rect 21180 16788 21232 16794
rect 21180 16730 21232 16736
rect 21270 16688 21326 16697
rect 21270 16623 21326 16632
rect 21284 16454 21312 16623
rect 21272 16448 21324 16454
rect 21272 16390 21324 16396
rect 21180 16108 21232 16114
rect 21180 16050 21232 16056
rect 21192 14550 21220 16050
rect 21284 16046 21312 16390
rect 21272 16040 21324 16046
rect 21272 15982 21324 15988
rect 21180 14544 21232 14550
rect 21180 14486 21232 14492
rect 21192 13938 21220 14486
rect 21180 13932 21232 13938
rect 21180 13874 21232 13880
rect 20996 13796 21048 13802
rect 20996 13738 21048 13744
rect 21008 13530 21036 13738
rect 20996 13524 21048 13530
rect 21180 13524 21232 13530
rect 21048 13484 21128 13512
rect 20996 13466 21048 13472
rect 20902 13424 20958 13433
rect 20902 13359 20958 13368
rect 20534 13152 20590 13161
rect 20534 13087 20590 13096
rect 20352 12980 20404 12986
rect 20352 12922 20404 12928
rect 20444 12912 20496 12918
rect 20272 12838 20392 12866
rect 20444 12854 20496 12860
rect 19996 12566 20116 12594
rect 20168 12640 20220 12646
rect 20168 12582 20220 12588
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19996 11268 20024 12566
rect 20074 12472 20130 12481
rect 20074 12407 20130 12416
rect 20088 12374 20116 12407
rect 20076 12368 20128 12374
rect 20076 12310 20128 12316
rect 20260 12232 20312 12238
rect 20260 12174 20312 12180
rect 19904 11240 20024 11268
rect 19904 10810 19932 11240
rect 19892 10804 19944 10810
rect 19892 10746 19944 10752
rect 20168 10804 20220 10810
rect 20168 10746 20220 10752
rect 20074 10704 20130 10713
rect 19984 10668 20036 10674
rect 20074 10639 20130 10648
rect 19984 10610 20036 10616
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19996 8922 20024 10610
rect 19628 8894 20024 8922
rect 19524 8628 19576 8634
rect 19524 8570 19576 8576
rect 19628 8378 19656 8894
rect 19984 8832 20036 8838
rect 19984 8774 20036 8780
rect 19536 8350 19656 8378
rect 19432 7540 19484 7546
rect 19432 7482 19484 7488
rect 19430 7032 19486 7041
rect 19340 6996 19392 7002
rect 19536 7018 19564 8350
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19800 8016 19852 8022
rect 19800 7958 19852 7964
rect 19812 7274 19840 7958
rect 19996 7954 20024 8774
rect 19984 7948 20036 7954
rect 19984 7890 20036 7896
rect 19800 7268 19852 7274
rect 19800 7210 19852 7216
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19486 6990 19564 7018
rect 19996 7002 20024 7890
rect 20088 7449 20116 10639
rect 20180 7585 20208 10746
rect 20166 7576 20222 7585
rect 20166 7511 20222 7520
rect 20168 7472 20220 7478
rect 20074 7440 20130 7449
rect 20168 7414 20220 7420
rect 20074 7375 20130 7384
rect 20076 7200 20128 7206
rect 20076 7142 20128 7148
rect 19984 6996 20036 7002
rect 19430 6967 19486 6976
rect 19340 6938 19392 6944
rect 19984 6938 20036 6944
rect 19248 6928 19300 6934
rect 19248 6870 19300 6876
rect 19156 6792 19208 6798
rect 19156 6734 19208 6740
rect 19168 6458 19196 6734
rect 19156 6452 19208 6458
rect 19156 6394 19208 6400
rect 19168 5846 19196 6394
rect 19260 5914 19288 6870
rect 19982 6760 20038 6769
rect 19982 6695 20038 6704
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19996 5914 20024 6695
rect 19248 5908 19300 5914
rect 19248 5850 19300 5856
rect 19984 5908 20036 5914
rect 19984 5850 20036 5856
rect 19156 5840 19208 5846
rect 20088 5817 20116 7142
rect 19156 5782 19208 5788
rect 20074 5808 20130 5817
rect 19800 5772 19852 5778
rect 20074 5743 20130 5752
rect 19800 5714 19852 5720
rect 19430 5536 19486 5545
rect 19430 5471 19486 5480
rect 18880 5160 18932 5166
rect 18878 5128 18880 5137
rect 18932 5128 18934 5137
rect 18878 5063 18934 5072
rect 18880 3936 18932 3942
rect 18880 3878 18932 3884
rect 18340 3602 18460 3618
rect 17224 3596 17276 3602
rect 17224 3538 17276 3544
rect 18328 3596 18460 3602
rect 18380 3590 18460 3596
rect 18328 3538 18380 3544
rect 17236 3194 17264 3538
rect 18326 3496 18382 3505
rect 18326 3431 18382 3440
rect 17592 3392 17644 3398
rect 17592 3334 17644 3340
rect 16672 3188 16724 3194
rect 16672 3130 16724 3136
rect 17224 3188 17276 3194
rect 17224 3130 17276 3136
rect 16684 2990 16712 3130
rect 16672 2984 16724 2990
rect 16672 2926 16724 2932
rect 17040 2848 17092 2854
rect 16210 2816 16266 2825
rect 16210 2751 16266 2760
rect 17038 2816 17040 2825
rect 17092 2816 17094 2825
rect 17038 2751 17094 2760
rect 16224 2650 16252 2751
rect 16212 2644 16264 2650
rect 16212 2586 16264 2592
rect 16856 2372 16908 2378
rect 16856 2314 16908 2320
rect 16132 1958 16252 1986
rect 16224 480 16252 1958
rect 16868 480 16896 2314
rect 17604 480 17632 3334
rect 17866 3224 17922 3233
rect 18340 3194 18368 3431
rect 18432 3194 18460 3590
rect 18708 3590 18828 3618
rect 17866 3159 17922 3168
rect 18328 3188 18380 3194
rect 17774 2952 17830 2961
rect 17774 2887 17776 2896
rect 17828 2887 17830 2896
rect 17776 2858 17828 2864
rect 17880 2650 17908 3159
rect 18328 3130 18380 3136
rect 18420 3188 18472 3194
rect 18420 3130 18472 3136
rect 18234 2680 18290 2689
rect 17868 2644 17920 2650
rect 18234 2615 18290 2624
rect 17868 2586 17920 2592
rect 18248 480 18276 2615
rect 18708 2514 18736 3590
rect 18892 3369 18920 3878
rect 18878 3360 18934 3369
rect 18878 3295 18934 3304
rect 19444 3194 19472 5471
rect 19812 5302 19840 5714
rect 19800 5296 19852 5302
rect 19798 5264 19800 5273
rect 19852 5264 19854 5273
rect 19798 5199 19854 5208
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19798 4720 19854 4729
rect 19798 4655 19800 4664
rect 19852 4655 19854 4664
rect 19800 4626 19852 4632
rect 19798 4448 19854 4457
rect 19798 4383 19854 4392
rect 19812 4078 19840 4383
rect 19982 4312 20038 4321
rect 19982 4247 20038 4256
rect 19800 4072 19852 4078
rect 19800 4014 19852 4020
rect 19996 3942 20024 4247
rect 20180 4146 20208 7414
rect 20272 7410 20300 12174
rect 20364 11626 20392 12838
rect 20352 11620 20404 11626
rect 20352 11562 20404 11568
rect 20350 11112 20406 11121
rect 20350 11047 20406 11056
rect 20364 9432 20392 11047
rect 20456 10266 20484 12854
rect 20640 12850 20760 12866
rect 20640 12844 20772 12850
rect 20640 12838 20720 12844
rect 20536 12640 20588 12646
rect 20536 12582 20588 12588
rect 20548 10810 20576 12582
rect 20640 11762 20668 12838
rect 20720 12786 20772 12792
rect 20812 12776 20864 12782
rect 20812 12718 20864 12724
rect 20720 12708 20772 12714
rect 20720 12650 20772 12656
rect 20732 12442 20760 12650
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 20720 12300 20772 12306
rect 20720 12242 20772 12248
rect 20732 11898 20760 12242
rect 20824 12170 20852 12718
rect 20916 12238 20944 13359
rect 21100 12714 21128 13484
rect 21180 13466 21232 13472
rect 21192 12918 21220 13466
rect 21180 12912 21232 12918
rect 21180 12854 21232 12860
rect 21088 12708 21140 12714
rect 21088 12650 21140 12656
rect 21180 12436 21232 12442
rect 21180 12378 21232 12384
rect 20996 12368 21048 12374
rect 20996 12310 21048 12316
rect 20904 12232 20956 12238
rect 20904 12174 20956 12180
rect 20812 12164 20864 12170
rect 20812 12106 20864 12112
rect 21008 11898 21036 12310
rect 21192 12102 21220 12378
rect 21284 12306 21312 15982
rect 21376 13841 21404 19110
rect 21560 17218 21588 21830
rect 21468 17190 21588 17218
rect 21362 13832 21418 13841
rect 21362 13767 21418 13776
rect 21364 13320 21416 13326
rect 21364 13262 21416 13268
rect 21376 12850 21404 13262
rect 21364 12844 21416 12850
rect 21364 12786 21416 12792
rect 21364 12708 21416 12714
rect 21364 12650 21416 12656
rect 21272 12300 21324 12306
rect 21272 12242 21324 12248
rect 21180 12096 21232 12102
rect 21180 12038 21232 12044
rect 20720 11892 20772 11898
rect 20720 11834 20772 11840
rect 20996 11892 21048 11898
rect 20996 11834 21048 11840
rect 20628 11756 20680 11762
rect 20628 11698 20680 11704
rect 20904 11688 20956 11694
rect 20904 11630 20956 11636
rect 20628 11620 20680 11626
rect 20628 11562 20680 11568
rect 20536 10804 20588 10810
rect 20536 10746 20588 10752
rect 20534 10568 20590 10577
rect 20534 10503 20590 10512
rect 20444 10260 20496 10266
rect 20444 10202 20496 10208
rect 20456 9586 20484 10202
rect 20444 9580 20496 9586
rect 20444 9522 20496 9528
rect 20364 9404 20484 9432
rect 20350 9344 20406 9353
rect 20350 9279 20406 9288
rect 20364 9178 20392 9279
rect 20352 9172 20404 9178
rect 20352 9114 20404 9120
rect 20456 8945 20484 9404
rect 20442 8936 20498 8945
rect 20442 8871 20498 8880
rect 20548 8838 20576 10503
rect 20352 8832 20404 8838
rect 20352 8774 20404 8780
rect 20536 8832 20588 8838
rect 20536 8774 20588 8780
rect 20364 7478 20392 8774
rect 20442 8664 20498 8673
rect 20442 8599 20498 8608
rect 20352 7472 20404 7478
rect 20352 7414 20404 7420
rect 20260 7404 20312 7410
rect 20260 7346 20312 7352
rect 20260 7200 20312 7206
rect 20260 7142 20312 7148
rect 20168 4140 20220 4146
rect 20168 4082 20220 4088
rect 19984 3936 20036 3942
rect 19984 3878 20036 3884
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19616 3528 19668 3534
rect 19616 3470 19668 3476
rect 19628 3233 19656 3470
rect 20166 3360 20222 3369
rect 20166 3295 20222 3304
rect 19614 3224 19670 3233
rect 19432 3188 19484 3194
rect 19614 3159 19670 3168
rect 19432 3130 19484 3136
rect 19246 3088 19302 3097
rect 19246 3023 19302 3032
rect 19260 2990 19288 3023
rect 19248 2984 19300 2990
rect 18786 2952 18842 2961
rect 19248 2926 19300 2932
rect 18786 2887 18842 2896
rect 18800 2650 18828 2887
rect 18878 2816 18934 2825
rect 18878 2751 18934 2760
rect 18788 2644 18840 2650
rect 18788 2586 18840 2592
rect 18696 2508 18748 2514
rect 18696 2450 18748 2456
rect 18892 480 18920 2751
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19524 2372 19576 2378
rect 19524 2314 19576 2320
rect 19536 480 19564 2314
rect 20180 1986 20208 3295
rect 20272 2650 20300 7142
rect 20350 7032 20406 7041
rect 20350 6967 20406 6976
rect 20364 3602 20392 6967
rect 20456 4078 20484 8599
rect 20536 8560 20588 8566
rect 20536 8502 20588 8508
rect 20548 7274 20576 8502
rect 20640 8378 20668 11562
rect 20812 11280 20864 11286
rect 20812 11222 20864 11228
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 20732 9654 20760 11086
rect 20824 10742 20852 11222
rect 20916 11218 20944 11630
rect 21192 11626 21220 12038
rect 21180 11620 21232 11626
rect 21180 11562 21232 11568
rect 20904 11212 20956 11218
rect 20904 11154 20956 11160
rect 21270 10840 21326 10849
rect 21270 10775 21326 10784
rect 21284 10742 21312 10775
rect 20812 10736 20864 10742
rect 20812 10678 20864 10684
rect 21272 10736 21324 10742
rect 21272 10678 21324 10684
rect 20824 10198 20852 10678
rect 21376 10674 21404 12650
rect 21468 11801 21496 17190
rect 21548 16176 21600 16182
rect 21548 16118 21600 16124
rect 21560 15638 21588 16118
rect 21548 15632 21600 15638
rect 21548 15574 21600 15580
rect 21546 13152 21602 13161
rect 21546 13087 21602 13096
rect 21560 12617 21588 13087
rect 21546 12608 21602 12617
rect 21546 12543 21602 12552
rect 21560 12374 21588 12543
rect 21548 12368 21600 12374
rect 21548 12310 21600 12316
rect 21548 12232 21600 12238
rect 21548 12174 21600 12180
rect 21454 11792 21510 11801
rect 21454 11727 21510 11736
rect 21560 11286 21588 12174
rect 21548 11280 21600 11286
rect 21548 11222 21600 11228
rect 21548 11008 21600 11014
rect 21548 10950 21600 10956
rect 21364 10668 21416 10674
rect 21364 10610 21416 10616
rect 20902 10568 20958 10577
rect 20902 10503 20904 10512
rect 20956 10503 20958 10512
rect 21362 10568 21418 10577
rect 21362 10503 21418 10512
rect 20904 10474 20956 10480
rect 20812 10192 20864 10198
rect 20812 10134 20864 10140
rect 20996 10056 21048 10062
rect 20996 9998 21048 10004
rect 20812 9920 20864 9926
rect 20812 9862 20864 9868
rect 20720 9648 20772 9654
rect 20720 9590 20772 9596
rect 20640 8350 20760 8378
rect 20628 8288 20680 8294
rect 20628 8230 20680 8236
rect 20640 7954 20668 8230
rect 20732 8022 20760 8350
rect 20720 8016 20772 8022
rect 20720 7958 20772 7964
rect 20628 7948 20680 7954
rect 20628 7890 20680 7896
rect 20720 7880 20772 7886
rect 20720 7822 20772 7828
rect 20732 7546 20760 7822
rect 20720 7540 20772 7546
rect 20720 7482 20772 7488
rect 20628 7472 20680 7478
rect 20628 7414 20680 7420
rect 20536 7268 20588 7274
rect 20536 7210 20588 7216
rect 20548 6866 20576 7210
rect 20536 6860 20588 6866
rect 20536 6802 20588 6808
rect 20536 6248 20588 6254
rect 20536 6190 20588 6196
rect 20548 5778 20576 6190
rect 20536 5772 20588 5778
rect 20536 5714 20588 5720
rect 20548 5370 20576 5714
rect 20536 5364 20588 5370
rect 20536 5306 20588 5312
rect 20640 5166 20668 7414
rect 20732 5778 20760 7482
rect 20824 7041 20852 9862
rect 21008 9722 21036 9998
rect 20996 9716 21048 9722
rect 20996 9658 21048 9664
rect 20996 9376 21048 9382
rect 20996 9318 21048 9324
rect 21008 9217 21036 9318
rect 20994 9208 21050 9217
rect 20994 9143 21050 9152
rect 21272 9036 21324 9042
rect 21272 8978 21324 8984
rect 21180 8832 21232 8838
rect 21180 8774 21232 8780
rect 20996 8424 21048 8430
rect 20996 8366 21048 8372
rect 20904 8288 20956 8294
rect 20904 8230 20956 8236
rect 20916 7886 20944 8230
rect 20904 7880 20956 7886
rect 20904 7822 20956 7828
rect 20904 7744 20956 7750
rect 20904 7686 20956 7692
rect 20916 7342 20944 7686
rect 20904 7336 20956 7342
rect 20904 7278 20956 7284
rect 21008 7290 21036 8366
rect 21192 8362 21220 8774
rect 21180 8356 21232 8362
rect 21180 8298 21232 8304
rect 21192 7750 21220 8298
rect 21284 7857 21312 8978
rect 21270 7848 21326 7857
rect 21270 7783 21326 7792
rect 21180 7744 21232 7750
rect 21180 7686 21232 7692
rect 21192 7410 21220 7686
rect 21180 7404 21232 7410
rect 21180 7346 21232 7352
rect 21008 7262 21220 7290
rect 20994 7168 21050 7177
rect 20994 7103 21050 7112
rect 20810 7032 20866 7041
rect 20810 6967 20866 6976
rect 20904 6860 20956 6866
rect 20904 6802 20956 6808
rect 20916 6458 20944 6802
rect 20904 6452 20956 6458
rect 20904 6394 20956 6400
rect 20812 6180 20864 6186
rect 20812 6122 20864 6128
rect 20824 5914 20852 6122
rect 20812 5908 20864 5914
rect 20812 5850 20864 5856
rect 20720 5772 20772 5778
rect 20720 5714 20772 5720
rect 21008 5234 21036 7103
rect 21088 6656 21140 6662
rect 21088 6598 21140 6604
rect 21100 5681 21128 6598
rect 21086 5672 21142 5681
rect 21086 5607 21142 5616
rect 20996 5228 21048 5234
rect 20996 5170 21048 5176
rect 20628 5160 20680 5166
rect 20628 5102 20680 5108
rect 20444 4072 20496 4078
rect 20444 4014 20496 4020
rect 21088 3936 21140 3942
rect 21088 3878 21140 3884
rect 20442 3768 20498 3777
rect 20442 3703 20444 3712
rect 20496 3703 20498 3712
rect 20444 3674 20496 3680
rect 20352 3596 20404 3602
rect 20352 3538 20404 3544
rect 20364 3194 20392 3538
rect 20352 3188 20404 3194
rect 20352 3130 20404 3136
rect 20456 2990 20484 3674
rect 21100 3505 21128 3878
rect 21192 3602 21220 7262
rect 21284 6866 21312 7783
rect 21272 6860 21324 6866
rect 21272 6802 21324 6808
rect 21376 6361 21404 10503
rect 21560 10198 21588 10950
rect 21548 10192 21600 10198
rect 21548 10134 21600 10140
rect 21560 9722 21588 10134
rect 21548 9716 21600 9722
rect 21548 9658 21600 9664
rect 21456 8832 21508 8838
rect 21456 8774 21508 8780
rect 21468 8401 21496 8774
rect 21454 8392 21510 8401
rect 21454 8327 21510 8336
rect 21362 6352 21418 6361
rect 21362 6287 21418 6296
rect 21548 5772 21600 5778
rect 21548 5714 21600 5720
rect 21560 5030 21588 5714
rect 21548 5024 21600 5030
rect 21548 4966 21600 4972
rect 21560 4185 21588 4966
rect 21546 4176 21602 4185
rect 21546 4111 21602 4120
rect 21652 3777 21680 22646
rect 21914 22607 21970 22616
rect 21732 21616 21784 21622
rect 21732 21558 21784 21564
rect 21744 19310 21772 21558
rect 21822 21040 21878 21049
rect 21822 20975 21878 20984
rect 21732 19304 21784 19310
rect 21732 19246 21784 19252
rect 21744 18902 21772 19246
rect 21732 18896 21784 18902
rect 21732 18838 21784 18844
rect 21730 18728 21786 18737
rect 21730 18663 21786 18672
rect 21744 17338 21772 18663
rect 21732 17332 21784 17338
rect 21732 17274 21784 17280
rect 21730 16552 21786 16561
rect 21730 16487 21786 16496
rect 21744 15638 21772 16487
rect 21836 15978 21864 20975
rect 21928 20942 21956 22607
rect 22008 21344 22060 21350
rect 22008 21286 22060 21292
rect 22020 21146 22048 21286
rect 22008 21140 22060 21146
rect 22008 21082 22060 21088
rect 21916 20936 21968 20942
rect 22112 20913 22140 23718
rect 22192 22160 22244 22166
rect 22192 22102 22244 22108
rect 22204 21146 22232 22102
rect 22192 21140 22244 21146
rect 22192 21082 22244 21088
rect 21916 20878 21968 20884
rect 22098 20904 22154 20913
rect 22008 20868 22060 20874
rect 22098 20839 22154 20848
rect 22008 20810 22060 20816
rect 22020 20074 22048 20810
rect 22204 20806 22232 21082
rect 22192 20800 22244 20806
rect 22192 20742 22244 20748
rect 22296 20369 22324 24686
rect 22376 22024 22428 22030
rect 22376 21966 22428 21972
rect 22282 20360 22338 20369
rect 22282 20295 22338 20304
rect 21928 20058 22140 20074
rect 21928 20052 22152 20058
rect 21928 20046 22100 20052
rect 21928 19174 21956 20046
rect 22100 19994 22152 20000
rect 22388 19718 22416 21966
rect 22480 21554 22508 24754
rect 22756 24410 22784 27520
rect 23294 27160 23350 27169
rect 23294 27095 23350 27104
rect 22744 24404 22796 24410
rect 22744 24346 22796 24352
rect 22560 24268 22612 24274
rect 22560 24210 22612 24216
rect 22572 23322 22600 24210
rect 23308 23798 23336 27095
rect 23492 24834 23520 27520
rect 24030 26616 24086 26625
rect 24030 26551 24086 26560
rect 23570 25936 23626 25945
rect 23570 25871 23626 25880
rect 23584 24886 23612 25871
rect 23400 24806 23520 24834
rect 23572 24880 23624 24886
rect 23572 24822 23624 24828
rect 23754 24848 23810 24857
rect 23400 24682 23428 24806
rect 23754 24783 23810 24792
rect 23388 24676 23440 24682
rect 23388 24618 23440 24624
rect 23296 23792 23348 23798
rect 23296 23734 23348 23740
rect 23112 23520 23164 23526
rect 23112 23462 23164 23468
rect 23480 23520 23532 23526
rect 23480 23462 23532 23468
rect 22560 23316 22612 23322
rect 22560 23258 22612 23264
rect 22836 23316 22888 23322
rect 22836 23258 22888 23264
rect 22468 21548 22520 21554
rect 22468 21490 22520 21496
rect 22560 21412 22612 21418
rect 22560 21354 22612 21360
rect 22744 21412 22796 21418
rect 22744 21354 22796 21360
rect 22572 21146 22600 21354
rect 22560 21140 22612 21146
rect 22560 21082 22612 21088
rect 22468 21004 22520 21010
rect 22468 20946 22520 20952
rect 22480 20262 22508 20946
rect 22572 20505 22600 21082
rect 22650 20904 22706 20913
rect 22650 20839 22706 20848
rect 22558 20496 22614 20505
rect 22558 20431 22614 20440
rect 22468 20256 22520 20262
rect 22468 20198 22520 20204
rect 22480 19922 22508 20198
rect 22572 19990 22600 20431
rect 22560 19984 22612 19990
rect 22560 19926 22612 19932
rect 22468 19916 22520 19922
rect 22468 19858 22520 19864
rect 22376 19712 22428 19718
rect 22376 19654 22428 19660
rect 22480 19242 22508 19858
rect 22008 19236 22060 19242
rect 22008 19178 22060 19184
rect 22468 19236 22520 19242
rect 22468 19178 22520 19184
rect 21916 19168 21968 19174
rect 21916 19110 21968 19116
rect 22020 18970 22048 19178
rect 22008 18964 22060 18970
rect 22008 18906 22060 18912
rect 22376 18896 22428 18902
rect 22376 18838 22428 18844
rect 22192 18828 22244 18834
rect 22192 18770 22244 18776
rect 22100 18692 22152 18698
rect 22100 18634 22152 18640
rect 22112 18222 22140 18634
rect 22100 18216 22152 18222
rect 22100 18158 22152 18164
rect 21916 16992 21968 16998
rect 21916 16934 21968 16940
rect 21928 16658 21956 16934
rect 21916 16652 21968 16658
rect 21916 16594 21968 16600
rect 21928 16266 21956 16594
rect 21928 16250 22140 16266
rect 21928 16244 22152 16250
rect 21928 16238 22100 16244
rect 21824 15972 21876 15978
rect 21824 15914 21876 15920
rect 21732 15632 21784 15638
rect 21730 15600 21732 15609
rect 21784 15600 21786 15609
rect 21730 15535 21786 15544
rect 21836 13530 21864 15914
rect 21928 14074 21956 16238
rect 22100 16186 22152 16192
rect 22008 15496 22060 15502
rect 22060 15444 22140 15450
rect 22008 15438 22140 15444
rect 22020 15422 22140 15438
rect 22204 15434 22232 18770
rect 22388 17882 22416 18838
rect 22468 18760 22520 18766
rect 22468 18702 22520 18708
rect 22480 18086 22508 18702
rect 22468 18080 22520 18086
rect 22468 18022 22520 18028
rect 22376 17876 22428 17882
rect 22376 17818 22428 17824
rect 22284 17536 22336 17542
rect 22284 17478 22336 17484
rect 22296 16726 22324 17478
rect 22388 17338 22416 17818
rect 22468 17536 22520 17542
rect 22468 17478 22520 17484
rect 22376 17332 22428 17338
rect 22376 17274 22428 17280
rect 22480 17105 22508 17478
rect 22466 17096 22522 17105
rect 22466 17031 22468 17040
rect 22520 17031 22522 17040
rect 22468 17002 22520 17008
rect 22480 16971 22508 17002
rect 22284 16720 22336 16726
rect 22284 16662 22336 16668
rect 22296 16561 22324 16662
rect 22282 16552 22338 16561
rect 22282 16487 22338 16496
rect 22112 14618 22140 15422
rect 22192 15428 22244 15434
rect 22192 15370 22244 15376
rect 22664 15314 22692 20839
rect 22756 20806 22784 21354
rect 22744 20800 22796 20806
rect 22744 20742 22796 20748
rect 22756 20398 22784 20742
rect 22744 20392 22796 20398
rect 22744 20334 22796 20340
rect 22744 20052 22796 20058
rect 22744 19994 22796 20000
rect 22204 15286 22692 15314
rect 22100 14612 22152 14618
rect 22100 14554 22152 14560
rect 21916 14068 21968 14074
rect 21916 14010 21968 14016
rect 21824 13524 21876 13530
rect 21824 13466 21876 13472
rect 21732 13184 21784 13190
rect 21732 13126 21784 13132
rect 21744 10062 21772 13126
rect 21928 12102 21956 14010
rect 22100 13728 22152 13734
rect 22100 13670 22152 13676
rect 22112 13530 22140 13670
rect 22100 13524 22152 13530
rect 22100 13466 22152 13472
rect 21916 12096 21968 12102
rect 21916 12038 21968 12044
rect 21928 11694 21956 12038
rect 21916 11688 21968 11694
rect 21822 11656 21878 11665
rect 21916 11630 21968 11636
rect 21822 11591 21878 11600
rect 21732 10056 21784 10062
rect 21732 9998 21784 10004
rect 21732 9036 21784 9042
rect 21732 8978 21784 8984
rect 21744 8430 21772 8978
rect 21732 8424 21784 8430
rect 21732 8366 21784 8372
rect 21836 5409 21864 11591
rect 21928 11098 21956 11630
rect 21928 11070 22140 11098
rect 22112 10810 22140 11070
rect 22204 10826 22232 15286
rect 22756 15201 22784 19994
rect 22848 18290 22876 23258
rect 23020 22092 23072 22098
rect 23020 22034 23072 22040
rect 23032 21350 23060 22034
rect 23020 21344 23072 21350
rect 23020 21286 23072 21292
rect 23032 21146 23060 21286
rect 23020 21140 23072 21146
rect 23020 21082 23072 21088
rect 22928 21072 22980 21078
rect 22928 21014 22980 21020
rect 22940 20346 22968 21014
rect 22940 20318 23060 20346
rect 22928 19984 22980 19990
rect 22928 19926 22980 19932
rect 22940 19786 22968 19926
rect 22928 19780 22980 19786
rect 22928 19722 22980 19728
rect 22940 18970 22968 19722
rect 22928 18964 22980 18970
rect 22928 18906 22980 18912
rect 23032 18465 23060 20318
rect 23124 19961 23152 23462
rect 23204 22024 23256 22030
rect 23204 21966 23256 21972
rect 23492 21978 23520 23462
rect 23662 22536 23718 22545
rect 23662 22471 23718 22480
rect 23216 21418 23244 21966
rect 23492 21950 23612 21978
rect 23480 21888 23532 21894
rect 23480 21830 23532 21836
rect 23492 21729 23520 21830
rect 23478 21720 23534 21729
rect 23478 21655 23534 21664
rect 23204 21412 23256 21418
rect 23204 21354 23256 21360
rect 23478 21312 23534 21321
rect 23478 21247 23534 21256
rect 23294 20904 23350 20913
rect 23294 20839 23350 20848
rect 23110 19952 23166 19961
rect 23110 19887 23166 19896
rect 23308 19854 23336 20839
rect 23388 20256 23440 20262
rect 23388 20198 23440 20204
rect 23400 19922 23428 20198
rect 23492 20058 23520 21247
rect 23480 20052 23532 20058
rect 23480 19994 23532 20000
rect 23478 19952 23534 19961
rect 23388 19916 23440 19922
rect 23478 19887 23534 19896
rect 23388 19858 23440 19864
rect 23296 19848 23348 19854
rect 23296 19790 23348 19796
rect 23308 19514 23336 19790
rect 23296 19508 23348 19514
rect 23296 19450 23348 19456
rect 23492 18970 23520 19887
rect 23480 18964 23532 18970
rect 23480 18906 23532 18912
rect 23018 18456 23074 18465
rect 23018 18391 23074 18400
rect 22836 18284 22888 18290
rect 22836 18226 22888 18232
rect 22834 17640 22890 17649
rect 22834 17575 22890 17584
rect 22848 15638 22876 17575
rect 22836 15632 22888 15638
rect 22836 15574 22888 15580
rect 22742 15192 22798 15201
rect 22848 15162 22876 15574
rect 22742 15127 22798 15136
rect 22836 15156 22888 15162
rect 22836 15098 22888 15104
rect 22560 15088 22612 15094
rect 22560 15030 22612 15036
rect 22284 13864 22336 13870
rect 22336 13812 22416 13818
rect 22284 13806 22416 13812
rect 22296 13790 22416 13806
rect 22284 13320 22336 13326
rect 22284 13262 22336 13268
rect 22296 12646 22324 13262
rect 22284 12640 22336 12646
rect 22284 12582 22336 12588
rect 22296 11626 22324 12582
rect 22284 11620 22336 11626
rect 22284 11562 22336 11568
rect 22296 11354 22324 11562
rect 22284 11348 22336 11354
rect 22284 11290 22336 11296
rect 22100 10804 22152 10810
rect 22204 10798 22324 10826
rect 22100 10746 22152 10752
rect 22008 10668 22060 10674
rect 22112 10656 22140 10746
rect 22112 10628 22232 10656
rect 22008 10610 22060 10616
rect 21916 9376 21968 9382
rect 21916 9318 21968 9324
rect 21928 9178 21956 9318
rect 21916 9172 21968 9178
rect 21916 9114 21968 9120
rect 21916 7948 21968 7954
rect 21916 7890 21968 7896
rect 21928 7546 21956 7890
rect 21916 7540 21968 7546
rect 21916 7482 21968 7488
rect 21914 7304 21970 7313
rect 21914 7239 21970 7248
rect 21928 6458 21956 7239
rect 22020 6905 22048 10610
rect 22100 10532 22152 10538
rect 22100 10474 22152 10480
rect 22112 10266 22140 10474
rect 22100 10260 22152 10266
rect 22100 10202 22152 10208
rect 22100 9648 22152 9654
rect 22100 9590 22152 9596
rect 22006 6896 22062 6905
rect 22112 6866 22140 9590
rect 22204 9042 22232 10628
rect 22192 9036 22244 9042
rect 22192 8978 22244 8984
rect 22204 8566 22232 8978
rect 22192 8560 22244 8566
rect 22192 8502 22244 8508
rect 22006 6831 22062 6840
rect 22100 6860 22152 6866
rect 22100 6802 22152 6808
rect 22296 6798 22324 10798
rect 22284 6792 22336 6798
rect 22284 6734 22336 6740
rect 22296 6458 22324 6734
rect 21916 6452 21968 6458
rect 21916 6394 21968 6400
rect 22284 6452 22336 6458
rect 22284 6394 22336 6400
rect 22388 5914 22416 13790
rect 22468 13796 22520 13802
rect 22468 13738 22520 13744
rect 22480 13326 22508 13738
rect 22468 13320 22520 13326
rect 22468 13262 22520 13268
rect 22572 11665 22600 15030
rect 22664 13462 22692 13493
rect 22652 13456 22704 13462
rect 22650 13424 22652 13433
rect 22704 13424 22706 13433
rect 22650 13359 22706 13368
rect 22664 12986 22692 13359
rect 22652 12980 22704 12986
rect 22652 12922 22704 12928
rect 22744 12300 22796 12306
rect 22744 12242 22796 12248
rect 22756 11898 22784 12242
rect 22744 11892 22796 11898
rect 22744 11834 22796 11840
rect 22558 11656 22614 11665
rect 22558 11591 22614 11600
rect 22756 11354 22784 11834
rect 22926 11792 22982 11801
rect 22926 11727 22982 11736
rect 22744 11348 22796 11354
rect 22744 11290 22796 11296
rect 22756 11082 22784 11290
rect 22744 11076 22796 11082
rect 22744 11018 22796 11024
rect 22836 10124 22888 10130
rect 22836 10066 22888 10072
rect 22560 9920 22612 9926
rect 22560 9862 22612 9868
rect 22572 9586 22600 9862
rect 22848 9722 22876 10066
rect 22836 9716 22888 9722
rect 22836 9658 22888 9664
rect 22560 9580 22612 9586
rect 22560 9522 22612 9528
rect 22572 9353 22600 9522
rect 22652 9444 22704 9450
rect 22652 9386 22704 9392
rect 22558 9344 22614 9353
rect 22558 9279 22614 9288
rect 22664 9178 22692 9386
rect 22652 9172 22704 9178
rect 22652 9114 22704 9120
rect 22558 9072 22614 9081
rect 22468 9036 22520 9042
rect 22558 9007 22614 9016
rect 22468 8978 22520 8984
rect 22480 8634 22508 8978
rect 22468 8628 22520 8634
rect 22468 8570 22520 8576
rect 22480 8090 22508 8570
rect 22468 8084 22520 8090
rect 22468 8026 22520 8032
rect 22466 6216 22522 6225
rect 22466 6151 22522 6160
rect 22100 5908 22152 5914
rect 22100 5850 22152 5856
rect 22376 5908 22428 5914
rect 22376 5850 22428 5856
rect 21822 5400 21878 5409
rect 22112 5370 22140 5850
rect 21822 5335 21878 5344
rect 22100 5364 22152 5370
rect 22100 5306 22152 5312
rect 22282 5128 22338 5137
rect 22282 5063 22284 5072
rect 22336 5063 22338 5072
rect 22284 5034 22336 5040
rect 21824 4684 21876 4690
rect 21824 4626 21876 4632
rect 21836 4282 21864 4626
rect 22100 4480 22152 4486
rect 22100 4422 22152 4428
rect 21824 4276 21876 4282
rect 21824 4218 21876 4224
rect 21836 3942 21864 4218
rect 21824 3936 21876 3942
rect 21824 3878 21876 3884
rect 21638 3768 21694 3777
rect 21638 3703 21694 3712
rect 21180 3596 21232 3602
rect 21180 3538 21232 3544
rect 22008 3596 22060 3602
rect 22008 3538 22060 3544
rect 21086 3496 21142 3505
rect 21086 3431 21142 3440
rect 21088 3392 21140 3398
rect 21088 3334 21140 3340
rect 21100 3097 21128 3334
rect 21192 3194 21220 3538
rect 21180 3188 21232 3194
rect 21180 3130 21232 3136
rect 21086 3088 21142 3097
rect 21086 3023 21142 3032
rect 20444 2984 20496 2990
rect 20444 2926 20496 2932
rect 21546 2952 21602 2961
rect 20628 2916 20680 2922
rect 22020 2922 22048 3538
rect 21546 2887 21602 2896
rect 22008 2916 22060 2922
rect 20628 2858 20680 2864
rect 20260 2644 20312 2650
rect 20260 2586 20312 2592
rect 20640 2553 20668 2858
rect 20626 2544 20682 2553
rect 20626 2479 20682 2488
rect 20904 2372 20956 2378
rect 20904 2314 20956 2320
rect 20180 1958 20300 1986
rect 20272 480 20300 1958
rect 20916 480 20944 2314
rect 21560 480 21588 2887
rect 22008 2858 22060 2864
rect 22112 2802 22140 4422
rect 22192 3936 22244 3942
rect 22480 3924 22508 6151
rect 22572 4078 22600 9007
rect 22652 5024 22704 5030
rect 22652 4966 22704 4972
rect 22664 4593 22692 4966
rect 22650 4584 22706 4593
rect 22650 4519 22706 4528
rect 22560 4072 22612 4078
rect 22560 4014 22612 4020
rect 22652 3936 22704 3942
rect 22480 3896 22600 3924
rect 22192 3878 22244 3884
rect 22204 2922 22232 3878
rect 22192 2916 22244 2922
rect 22192 2858 22244 2864
rect 22112 2774 22232 2802
rect 21916 2304 21968 2310
rect 21916 2246 21968 2252
rect 21928 1601 21956 2246
rect 21914 1592 21970 1601
rect 21914 1527 21970 1536
rect 22204 480 22232 2774
rect 22572 2650 22600 3896
rect 22652 3878 22704 3884
rect 22664 3641 22692 3878
rect 22650 3632 22706 3641
rect 22940 3602 22968 11727
rect 23032 4826 23060 18391
rect 23492 18358 23520 18906
rect 23480 18352 23532 18358
rect 23480 18294 23532 18300
rect 23480 18148 23532 18154
rect 23480 18090 23532 18096
rect 23112 16992 23164 16998
rect 23112 16934 23164 16940
rect 23296 16992 23348 16998
rect 23296 16934 23348 16940
rect 23124 16454 23152 16934
rect 23112 16448 23164 16454
rect 23112 16390 23164 16396
rect 23124 15502 23152 16390
rect 23308 16250 23336 16934
rect 23492 16250 23520 18090
rect 23584 17882 23612 21950
rect 23676 19281 23704 22471
rect 23768 21486 23796 24783
rect 23940 23588 23992 23594
rect 23940 23530 23992 23536
rect 23848 23520 23900 23526
rect 23848 23462 23900 23468
rect 23756 21480 23808 21486
rect 23756 21422 23808 21428
rect 23860 21078 23888 23462
rect 23848 21072 23900 21078
rect 23848 21014 23900 21020
rect 23952 20754 23980 23530
rect 24044 21706 24072 26551
rect 24136 24410 24164 27520
rect 24596 26314 24624 27639
rect 24766 27520 24822 28000
rect 25502 27520 25558 28000
rect 26146 27520 26202 28000
rect 26882 27520 26938 28000
rect 27526 27520 27582 28000
rect 24584 26308 24636 26314
rect 24584 26250 24636 26256
rect 24780 25514 24808 27520
rect 24688 25486 24808 25514
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24124 24404 24176 24410
rect 24124 24346 24176 24352
rect 24216 24268 24268 24274
rect 24216 24210 24268 24216
rect 24228 23662 24256 24210
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24688 23866 24716 25486
rect 24766 25392 24822 25401
rect 24766 25327 24768 25336
rect 24820 25327 24822 25336
rect 24768 25298 24820 25304
rect 24860 24268 24912 24274
rect 24860 24210 24912 24216
rect 24676 23860 24728 23866
rect 24676 23802 24728 23808
rect 24216 23656 24268 23662
rect 24214 23624 24216 23633
rect 24268 23624 24270 23633
rect 24214 23559 24270 23568
rect 24674 23624 24730 23633
rect 24674 23559 24730 23568
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24688 22778 24716 23559
rect 24872 23526 24900 24210
rect 24950 23896 25006 23905
rect 24950 23831 24952 23840
rect 25004 23831 25006 23840
rect 24952 23802 25004 23808
rect 25516 23633 25544 27520
rect 25502 23624 25558 23633
rect 25502 23559 25558 23568
rect 24860 23520 24912 23526
rect 24766 23488 24822 23497
rect 26160 23497 26188 27520
rect 26896 24410 26924 27520
rect 26884 24404 26936 24410
rect 26884 24346 26936 24352
rect 27540 23905 27568 27520
rect 27526 23896 27582 23905
rect 27526 23831 27582 23840
rect 24860 23462 24912 23468
rect 26146 23488 26202 23497
rect 24766 23423 24822 23432
rect 26146 23423 26202 23432
rect 24780 23322 24808 23423
rect 24768 23316 24820 23322
rect 24768 23258 24820 23264
rect 24860 23180 24912 23186
rect 24860 23122 24912 23128
rect 24676 22772 24728 22778
rect 24676 22714 24728 22720
rect 24872 22438 24900 23122
rect 24216 22432 24268 22438
rect 24216 22374 24268 22380
rect 24860 22432 24912 22438
rect 24860 22374 24912 22380
rect 25780 22432 25832 22438
rect 25780 22374 25832 22380
rect 24044 21678 24164 21706
rect 24030 21584 24086 21593
rect 24030 21519 24086 21528
rect 23768 20726 23980 20754
rect 23662 19272 23718 19281
rect 23662 19207 23718 19216
rect 23572 17876 23624 17882
rect 23572 17818 23624 17824
rect 23768 17762 23796 20726
rect 23940 20392 23992 20398
rect 23940 20334 23992 20340
rect 23848 19712 23900 19718
rect 23848 19654 23900 19660
rect 23860 19242 23888 19654
rect 23952 19446 23980 20334
rect 23940 19440 23992 19446
rect 23940 19382 23992 19388
rect 23848 19236 23900 19242
rect 23848 19178 23900 19184
rect 24044 18306 24072 21519
rect 24136 21434 24164 21678
rect 24228 21554 24256 22374
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24216 21548 24268 21554
rect 24216 21490 24268 21496
rect 24676 21480 24728 21486
rect 24136 21406 24256 21434
rect 24676 21422 24728 21428
rect 24228 21185 24256 21406
rect 24214 21176 24270 21185
rect 24214 21111 24270 21120
rect 24124 20256 24176 20262
rect 24124 20198 24176 20204
rect 24136 19922 24164 20198
rect 24124 19916 24176 19922
rect 24124 19858 24176 19864
rect 24136 19718 24164 19858
rect 24124 19712 24176 19718
rect 24124 19654 24176 19660
rect 24136 19514 24164 19654
rect 24124 19508 24176 19514
rect 24124 19450 24176 19456
rect 24228 19394 24256 21111
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24688 19786 24716 21422
rect 24860 20936 24912 20942
rect 24766 20904 24822 20913
rect 24822 20884 24860 20890
rect 24822 20878 24912 20884
rect 24822 20862 24900 20878
rect 24766 20839 24822 20848
rect 25504 20528 25556 20534
rect 25502 20496 25504 20505
rect 25556 20496 25558 20505
rect 25502 20431 25558 20440
rect 24860 19984 24912 19990
rect 24860 19926 24912 19932
rect 24768 19848 24820 19854
rect 24768 19790 24820 19796
rect 24676 19780 24728 19786
rect 24676 19722 24728 19728
rect 24674 19680 24730 19689
rect 24289 19612 24585 19632
rect 24674 19615 24730 19624
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24582 19408 24638 19417
rect 24228 19366 24440 19394
rect 24122 19000 24178 19009
rect 24122 18935 24178 18944
rect 23952 18278 24072 18306
rect 23848 17876 23900 17882
rect 23848 17818 23900 17824
rect 23584 17734 23796 17762
rect 23296 16244 23348 16250
rect 23296 16186 23348 16192
rect 23480 16244 23532 16250
rect 23480 16186 23532 16192
rect 23202 16144 23258 16153
rect 23202 16079 23258 16088
rect 23216 15858 23244 16079
rect 23308 16046 23336 16186
rect 23296 16040 23348 16046
rect 23296 15982 23348 15988
rect 23584 15960 23612 17734
rect 23664 17672 23716 17678
rect 23664 17614 23716 17620
rect 23676 17134 23704 17614
rect 23756 17536 23808 17542
rect 23756 17478 23808 17484
rect 23664 17128 23716 17134
rect 23664 17070 23716 17076
rect 23676 16998 23704 17070
rect 23768 17066 23796 17478
rect 23756 17060 23808 17066
rect 23756 17002 23808 17008
rect 23664 16992 23716 16998
rect 23664 16934 23716 16940
rect 23676 16794 23704 16934
rect 23664 16788 23716 16794
rect 23664 16730 23716 16736
rect 23860 16153 23888 17818
rect 23952 17513 23980 18278
rect 24032 18216 24084 18222
rect 24032 18158 24084 18164
rect 23938 17504 23994 17513
rect 23938 17439 23994 17448
rect 23846 16144 23902 16153
rect 24044 16130 24072 18158
rect 24136 17377 24164 18935
rect 24216 18828 24268 18834
rect 24216 18770 24268 18776
rect 24228 18426 24256 18770
rect 24412 18737 24440 19366
rect 24582 19343 24638 19352
rect 24492 19236 24544 19242
rect 24492 19178 24544 19184
rect 24504 18902 24532 19178
rect 24492 18896 24544 18902
rect 24492 18838 24544 18844
rect 24596 18766 24624 19343
rect 24584 18760 24636 18766
rect 24398 18728 24454 18737
rect 24584 18702 24636 18708
rect 24398 18663 24454 18672
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24216 18420 24268 18426
rect 24216 18362 24268 18368
rect 24688 18222 24716 19615
rect 24780 18698 24808 19790
rect 24872 19242 24900 19926
rect 24860 19236 24912 19242
rect 24860 19178 24912 19184
rect 24768 18692 24820 18698
rect 24768 18634 24820 18640
rect 24872 18426 24900 19178
rect 24952 18896 25004 18902
rect 24952 18838 25004 18844
rect 24860 18420 24912 18426
rect 24860 18362 24912 18368
rect 24964 18290 24992 18838
rect 25044 18760 25096 18766
rect 25044 18702 25096 18708
rect 24952 18284 25004 18290
rect 24952 18226 25004 18232
rect 24676 18216 24728 18222
rect 24676 18158 24728 18164
rect 24768 18148 24820 18154
rect 24768 18090 24820 18096
rect 24216 17740 24268 17746
rect 24216 17682 24268 17688
rect 24122 17368 24178 17377
rect 24122 17303 24178 17312
rect 24228 16794 24256 17682
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24676 16992 24728 16998
rect 24676 16934 24728 16940
rect 24216 16788 24268 16794
rect 24216 16730 24268 16736
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24044 16102 24164 16130
rect 23846 16079 23902 16088
rect 24032 16040 24084 16046
rect 24032 15982 24084 15988
rect 23400 15932 23612 15960
rect 23216 15830 23336 15858
rect 23112 15496 23164 15502
rect 23112 15438 23164 15444
rect 23124 14618 23152 15438
rect 23112 14612 23164 14618
rect 23112 14554 23164 14560
rect 23112 14068 23164 14074
rect 23112 14010 23164 14016
rect 23124 13530 23152 14010
rect 23204 14000 23256 14006
rect 23204 13942 23256 13948
rect 23112 13524 23164 13530
rect 23112 13466 23164 13472
rect 23112 13388 23164 13394
rect 23112 13330 23164 13336
rect 23124 12646 23152 13330
rect 23112 12640 23164 12646
rect 23112 12582 23164 12588
rect 23124 12481 23152 12582
rect 23110 12472 23166 12481
rect 23110 12407 23166 12416
rect 23112 10056 23164 10062
rect 23112 9998 23164 10004
rect 23124 9450 23152 9998
rect 23112 9444 23164 9450
rect 23112 9386 23164 9392
rect 23124 9042 23152 9386
rect 23112 9036 23164 9042
rect 23112 8978 23164 8984
rect 23216 7562 23244 13942
rect 23308 10266 23336 15830
rect 23400 15706 23428 15932
rect 24044 15706 24072 15982
rect 23388 15700 23440 15706
rect 23388 15642 23440 15648
rect 24032 15700 24084 15706
rect 24032 15642 24084 15648
rect 23400 15094 23428 15642
rect 23662 15464 23718 15473
rect 24044 15450 24072 15642
rect 23662 15399 23718 15408
rect 23860 15422 24072 15450
rect 23388 15088 23440 15094
rect 23388 15030 23440 15036
rect 23480 14816 23532 14822
rect 23480 14758 23532 14764
rect 23492 14278 23520 14758
rect 23480 14272 23532 14278
rect 23480 14214 23532 14220
rect 23492 13258 23520 14214
rect 23572 14000 23624 14006
rect 23572 13942 23624 13948
rect 23480 13252 23532 13258
rect 23480 13194 23532 13200
rect 23584 11898 23612 13942
rect 23676 13546 23704 15399
rect 23756 15088 23808 15094
rect 23756 15030 23808 15036
rect 23768 13870 23796 15030
rect 23860 14482 23888 15422
rect 23940 15360 23992 15366
rect 23940 15302 23992 15308
rect 23952 14958 23980 15302
rect 24032 15156 24084 15162
rect 24032 15098 24084 15104
rect 23940 14952 23992 14958
rect 23940 14894 23992 14900
rect 23848 14476 23900 14482
rect 23848 14418 23900 14424
rect 23860 13938 23888 14418
rect 23952 14278 23980 14894
rect 24044 14550 24072 15098
rect 24032 14544 24084 14550
rect 24032 14486 24084 14492
rect 23940 14272 23992 14278
rect 23940 14214 23992 14220
rect 23952 13938 23980 14214
rect 24044 14074 24072 14486
rect 24032 14068 24084 14074
rect 24032 14010 24084 14016
rect 23848 13932 23900 13938
rect 23848 13874 23900 13880
rect 23940 13932 23992 13938
rect 23940 13874 23992 13880
rect 23756 13864 23808 13870
rect 23756 13806 23808 13812
rect 23676 13518 24072 13546
rect 23848 13456 23900 13462
rect 23848 13398 23900 13404
rect 23756 12912 23808 12918
rect 23756 12854 23808 12860
rect 23664 12096 23716 12102
rect 23664 12038 23716 12044
rect 23572 11892 23624 11898
rect 23572 11834 23624 11840
rect 23676 11014 23704 12038
rect 23664 11008 23716 11014
rect 23664 10950 23716 10956
rect 23676 10810 23704 10950
rect 23664 10804 23716 10810
rect 23664 10746 23716 10752
rect 23676 10606 23704 10746
rect 23664 10600 23716 10606
rect 23664 10542 23716 10548
rect 23664 10464 23716 10470
rect 23664 10406 23716 10412
rect 23296 10260 23348 10266
rect 23296 10202 23348 10208
rect 23308 9722 23336 10202
rect 23676 10198 23704 10406
rect 23768 10198 23796 12854
rect 23860 12442 23888 13398
rect 24044 13274 24072 13518
rect 24136 13394 24164 16102
rect 24688 16046 24716 16934
rect 24780 16794 24808 18090
rect 24768 16788 24820 16794
rect 24768 16730 24820 16736
rect 24860 16720 24912 16726
rect 24860 16662 24912 16668
rect 24676 16040 24728 16046
rect 24676 15982 24728 15988
rect 24676 15904 24728 15910
rect 24676 15846 24728 15852
rect 24688 15620 24716 15846
rect 24768 15632 24820 15638
rect 24688 15592 24768 15620
rect 24216 15360 24268 15366
rect 24216 15302 24268 15308
rect 24228 15026 24256 15302
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24216 15020 24268 15026
rect 24216 14962 24268 14968
rect 24228 14618 24256 14962
rect 24688 14822 24716 15592
rect 24872 15620 24900 16662
rect 25056 16017 25084 18702
rect 25320 18284 25372 18290
rect 25320 18226 25372 18232
rect 25332 17882 25360 18226
rect 25320 17876 25372 17882
rect 25320 17818 25372 17824
rect 25412 16652 25464 16658
rect 25412 16594 25464 16600
rect 25320 16584 25372 16590
rect 25320 16526 25372 16532
rect 25042 16008 25098 16017
rect 25332 15994 25360 16526
rect 25424 16250 25452 16594
rect 25412 16244 25464 16250
rect 25412 16186 25464 16192
rect 25410 16008 25466 16017
rect 25332 15966 25410 15994
rect 25042 15943 25098 15952
rect 25410 15943 25466 15952
rect 24820 15592 24900 15620
rect 24768 15574 24820 15580
rect 24860 15496 24912 15502
rect 24860 15438 24912 15444
rect 24872 15178 24900 15438
rect 24780 15162 24900 15178
rect 24768 15156 24900 15162
rect 24820 15150 24900 15156
rect 24768 15098 24820 15104
rect 24676 14816 24728 14822
rect 24676 14758 24728 14764
rect 24216 14612 24268 14618
rect 24216 14554 24268 14560
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24400 13864 24452 13870
rect 24400 13806 24452 13812
rect 24412 13530 24440 13806
rect 24400 13524 24452 13530
rect 24400 13466 24452 13472
rect 24124 13388 24176 13394
rect 24124 13330 24176 13336
rect 24044 13246 24164 13274
rect 24030 13152 24086 13161
rect 24030 13087 24086 13096
rect 23848 12436 23900 12442
rect 23848 12378 23900 12384
rect 23940 11688 23992 11694
rect 23940 11630 23992 11636
rect 23952 11218 23980 11630
rect 23940 11212 23992 11218
rect 23940 11154 23992 11160
rect 23952 10810 23980 11154
rect 23940 10804 23992 10810
rect 23940 10746 23992 10752
rect 23664 10192 23716 10198
rect 23662 10160 23664 10169
rect 23756 10192 23808 10198
rect 23716 10160 23718 10169
rect 23756 10134 23808 10140
rect 23662 10095 23718 10104
rect 23940 10056 23992 10062
rect 23570 10024 23626 10033
rect 23940 9998 23992 10004
rect 23570 9959 23626 9968
rect 23296 9716 23348 9722
rect 23296 9658 23348 9664
rect 23386 9480 23442 9489
rect 23386 9415 23442 9424
rect 23124 7534 23244 7562
rect 23020 4820 23072 4826
rect 23020 4762 23072 4768
rect 23032 4146 23060 4762
rect 23020 4140 23072 4146
rect 23020 4082 23072 4088
rect 22650 3567 22706 3576
rect 22928 3596 22980 3602
rect 22928 3538 22980 3544
rect 22926 3496 22982 3505
rect 22926 3431 22982 3440
rect 22560 2644 22612 2650
rect 22560 2586 22612 2592
rect 22836 2508 22888 2514
rect 22836 2450 22888 2456
rect 22848 1737 22876 2450
rect 22834 1728 22890 1737
rect 22834 1663 22890 1672
rect 22940 480 22968 3431
rect 23124 3194 23152 7534
rect 23204 7472 23256 7478
rect 23204 7414 23256 7420
rect 23216 7342 23244 7414
rect 23400 7410 23428 9415
rect 23480 9376 23532 9382
rect 23480 9318 23532 9324
rect 23492 9081 23520 9318
rect 23478 9072 23534 9081
rect 23478 9007 23534 9016
rect 23388 7404 23440 7410
rect 23388 7346 23440 7352
rect 23204 7336 23256 7342
rect 23204 7278 23256 7284
rect 23216 7002 23244 7278
rect 23204 6996 23256 7002
rect 23204 6938 23256 6944
rect 23294 6896 23350 6905
rect 23294 6831 23296 6840
rect 23348 6831 23350 6840
rect 23296 6802 23348 6808
rect 23308 6458 23336 6802
rect 23480 6656 23532 6662
rect 23480 6598 23532 6604
rect 23296 6452 23348 6458
rect 23296 6394 23348 6400
rect 23492 5030 23520 6598
rect 23584 6474 23612 9959
rect 23952 9586 23980 9998
rect 23940 9580 23992 9586
rect 23940 9522 23992 9528
rect 23756 9172 23808 9178
rect 23756 9114 23808 9120
rect 23664 8492 23716 8498
rect 23664 8434 23716 8440
rect 23676 7954 23704 8434
rect 23768 8430 23796 9114
rect 23846 9072 23902 9081
rect 23846 9007 23902 9016
rect 23756 8424 23808 8430
rect 23756 8366 23808 8372
rect 23768 8090 23796 8366
rect 23756 8084 23808 8090
rect 23756 8026 23808 8032
rect 23664 7948 23716 7954
rect 23664 7890 23716 7896
rect 23676 7546 23704 7890
rect 23664 7540 23716 7546
rect 23664 7482 23716 7488
rect 23584 6446 23704 6474
rect 23572 6384 23624 6390
rect 23572 6326 23624 6332
rect 23584 6225 23612 6326
rect 23570 6216 23626 6225
rect 23570 6151 23626 6160
rect 23572 5840 23624 5846
rect 23572 5782 23624 5788
rect 23584 5302 23612 5782
rect 23572 5296 23624 5302
rect 23572 5238 23624 5244
rect 23480 5024 23532 5030
rect 23480 4966 23532 4972
rect 23676 4842 23704 6446
rect 23756 6452 23808 6458
rect 23756 6394 23808 6400
rect 23584 4814 23704 4842
rect 23584 4321 23612 4814
rect 23662 4720 23718 4729
rect 23662 4655 23664 4664
rect 23716 4655 23718 4664
rect 23664 4626 23716 4632
rect 23570 4312 23626 4321
rect 23676 4282 23704 4626
rect 23570 4247 23626 4256
rect 23664 4276 23716 4282
rect 23664 4218 23716 4224
rect 23204 4140 23256 4146
rect 23204 4082 23256 4088
rect 23112 3188 23164 3194
rect 23112 3130 23164 3136
rect 23124 2990 23152 3130
rect 23112 2984 23164 2990
rect 23112 2926 23164 2932
rect 23018 2680 23074 2689
rect 23018 2615 23020 2624
rect 23072 2615 23074 2624
rect 23020 2586 23072 2592
rect 23216 1873 23244 4082
rect 23768 4078 23796 6394
rect 23860 5545 23888 9007
rect 23952 7993 23980 9522
rect 24044 9518 24072 13087
rect 24136 10674 24164 13246
rect 24216 13184 24268 13190
rect 24216 13126 24268 13132
rect 24228 12850 24256 13126
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24216 12844 24268 12850
rect 24216 12786 24268 12792
rect 24308 12708 24360 12714
rect 24308 12650 24360 12656
rect 24320 12170 24348 12650
rect 24308 12164 24360 12170
rect 24308 12106 24360 12112
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24688 11937 24716 14758
rect 24860 13388 24912 13394
rect 24860 13330 24912 13336
rect 24872 12986 24900 13330
rect 24860 12980 24912 12986
rect 24860 12922 24912 12928
rect 25056 12646 25084 15943
rect 25424 15706 25452 15943
rect 25412 15700 25464 15706
rect 25412 15642 25464 15648
rect 25424 15162 25452 15642
rect 25412 15156 25464 15162
rect 25412 15098 25464 15104
rect 25228 14816 25280 14822
rect 25228 14758 25280 14764
rect 25240 13462 25268 14758
rect 25228 13456 25280 13462
rect 25228 13398 25280 13404
rect 25688 13456 25740 13462
rect 25688 13398 25740 13404
rect 25044 12640 25096 12646
rect 25044 12582 25096 12588
rect 25240 12442 25268 13398
rect 25700 12986 25728 13398
rect 25688 12980 25740 12986
rect 25688 12922 25740 12928
rect 25228 12436 25280 12442
rect 25228 12378 25280 12384
rect 25792 12209 25820 22374
rect 25870 13832 25926 13841
rect 25870 13767 25926 13776
rect 25778 12200 25834 12209
rect 25778 12135 25834 12144
rect 24860 12096 24912 12102
rect 24860 12038 24912 12044
rect 25136 12096 25188 12102
rect 25136 12038 25188 12044
rect 24674 11928 24730 11937
rect 24872 11898 24900 12038
rect 24674 11863 24730 11872
rect 24860 11892 24912 11898
rect 24860 11834 24912 11840
rect 25148 11393 25176 12038
rect 25134 11384 25190 11393
rect 25134 11319 25190 11328
rect 24952 11076 25004 11082
rect 24952 11018 25004 11024
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24676 10736 24728 10742
rect 24676 10678 24728 10684
rect 24124 10668 24176 10674
rect 24124 10610 24176 10616
rect 24688 10198 24716 10678
rect 24768 10464 24820 10470
rect 24768 10406 24820 10412
rect 24216 10192 24268 10198
rect 24216 10134 24268 10140
rect 24676 10192 24728 10198
rect 24676 10134 24728 10140
rect 24124 9920 24176 9926
rect 24124 9862 24176 9868
rect 24032 9512 24084 9518
rect 24032 9454 24084 9460
rect 24044 9178 24072 9454
rect 24032 9172 24084 9178
rect 24032 9114 24084 9120
rect 24136 8650 24164 9862
rect 24228 9722 24256 10134
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24216 9716 24268 9722
rect 24216 9658 24268 9664
rect 24582 9616 24638 9625
rect 24582 9551 24638 9560
rect 24596 8922 24624 9551
rect 24688 9178 24716 10134
rect 24676 9172 24728 9178
rect 24676 9114 24728 9120
rect 24596 8894 24716 8922
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24044 8622 24164 8650
rect 23938 7984 23994 7993
rect 23938 7919 23994 7928
rect 23940 6792 23992 6798
rect 23940 6734 23992 6740
rect 23952 6254 23980 6734
rect 23940 6248 23992 6254
rect 23940 6190 23992 6196
rect 23952 5778 23980 6190
rect 23940 5772 23992 5778
rect 23940 5714 23992 5720
rect 23846 5536 23902 5545
rect 23846 5471 23902 5480
rect 23848 5228 23900 5234
rect 23848 5170 23900 5176
rect 23860 4554 23888 5170
rect 23952 4758 23980 5714
rect 23940 4752 23992 4758
rect 23940 4694 23992 4700
rect 23848 4548 23900 4554
rect 23848 4490 23900 4496
rect 23756 4072 23808 4078
rect 23756 4014 23808 4020
rect 23952 3738 23980 4694
rect 23940 3732 23992 3738
rect 23940 3674 23992 3680
rect 23296 3596 23348 3602
rect 23296 3538 23348 3544
rect 23308 3194 23336 3538
rect 23388 3392 23440 3398
rect 23388 3334 23440 3340
rect 23296 3188 23348 3194
rect 23296 3130 23348 3136
rect 23400 2961 23428 3334
rect 24044 3194 24072 8622
rect 24122 8528 24178 8537
rect 24122 8463 24178 8472
rect 24136 7721 24164 8463
rect 24688 8242 24716 8894
rect 24320 8214 24716 8242
rect 24320 7834 24348 8214
rect 24780 8106 24808 10406
rect 24964 10062 24992 11018
rect 25228 10600 25280 10606
rect 25226 10568 25228 10577
rect 25280 10568 25282 10577
rect 25226 10503 25282 10512
rect 24952 10056 25004 10062
rect 24952 9998 25004 10004
rect 25228 9920 25280 9926
rect 25228 9862 25280 9868
rect 25240 9518 25268 9862
rect 25228 9512 25280 9518
rect 25226 9480 25228 9489
rect 25280 9480 25282 9489
rect 25226 9415 25282 9424
rect 25412 9376 25464 9382
rect 25412 9318 25464 9324
rect 25226 9208 25282 9217
rect 25226 9143 25282 9152
rect 25240 9110 25268 9143
rect 25228 9104 25280 9110
rect 25228 9046 25280 9052
rect 24860 8832 24912 8838
rect 24860 8774 24912 8780
rect 24228 7806 24348 7834
rect 24688 8078 24808 8106
rect 24122 7712 24178 7721
rect 24122 7647 24178 7656
rect 24124 6656 24176 6662
rect 24124 6598 24176 6604
rect 24136 6322 24164 6598
rect 24124 6316 24176 6322
rect 24124 6258 24176 6264
rect 24136 5846 24164 6258
rect 24124 5840 24176 5846
rect 24124 5782 24176 5788
rect 24228 5250 24256 7806
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24584 7336 24636 7342
rect 24688 7313 24716 8078
rect 24768 8016 24820 8022
rect 24872 7970 24900 8774
rect 25240 8634 25268 9046
rect 25228 8628 25280 8634
rect 25228 8570 25280 8576
rect 25136 8288 25188 8294
rect 25136 8230 25188 8236
rect 24820 7964 24900 7970
rect 24768 7958 24900 7964
rect 24780 7942 24900 7958
rect 25148 7954 25176 8230
rect 24872 7426 24900 7942
rect 25136 7948 25188 7954
rect 25136 7890 25188 7896
rect 24780 7410 24900 7426
rect 25148 7410 25176 7890
rect 25320 7744 25372 7750
rect 25320 7686 25372 7692
rect 24768 7404 24900 7410
rect 24820 7398 24900 7404
rect 25136 7404 25188 7410
rect 24768 7346 24820 7352
rect 25136 7346 25188 7352
rect 24584 7278 24636 7284
rect 24674 7304 24730 7313
rect 24596 7002 24624 7278
rect 24674 7239 24730 7248
rect 25044 7200 25096 7206
rect 25044 7142 25096 7148
rect 24584 6996 24636 7002
rect 24584 6938 24636 6944
rect 24596 6746 24624 6938
rect 24768 6860 24820 6866
rect 24768 6802 24820 6808
rect 24596 6718 24716 6746
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24688 6254 24716 6718
rect 24780 6458 24808 6802
rect 25056 6730 25084 7142
rect 25148 6798 25176 7346
rect 25332 7342 25360 7686
rect 25320 7336 25372 7342
rect 25320 7278 25372 7284
rect 25320 6860 25372 6866
rect 25320 6802 25372 6808
rect 25136 6792 25188 6798
rect 25136 6734 25188 6740
rect 25044 6724 25096 6730
rect 25044 6666 25096 6672
rect 24768 6452 24820 6458
rect 24768 6394 24820 6400
rect 24676 6248 24728 6254
rect 24676 6190 24728 6196
rect 24676 6112 24728 6118
rect 24676 6054 24728 6060
rect 24688 5778 24716 6054
rect 25332 5914 25360 6802
rect 25424 6089 25452 9318
rect 25792 9178 25820 12135
rect 25780 9172 25832 9178
rect 25780 9114 25832 9120
rect 25504 8968 25556 8974
rect 25504 8910 25556 8916
rect 25516 8362 25544 8910
rect 25792 8566 25820 9114
rect 25780 8560 25832 8566
rect 25780 8502 25832 8508
rect 25504 8356 25556 8362
rect 25504 8298 25556 8304
rect 25504 7336 25556 7342
rect 25504 7278 25556 7284
rect 25516 7177 25544 7278
rect 25688 7200 25740 7206
rect 25502 7168 25558 7177
rect 25688 7142 25740 7148
rect 25502 7103 25558 7112
rect 25504 6792 25556 6798
rect 25504 6734 25556 6740
rect 25516 6458 25544 6734
rect 25504 6452 25556 6458
rect 25504 6394 25556 6400
rect 25410 6080 25466 6089
rect 25410 6015 25466 6024
rect 25320 5908 25372 5914
rect 25320 5850 25372 5856
rect 24676 5772 24728 5778
rect 24676 5714 24728 5720
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24688 5302 24716 5714
rect 24768 5568 24820 5574
rect 24768 5510 24820 5516
rect 24780 5370 24808 5510
rect 24768 5364 24820 5370
rect 24768 5306 24820 5312
rect 24136 5222 24256 5250
rect 24308 5296 24360 5302
rect 24308 5238 24360 5244
rect 24676 5296 24728 5302
rect 24676 5238 24728 5244
rect 25410 5264 25466 5273
rect 24136 3505 24164 5222
rect 24320 5098 24348 5238
rect 25410 5199 25412 5208
rect 25464 5199 25466 5208
rect 25412 5170 25464 5176
rect 24308 5092 24360 5098
rect 24308 5034 24360 5040
rect 24216 5024 24268 5030
rect 25700 5001 25728 7142
rect 25884 6866 25912 13767
rect 25962 12472 26018 12481
rect 25962 12407 26018 12416
rect 25872 6860 25924 6866
rect 25872 6802 25924 6808
rect 24216 4966 24268 4972
rect 25686 4992 25742 5001
rect 24228 4826 24256 4966
rect 25686 4927 25742 4936
rect 24216 4820 24268 4826
rect 24216 4762 24268 4768
rect 25228 4684 25280 4690
rect 25228 4626 25280 4632
rect 25044 4480 25096 4486
rect 25044 4422 25096 4428
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24492 3936 24544 3942
rect 24492 3878 24544 3884
rect 24214 3632 24270 3641
rect 24214 3567 24270 3576
rect 24122 3496 24178 3505
rect 24122 3431 24178 3440
rect 24124 3392 24176 3398
rect 24124 3334 24176 3340
rect 24032 3188 24084 3194
rect 24032 3130 24084 3136
rect 23570 3088 23626 3097
rect 23570 3023 23626 3032
rect 23754 3088 23810 3097
rect 23754 3023 23810 3032
rect 23386 2952 23442 2961
rect 23386 2887 23442 2896
rect 23202 1864 23258 1873
rect 23202 1799 23258 1808
rect 23584 480 23612 3023
rect 23768 1465 23796 3023
rect 24044 2990 24072 3130
rect 24032 2984 24084 2990
rect 24032 2926 24084 2932
rect 23754 1456 23810 1465
rect 23754 1391 23810 1400
rect 294 0 350 480
rect 938 0 994 480
rect 1582 0 1638 480
rect 2226 0 2282 480
rect 2870 0 2926 480
rect 3606 0 3662 480
rect 4250 0 4306 480
rect 4894 0 4950 480
rect 5538 0 5594 480
rect 6274 0 6330 480
rect 6918 0 6974 480
rect 7562 0 7618 480
rect 8206 0 8262 480
rect 8942 0 8998 480
rect 9586 0 9642 480
rect 10230 0 10286 480
rect 10874 0 10930 480
rect 11610 0 11666 480
rect 12254 0 12310 480
rect 12898 0 12954 480
rect 13542 0 13598 480
rect 14278 0 14334 480
rect 14922 0 14978 480
rect 15566 0 15622 480
rect 16210 0 16266 480
rect 16854 0 16910 480
rect 17590 0 17646 480
rect 18234 0 18290 480
rect 18878 0 18934 480
rect 19522 0 19578 480
rect 20258 0 20314 480
rect 20902 0 20958 480
rect 21546 0 21602 480
rect 22190 0 22246 480
rect 22926 0 22982 480
rect 23570 0 23626 480
rect 24136 377 24164 3334
rect 24228 480 24256 3567
rect 24504 3505 24532 3878
rect 25056 3777 25084 4422
rect 25240 4078 25268 4626
rect 25976 4146 26004 12407
rect 27526 4176 27582 4185
rect 25964 4140 26016 4146
rect 27526 4111 27582 4120
rect 25964 4082 26016 4088
rect 25228 4072 25280 4078
rect 25226 4040 25228 4049
rect 25280 4040 25282 4049
rect 25226 3975 25282 3984
rect 26884 4004 26936 4010
rect 26884 3946 26936 3952
rect 24858 3768 24914 3777
rect 24858 3703 24914 3712
rect 25042 3768 25098 3777
rect 25042 3703 25098 3712
rect 24768 3596 24820 3602
rect 24768 3538 24820 3544
rect 24490 3496 24546 3505
rect 24490 3431 24546 3440
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24780 3194 24808 3538
rect 24768 3188 24820 3194
rect 24768 3130 24820 3136
rect 24872 2990 24900 3703
rect 26238 3496 26294 3505
rect 26238 3431 26294 3440
rect 24860 2984 24912 2990
rect 24860 2926 24912 2932
rect 24950 2952 25006 2961
rect 24950 2887 25006 2896
rect 24860 2848 24912 2854
rect 24688 2796 24860 2802
rect 24688 2790 24912 2796
rect 24688 2774 24900 2790
rect 24582 2544 24638 2553
rect 24582 2479 24584 2488
rect 24636 2479 24638 2488
rect 24584 2450 24636 2456
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24688 1465 24716 2774
rect 24768 2304 24820 2310
rect 24768 2246 24820 2252
rect 24674 1456 24730 1465
rect 24674 1391 24730 1400
rect 24780 921 24808 2246
rect 24964 1714 24992 2887
rect 24872 1686 24992 1714
rect 24766 912 24822 921
rect 24766 847 24822 856
rect 24872 480 24900 1686
rect 25594 1592 25650 1601
rect 25594 1527 25650 1536
rect 25608 480 25636 1527
rect 26252 480 26280 3431
rect 26896 480 26924 3946
rect 27540 480 27568 4111
rect 24122 368 24178 377
rect 24122 303 24178 312
rect 24214 0 24270 480
rect 24858 0 24914 480
rect 25594 0 25650 480
rect 26238 0 26294 480
rect 26882 0 26938 480
rect 27526 0 27582 480
<< via2 >>
rect 24582 27648 24638 27704
rect 1582 24384 1638 24440
rect 938 23568 994 23624
rect 2962 24792 3018 24848
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 4986 24656 5042 24712
rect 4342 24112 4398 24168
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 3698 23704 3754 23760
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 6642 22228 6698 22264
rect 6642 22208 6644 22228
rect 6644 22208 6696 22228
rect 6696 22208 6698 22228
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 2318 20440 2374 20496
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 294 19216 350 19272
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5446 15408 5502 15464
rect 5354 15000 5410 15056
rect 3606 8880 3662 8936
rect 2226 7928 2282 7984
rect 294 5208 350 5264
rect 1674 4664 1730 4720
rect 1582 3984 1638 4040
rect 938 3712 994 3768
rect 1674 3712 1730 3768
rect 2870 2896 2926 2952
rect 4066 7928 4122 7984
rect 4066 6976 4122 7032
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 7286 21120 7342 21176
rect 8206 23296 8262 23352
rect 8114 22752 8170 22808
rect 7746 21936 7802 21992
rect 7654 20984 7710 21040
rect 7194 13368 7250 13424
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 6274 6296 6330 6352
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5538 3032 5594 3088
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 7562 5616 7618 5672
rect 6918 3984 6974 4040
rect 8206 22480 8262 22536
rect 9954 24828 9956 24848
rect 9956 24828 10008 24848
rect 10008 24828 10010 24848
rect 9954 24792 10010 24828
rect 9954 24656 10010 24712
rect 9126 21664 9182 21720
rect 8482 21120 8538 21176
rect 8758 20984 8814 21040
rect 9770 21936 9826 21992
rect 9678 20984 9734 21040
rect 10046 24384 10102 24440
rect 9954 21936 10010 21992
rect 8482 19760 8538 19816
rect 8942 7520 8998 7576
rect 8206 6724 8262 6760
rect 8206 6704 8208 6724
rect 8208 6704 8260 6724
rect 8260 6704 8262 6724
rect 8022 3576 8078 3632
rect 9770 15000 9826 15056
rect 9954 14864 10010 14920
rect 9494 5752 9550 5808
rect 9310 3984 9366 4040
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10322 24656 10378 24712
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10138 23296 10194 23352
rect 10322 22480 10378 22536
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10138 22228 10194 22264
rect 10138 22208 10140 22228
rect 10140 22208 10192 22228
rect 10192 22208 10194 22228
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10782 22380 10784 22400
rect 10784 22380 10836 22400
rect 10836 22380 10838 22400
rect 10782 22344 10838 22380
rect 11426 23976 11482 24032
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10690 18672 10746 18728
rect 10598 18420 10654 18456
rect 10598 18400 10600 18420
rect 10600 18400 10652 18420
rect 10652 18400 10654 18420
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10138 17040 10194 17096
rect 10782 16904 10838 16960
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10966 18264 11022 18320
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10598 10548 10600 10568
rect 10600 10548 10652 10568
rect 10652 10548 10654 10568
rect 10598 10512 10654 10548
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10230 3596 10286 3632
rect 10230 3576 10232 3596
rect 10232 3576 10284 3596
rect 10284 3576 10286 3596
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 9586 1672 9642 1728
rect 10782 15428 10838 15464
rect 10782 15408 10784 15428
rect 10784 15408 10836 15428
rect 10836 15408 10838 15428
rect 11150 16088 11206 16144
rect 11242 12144 11298 12200
rect 11886 23024 11942 23080
rect 11702 22092 11758 22128
rect 11702 22072 11704 22092
rect 11704 22072 11756 22092
rect 11756 22072 11758 22092
rect 12622 24112 12678 24168
rect 11426 15952 11482 16008
rect 11610 13368 11666 13424
rect 10966 9696 11022 9752
rect 11610 10376 11666 10432
rect 12806 22208 12862 22264
rect 12806 20848 12862 20904
rect 12070 19216 12126 19272
rect 12162 18164 12164 18184
rect 12164 18164 12216 18184
rect 12216 18164 12218 18184
rect 12162 18128 12218 18164
rect 12622 18944 12678 19000
rect 12622 18400 12678 18456
rect 11978 13368 12034 13424
rect 12254 13232 12310 13288
rect 12162 12280 12218 12336
rect 11794 10512 11850 10568
rect 11702 9152 11758 9208
rect 10874 7112 10930 7168
rect 11058 6296 11114 6352
rect 11334 1536 11390 1592
rect 13450 24656 13506 24712
rect 13082 23976 13138 24032
rect 13266 23316 13322 23352
rect 13266 23296 13268 23316
rect 13268 23296 13320 23316
rect 13320 23296 13322 23316
rect 13082 22636 13138 22672
rect 13082 22616 13084 22636
rect 13084 22616 13136 22636
rect 13136 22616 13138 22636
rect 13082 20168 13138 20224
rect 12990 16940 12992 16960
rect 12992 16940 13044 16960
rect 13044 16940 13046 16960
rect 12990 16904 13046 16940
rect 12898 16496 12954 16552
rect 12622 7792 12678 7848
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 15290 24112 15346 24168
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 14002 22752 14058 22808
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14186 22072 14242 22128
rect 14186 21428 14188 21448
rect 14188 21428 14240 21448
rect 14240 21428 14242 21448
rect 14186 21392 14242 21428
rect 13726 20052 13782 20088
rect 13726 20032 13728 20052
rect 13728 20032 13780 20052
rect 13780 20032 13782 20052
rect 14186 19760 14242 19816
rect 13634 18944 13690 19000
rect 13450 18400 13506 18456
rect 13726 17992 13782 18048
rect 14094 17040 14150 17096
rect 13266 15544 13322 15600
rect 13634 15544 13690 15600
rect 13174 12824 13230 12880
rect 12898 5616 12954 5672
rect 12898 4936 12954 4992
rect 12806 2372 12862 2408
rect 12806 2352 12808 2372
rect 12808 2352 12860 2372
rect 12860 2352 12862 2372
rect 12254 1808 12310 1864
rect 13174 5208 13230 5264
rect 14370 17720 14426 17776
rect 14002 14864 14058 14920
rect 14370 14592 14426 14648
rect 13818 12416 13874 12472
rect 13726 11620 13782 11656
rect 13726 11600 13728 11620
rect 13728 11600 13780 11620
rect 13780 11600 13782 11620
rect 13542 9696 13598 9752
rect 14370 12824 14426 12880
rect 14370 12416 14426 12472
rect 14002 9288 14058 9344
rect 13542 9016 13598 9072
rect 13450 8336 13506 8392
rect 14646 22480 14702 22536
rect 14554 9968 14610 10024
rect 13634 6316 13690 6352
rect 13634 6296 13636 6316
rect 13636 6296 13688 6316
rect 13688 6296 13690 6316
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14738 21684 14794 21720
rect 14738 21664 14740 21684
rect 14740 21664 14792 21684
rect 14792 21664 14794 21684
rect 15842 24112 15898 24168
rect 16118 23588 16174 23624
rect 16118 23568 16120 23588
rect 16120 23568 16172 23588
rect 16172 23568 16174 23588
rect 16302 24556 16304 24576
rect 16304 24556 16356 24576
rect 16356 24556 16358 24576
rect 16302 24520 16358 24556
rect 18602 24792 18658 24848
rect 16486 24248 16542 24304
rect 16394 23724 16450 23760
rect 16394 23704 16396 23724
rect 16396 23704 16448 23724
rect 16448 23704 16450 23724
rect 16394 22888 16450 22944
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 15658 20712 15714 20768
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14830 18264 14886 18320
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14830 17196 14886 17232
rect 14830 17176 14832 17196
rect 14832 17176 14884 17196
rect 14884 17176 14886 17196
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14738 13504 14794 13560
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 15290 12552 15346 12608
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 13542 4120 13598 4176
rect 13634 4004 13690 4040
rect 13634 3984 13636 4004
rect 13636 3984 13688 4004
rect 13688 3984 13690 4004
rect 13634 3848 13690 3904
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 15198 4936 15254 4992
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14830 4120 14886 4176
rect 15934 20848 15990 20904
rect 15750 20168 15806 20224
rect 15750 19236 15806 19272
rect 15750 19216 15752 19236
rect 15752 19216 15804 19236
rect 15804 19216 15806 19236
rect 15842 19116 15844 19136
rect 15844 19116 15896 19136
rect 15896 19116 15898 19136
rect 15658 18128 15714 18184
rect 15842 19080 15898 19116
rect 15842 17992 15898 18048
rect 15658 14592 15714 14648
rect 15474 8336 15530 8392
rect 15566 7268 15622 7304
rect 15566 7248 15568 7268
rect 15568 7248 15620 7268
rect 15620 7248 15622 7268
rect 15934 14884 15990 14920
rect 15934 14864 15936 14884
rect 15936 14864 15988 14884
rect 15988 14864 15990 14884
rect 16946 23432 17002 23488
rect 17590 23024 17646 23080
rect 17958 24520 18014 24576
rect 18326 23296 18382 23352
rect 17958 22752 18014 22808
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 20718 24792 20774 24848
rect 19430 24656 19486 24712
rect 18694 23432 18750 23488
rect 18878 22616 18934 22672
rect 18602 22344 18658 22400
rect 18142 22208 18198 22264
rect 17314 21936 17370 21992
rect 16670 19080 16726 19136
rect 16762 17176 16818 17232
rect 16946 16940 16948 16960
rect 16948 16940 17000 16960
rect 17000 16940 17002 16960
rect 16946 16904 17002 16940
rect 16854 16496 16910 16552
rect 16118 15952 16174 16008
rect 16026 14592 16082 14648
rect 15842 14320 15898 14376
rect 15934 10512 15990 10568
rect 15842 9968 15898 10024
rect 15750 7792 15806 7848
rect 14922 3440 14978 3496
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 15658 3884 15660 3904
rect 15660 3884 15712 3904
rect 15712 3884 15714 3904
rect 15658 3848 15714 3884
rect 15750 3712 15806 3768
rect 17774 20712 17830 20768
rect 17406 20440 17462 20496
rect 16854 10784 16910 10840
rect 16302 9152 16358 9208
rect 16210 8880 16266 8936
rect 16210 7148 16212 7168
rect 16212 7148 16264 7168
rect 16264 7148 16266 7168
rect 16210 7112 16266 7148
rect 16118 3576 16174 3632
rect 16486 5364 16542 5400
rect 16486 5344 16488 5364
rect 16488 5344 16540 5364
rect 16540 5344 16542 5364
rect 16118 3440 16174 3496
rect 17774 17992 17830 18048
rect 17498 16632 17554 16688
rect 17498 13368 17554 13424
rect 17682 12588 17684 12608
rect 17684 12588 17736 12608
rect 17736 12588 17738 12608
rect 17682 12552 17738 12588
rect 18878 22072 18934 22128
rect 19246 23160 19302 23216
rect 19246 23024 19302 23080
rect 19154 22480 19210 22536
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19614 24284 19616 24304
rect 19616 24284 19668 24304
rect 19668 24284 19670 24304
rect 19614 24248 19670 24284
rect 20074 24248 20130 24304
rect 20258 23568 20314 23624
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19522 23160 19578 23216
rect 19338 22208 19394 22264
rect 18234 17992 18290 18048
rect 18602 18400 18658 18456
rect 18418 17040 18474 17096
rect 18786 16904 18842 16960
rect 18234 15136 18290 15192
rect 17774 11600 17830 11656
rect 17498 9696 17554 9752
rect 18694 15972 18750 16008
rect 18694 15952 18696 15972
rect 18696 15952 18748 15972
rect 18748 15952 18750 15972
rect 18602 12824 18658 12880
rect 18418 12552 18474 12608
rect 18970 17176 19026 17232
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 20074 21120 20130 21176
rect 20074 20984 20130 21040
rect 19982 20848 20038 20904
rect 19338 20304 19394 20360
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 18970 15544 19026 15600
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19246 16668 19248 16688
rect 19248 16668 19300 16688
rect 19300 16668 19302 16688
rect 19246 16632 19302 16668
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19430 15408 19486 15464
rect 19982 14864 20038 14920
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 20718 22924 20720 22944
rect 20720 22924 20772 22944
rect 20772 22924 20774 22944
rect 20718 22888 20774 22924
rect 20534 22752 20590 22808
rect 20350 21684 20406 21720
rect 20350 21664 20352 21684
rect 20352 21664 20404 21684
rect 20404 21664 20406 21684
rect 20718 21428 20720 21448
rect 20720 21428 20772 21448
rect 20772 21428 20774 21448
rect 20718 21392 20774 21428
rect 20810 20460 20866 20496
rect 20810 20440 20812 20460
rect 20812 20440 20864 20460
rect 20864 20440 20866 20460
rect 21086 24132 21142 24168
rect 21086 24112 21088 24132
rect 21088 24112 21140 24132
rect 21140 24112 21142 24132
rect 21362 22072 21418 22128
rect 21178 20984 21234 21040
rect 21914 23296 21970 23352
rect 21546 22500 21602 22536
rect 21546 22480 21548 22500
rect 21548 22480 21600 22500
rect 21600 22480 21602 22500
rect 20902 18672 20958 18728
rect 20626 17584 20682 17640
rect 20626 17312 20682 17368
rect 20258 14592 20314 14648
rect 18878 12688 18934 12744
rect 18602 11056 18658 11112
rect 19430 12416 19486 12472
rect 18786 10104 18842 10160
rect 18786 9696 18842 9752
rect 18234 7828 18236 7848
rect 18236 7828 18288 7848
rect 18288 7828 18290 7848
rect 17958 7656 18014 7712
rect 18234 7792 18290 7828
rect 17958 6704 18014 6760
rect 16762 6160 16818 6216
rect 18694 7384 18750 7440
rect 18326 4664 18382 4720
rect 17222 3712 17278 3768
rect 19338 9288 19394 9344
rect 20626 14864 20682 14920
rect 21270 16632 21326 16688
rect 20902 13368 20958 13424
rect 20534 13096 20590 13152
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 20074 12416 20130 12472
rect 20074 10648 20130 10704
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19430 6976 19486 7032
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 20166 7520 20222 7576
rect 20074 7384 20130 7440
rect 19982 6704 20038 6760
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 20074 5752 20130 5808
rect 19430 5480 19486 5536
rect 18878 5108 18880 5128
rect 18880 5108 18932 5128
rect 18932 5108 18934 5128
rect 18878 5072 18934 5108
rect 18326 3440 18382 3496
rect 16210 2760 16266 2816
rect 17038 2796 17040 2816
rect 17040 2796 17092 2816
rect 17092 2796 17094 2816
rect 17038 2760 17094 2796
rect 17866 3168 17922 3224
rect 17774 2916 17830 2952
rect 17774 2896 17776 2916
rect 17776 2896 17828 2916
rect 17828 2896 17830 2916
rect 18234 2624 18290 2680
rect 18878 3304 18934 3360
rect 19798 5244 19800 5264
rect 19800 5244 19852 5264
rect 19852 5244 19854 5264
rect 19798 5208 19854 5244
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19798 4684 19854 4720
rect 19798 4664 19800 4684
rect 19800 4664 19852 4684
rect 19852 4664 19854 4684
rect 19798 4392 19854 4448
rect 19982 4256 20038 4312
rect 20350 11056 20406 11112
rect 21362 13776 21418 13832
rect 20534 10512 20590 10568
rect 20350 9288 20406 9344
rect 20442 8880 20498 8936
rect 20442 8608 20498 8664
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 20166 3304 20222 3360
rect 19614 3168 19670 3224
rect 19246 3032 19302 3088
rect 18786 2896 18842 2952
rect 18878 2760 18934 2816
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 20350 6976 20406 7032
rect 21270 10784 21326 10840
rect 21546 13096 21602 13152
rect 21546 12552 21602 12608
rect 21454 11736 21510 11792
rect 20902 10532 20958 10568
rect 20902 10512 20904 10532
rect 20904 10512 20956 10532
rect 20956 10512 20958 10532
rect 21362 10512 21418 10568
rect 20994 9152 21050 9208
rect 21270 7792 21326 7848
rect 20994 7112 21050 7168
rect 20810 6976 20866 7032
rect 21086 5616 21142 5672
rect 20442 3732 20498 3768
rect 20442 3712 20444 3732
rect 20444 3712 20496 3732
rect 20496 3712 20498 3732
rect 21454 8336 21510 8392
rect 21362 6296 21418 6352
rect 21546 4120 21602 4176
rect 21914 22616 21970 22672
rect 21822 20984 21878 21040
rect 21730 18672 21786 18728
rect 21730 16496 21786 16552
rect 22098 20848 22154 20904
rect 22282 20304 22338 20360
rect 23294 27104 23350 27160
rect 24030 26560 24086 26616
rect 23570 25880 23626 25936
rect 23754 24792 23810 24848
rect 22650 20848 22706 20904
rect 22558 20440 22614 20496
rect 21730 15580 21732 15600
rect 21732 15580 21784 15600
rect 21784 15580 21786 15600
rect 21730 15544 21786 15580
rect 22466 17060 22522 17096
rect 22466 17040 22468 17060
rect 22468 17040 22520 17060
rect 22520 17040 22522 17060
rect 22282 16496 22338 16552
rect 21822 11600 21878 11656
rect 23662 22480 23718 22536
rect 23478 21664 23534 21720
rect 23478 21256 23534 21312
rect 23294 20848 23350 20904
rect 23110 19896 23166 19952
rect 23478 19896 23534 19952
rect 23018 18400 23074 18456
rect 22834 17584 22890 17640
rect 22742 15136 22798 15192
rect 21914 7248 21970 7304
rect 22006 6840 22062 6896
rect 22650 13404 22652 13424
rect 22652 13404 22704 13424
rect 22704 13404 22706 13424
rect 22650 13368 22706 13404
rect 22558 11600 22614 11656
rect 22926 11736 22982 11792
rect 22558 9288 22614 9344
rect 22558 9016 22614 9072
rect 22466 6160 22522 6216
rect 21822 5344 21878 5400
rect 22282 5092 22338 5128
rect 22282 5072 22284 5092
rect 22284 5072 22336 5092
rect 22336 5072 22338 5092
rect 21638 3712 21694 3768
rect 21086 3440 21142 3496
rect 21086 3032 21142 3088
rect 21546 2896 21602 2952
rect 20626 2488 20682 2544
rect 22650 4528 22706 4584
rect 21914 1536 21970 1592
rect 22650 3576 22706 3632
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24766 25356 24822 25392
rect 24766 25336 24768 25356
rect 24768 25336 24820 25356
rect 24820 25336 24822 25356
rect 24214 23604 24216 23624
rect 24216 23604 24268 23624
rect 24268 23604 24270 23624
rect 24214 23568 24270 23604
rect 24674 23568 24730 23624
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24950 23860 25006 23896
rect 24950 23840 24952 23860
rect 24952 23840 25004 23860
rect 25004 23840 25006 23860
rect 25502 23568 25558 23624
rect 24766 23432 24822 23488
rect 27526 23840 27582 23896
rect 26146 23432 26202 23488
rect 24030 21528 24086 21584
rect 23662 19216 23718 19272
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24214 21120 24270 21176
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24766 20848 24822 20904
rect 25502 20476 25504 20496
rect 25504 20476 25556 20496
rect 25556 20476 25558 20496
rect 25502 20440 25558 20476
rect 24674 19624 24730 19680
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24122 18944 24178 19000
rect 23202 16088 23258 16144
rect 23938 17448 23994 17504
rect 23846 16088 23902 16144
rect 24582 19352 24638 19408
rect 24398 18672 24454 18728
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24122 17312 24178 17368
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 23110 12416 23166 12472
rect 23662 15408 23718 15464
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 25042 15952 25098 16008
rect 25410 15952 25466 16008
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24030 13096 24086 13152
rect 23662 10140 23664 10160
rect 23664 10140 23716 10160
rect 23716 10140 23718 10160
rect 23662 10104 23718 10140
rect 23570 9968 23626 10024
rect 23386 9424 23442 9480
rect 22926 3440 22982 3496
rect 22834 1672 22890 1728
rect 23478 9016 23534 9072
rect 23294 6860 23350 6896
rect 23294 6840 23296 6860
rect 23296 6840 23348 6860
rect 23348 6840 23350 6860
rect 23846 9016 23902 9072
rect 23570 6160 23626 6216
rect 23662 4684 23718 4720
rect 23662 4664 23664 4684
rect 23664 4664 23716 4684
rect 23716 4664 23718 4684
rect 23570 4256 23626 4312
rect 23018 2644 23074 2680
rect 23018 2624 23020 2644
rect 23020 2624 23072 2644
rect 23072 2624 23074 2644
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 25870 13776 25926 13832
rect 25778 12144 25834 12200
rect 24674 11872 24730 11928
rect 25134 11328 25190 11384
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24582 9560 24638 9616
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 23938 7928 23994 7984
rect 23846 5480 23902 5536
rect 24122 8472 24178 8528
rect 25226 10548 25228 10568
rect 25228 10548 25280 10568
rect 25280 10548 25282 10568
rect 25226 10512 25282 10548
rect 25226 9460 25228 9480
rect 25228 9460 25280 9480
rect 25280 9460 25282 9480
rect 25226 9424 25282 9460
rect 25226 9152 25282 9208
rect 24122 7656 24178 7712
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24674 7248 24730 7304
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 25502 7112 25558 7168
rect 25410 6024 25466 6080
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 25410 5228 25466 5264
rect 25410 5208 25412 5228
rect 25412 5208 25464 5228
rect 25464 5208 25466 5228
rect 25962 12416 26018 12472
rect 25686 4936 25742 4992
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24214 3576 24270 3632
rect 24122 3440 24178 3496
rect 23570 3032 23626 3088
rect 23754 3032 23810 3088
rect 23386 2896 23442 2952
rect 23202 1808 23258 1864
rect 23754 1400 23810 1456
rect 27526 4120 27582 4176
rect 25226 4020 25228 4040
rect 25228 4020 25280 4040
rect 25280 4020 25282 4040
rect 25226 3984 25282 4020
rect 24858 3712 24914 3768
rect 25042 3712 25098 3768
rect 24490 3440 24546 3496
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 26238 3440 26294 3496
rect 24950 2896 25006 2952
rect 24582 2508 24638 2544
rect 24582 2488 24584 2508
rect 24584 2488 24636 2508
rect 24636 2488 24638 2508
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 24674 1400 24730 1456
rect 24766 856 24822 912
rect 25594 1536 25650 1592
rect 24122 312 24178 368
<< metal3 >>
rect 24577 27706 24643 27709
rect 27520 27706 28000 27736
rect 24577 27704 28000 27706
rect 24577 27648 24582 27704
rect 24638 27648 28000 27704
rect 24577 27646 28000 27648
rect 24577 27643 24643 27646
rect 27520 27616 28000 27646
rect 23289 27162 23355 27165
rect 27520 27162 28000 27192
rect 23289 27160 28000 27162
rect 23289 27104 23294 27160
rect 23350 27104 28000 27160
rect 23289 27102 28000 27104
rect 23289 27099 23355 27102
rect 27520 27072 28000 27102
rect 24025 26618 24091 26621
rect 27520 26618 28000 26648
rect 24025 26616 28000 26618
rect 24025 26560 24030 26616
rect 24086 26560 28000 26616
rect 24025 26558 28000 26560
rect 24025 26555 24091 26558
rect 27520 26528 28000 26558
rect 23565 25938 23631 25941
rect 27520 25938 28000 25968
rect 23565 25936 28000 25938
rect 23565 25880 23570 25936
rect 23626 25880 28000 25936
rect 23565 25878 28000 25880
rect 23565 25875 23631 25878
rect 27520 25848 28000 25878
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 24761 25394 24827 25397
rect 27520 25394 28000 25424
rect 24761 25392 28000 25394
rect 24761 25336 24766 25392
rect 24822 25336 28000 25392
rect 24761 25334 28000 25336
rect 24761 25331 24827 25334
rect 27520 25304 28000 25334
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 2957 24850 3023 24853
rect 9949 24850 10015 24853
rect 2957 24848 10015 24850
rect 2957 24792 2962 24848
rect 3018 24792 9954 24848
rect 10010 24792 10015 24848
rect 2957 24790 10015 24792
rect 2957 24787 3023 24790
rect 9949 24787 10015 24790
rect 18597 24850 18663 24853
rect 20713 24850 20779 24853
rect 18597 24848 20779 24850
rect 18597 24792 18602 24848
rect 18658 24792 20718 24848
rect 20774 24792 20779 24848
rect 18597 24790 20779 24792
rect 18597 24787 18663 24790
rect 20713 24787 20779 24790
rect 23749 24850 23815 24853
rect 27520 24850 28000 24880
rect 23749 24848 28000 24850
rect 23749 24792 23754 24848
rect 23810 24792 28000 24848
rect 23749 24790 28000 24792
rect 23749 24787 23815 24790
rect 27520 24760 28000 24790
rect 4981 24714 5047 24717
rect 9949 24714 10015 24717
rect 10317 24714 10383 24717
rect 4981 24712 10383 24714
rect 4981 24656 4986 24712
rect 5042 24656 9954 24712
rect 10010 24656 10322 24712
rect 10378 24656 10383 24712
rect 4981 24654 10383 24656
rect 4981 24651 5047 24654
rect 9949 24651 10015 24654
rect 10317 24651 10383 24654
rect 13445 24714 13511 24717
rect 19425 24714 19491 24717
rect 13445 24712 19491 24714
rect 13445 24656 13450 24712
rect 13506 24656 19430 24712
rect 19486 24656 19491 24712
rect 13445 24654 19491 24656
rect 13445 24651 13511 24654
rect 19425 24651 19491 24654
rect 16297 24578 16363 24581
rect 17953 24578 18019 24581
rect 16297 24576 18019 24578
rect 16297 24520 16302 24576
rect 16358 24520 17958 24576
rect 18014 24520 18019 24576
rect 16297 24518 18019 24520
rect 16297 24515 16363 24518
rect 17953 24515 18019 24518
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 1577 24442 1643 24445
rect 10041 24442 10107 24445
rect 1577 24440 10107 24442
rect 1577 24384 1582 24440
rect 1638 24384 10046 24440
rect 10102 24384 10107 24440
rect 1577 24382 10107 24384
rect 1577 24379 1643 24382
rect 10041 24379 10107 24382
rect 16481 24306 16547 24309
rect 19609 24306 19675 24309
rect 16481 24304 19675 24306
rect 16481 24248 16486 24304
rect 16542 24248 19614 24304
rect 19670 24248 19675 24304
rect 16481 24246 19675 24248
rect 16481 24243 16547 24246
rect 19609 24243 19675 24246
rect 20069 24306 20135 24309
rect 20069 24304 27538 24306
rect 20069 24248 20074 24304
rect 20130 24248 27538 24304
rect 20069 24246 27538 24248
rect 20069 24243 20135 24246
rect 27478 24200 27538 24246
rect 4337 24170 4403 24173
rect 12617 24170 12683 24173
rect 15285 24170 15351 24173
rect 4337 24168 9506 24170
rect 4337 24112 4342 24168
rect 4398 24112 9506 24168
rect 4337 24110 9506 24112
rect 4337 24107 4403 24110
rect 9446 24034 9506 24110
rect 12617 24168 15351 24170
rect 12617 24112 12622 24168
rect 12678 24112 15290 24168
rect 15346 24112 15351 24168
rect 12617 24110 15351 24112
rect 12617 24107 12683 24110
rect 15285 24107 15351 24110
rect 15837 24170 15903 24173
rect 21081 24170 21147 24173
rect 15837 24168 21147 24170
rect 15837 24112 15842 24168
rect 15898 24112 21086 24168
rect 21142 24112 21147 24168
rect 15837 24110 21147 24112
rect 27478 24110 28000 24200
rect 15837 24107 15903 24110
rect 21081 24107 21147 24110
rect 27520 24080 28000 24110
rect 11421 24034 11487 24037
rect 13077 24034 13143 24037
rect 9446 24032 13143 24034
rect 9446 23976 11426 24032
rect 11482 23976 13082 24032
rect 13138 23976 13143 24032
rect 9446 23974 13143 23976
rect 11421 23971 11487 23974
rect 13077 23971 13143 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 24945 23898 25011 23901
rect 27521 23898 27587 23901
rect 24945 23896 27587 23898
rect 24945 23840 24950 23896
rect 25006 23840 27526 23896
rect 27582 23840 27587 23896
rect 24945 23838 27587 23840
rect 24945 23835 25011 23838
rect 27521 23835 27587 23838
rect 3693 23762 3759 23765
rect 16389 23762 16455 23765
rect 3693 23760 16455 23762
rect 3693 23704 3698 23760
rect 3754 23704 16394 23760
rect 16450 23704 16455 23760
rect 3693 23702 16455 23704
rect 3693 23699 3759 23702
rect 16389 23699 16455 23702
rect 24534 23702 25698 23762
rect 933 23626 999 23629
rect 16113 23626 16179 23629
rect 933 23624 16179 23626
rect 933 23568 938 23624
rect 994 23568 16118 23624
rect 16174 23568 16179 23624
rect 933 23566 16179 23568
rect 933 23563 999 23566
rect 16113 23563 16179 23566
rect 20253 23626 20319 23629
rect 24209 23626 24275 23629
rect 20253 23624 24275 23626
rect 20253 23568 20258 23624
rect 20314 23568 24214 23624
rect 24270 23568 24275 23624
rect 20253 23566 24275 23568
rect 20253 23563 20319 23566
rect 24209 23563 24275 23566
rect 16941 23490 17007 23493
rect 18689 23490 18755 23493
rect 16941 23488 18755 23490
rect 16941 23432 16946 23488
rect 17002 23432 18694 23488
rect 18750 23432 18755 23488
rect 16941 23430 18755 23432
rect 16941 23427 17007 23430
rect 18689 23427 18755 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 8201 23354 8267 23357
rect 10133 23354 10199 23357
rect 8201 23352 10199 23354
rect 8201 23296 8206 23352
rect 8262 23296 10138 23352
rect 10194 23296 10199 23352
rect 8201 23294 10199 23296
rect 8201 23291 8267 23294
rect 10133 23291 10199 23294
rect 13261 23354 13327 23357
rect 18321 23354 18387 23357
rect 13261 23352 18387 23354
rect 13261 23296 13266 23352
rect 13322 23296 18326 23352
rect 18382 23296 18387 23352
rect 13261 23294 18387 23296
rect 13261 23291 13327 23294
rect 18321 23291 18387 23294
rect 21909 23354 21975 23357
rect 24534 23354 24594 23702
rect 24669 23626 24735 23629
rect 25497 23626 25563 23629
rect 24669 23624 25563 23626
rect 24669 23568 24674 23624
rect 24730 23568 25502 23624
rect 25558 23568 25563 23624
rect 24669 23566 25563 23568
rect 25638 23626 25698 23702
rect 27520 23626 28000 23656
rect 25638 23566 28000 23626
rect 24669 23563 24735 23566
rect 25497 23563 25563 23566
rect 27520 23536 28000 23566
rect 24761 23490 24827 23493
rect 26141 23490 26207 23493
rect 24761 23488 26207 23490
rect 24761 23432 24766 23488
rect 24822 23432 26146 23488
rect 26202 23432 26207 23488
rect 24761 23430 26207 23432
rect 24761 23427 24827 23430
rect 26141 23427 26207 23430
rect 21909 23352 24594 23354
rect 21909 23296 21914 23352
rect 21970 23296 24594 23352
rect 21909 23294 24594 23296
rect 21909 23291 21975 23294
rect 19241 23218 19307 23221
rect 19517 23218 19583 23221
rect 19241 23216 19583 23218
rect 19241 23160 19246 23216
rect 19302 23160 19522 23216
rect 19578 23160 19583 23216
rect 19241 23158 19583 23160
rect 19241 23155 19307 23158
rect 19517 23155 19583 23158
rect 11881 23082 11947 23085
rect 17585 23082 17651 23085
rect 11881 23080 17651 23082
rect 11881 23024 11886 23080
rect 11942 23024 17590 23080
rect 17646 23024 17651 23080
rect 11881 23022 17651 23024
rect 11881 23019 11947 23022
rect 17585 23019 17651 23022
rect 19241 23082 19307 23085
rect 27520 23082 28000 23112
rect 19241 23080 28000 23082
rect 19241 23024 19246 23080
rect 19302 23024 28000 23080
rect 19241 23022 28000 23024
rect 19241 23019 19307 23022
rect 27520 22992 28000 23022
rect 16389 22946 16455 22949
rect 20713 22946 20779 22949
rect 16389 22944 20779 22946
rect 16389 22888 16394 22944
rect 16450 22888 20718 22944
rect 20774 22888 20779 22944
rect 16389 22886 20779 22888
rect 16389 22883 16455 22886
rect 20713 22883 20779 22886
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 8109 22810 8175 22813
rect 13997 22810 14063 22813
rect 8109 22808 14063 22810
rect 8109 22752 8114 22808
rect 8170 22752 14002 22808
rect 14058 22752 14063 22808
rect 8109 22750 14063 22752
rect 8109 22747 8175 22750
rect 13997 22747 14063 22750
rect 17953 22810 18019 22813
rect 20529 22810 20595 22813
rect 17953 22808 20595 22810
rect 17953 22752 17958 22808
rect 18014 22752 20534 22808
rect 20590 22752 20595 22808
rect 17953 22750 20595 22752
rect 17953 22747 18019 22750
rect 20529 22747 20595 22750
rect 13077 22674 13143 22677
rect 18873 22674 18939 22677
rect 21909 22674 21975 22677
rect 13077 22672 18939 22674
rect 13077 22616 13082 22672
rect 13138 22616 18878 22672
rect 18934 22616 18939 22672
rect 13077 22614 18939 22616
rect 13077 22611 13143 22614
rect 18873 22611 18939 22614
rect 19014 22672 21975 22674
rect 19014 22616 21914 22672
rect 21970 22616 21975 22672
rect 19014 22614 21975 22616
rect 8201 22538 8267 22541
rect 10317 22538 10383 22541
rect 8201 22536 10383 22538
rect 8201 22480 8206 22536
rect 8262 22480 10322 22536
rect 10378 22480 10383 22536
rect 8201 22478 10383 22480
rect 8201 22475 8267 22478
rect 10317 22475 10383 22478
rect 14641 22538 14707 22541
rect 19014 22538 19074 22614
rect 21909 22611 21975 22614
rect 14641 22536 19074 22538
rect 14641 22480 14646 22536
rect 14702 22480 19074 22536
rect 14641 22478 19074 22480
rect 19149 22538 19215 22541
rect 21541 22538 21607 22541
rect 19149 22536 21607 22538
rect 19149 22480 19154 22536
rect 19210 22480 21546 22536
rect 21602 22480 21607 22536
rect 19149 22478 21607 22480
rect 14641 22475 14707 22478
rect 19149 22475 19215 22478
rect 21541 22475 21607 22478
rect 23657 22538 23723 22541
rect 27520 22538 28000 22568
rect 23657 22536 28000 22538
rect 23657 22480 23662 22536
rect 23718 22480 28000 22536
rect 23657 22478 28000 22480
rect 23657 22475 23723 22478
rect 27520 22448 28000 22478
rect 10777 22402 10843 22405
rect 18597 22402 18663 22405
rect 10777 22400 18663 22402
rect 10777 22344 10782 22400
rect 10838 22344 18602 22400
rect 18658 22344 18663 22400
rect 10777 22342 18663 22344
rect 10777 22339 10843 22342
rect 18597 22339 18663 22342
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 6637 22266 6703 22269
rect 10133 22266 10199 22269
rect 6637 22264 10199 22266
rect 6637 22208 6642 22264
rect 6698 22208 10138 22264
rect 10194 22208 10199 22264
rect 6637 22206 10199 22208
rect 6637 22203 6703 22206
rect 10133 22203 10199 22206
rect 12801 22266 12867 22269
rect 18137 22266 18203 22269
rect 19333 22266 19399 22269
rect 12801 22264 19399 22266
rect 12801 22208 12806 22264
rect 12862 22208 18142 22264
rect 18198 22208 19338 22264
rect 19394 22208 19399 22264
rect 12801 22206 19399 22208
rect 12801 22203 12867 22206
rect 18137 22203 18203 22206
rect 19333 22203 19399 22206
rect 11697 22130 11763 22133
rect 14181 22130 14247 22133
rect 11697 22128 14247 22130
rect 11697 22072 11702 22128
rect 11758 22072 14186 22128
rect 14242 22072 14247 22128
rect 11697 22070 14247 22072
rect 11697 22067 11763 22070
rect 14181 22067 14247 22070
rect 18873 22130 18939 22133
rect 21357 22130 21423 22133
rect 18873 22128 21423 22130
rect 18873 22072 18878 22128
rect 18934 22072 21362 22128
rect 21418 22072 21423 22128
rect 18873 22070 21423 22072
rect 18873 22067 18939 22070
rect 21357 22067 21423 22070
rect 7741 21994 7807 21997
rect 9765 21994 9831 21997
rect 7741 21992 9831 21994
rect 7741 21936 7746 21992
rect 7802 21936 9770 21992
rect 9826 21936 9831 21992
rect 7741 21934 9831 21936
rect 7741 21931 7807 21934
rect 9765 21931 9831 21934
rect 9949 21994 10015 21997
rect 17309 21994 17375 21997
rect 9949 21992 17375 21994
rect 9949 21936 9954 21992
rect 10010 21936 17314 21992
rect 17370 21936 17375 21992
rect 9949 21934 17375 21936
rect 9949 21931 10015 21934
rect 17309 21931 17375 21934
rect 27520 21858 28000 21888
rect 24718 21798 28000 21858
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 9121 21722 9187 21725
rect 14733 21722 14799 21725
rect 9121 21720 14799 21722
rect 9121 21664 9126 21720
rect 9182 21664 14738 21720
rect 14794 21664 14799 21720
rect 9121 21662 14799 21664
rect 9121 21659 9187 21662
rect 14733 21659 14799 21662
rect 20345 21722 20411 21725
rect 23473 21722 23539 21725
rect 20345 21720 23539 21722
rect 20345 21664 20350 21720
rect 20406 21664 23478 21720
rect 23534 21664 23539 21720
rect 20345 21662 23539 21664
rect 20345 21659 20411 21662
rect 23473 21659 23539 21662
rect 24025 21586 24091 21589
rect 24718 21586 24778 21798
rect 27520 21768 28000 21798
rect 24025 21584 24778 21586
rect 24025 21528 24030 21584
rect 24086 21528 24778 21584
rect 24025 21526 24778 21528
rect 24025 21523 24091 21526
rect 14181 21450 14247 21453
rect 20713 21450 20779 21453
rect 14181 21448 20779 21450
rect 14181 21392 14186 21448
rect 14242 21392 20718 21448
rect 20774 21392 20779 21448
rect 14181 21390 20779 21392
rect 14181 21387 14247 21390
rect 20713 21387 20779 21390
rect 23473 21314 23539 21317
rect 27520 21314 28000 21344
rect 23473 21312 28000 21314
rect 23473 21256 23478 21312
rect 23534 21256 28000 21312
rect 23473 21254 28000 21256
rect 23473 21251 23539 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 27520 21224 28000 21254
rect 19610 21183 19930 21184
rect 7281 21178 7347 21181
rect 8477 21178 8543 21181
rect 7281 21176 8543 21178
rect 7281 21120 7286 21176
rect 7342 21120 8482 21176
rect 8538 21120 8543 21176
rect 7281 21118 8543 21120
rect 7281 21115 7347 21118
rect 8477 21115 8543 21118
rect 20069 21178 20135 21181
rect 24209 21178 24275 21181
rect 20069 21176 24275 21178
rect 20069 21120 20074 21176
rect 20130 21120 24214 21176
rect 24270 21120 24275 21176
rect 20069 21118 24275 21120
rect 20069 21115 20135 21118
rect 24209 21115 24275 21118
rect 0 21042 480 21072
rect 7649 21042 7715 21045
rect 8753 21042 8819 21045
rect 9673 21042 9739 21045
rect 0 21040 9739 21042
rect 0 20984 7654 21040
rect 7710 20984 8758 21040
rect 8814 20984 9678 21040
rect 9734 20984 9739 21040
rect 0 20982 9739 20984
rect 0 20952 480 20982
rect 7649 20979 7715 20982
rect 8753 20979 8819 20982
rect 9673 20979 9739 20982
rect 20069 21042 20135 21045
rect 21173 21042 21239 21045
rect 20069 21040 21239 21042
rect 20069 20984 20074 21040
rect 20130 20984 21178 21040
rect 21234 20984 21239 21040
rect 20069 20982 21239 20984
rect 20069 20979 20135 20982
rect 21173 20979 21239 20982
rect 21817 21042 21883 21045
rect 21817 21040 24962 21042
rect 21817 20984 21822 21040
rect 21878 20984 24962 21040
rect 21817 20982 24962 20984
rect 21817 20979 21883 20982
rect 12801 20906 12867 20909
rect 15929 20906 15995 20909
rect 12801 20904 15995 20906
rect 12801 20848 12806 20904
rect 12862 20848 15934 20904
rect 15990 20848 15995 20904
rect 12801 20846 15995 20848
rect 12801 20843 12867 20846
rect 15929 20843 15995 20846
rect 19977 20906 20043 20909
rect 22093 20906 22159 20909
rect 22645 20906 22711 20909
rect 19977 20904 22711 20906
rect 19977 20848 19982 20904
rect 20038 20848 22098 20904
rect 22154 20848 22650 20904
rect 22706 20848 22711 20904
rect 19977 20846 22711 20848
rect 19977 20843 20043 20846
rect 22093 20843 22159 20846
rect 22645 20843 22711 20846
rect 23289 20906 23355 20909
rect 24761 20906 24827 20909
rect 23289 20904 24827 20906
rect 23289 20848 23294 20904
rect 23350 20848 24766 20904
rect 24822 20848 24827 20904
rect 23289 20846 24827 20848
rect 23289 20843 23355 20846
rect 24761 20843 24827 20846
rect 15653 20770 15719 20773
rect 17769 20770 17835 20773
rect 15653 20768 17835 20770
rect 15653 20712 15658 20768
rect 15714 20712 17774 20768
rect 17830 20712 17835 20768
rect 15653 20710 17835 20712
rect 24902 20770 24962 20982
rect 27520 20770 28000 20800
rect 24902 20710 28000 20770
rect 15653 20707 15719 20710
rect 17769 20707 17835 20710
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 27520 20680 28000 20710
rect 24277 20639 24597 20640
rect 2313 20498 2379 20501
rect 17401 20498 17467 20501
rect 20805 20498 20871 20501
rect 2313 20496 20871 20498
rect 2313 20440 2318 20496
rect 2374 20440 17406 20496
rect 17462 20440 20810 20496
rect 20866 20440 20871 20496
rect 2313 20438 20871 20440
rect 2313 20435 2379 20438
rect 17401 20435 17467 20438
rect 20805 20435 20871 20438
rect 22553 20498 22619 20501
rect 25497 20498 25563 20501
rect 22553 20496 25563 20498
rect 22553 20440 22558 20496
rect 22614 20440 25502 20496
rect 25558 20440 25563 20496
rect 22553 20438 25563 20440
rect 22553 20435 22619 20438
rect 25497 20435 25563 20438
rect 19333 20362 19399 20365
rect 22277 20362 22343 20365
rect 19333 20360 22343 20362
rect 19333 20304 19338 20360
rect 19394 20304 22282 20360
rect 22338 20304 22343 20360
rect 19333 20302 22343 20304
rect 19333 20299 19399 20302
rect 22277 20299 22343 20302
rect 13077 20226 13143 20229
rect 15745 20226 15811 20229
rect 13077 20224 15811 20226
rect 13077 20168 13082 20224
rect 13138 20168 15750 20224
rect 15806 20168 15811 20224
rect 13077 20166 15811 20168
rect 13077 20163 13143 20166
rect 15745 20163 15811 20166
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 13721 20090 13787 20093
rect 27520 20090 28000 20120
rect 13721 20088 13922 20090
rect 13721 20032 13726 20088
rect 13782 20032 13922 20088
rect 13721 20030 13922 20032
rect 13721 20027 13787 20030
rect 13862 19954 13922 20030
rect 24902 20030 28000 20090
rect 23105 19954 23171 19957
rect 23473 19954 23539 19957
rect 13862 19952 23539 19954
rect 13862 19896 23110 19952
rect 23166 19896 23478 19952
rect 23534 19896 23539 19952
rect 13862 19894 23539 19896
rect 23105 19891 23171 19894
rect 23473 19891 23539 19894
rect 8477 19818 8543 19821
rect 14181 19818 14247 19821
rect 8477 19816 14247 19818
rect 8477 19760 8482 19816
rect 8538 19760 14186 19816
rect 14242 19760 14247 19816
rect 8477 19758 14247 19760
rect 8477 19755 8543 19758
rect 14181 19755 14247 19758
rect 24669 19682 24735 19685
rect 24902 19682 24962 20030
rect 27520 20000 28000 20030
rect 24669 19680 24962 19682
rect 24669 19624 24674 19680
rect 24730 19624 24962 19680
rect 24669 19622 24962 19624
rect 24669 19619 24735 19622
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 27520 19546 28000 19576
rect 24718 19486 28000 19546
rect 24577 19410 24643 19413
rect 24718 19410 24778 19486
rect 27520 19456 28000 19486
rect 24577 19408 24778 19410
rect 24577 19352 24582 19408
rect 24638 19352 24778 19408
rect 24577 19350 24778 19352
rect 24577 19347 24643 19350
rect 289 19274 355 19277
rect 12065 19274 12131 19277
rect 15745 19274 15811 19277
rect 23657 19274 23723 19277
rect 289 19272 15811 19274
rect 289 19216 294 19272
rect 350 19216 12070 19272
rect 12126 19216 15750 19272
rect 15806 19216 15811 19272
rect 289 19214 15811 19216
rect 289 19211 355 19214
rect 12065 19211 12131 19214
rect 15745 19211 15811 19214
rect 16806 19272 23723 19274
rect 16806 19216 23662 19272
rect 23718 19216 23723 19272
rect 16806 19214 23723 19216
rect 15837 19138 15903 19141
rect 16665 19138 16731 19141
rect 15837 19136 16731 19138
rect 15837 19080 15842 19136
rect 15898 19080 16670 19136
rect 16726 19080 16731 19136
rect 15837 19078 16731 19080
rect 15837 19075 15903 19078
rect 16665 19075 16731 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 12617 19002 12683 19005
rect 13629 19002 13695 19005
rect 16806 19002 16866 19214
rect 23657 19211 23723 19214
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 12617 19000 16866 19002
rect 12617 18944 12622 19000
rect 12678 18944 13634 19000
rect 13690 18944 16866 19000
rect 12617 18942 16866 18944
rect 24117 19002 24183 19005
rect 27520 19002 28000 19032
rect 24117 19000 28000 19002
rect 24117 18944 24122 19000
rect 24178 18944 28000 19000
rect 24117 18942 28000 18944
rect 12617 18939 12683 18942
rect 13629 18939 13695 18942
rect 24117 18939 24183 18942
rect 27520 18912 28000 18942
rect 10685 18730 10751 18733
rect 20897 18730 20963 18733
rect 21725 18730 21791 18733
rect 10685 18728 21791 18730
rect 10685 18672 10690 18728
rect 10746 18672 20902 18728
rect 20958 18672 21730 18728
rect 21786 18672 21791 18728
rect 10685 18670 21791 18672
rect 10685 18667 10751 18670
rect 20897 18667 20963 18670
rect 21725 18667 21791 18670
rect 23974 18668 23980 18732
rect 24044 18730 24050 18732
rect 24393 18730 24459 18733
rect 24044 18728 24459 18730
rect 24044 18672 24398 18728
rect 24454 18672 24459 18728
rect 24044 18670 24459 18672
rect 24044 18668 24050 18670
rect 24393 18667 24459 18670
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 10593 18458 10659 18461
rect 12617 18458 12683 18461
rect 13445 18458 13511 18461
rect 10593 18456 13511 18458
rect 10593 18400 10598 18456
rect 10654 18400 12622 18456
rect 12678 18400 13450 18456
rect 13506 18400 13511 18456
rect 10593 18398 13511 18400
rect 10593 18395 10659 18398
rect 12617 18395 12683 18398
rect 13445 18395 13511 18398
rect 18597 18458 18663 18461
rect 23013 18458 23079 18461
rect 27520 18458 28000 18488
rect 18597 18456 23079 18458
rect 18597 18400 18602 18456
rect 18658 18400 23018 18456
rect 23074 18400 23079 18456
rect 18597 18398 23079 18400
rect 18597 18395 18663 18398
rect 23013 18395 23079 18398
rect 24902 18398 28000 18458
rect 10961 18322 11027 18325
rect 14825 18322 14891 18325
rect 10961 18320 14891 18322
rect 10961 18264 10966 18320
rect 11022 18264 14830 18320
rect 14886 18264 14891 18320
rect 10961 18262 14891 18264
rect 10961 18259 11027 18262
rect 14825 18259 14891 18262
rect 12157 18186 12223 18189
rect 15653 18186 15719 18189
rect 24902 18186 24962 18398
rect 27520 18368 28000 18398
rect 12157 18184 24962 18186
rect 12157 18128 12162 18184
rect 12218 18128 15658 18184
rect 15714 18128 24962 18184
rect 12157 18126 24962 18128
rect 12157 18123 12223 18126
rect 15653 18123 15719 18126
rect 13721 18050 13787 18053
rect 15837 18050 15903 18053
rect 13721 18048 15903 18050
rect 13721 17992 13726 18048
rect 13782 17992 15842 18048
rect 15898 17992 15903 18048
rect 13721 17990 15903 17992
rect 13721 17987 13787 17990
rect 15837 17987 15903 17990
rect 17769 18050 17835 18053
rect 18229 18050 18295 18053
rect 17769 18048 18295 18050
rect 17769 17992 17774 18048
rect 17830 17992 18234 18048
rect 18290 17992 18295 18048
rect 17769 17990 18295 17992
rect 17769 17987 17835 17990
rect 18229 17987 18295 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 14365 17778 14431 17781
rect 27520 17778 28000 17808
rect 14365 17776 28000 17778
rect 14365 17720 14370 17776
rect 14426 17720 28000 17776
rect 14365 17718 28000 17720
rect 14365 17715 14431 17718
rect 27520 17688 28000 17718
rect 20621 17642 20687 17645
rect 22829 17642 22895 17645
rect 20621 17640 22895 17642
rect 20621 17584 20626 17640
rect 20682 17584 22834 17640
rect 22890 17584 22895 17640
rect 20621 17582 22895 17584
rect 20621 17579 20687 17582
rect 22829 17579 22895 17582
rect 23933 17506 23999 17509
rect 15886 17504 23999 17506
rect 15886 17448 23938 17504
rect 23994 17448 23999 17504
rect 15886 17446 23999 17448
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 14825 17234 14891 17237
rect 15886 17234 15946 17446
rect 23933 17443 23999 17446
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 20621 17370 20687 17373
rect 24117 17370 24183 17373
rect 20621 17368 24183 17370
rect 20621 17312 20626 17368
rect 20682 17312 24122 17368
rect 24178 17312 24183 17368
rect 20621 17310 24183 17312
rect 20621 17307 20687 17310
rect 24117 17307 24183 17310
rect 14825 17232 15946 17234
rect 14825 17176 14830 17232
rect 14886 17176 15946 17232
rect 14825 17174 15946 17176
rect 16757 17234 16823 17237
rect 18965 17234 19031 17237
rect 27520 17234 28000 17264
rect 16757 17232 28000 17234
rect 16757 17176 16762 17232
rect 16818 17176 18970 17232
rect 19026 17176 28000 17232
rect 16757 17174 28000 17176
rect 14825 17171 14891 17174
rect 16757 17171 16823 17174
rect 18965 17171 19031 17174
rect 27520 17144 28000 17174
rect 10133 17098 10199 17101
rect 14089 17098 14155 17101
rect 10133 17096 14155 17098
rect 10133 17040 10138 17096
rect 10194 17040 14094 17096
rect 14150 17040 14155 17096
rect 10133 17038 14155 17040
rect 10133 17035 10199 17038
rect 14089 17035 14155 17038
rect 18413 17098 18479 17101
rect 22461 17098 22527 17101
rect 18413 17096 22527 17098
rect 18413 17040 18418 17096
rect 18474 17040 22466 17096
rect 22522 17040 22527 17096
rect 18413 17038 22527 17040
rect 18413 17035 18479 17038
rect 22461 17035 22527 17038
rect 10777 16962 10843 16965
rect 12985 16962 13051 16965
rect 10777 16960 13051 16962
rect 10777 16904 10782 16960
rect 10838 16904 12990 16960
rect 13046 16904 13051 16960
rect 10777 16902 13051 16904
rect 10777 16899 10843 16902
rect 12985 16899 13051 16902
rect 16941 16962 17007 16965
rect 18781 16962 18847 16965
rect 16941 16960 18847 16962
rect 16941 16904 16946 16960
rect 17002 16904 18786 16960
rect 18842 16904 18847 16960
rect 16941 16902 18847 16904
rect 16941 16899 17007 16902
rect 18781 16899 18847 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 17493 16690 17559 16693
rect 19241 16690 19307 16693
rect 17493 16688 19307 16690
rect 17493 16632 17498 16688
rect 17554 16632 19246 16688
rect 19302 16632 19307 16688
rect 17493 16630 19307 16632
rect 17493 16627 17559 16630
rect 19241 16627 19307 16630
rect 21265 16690 21331 16693
rect 27520 16690 28000 16720
rect 21265 16688 28000 16690
rect 21265 16632 21270 16688
rect 21326 16632 28000 16688
rect 21265 16630 28000 16632
rect 21265 16627 21331 16630
rect 27520 16600 28000 16630
rect 12893 16554 12959 16557
rect 16849 16554 16915 16557
rect 12893 16552 16915 16554
rect 12893 16496 12898 16552
rect 12954 16496 16854 16552
rect 16910 16496 16915 16552
rect 12893 16494 16915 16496
rect 12893 16491 12959 16494
rect 16849 16491 16915 16494
rect 21725 16554 21791 16557
rect 22277 16554 22343 16557
rect 21725 16552 22343 16554
rect 21725 16496 21730 16552
rect 21786 16496 22282 16552
rect 22338 16496 22343 16552
rect 21725 16494 22343 16496
rect 21725 16491 21791 16494
rect 22277 16491 22343 16494
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 11145 16146 11211 16149
rect 23197 16146 23263 16149
rect 23841 16146 23907 16149
rect 11145 16144 23907 16146
rect 11145 16088 11150 16144
rect 11206 16088 23202 16144
rect 23258 16088 23846 16144
rect 23902 16088 23907 16144
rect 11145 16086 23907 16088
rect 11145 16083 11211 16086
rect 23197 16083 23263 16086
rect 23841 16083 23907 16086
rect 11421 16010 11487 16013
rect 16113 16010 16179 16013
rect 11421 16008 16179 16010
rect 11421 15952 11426 16008
rect 11482 15952 16118 16008
rect 16174 15952 16179 16008
rect 11421 15950 16179 15952
rect 11421 15947 11487 15950
rect 16113 15947 16179 15950
rect 18689 16010 18755 16013
rect 25037 16010 25103 16013
rect 18689 16008 25103 16010
rect 18689 15952 18694 16008
rect 18750 15952 25042 16008
rect 25098 15952 25103 16008
rect 18689 15950 25103 15952
rect 18689 15947 18755 15950
rect 25037 15947 25103 15950
rect 25405 16010 25471 16013
rect 27520 16010 28000 16040
rect 25405 16008 28000 16010
rect 25405 15952 25410 16008
rect 25466 15952 28000 16008
rect 25405 15950 28000 15952
rect 25405 15947 25471 15950
rect 27520 15920 28000 15950
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 13261 15602 13327 15605
rect 13629 15602 13695 15605
rect 13261 15600 13695 15602
rect 13261 15544 13266 15600
rect 13322 15544 13634 15600
rect 13690 15544 13695 15600
rect 13261 15542 13695 15544
rect 13261 15539 13327 15542
rect 13629 15539 13695 15542
rect 18965 15602 19031 15605
rect 21725 15602 21791 15605
rect 18965 15600 21791 15602
rect 18965 15544 18970 15600
rect 19026 15544 21730 15600
rect 21786 15544 21791 15600
rect 18965 15542 21791 15544
rect 18965 15539 19031 15542
rect 21725 15539 21791 15542
rect 5441 15466 5507 15469
rect 10777 15466 10843 15469
rect 5441 15464 10843 15466
rect 5441 15408 5446 15464
rect 5502 15408 10782 15464
rect 10838 15408 10843 15464
rect 5441 15406 10843 15408
rect 5441 15403 5507 15406
rect 10777 15403 10843 15406
rect 19425 15466 19491 15469
rect 23657 15466 23723 15469
rect 27520 15466 28000 15496
rect 19425 15464 28000 15466
rect 19425 15408 19430 15464
rect 19486 15408 23662 15464
rect 23718 15408 28000 15464
rect 19425 15406 28000 15408
rect 19425 15403 19491 15406
rect 23657 15403 23723 15406
rect 27520 15376 28000 15406
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 18229 15194 18295 15197
rect 22737 15194 22803 15197
rect 18229 15192 22803 15194
rect 18229 15136 18234 15192
rect 18290 15136 22742 15192
rect 22798 15136 22803 15192
rect 18229 15134 22803 15136
rect 18229 15131 18295 15134
rect 22737 15131 22803 15134
rect 5349 15058 5415 15061
rect 9765 15058 9831 15061
rect 5349 15056 9831 15058
rect 5349 15000 5354 15056
rect 5410 15000 9770 15056
rect 9826 15000 9831 15056
rect 5349 14998 9831 15000
rect 5349 14995 5415 14998
rect 9765 14995 9831 14998
rect 9949 14922 10015 14925
rect 13997 14922 14063 14925
rect 9949 14920 14063 14922
rect 9949 14864 9954 14920
rect 10010 14864 14002 14920
rect 14058 14864 14063 14920
rect 9949 14862 14063 14864
rect 9949 14859 10015 14862
rect 13997 14859 14063 14862
rect 15929 14922 15995 14925
rect 19977 14922 20043 14925
rect 20621 14922 20687 14925
rect 27520 14922 28000 14952
rect 15929 14920 20178 14922
rect 15929 14864 15934 14920
rect 15990 14864 19982 14920
rect 20038 14864 20178 14920
rect 15929 14862 20178 14864
rect 15929 14859 15995 14862
rect 19977 14859 20043 14862
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 14365 14650 14431 14653
rect 15653 14650 15719 14653
rect 16021 14650 16087 14653
rect 14365 14648 16087 14650
rect 14365 14592 14370 14648
rect 14426 14592 15658 14648
rect 15714 14592 16026 14648
rect 16082 14592 16087 14648
rect 14365 14590 16087 14592
rect 20118 14650 20178 14862
rect 20621 14920 28000 14922
rect 20621 14864 20626 14920
rect 20682 14864 28000 14920
rect 20621 14862 28000 14864
rect 20621 14859 20687 14862
rect 27520 14832 28000 14862
rect 20253 14650 20319 14653
rect 20118 14648 20319 14650
rect 20118 14592 20258 14648
rect 20314 14592 20319 14648
rect 20118 14590 20319 14592
rect 14365 14587 14431 14590
rect 15653 14587 15719 14590
rect 16021 14587 16087 14590
rect 20253 14587 20319 14590
rect 15837 14378 15903 14381
rect 27520 14378 28000 14408
rect 15837 14376 28000 14378
rect 15837 14320 15842 14376
rect 15898 14320 28000 14376
rect 15837 14318 28000 14320
rect 15837 14315 15903 14318
rect 27520 14288 28000 14318
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 21357 13834 21423 13837
rect 25865 13834 25931 13837
rect 21357 13832 25931 13834
rect 21357 13776 21362 13832
rect 21418 13776 25870 13832
rect 25926 13776 25931 13832
rect 21357 13774 25931 13776
rect 21357 13771 21423 13774
rect 25865 13771 25931 13774
rect 27520 13698 28000 13728
rect 23476 13638 28000 13698
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 14733 13562 14799 13565
rect 14733 13560 18522 13562
rect 14733 13504 14738 13560
rect 14794 13504 18522 13560
rect 14733 13502 18522 13504
rect 14733 13499 14799 13502
rect 7189 13426 7255 13429
rect 11605 13426 11671 13429
rect 7189 13424 11671 13426
rect 7189 13368 7194 13424
rect 7250 13368 11610 13424
rect 11666 13368 11671 13424
rect 7189 13366 11671 13368
rect 7189 13363 7255 13366
rect 11605 13363 11671 13366
rect 11973 13426 12039 13429
rect 17493 13426 17559 13429
rect 11973 13424 17559 13426
rect 11973 13368 11978 13424
rect 12034 13368 17498 13424
rect 17554 13368 17559 13424
rect 11973 13366 17559 13368
rect 18462 13426 18522 13502
rect 20897 13426 20963 13429
rect 22645 13426 22711 13429
rect 18462 13424 22711 13426
rect 18462 13368 20902 13424
rect 20958 13368 22650 13424
rect 22706 13368 22711 13424
rect 18462 13366 22711 13368
rect 11973 13363 12039 13366
rect 17493 13363 17559 13366
rect 20897 13363 20963 13366
rect 22645 13363 22711 13366
rect 12249 13290 12315 13293
rect 23476 13290 23536 13638
rect 27520 13608 28000 13638
rect 12249 13288 23536 13290
rect 12249 13232 12254 13288
rect 12310 13232 23536 13288
rect 12249 13230 23536 13232
rect 12249 13227 12315 13230
rect 20529 13154 20595 13157
rect 21541 13154 21607 13157
rect 24025 13156 24091 13157
rect 20529 13152 21607 13154
rect 20529 13096 20534 13152
rect 20590 13096 21546 13152
rect 21602 13096 21607 13152
rect 20529 13094 21607 13096
rect 20529 13091 20595 13094
rect 21541 13091 21607 13094
rect 23974 13092 23980 13156
rect 24044 13154 24091 13156
rect 27520 13154 28000 13184
rect 24044 13152 24136 13154
rect 24086 13096 24136 13152
rect 24044 13094 24136 13096
rect 24902 13094 28000 13154
rect 24044 13092 24091 13094
rect 24025 13091 24091 13092
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 13169 12882 13235 12885
rect 14365 12882 14431 12885
rect 18597 12882 18663 12885
rect 13169 12880 14431 12882
rect 13169 12824 13174 12880
rect 13230 12824 14370 12880
rect 14426 12824 14431 12880
rect 13169 12822 14431 12824
rect 13169 12819 13235 12822
rect 14365 12819 14431 12822
rect 18416 12880 18663 12882
rect 18416 12824 18602 12880
rect 18658 12824 18663 12880
rect 18416 12822 18663 12824
rect 18416 12613 18476 12822
rect 18597 12819 18663 12822
rect 18873 12746 18939 12749
rect 24902 12746 24962 13094
rect 27520 13064 28000 13094
rect 18873 12744 24962 12746
rect 18873 12688 18878 12744
rect 18934 12688 24962 12744
rect 18873 12686 24962 12688
rect 18873 12683 18939 12686
rect 15285 12610 15351 12613
rect 17677 12610 17743 12613
rect 15285 12608 17743 12610
rect 15285 12552 15290 12608
rect 15346 12552 17682 12608
rect 17738 12552 17743 12608
rect 15285 12550 17743 12552
rect 15285 12547 15351 12550
rect 17677 12547 17743 12550
rect 18413 12608 18479 12613
rect 18413 12552 18418 12608
rect 18474 12552 18479 12608
rect 18413 12547 18479 12552
rect 21541 12610 21607 12613
rect 27520 12610 28000 12640
rect 21541 12608 28000 12610
rect 21541 12552 21546 12608
rect 21602 12552 28000 12608
rect 21541 12550 28000 12552
rect 21541 12547 21607 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 27520 12520 28000 12550
rect 19610 12479 19930 12480
rect 13813 12474 13879 12477
rect 12758 12472 13879 12474
rect 12758 12416 13818 12472
rect 13874 12416 13879 12472
rect 12758 12414 13879 12416
rect 12157 12338 12223 12341
rect 12758 12338 12818 12414
rect 13813 12411 13879 12414
rect 14365 12474 14431 12477
rect 19425 12474 19491 12477
rect 14365 12472 19491 12474
rect 14365 12416 14370 12472
rect 14426 12416 19430 12472
rect 19486 12416 19491 12472
rect 14365 12414 19491 12416
rect 14365 12411 14431 12414
rect 19425 12411 19491 12414
rect 20069 12474 20135 12477
rect 23105 12474 23171 12477
rect 25957 12474 26023 12477
rect 20069 12472 26023 12474
rect 20069 12416 20074 12472
rect 20130 12416 23110 12472
rect 23166 12416 25962 12472
rect 26018 12416 26023 12472
rect 20069 12414 26023 12416
rect 20069 12411 20135 12414
rect 23105 12411 23171 12414
rect 25957 12411 26023 12414
rect 12157 12336 12818 12338
rect 12157 12280 12162 12336
rect 12218 12280 12818 12336
rect 12157 12278 12818 12280
rect 12157 12275 12223 12278
rect 11237 12202 11303 12205
rect 25773 12202 25839 12205
rect 11237 12200 25839 12202
rect 11237 12144 11242 12200
rect 11298 12144 25778 12200
rect 25834 12144 25839 12200
rect 11237 12142 25839 12144
rect 11237 12139 11303 12142
rect 25773 12139 25839 12142
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 24669 11930 24735 11933
rect 27520 11930 28000 11960
rect 24669 11928 28000 11930
rect 24669 11872 24674 11928
rect 24730 11872 28000 11928
rect 24669 11870 28000 11872
rect 24669 11867 24735 11870
rect 27520 11840 28000 11870
rect 21449 11794 21515 11797
rect 22921 11794 22987 11797
rect 21449 11792 22987 11794
rect 21449 11736 21454 11792
rect 21510 11736 22926 11792
rect 22982 11736 22987 11792
rect 21449 11734 22987 11736
rect 21449 11731 21515 11734
rect 22921 11731 22987 11734
rect 13721 11658 13787 11661
rect 17769 11658 17835 11661
rect 13721 11656 17835 11658
rect 13721 11600 13726 11656
rect 13782 11600 17774 11656
rect 17830 11600 17835 11656
rect 13721 11598 17835 11600
rect 13721 11595 13787 11598
rect 17769 11595 17835 11598
rect 21817 11658 21883 11661
rect 22553 11658 22619 11661
rect 21817 11656 22619 11658
rect 21817 11600 21822 11656
rect 21878 11600 22558 11656
rect 22614 11600 22619 11656
rect 21817 11598 22619 11600
rect 21817 11595 21883 11598
rect 22553 11595 22619 11598
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 25129 11386 25195 11389
rect 27520 11386 28000 11416
rect 25129 11384 28000 11386
rect 25129 11328 25134 11384
rect 25190 11328 28000 11384
rect 25129 11326 28000 11328
rect 25129 11323 25195 11326
rect 27520 11296 28000 11326
rect 18597 11114 18663 11117
rect 20345 11114 20411 11117
rect 18597 11112 20411 11114
rect 18597 11056 18602 11112
rect 18658 11056 20350 11112
rect 20406 11056 20411 11112
rect 18597 11054 20411 11056
rect 18597 11051 18663 11054
rect 20345 11051 20411 11054
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 16849 10842 16915 10845
rect 21265 10842 21331 10845
rect 27520 10842 28000 10872
rect 16849 10840 21331 10842
rect 16849 10784 16854 10840
rect 16910 10784 21270 10840
rect 21326 10784 21331 10840
rect 16849 10782 21331 10784
rect 16849 10779 16915 10782
rect 21265 10779 21331 10782
rect 24902 10782 28000 10842
rect 20069 10706 20135 10709
rect 24902 10706 24962 10782
rect 27520 10752 28000 10782
rect 20069 10704 24962 10706
rect 20069 10648 20074 10704
rect 20130 10648 24962 10704
rect 20069 10646 24962 10648
rect 20069 10643 20135 10646
rect 10593 10570 10659 10573
rect 11789 10570 11855 10573
rect 15929 10570 15995 10573
rect 20529 10570 20595 10573
rect 20897 10570 20963 10573
rect 10593 10568 15995 10570
rect 10593 10512 10598 10568
rect 10654 10512 11794 10568
rect 11850 10512 15934 10568
rect 15990 10512 15995 10568
rect 10593 10510 15995 10512
rect 10593 10507 10659 10510
rect 11789 10507 11855 10510
rect 15929 10507 15995 10510
rect 18646 10568 20963 10570
rect 18646 10512 20534 10568
rect 20590 10512 20902 10568
rect 20958 10512 20963 10568
rect 18646 10510 20963 10512
rect 11605 10434 11671 10437
rect 18646 10434 18706 10510
rect 20529 10507 20595 10510
rect 20897 10507 20963 10510
rect 21357 10570 21423 10573
rect 25221 10570 25287 10573
rect 21357 10568 25287 10570
rect 21357 10512 21362 10568
rect 21418 10512 25226 10568
rect 25282 10512 25287 10568
rect 21357 10510 25287 10512
rect 21357 10507 21423 10510
rect 25221 10507 25287 10510
rect 11605 10432 18706 10434
rect 11605 10376 11610 10432
rect 11666 10376 18706 10432
rect 11605 10374 18706 10376
rect 11605 10371 11671 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 18781 10162 18847 10165
rect 23657 10162 23723 10165
rect 27520 10162 28000 10192
rect 18781 10160 23723 10162
rect 18781 10104 18786 10160
rect 18842 10104 23662 10160
rect 23718 10104 23723 10160
rect 18781 10102 23723 10104
rect 18781 10099 18847 10102
rect 23657 10099 23723 10102
rect 23798 10102 28000 10162
rect 14549 10026 14615 10029
rect 15837 10026 15903 10029
rect 14549 10024 15903 10026
rect 14549 9968 14554 10024
rect 14610 9968 15842 10024
rect 15898 9968 15903 10024
rect 14549 9966 15903 9968
rect 14549 9963 14615 9966
rect 15837 9963 15903 9966
rect 23565 10026 23631 10029
rect 23798 10026 23858 10102
rect 27520 10072 28000 10102
rect 23565 10024 23858 10026
rect 23565 9968 23570 10024
rect 23626 9968 23858 10024
rect 23565 9966 23858 9968
rect 23565 9963 23631 9966
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 10961 9754 11027 9757
rect 13537 9754 13603 9757
rect 10961 9752 13603 9754
rect 10961 9696 10966 9752
rect 11022 9696 13542 9752
rect 13598 9696 13603 9752
rect 10961 9694 13603 9696
rect 10961 9691 11027 9694
rect 13537 9691 13603 9694
rect 17493 9754 17559 9757
rect 18781 9754 18847 9757
rect 17493 9752 18847 9754
rect 17493 9696 17498 9752
rect 17554 9696 18786 9752
rect 18842 9696 18847 9752
rect 17493 9694 18847 9696
rect 17493 9691 17559 9694
rect 18781 9691 18847 9694
rect 24577 9618 24643 9621
rect 27520 9618 28000 9648
rect 24577 9616 28000 9618
rect 24577 9560 24582 9616
rect 24638 9560 28000 9616
rect 24577 9558 28000 9560
rect 24577 9555 24643 9558
rect 27520 9528 28000 9558
rect 23381 9482 23447 9485
rect 25221 9482 25287 9485
rect 23381 9480 25287 9482
rect 23381 9424 23386 9480
rect 23442 9424 25226 9480
rect 25282 9424 25287 9480
rect 23381 9422 25287 9424
rect 23381 9419 23447 9422
rect 25221 9419 25287 9422
rect 13997 9346 14063 9349
rect 19333 9346 19399 9349
rect 13997 9344 19399 9346
rect 13997 9288 14002 9344
rect 14058 9288 19338 9344
rect 19394 9288 19399 9344
rect 13997 9286 19399 9288
rect 13997 9283 14063 9286
rect 19333 9283 19399 9286
rect 20345 9346 20411 9349
rect 22553 9346 22619 9349
rect 20345 9344 22619 9346
rect 20345 9288 20350 9344
rect 20406 9288 22558 9344
rect 22614 9288 22619 9344
rect 20345 9286 22619 9288
rect 20345 9283 20411 9286
rect 22553 9283 22619 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 11697 9210 11763 9213
rect 16297 9210 16363 9213
rect 11697 9208 16363 9210
rect 11697 9152 11702 9208
rect 11758 9152 16302 9208
rect 16358 9152 16363 9208
rect 11697 9150 16363 9152
rect 11697 9147 11763 9150
rect 16297 9147 16363 9150
rect 20989 9210 21055 9213
rect 25221 9210 25287 9213
rect 20989 9208 25287 9210
rect 20989 9152 20994 9208
rect 21050 9152 25226 9208
rect 25282 9152 25287 9208
rect 20989 9150 25287 9152
rect 20989 9147 21055 9150
rect 25221 9147 25287 9150
rect 13537 9074 13603 9077
rect 22553 9074 22619 9077
rect 23473 9074 23539 9077
rect 13537 9072 23539 9074
rect 13537 9016 13542 9072
rect 13598 9016 22558 9072
rect 22614 9016 23478 9072
rect 23534 9016 23539 9072
rect 13537 9014 23539 9016
rect 13537 9011 13603 9014
rect 22553 9011 22619 9014
rect 23473 9011 23539 9014
rect 23841 9074 23907 9077
rect 27520 9074 28000 9104
rect 23841 9072 28000 9074
rect 23841 9016 23846 9072
rect 23902 9016 28000 9072
rect 23841 9014 28000 9016
rect 23841 9011 23907 9014
rect 27520 8984 28000 9014
rect 3601 8938 3667 8941
rect 16205 8938 16271 8941
rect 3601 8936 16271 8938
rect 3601 8880 3606 8936
rect 3662 8880 16210 8936
rect 16266 8880 16271 8936
rect 3601 8878 16271 8880
rect 3601 8875 3667 8878
rect 16205 8875 16271 8878
rect 20437 8936 20503 8941
rect 20437 8880 20442 8936
rect 20498 8880 20503 8936
rect 20437 8875 20503 8880
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 20440 8669 20500 8875
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 20437 8664 20503 8669
rect 20437 8608 20442 8664
rect 20498 8608 20503 8664
rect 20437 8603 20503 8608
rect 24117 8530 24183 8533
rect 27520 8530 28000 8560
rect 24117 8528 28000 8530
rect 24117 8472 24122 8528
rect 24178 8472 28000 8528
rect 24117 8470 28000 8472
rect 24117 8467 24183 8470
rect 27520 8440 28000 8470
rect 13445 8394 13511 8397
rect 15469 8394 15535 8397
rect 13445 8392 15535 8394
rect 13445 8336 13450 8392
rect 13506 8336 15474 8392
rect 15530 8336 15535 8392
rect 13445 8334 15535 8336
rect 13445 8331 13511 8334
rect 15469 8331 15535 8334
rect 21449 8394 21515 8397
rect 21449 8392 24778 8394
rect 21449 8336 21454 8392
rect 21510 8336 24778 8392
rect 21449 8334 24778 8336
rect 21449 8331 21515 8334
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 2221 7986 2287 7989
rect 4061 7986 4127 7989
rect 23933 7986 23999 7989
rect 2221 7984 3986 7986
rect 2221 7928 2226 7984
rect 2282 7928 3986 7984
rect 2221 7926 3986 7928
rect 2221 7923 2287 7926
rect 3926 7306 3986 7926
rect 4061 7984 23999 7986
rect 4061 7928 4066 7984
rect 4122 7928 23938 7984
rect 23994 7928 23999 7984
rect 4061 7926 23999 7928
rect 4061 7923 4127 7926
rect 23933 7923 23999 7926
rect 12617 7850 12683 7853
rect 15745 7850 15811 7853
rect 12617 7848 15811 7850
rect 12617 7792 12622 7848
rect 12678 7792 15750 7848
rect 15806 7792 15811 7848
rect 12617 7790 15811 7792
rect 12617 7787 12683 7790
rect 15745 7787 15811 7790
rect 18229 7850 18295 7853
rect 21265 7850 21331 7853
rect 18229 7848 21331 7850
rect 18229 7792 18234 7848
rect 18290 7792 21270 7848
rect 21326 7792 21331 7848
rect 18229 7790 21331 7792
rect 24718 7850 24778 8334
rect 27520 7850 28000 7880
rect 24718 7790 28000 7850
rect 18229 7787 18295 7790
rect 21265 7787 21331 7790
rect 27520 7760 28000 7790
rect 17953 7714 18019 7717
rect 24117 7714 24183 7717
rect 17953 7712 24183 7714
rect 17953 7656 17958 7712
rect 18014 7656 24122 7712
rect 24178 7656 24183 7712
rect 17953 7654 24183 7656
rect 17953 7651 18019 7654
rect 24117 7651 24183 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 8937 7578 9003 7581
rect 20161 7578 20227 7581
rect 8937 7576 12634 7578
rect 8937 7520 8942 7576
rect 8998 7520 12634 7576
rect 8937 7518 12634 7520
rect 8937 7515 9003 7518
rect 12574 7442 12634 7518
rect 15334 7576 20227 7578
rect 15334 7520 20166 7576
rect 20222 7520 20227 7576
rect 15334 7518 20227 7520
rect 15334 7442 15394 7518
rect 20161 7515 20227 7518
rect 12574 7382 15394 7442
rect 18689 7442 18755 7445
rect 20069 7442 20135 7445
rect 18689 7440 20135 7442
rect 18689 7384 18694 7440
rect 18750 7384 20074 7440
rect 20130 7384 20135 7440
rect 18689 7382 20135 7384
rect 18689 7379 18755 7382
rect 20069 7379 20135 7382
rect 15561 7306 15627 7309
rect 21909 7306 21975 7309
rect 3926 7246 10794 7306
rect 10277 7104 10597 7105
rect 0 7034 480 7064
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 4061 7034 4127 7037
rect 0 7032 4127 7034
rect 0 6976 4066 7032
rect 4122 6976 4127 7032
rect 0 6974 4127 6976
rect 10734 7034 10794 7246
rect 15561 7304 21975 7306
rect 15561 7248 15566 7304
rect 15622 7248 21914 7304
rect 21970 7248 21975 7304
rect 15561 7246 21975 7248
rect 15561 7243 15627 7246
rect 21909 7243 21975 7246
rect 24669 7306 24735 7309
rect 27520 7306 28000 7336
rect 24669 7304 28000 7306
rect 24669 7248 24674 7304
rect 24730 7248 28000 7304
rect 24669 7246 28000 7248
rect 24669 7243 24735 7246
rect 27520 7216 28000 7246
rect 10869 7170 10935 7173
rect 16205 7170 16271 7173
rect 10869 7168 16271 7170
rect 10869 7112 10874 7168
rect 10930 7112 16210 7168
rect 16266 7112 16271 7168
rect 10869 7110 16271 7112
rect 10869 7107 10935 7110
rect 16205 7107 16271 7110
rect 20989 7170 21055 7173
rect 25497 7170 25563 7173
rect 20989 7168 25563 7170
rect 20989 7112 20994 7168
rect 21050 7112 25502 7168
rect 25558 7112 25563 7168
rect 20989 7110 25563 7112
rect 20989 7107 21055 7110
rect 25497 7107 25563 7110
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 19425 7034 19491 7037
rect 10734 7032 19491 7034
rect 10734 6976 19430 7032
rect 19486 6976 19491 7032
rect 10734 6974 19491 6976
rect 0 6944 480 6974
rect 4061 6971 4127 6974
rect 19425 6971 19491 6974
rect 20345 7034 20411 7037
rect 20805 7034 20871 7037
rect 20345 7032 20871 7034
rect 20345 6976 20350 7032
rect 20406 6976 20810 7032
rect 20866 6976 20871 7032
rect 20345 6974 20871 6976
rect 20345 6971 20411 6974
rect 20805 6971 20871 6974
rect 22001 6898 22067 6901
rect 23289 6898 23355 6901
rect 22001 6896 23355 6898
rect 22001 6840 22006 6896
rect 22062 6840 23294 6896
rect 23350 6840 23355 6896
rect 22001 6838 23355 6840
rect 22001 6835 22067 6838
rect 23289 6835 23355 6838
rect 8201 6762 8267 6765
rect 17953 6762 18019 6765
rect 8201 6760 18019 6762
rect 8201 6704 8206 6760
rect 8262 6704 17958 6760
rect 18014 6704 18019 6760
rect 8201 6702 18019 6704
rect 8201 6699 8267 6702
rect 17953 6699 18019 6702
rect 19977 6762 20043 6765
rect 27520 6762 28000 6792
rect 19977 6760 28000 6762
rect 19977 6704 19982 6760
rect 20038 6704 28000 6760
rect 19977 6702 28000 6704
rect 19977 6699 20043 6702
rect 27520 6672 28000 6702
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 6269 6354 6335 6357
rect 11053 6354 11119 6357
rect 6269 6352 11119 6354
rect 6269 6296 6274 6352
rect 6330 6296 11058 6352
rect 11114 6296 11119 6352
rect 6269 6294 11119 6296
rect 6269 6291 6335 6294
rect 11053 6291 11119 6294
rect 13629 6354 13695 6357
rect 21357 6354 21423 6357
rect 13629 6352 21423 6354
rect 13629 6296 13634 6352
rect 13690 6296 21362 6352
rect 21418 6296 21423 6352
rect 13629 6294 21423 6296
rect 13629 6291 13695 6294
rect 21357 6291 21423 6294
rect 16757 6218 16823 6221
rect 22461 6218 22527 6221
rect 23565 6218 23631 6221
rect 16757 6216 23631 6218
rect 16757 6160 16762 6216
rect 16818 6160 22466 6216
rect 22522 6160 23570 6216
rect 23626 6160 23631 6216
rect 16757 6158 23631 6160
rect 16757 6155 16823 6158
rect 22461 6155 22527 6158
rect 23565 6155 23631 6158
rect 25405 6082 25471 6085
rect 27520 6082 28000 6112
rect 25405 6080 28000 6082
rect 25405 6024 25410 6080
rect 25466 6024 28000 6080
rect 25405 6022 28000 6024
rect 25405 6019 25471 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 27520 5992 28000 6022
rect 19610 5951 19930 5952
rect 9489 5810 9555 5813
rect 20069 5810 20135 5813
rect 9489 5808 20135 5810
rect 9489 5752 9494 5808
rect 9550 5752 20074 5808
rect 20130 5752 20135 5808
rect 9489 5750 20135 5752
rect 9489 5747 9555 5750
rect 20069 5747 20135 5750
rect 7557 5674 7623 5677
rect 12893 5674 12959 5677
rect 7557 5672 12959 5674
rect 7557 5616 7562 5672
rect 7618 5616 12898 5672
rect 12954 5616 12959 5672
rect 7557 5614 12959 5616
rect 7557 5611 7623 5614
rect 12893 5611 12959 5614
rect 21081 5674 21147 5677
rect 21081 5672 24778 5674
rect 21081 5616 21086 5672
rect 21142 5616 24778 5672
rect 21081 5614 24778 5616
rect 21081 5611 21147 5614
rect 19425 5538 19491 5541
rect 23841 5538 23907 5541
rect 19425 5536 23907 5538
rect 19425 5480 19430 5536
rect 19486 5480 23846 5536
rect 23902 5480 23907 5536
rect 19425 5478 23907 5480
rect 24718 5538 24778 5614
rect 27520 5538 28000 5568
rect 24718 5478 28000 5538
rect 19425 5475 19491 5478
rect 23841 5475 23907 5478
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 27520 5448 28000 5478
rect 24277 5407 24597 5408
rect 16481 5402 16547 5405
rect 21817 5402 21883 5405
rect 16481 5400 21883 5402
rect 16481 5344 16486 5400
rect 16542 5344 21822 5400
rect 21878 5344 21883 5400
rect 16481 5342 21883 5344
rect 16481 5339 16547 5342
rect 21817 5339 21883 5342
rect 289 5266 355 5269
rect 13169 5266 13235 5269
rect 289 5264 13235 5266
rect 289 5208 294 5264
rect 350 5208 13174 5264
rect 13230 5208 13235 5264
rect 289 5206 13235 5208
rect 289 5203 355 5206
rect 13169 5203 13235 5206
rect 19793 5266 19859 5269
rect 25405 5266 25471 5269
rect 19793 5264 25471 5266
rect 19793 5208 19798 5264
rect 19854 5208 25410 5264
rect 25466 5208 25471 5264
rect 19793 5206 25471 5208
rect 19793 5203 19859 5206
rect 25405 5203 25471 5206
rect 18873 5130 18939 5133
rect 22277 5130 22343 5133
rect 18873 5128 22343 5130
rect 18873 5072 18878 5128
rect 18934 5072 22282 5128
rect 22338 5072 22343 5128
rect 18873 5070 22343 5072
rect 18873 5067 18939 5070
rect 22277 5067 22343 5070
rect 12893 4994 12959 4997
rect 15193 4994 15259 4997
rect 12893 4992 15259 4994
rect 12893 4936 12898 4992
rect 12954 4936 15198 4992
rect 15254 4936 15259 4992
rect 12893 4934 15259 4936
rect 12893 4931 12959 4934
rect 15193 4931 15259 4934
rect 25681 4994 25747 4997
rect 27520 4994 28000 5024
rect 25681 4992 28000 4994
rect 25681 4936 25686 4992
rect 25742 4936 28000 4992
rect 25681 4934 28000 4936
rect 25681 4931 25747 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 27520 4904 28000 4934
rect 19610 4863 19930 4864
rect 1669 4722 1735 4725
rect 18321 4722 18387 4725
rect 1669 4720 18387 4722
rect 1669 4664 1674 4720
rect 1730 4664 18326 4720
rect 18382 4664 18387 4720
rect 1669 4662 18387 4664
rect 1669 4659 1735 4662
rect 18321 4659 18387 4662
rect 19793 4722 19859 4725
rect 23657 4722 23723 4725
rect 19793 4720 23723 4722
rect 19793 4664 19798 4720
rect 19854 4664 23662 4720
rect 23718 4664 23723 4720
rect 19793 4662 23723 4664
rect 19793 4659 19859 4662
rect 23657 4659 23723 4662
rect 22645 4586 22711 4589
rect 13310 4526 19396 4586
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 13310 4178 13370 4526
rect 19336 4484 19396 4526
rect 22645 4584 25146 4586
rect 22645 4528 22650 4584
rect 22706 4528 25146 4584
rect 22645 4526 25146 4528
rect 22645 4523 22711 4526
rect 19336 4450 19442 4484
rect 19793 4450 19859 4453
rect 19336 4448 19859 4450
rect 19336 4424 19798 4448
rect 19382 4392 19798 4424
rect 19854 4392 19859 4448
rect 19382 4390 19859 4392
rect 25086 4450 25146 4526
rect 27520 4450 28000 4480
rect 25086 4390 28000 4450
rect 19793 4387 19859 4390
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 27520 4360 28000 4390
rect 24277 4319 24597 4320
rect 19977 4314 20043 4317
rect 23565 4314 23631 4317
rect 19977 4312 23631 4314
rect 19977 4256 19982 4312
rect 20038 4256 23570 4312
rect 23626 4256 23631 4312
rect 19977 4254 23631 4256
rect 19977 4251 20043 4254
rect 23565 4251 23631 4254
rect 3926 4118 13370 4178
rect 13537 4178 13603 4181
rect 14825 4178 14891 4181
rect 13537 4176 14891 4178
rect 13537 4120 13542 4176
rect 13598 4120 14830 4176
rect 14886 4120 14891 4176
rect 13537 4118 14891 4120
rect 1577 4042 1643 4045
rect 3926 4042 3986 4118
rect 13537 4115 13603 4118
rect 14825 4115 14891 4118
rect 21541 4178 21607 4181
rect 27521 4178 27587 4181
rect 21541 4176 27587 4178
rect 21541 4120 21546 4176
rect 21602 4120 27526 4176
rect 27582 4120 27587 4176
rect 21541 4118 27587 4120
rect 21541 4115 21607 4118
rect 27521 4115 27587 4118
rect 1577 4040 3986 4042
rect 1577 3984 1582 4040
rect 1638 3984 3986 4040
rect 1577 3982 3986 3984
rect 6913 4042 6979 4045
rect 9305 4042 9371 4045
rect 6913 4040 9371 4042
rect 6913 3984 6918 4040
rect 6974 3984 9310 4040
rect 9366 3984 9371 4040
rect 6913 3982 9371 3984
rect 1577 3979 1643 3982
rect 6913 3979 6979 3982
rect 9305 3979 9371 3982
rect 13629 4042 13695 4045
rect 25221 4042 25287 4045
rect 13629 4040 25287 4042
rect 13629 3984 13634 4040
rect 13690 3984 25226 4040
rect 25282 3984 25287 4040
rect 13629 3982 25287 3984
rect 13629 3979 13695 3982
rect 25221 3979 25287 3982
rect 13629 3906 13695 3909
rect 15653 3906 15719 3909
rect 13629 3904 15719 3906
rect 13629 3848 13634 3904
rect 13690 3848 15658 3904
rect 15714 3848 15719 3904
rect 13629 3846 15719 3848
rect 13629 3843 13695 3846
rect 15653 3843 15719 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 933 3770 999 3773
rect 1669 3770 1735 3773
rect 933 3768 1735 3770
rect 933 3712 938 3768
rect 994 3712 1674 3768
rect 1730 3712 1735 3768
rect 933 3710 1735 3712
rect 933 3707 999 3710
rect 1669 3707 1735 3710
rect 15745 3770 15811 3773
rect 17217 3770 17283 3773
rect 15745 3768 17283 3770
rect 15745 3712 15750 3768
rect 15806 3712 17222 3768
rect 17278 3712 17283 3768
rect 15745 3710 17283 3712
rect 15745 3707 15811 3710
rect 17217 3707 17283 3710
rect 20437 3770 20503 3773
rect 21633 3770 21699 3773
rect 24853 3770 24919 3773
rect 20437 3768 21699 3770
rect 20437 3712 20442 3768
rect 20498 3712 21638 3768
rect 21694 3712 21699 3768
rect 20437 3710 21699 3712
rect 20437 3707 20503 3710
rect 21633 3707 21699 3710
rect 22510 3768 24919 3770
rect 22510 3712 24858 3768
rect 24914 3712 24919 3768
rect 22510 3710 24919 3712
rect 8017 3634 8083 3637
rect 10225 3634 10291 3637
rect 8017 3632 10291 3634
rect 8017 3576 8022 3632
rect 8078 3576 10230 3632
rect 10286 3576 10291 3632
rect 8017 3574 10291 3576
rect 8017 3571 8083 3574
rect 10225 3571 10291 3574
rect 16113 3634 16179 3637
rect 22510 3634 22570 3710
rect 24853 3707 24919 3710
rect 25037 3770 25103 3773
rect 27520 3770 28000 3800
rect 25037 3768 28000 3770
rect 25037 3712 25042 3768
rect 25098 3712 28000 3768
rect 25037 3710 28000 3712
rect 25037 3707 25103 3710
rect 27520 3680 28000 3710
rect 16113 3632 22570 3634
rect 16113 3576 16118 3632
rect 16174 3576 22570 3632
rect 16113 3574 22570 3576
rect 22645 3634 22711 3637
rect 24209 3634 24275 3637
rect 22645 3632 24275 3634
rect 22645 3576 22650 3632
rect 22706 3576 24214 3632
rect 24270 3576 24275 3632
rect 22645 3574 24275 3576
rect 16113 3571 16179 3574
rect 22645 3571 22711 3574
rect 24209 3571 24275 3574
rect 14917 3498 14983 3501
rect 16113 3498 16179 3501
rect 14917 3496 16179 3498
rect 14917 3440 14922 3496
rect 14978 3440 16118 3496
rect 16174 3440 16179 3496
rect 14917 3438 16179 3440
rect 14917 3435 14983 3438
rect 16113 3435 16179 3438
rect 18321 3498 18387 3501
rect 21081 3498 21147 3501
rect 22921 3498 22987 3501
rect 24117 3498 24183 3501
rect 18321 3496 20362 3498
rect 18321 3440 18326 3496
rect 18382 3440 20362 3496
rect 18321 3438 20362 3440
rect 18321 3435 18387 3438
rect 18873 3362 18939 3365
rect 20161 3362 20227 3365
rect 18873 3360 20227 3362
rect 18873 3304 18878 3360
rect 18934 3304 20166 3360
rect 20222 3304 20227 3360
rect 18873 3302 20227 3304
rect 20302 3362 20362 3438
rect 21081 3496 22987 3498
rect 21081 3440 21086 3496
rect 21142 3440 22926 3496
rect 22982 3440 22987 3496
rect 21081 3438 22987 3440
rect 21081 3435 21147 3438
rect 22921 3435 22987 3438
rect 23982 3496 24183 3498
rect 23982 3440 24122 3496
rect 24178 3440 24183 3496
rect 23982 3438 24183 3440
rect 23982 3362 24042 3438
rect 24117 3435 24183 3438
rect 24485 3498 24551 3501
rect 26233 3498 26299 3501
rect 24485 3496 26299 3498
rect 24485 3440 24490 3496
rect 24546 3440 26238 3496
rect 26294 3440 26299 3496
rect 24485 3438 26299 3440
rect 24485 3435 24551 3438
rect 26233 3435 26299 3438
rect 20302 3302 24042 3362
rect 18873 3299 18939 3302
rect 20161 3299 20227 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 17861 3226 17927 3229
rect 19609 3226 19675 3229
rect 27520 3226 28000 3256
rect 17861 3224 19675 3226
rect 17861 3168 17866 3224
rect 17922 3168 19614 3224
rect 19670 3168 19675 3224
rect 17861 3166 19675 3168
rect 17861 3163 17927 3166
rect 19609 3163 19675 3166
rect 25638 3166 28000 3226
rect 5533 3090 5599 3093
rect 19241 3090 19307 3093
rect 5533 3088 19307 3090
rect 5533 3032 5538 3088
rect 5594 3032 19246 3088
rect 19302 3032 19307 3088
rect 5533 3030 19307 3032
rect 5533 3027 5599 3030
rect 19241 3027 19307 3030
rect 21081 3090 21147 3093
rect 23565 3090 23631 3093
rect 21081 3088 23631 3090
rect 21081 3032 21086 3088
rect 21142 3032 23570 3088
rect 23626 3032 23631 3088
rect 21081 3030 23631 3032
rect 21081 3027 21147 3030
rect 23565 3027 23631 3030
rect 23749 3090 23815 3093
rect 25638 3090 25698 3166
rect 27520 3136 28000 3166
rect 23749 3088 25698 3090
rect 23749 3032 23754 3088
rect 23810 3032 25698 3088
rect 23749 3030 25698 3032
rect 23749 3027 23815 3030
rect 2865 2954 2931 2957
rect 17769 2954 17835 2957
rect 2865 2952 17835 2954
rect 2865 2896 2870 2952
rect 2926 2896 17774 2952
rect 17830 2896 17835 2952
rect 2865 2894 17835 2896
rect 2865 2891 2931 2894
rect 17769 2891 17835 2894
rect 18781 2954 18847 2957
rect 21541 2954 21607 2957
rect 18781 2952 21607 2954
rect 18781 2896 18786 2952
rect 18842 2896 21546 2952
rect 21602 2896 21607 2952
rect 18781 2894 21607 2896
rect 18781 2891 18847 2894
rect 21541 2891 21607 2894
rect 23381 2954 23447 2957
rect 24945 2954 25011 2957
rect 23381 2952 25011 2954
rect 23381 2896 23386 2952
rect 23442 2896 24950 2952
rect 25006 2896 25011 2952
rect 23381 2894 25011 2896
rect 23381 2891 23447 2894
rect 24945 2891 25011 2894
rect 16205 2818 16271 2821
rect 17033 2818 17099 2821
rect 18873 2818 18939 2821
rect 16205 2816 16866 2818
rect 16205 2760 16210 2816
rect 16266 2760 16866 2816
rect 16205 2758 16866 2760
rect 16205 2755 16271 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 16806 2682 16866 2758
rect 17033 2816 18939 2818
rect 17033 2760 17038 2816
rect 17094 2760 18878 2816
rect 18934 2760 18939 2816
rect 17033 2758 18939 2760
rect 17033 2755 17099 2758
rect 18873 2755 18939 2758
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 18229 2682 18295 2685
rect 16806 2680 18295 2682
rect 16806 2624 18234 2680
rect 18290 2624 18295 2680
rect 16806 2622 18295 2624
rect 18229 2619 18295 2622
rect 23013 2682 23079 2685
rect 27520 2682 28000 2712
rect 23013 2680 28000 2682
rect 23013 2624 23018 2680
rect 23074 2624 28000 2680
rect 23013 2622 28000 2624
rect 23013 2619 23079 2622
rect 27520 2592 28000 2622
rect 20621 2546 20687 2549
rect 24577 2546 24643 2549
rect 20621 2544 24643 2546
rect 20621 2488 20626 2544
rect 20682 2488 24582 2544
rect 24638 2488 24643 2544
rect 20621 2486 24643 2488
rect 20621 2483 20687 2486
rect 24577 2483 24643 2486
rect 12801 2410 12867 2413
rect 12801 2408 26986 2410
rect 12801 2352 12806 2408
rect 12862 2352 26986 2408
rect 12801 2350 26986 2352
rect 12801 2347 12867 2350
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 26926 2002 26986 2350
rect 27520 2002 28000 2032
rect 26926 1942 28000 2002
rect 27520 1912 28000 1942
rect 12249 1866 12315 1869
rect 23197 1866 23263 1869
rect 12249 1864 23263 1866
rect 12249 1808 12254 1864
rect 12310 1808 23202 1864
rect 23258 1808 23263 1864
rect 12249 1806 23263 1808
rect 12249 1803 12315 1806
rect 23197 1803 23263 1806
rect 9581 1730 9647 1733
rect 22829 1730 22895 1733
rect 9581 1728 22895 1730
rect 9581 1672 9586 1728
rect 9642 1672 22834 1728
rect 22890 1672 22895 1728
rect 9581 1670 22895 1672
rect 9581 1667 9647 1670
rect 22829 1667 22895 1670
rect 11329 1594 11395 1597
rect 21909 1594 21975 1597
rect 25589 1594 25655 1597
rect 11329 1592 21466 1594
rect 11329 1536 11334 1592
rect 11390 1536 21466 1592
rect 11329 1534 21466 1536
rect 11329 1531 11395 1534
rect 21406 1458 21466 1534
rect 21909 1592 25655 1594
rect 21909 1536 21914 1592
rect 21970 1536 25594 1592
rect 25650 1536 25655 1592
rect 21909 1534 25655 1536
rect 21909 1531 21975 1534
rect 25589 1531 25655 1534
rect 23749 1458 23815 1461
rect 21406 1456 23815 1458
rect 21406 1400 23754 1456
rect 23810 1400 23815 1456
rect 21406 1398 23815 1400
rect 23749 1395 23815 1398
rect 24669 1458 24735 1461
rect 27520 1458 28000 1488
rect 24669 1456 28000 1458
rect 24669 1400 24674 1456
rect 24730 1400 28000 1456
rect 24669 1398 28000 1400
rect 24669 1395 24735 1398
rect 27520 1368 28000 1398
rect 24761 914 24827 917
rect 27520 914 28000 944
rect 24761 912 28000 914
rect 24761 856 24766 912
rect 24822 856 28000 912
rect 24761 854 28000 856
rect 24761 851 24827 854
rect 27520 824 28000 854
rect 24117 370 24183 373
rect 27520 370 28000 400
rect 24117 368 28000 370
rect 24117 312 24122 368
rect 24178 312 28000 368
rect 24117 310 28000 312
rect 24117 307 24183 310
rect 27520 280 28000 310
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 23980 18668 24044 18732
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 23980 13152 24044 13156
rect 23980 13096 24030 13152
rect 24030 13096 24044 13152
rect 23980 13092 24044 13096
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 23979 18732 24045 18733
rect 23979 18668 23980 18732
rect 24044 18668 24045 18732
rect 23979 18667 24045 18668
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 23982 13157 24042 18667
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 23979 13156 24045 13157
rect 23979 13092 23980 13156
rect 24044 13092 24045 13156
rect 23979 13091 24045 13092
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_39
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_8  FILLER_1_51 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_59 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 774 592
use scs8hd_buf_4  mux_right_track_8.scs8hd_buf_4_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8648 0 1 2720
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.scs8hd_buf_4_0__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 9384 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_87
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_88
timestamp 1586364061
transform 1 0 9200 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_1_92
timestamp 1586364061
transform 1 0 9568 0 1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_1_98 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_105
timestamp 1586364061
transform 1 0 10764 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_101
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 314 592
use scs8hd_buf_4  mux_right_track_6.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 10856 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_112
timestamp 1586364061
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _070_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11132 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_6  FILLER_1_116
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 590 592
use scs8hd_decap_6  FILLER_0_117
timestamp 1586364061
transform 1 0 11868 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_113
timestamp 1586364061
transform 1 0 11500 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 11684 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_127
timestamp 1586364061
transform 1 0 12788 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_123
timestamp 1586364061
transform 1 0 12420 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 12604 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _072_
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_134
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_133
timestamp 1586364061
transform 1 0 13340 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_129
timestamp 1586364061
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_track_3.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 12880 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_138
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_1_142
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_141
timestamp 1586364061
transform 1 0 14076 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _091_
timestamp 1586364061
transform 1 0 14260 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_148
timestamp 1586364061
transform 1 0 14720 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_track_1.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 14812 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_155
timestamp 1586364061
transform 1 0 15364 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 15548 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_1_163
timestamp 1586364061
transform 1 0 16100 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 15916 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _089_
timestamp 1586364061
transform 1 0 16008 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_170
timestamp 1586364061
transform 1 0 16744 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_166
timestamp 1586364061
transform 1 0 16376 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 16652 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _088_
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_175
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_178
timestamp 1586364061
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _087_
timestamp 1586364061
transform 1 0 17112 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__A
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _059_
timestamp 1586364061
transform 1 0 18124 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_193
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_189
timestamp 1586364061
transform 1 0 18492 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__A
timestamp 1586364061
transform 1 0 18676 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _084_
timestamp 1586364061
transform 1 0 18584 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_194
timestamp 1586364061
transform 1 0 18952 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _060_
timestamp 1586364061
transform 1 0 19228 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_198
timestamp 1586364061
transform 1 0 19320 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_205
timestamp 1586364061
transform 1 0 19964 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_201
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__060__A
timestamp 1586364061
transform 1 0 19780 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _085_
timestamp 1586364061
transform 1 0 19688 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_6  FILLER_0_210
timestamp 1586364061
transform 1 0 20424 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_206
timestamp 1586364061
transform 1 0 20056 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20148 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 20240 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_4  mux_right_track_2.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 20332 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_215
timestamp 1586364061
transform 1 0 20884 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_0_216
timestamp 1586364061
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 21068 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_1_219
timestamp 1586364061
transform 1 0 21252 0 1 2720
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 21988 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _078_
timestamp 1586364061
transform 1 0 21712 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_229
timestamp 1586364061
transform 1 0 22172 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_232
timestamp 1586364061
transform 1 0 22448 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_228
timestamp 1586364061
transform 1 0 22080 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_track_25.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22264 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_236
timestamp 1586364061
transform 1 0 22816 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _071_
timestamp 1586364061
transform 1 0 22816 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_240
timestamp 1586364061
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_244
timestamp 1586364061
transform 1 0 23552 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_240
timestamp 1586364061
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_251
timestamp 1586364061
transform 1 0 24196 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_4  mux_bottom_track_33.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_255
timestamp 1586364061
transform 1 0 24564 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24380 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _074_
timestamp 1586364061
transform 1 0 24564 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_1_267
timestamp 1586364061
transform 1 0 25668 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_263
timestamp 1586364061
transform 1 0 25300 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_259
timestamp 1586364061
transform 1 0 24932 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 25484 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _073_
timestamp 1586364061
transform 1 0 24932 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_275
timestamp 1586364061
transform 1 0 26404 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_275
timestamp 1586364061
transform 1 0 26404 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_263
timestamp 1586364061
transform 1 0 25300 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_buf_4  mux_right_track_10.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 590 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 406 592
use scs8hd_buf_2  _095_
timestamp 1586364061
transform 1 0 12236 0 -1 3808
box -38 -48 406 592
use scs8hd_buf_4  mux_bottom_track_5.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 13340 0 -1 3808
box -38 -48 590 592
use scs8hd_decap_8  FILLER_2_125
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_139
timestamp 1586364061
transform 1 0 13892 0 -1 3808
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_2_151
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 590 592
use scs8hd_buf_2  _090_
timestamp 1586364061
transform 1 0 17204 0 -1 3808
box -38 -48 406 592
use scs8hd_buf_4  mux_bottom_track_9.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 15916 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_160
timestamp 1586364061
transform 1 0 15824 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_167
timestamp 1586364061
transform 1 0 16468 0 -1 3808
box -38 -48 774 592
use scs8hd_buf_2  _057_
timestamp 1586364061
transform 1 0 18308 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_2_179
timestamp 1586364061
transform 1 0 17572 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_8  FILLER_2_191
timestamp 1586364061
transform 1 0 18676 0 -1 3808
box -38 -48 774 592
use scs8hd_buf_2  _081_
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use scs8hd_buf_4  mux_bottom_track_17.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 19412 0 -1 3808
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20332 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_205
timestamp 1586364061
transform 1 0 19964 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_3  FILLER_2_211
timestamp 1586364061
transform 1 0 20516 0 -1 3808
box -38 -48 314 592
use scs8hd_buf_2  _079_
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_2_219
timestamp 1586364061
transform 1 0 21252 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_8  FILLER_2_231
timestamp 1586364061
transform 1 0 22356 0 -1 3808
box -38 -48 774 592
use scs8hd_buf_2  _075_
timestamp 1586364061
transform 1 0 24564 0 -1 3808
box -38 -48 406 592
use scs8hd_buf_4  mux_right_track_0.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 23828 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_245
timestamp 1586364061
transform 1 0 23644 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_249
timestamp 1586364061
transform 1 0 24012 0 -1 3808
box -38 -48 590 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_259
timestamp 1586364061
transform 1 0 24932 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_2_271
timestamp 1586364061
transform 1 0 26036 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_110
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use scs8hd_buf_4  mux_right_track_12.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 13340 0 1 3808
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 13156 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 774 592
use scs8hd_buf_2  _092_
timestamp 1586364061
transform 1 0 14720 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 14076 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 15640 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_139
timestamp 1586364061
transform 1 0 13892 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_143
timestamp 1586364061
transform 1 0 14260 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_152
timestamp 1586364061
transform 1 0 15088 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_156
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 222 592
use scs8hd_buf_4  mux_right_track_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 15824 0 1 3808
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 16560 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_166
timestamp 1586364061
transform 1 0 16376 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_170
timestamp 1586364061
transform 1 0 16744 0 1 3808
box -38 -48 1142 592
use scs8hd_buf_2  _086_
timestamp 1586364061
transform 1 0 18676 0 1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_182
timestamp 1586364061
transform 1 0 17848 0 1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_3_190
timestamp 1586364061
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_195
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _058_
timestamp 1586364061
transform 1 0 19780 0 1 3808
box -38 -48 406 592
use scs8hd_buf_2  _082_
timestamp 1586364061
transform 1 0 20884 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__058__A
timestamp 1586364061
transform 1 0 20332 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_199
timestamp 1586364061
transform 1 0 19412 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_207
timestamp 1586364061
transform 1 0 20148 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_211
timestamp 1586364061
transform 1 0 20516 0 1 3808
box -38 -48 406 592
use scs8hd_buf_2  _080_
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 21436 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 22264 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 21804 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_219
timestamp 1586364061
transform 1 0 21252 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_223
timestamp 1586364061
transform 1 0 21620 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_227
timestamp 1586364061
transform 1 0 21988 0 1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_3_236
timestamp 1586364061
transform 1 0 22816 0 1 3808
box -38 -48 406 592
use scs8hd_buf_2  _077_
timestamp 1586364061
transform 1 0 24288 0 1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 23276 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 23828 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_240
timestamp 1586364061
transform 1 0 23184 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_243
timestamp 1586364061
transform 1 0 23460 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_249
timestamp 1586364061
transform 1 0 24012 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_256
timestamp 1586364061
transform 1 0 24656 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _076_
timestamp 1586364061
transform 1 0 25392 0 1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 24840 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 25944 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 25208 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_260
timestamp 1586364061
transform 1 0 25024 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_268
timestamp 1586364061
transform 1 0 25760 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_272
timestamp 1586364061
transform 1 0 26128 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_276
timestamp 1586364061
transform 1 0 26496 0 1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_buf_2  _094_
timestamp 1586364061
transform 1 0 13340 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_4  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_6  FILLER_4_137
timestamp 1586364061
transform 1 0 13708 0 -1 4896
box -38 -48 590 592
use scs8hd_buf_2  _093_
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 14352 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 14720 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_143
timestamp 1586364061
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_146
timestamp 1586364061
transform 1 0 14536 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_150
timestamp 1586364061
transform 1 0 14904 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_158
timestamp 1586364061
transform 1 0 15640 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 15824 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 16192 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_162
timestamp 1586364061
transform 1 0 16008 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use scs8hd_conb_1  _030_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19780 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_206
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_8  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 774 592
use scs8hd_buf_2  _083_
timestamp 1586364061
transform 1 0 21804 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_223
timestamp 1586364061
transform 1 0 21620 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_229
timestamp 1586364061
transform 1 0 22172 0 -1 4896
box -38 -48 1142 592
use scs8hd_mux2_2  mux_right_track_22.mux_l1_in_1_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 23276 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 24288 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_250
timestamp 1586364061
transform 1 0 24104 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_254
timestamp 1586364061
transform 1 0 24472 0 -1 4896
box -38 -48 406 592
use scs8hd_buf_2  _069_
timestamp 1586364061
transform 1 0 24840 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_262
timestamp 1586364061
transform 1 0 25208 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_4_274
timestamp 1586364061
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use scs8hd_conb_1  _031_
timestamp 1586364061
transform 1 0 13340 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 13156 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_136
timestamp 1586364061
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_24.mux_l3_in_0_
timestamp 1586364061
transform 1 0 14352 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 15364 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 14168 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_140
timestamp 1586364061
transform 1 0 13984 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_153
timestamp 1586364061
transform 1 0 15180 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_157
timestamp 1586364061
transform 1 0 15548 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_24.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15916 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 16928 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_170
timestamp 1586364061
transform 1 0 16744 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_174
timestamp 1586364061
transform 1 0 17112 0 1 4896
box -38 -48 774 592
use scs8hd_buf_4  mux_right_track_14.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18584 0 1 4896
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 19320 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_182
timestamp 1586364061
transform 1 0 17848 0 1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 590 592
use scs8hd_fill_2  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 222 592
use scs8hd_buf_4  mux_right_track_16.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 20700 0 1 4896
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 20516 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20148 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 19688 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_200
timestamp 1586364061
transform 1 0 19504 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_204
timestamp 1586364061
transform 1 0 19872 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_209
timestamp 1586364061
transform 1 0 20332 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _068_
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 21436 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 22264 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_219
timestamp 1586364061
transform 1 0 21252 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_223
timestamp 1586364061
transform 1 0 21620 0 1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_5_229
timestamp 1586364061
transform 1 0 22172 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_236
timestamp 1586364061
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_22.mux_l2_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_22.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_22.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 24656 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_240
timestamp 1586364061
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_254
timestamp 1586364061
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use scs8hd_buf_4  mux_right_track_22.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 25208 0 1 4896
box -38 -48 590 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 25024 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 25944 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_258
timestamp 1586364061
transform 1 0 24840 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_268
timestamp 1586364061
transform 1 0 25760 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_272
timestamp 1586364061
transform 1 0 26128 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_276
timestamp 1586364061
transform 1 0 26496 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__061__A
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_77
timestamp 1586364061
transform 1 0 8188 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_89
timestamp 1586364061
transform 1 0 9292 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_101
timestamp 1586364061
transform 1 0 10396 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_113
timestamp 1586364061
transform 1 0 11500 0 1 5984
box -38 -48 774 592
use scs8hd_mux2_2  mux_right_track_24.mux_l2_in_1_
timestamp 1586364061
transform 1 0 13616 0 -1 5984
box -38 -48 866 592
use scs8hd_buf_4  mux_right_track_24.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 13340 0 1 5984
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_135
timestamp 1586364061
transform 1 0 13524 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_121
timestamp 1586364061
transform 1 0 12236 0 1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_131
timestamp 1586364061
transform 1 0 13156 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_143
timestamp 1586364061
transform 1 0 14260 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_139
timestamp 1586364061
transform 1 0 13892 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14076 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 14444 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_149
timestamp 1586364061
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_2_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_26.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 16560 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_26.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 16928 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_173
timestamp 1586364061
transform 1 0 17020 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_166
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_170
timestamp 1586364061
transform 1 0 16744 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_174
timestamp 1586364061
transform 1 0 17112 0 1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_180
timestamp 1586364061
transform 1 0 17664 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_6_186
timestamp 1586364061
transform 1 0 18216 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_6_181
timestamp 1586364061
transform 1 0 17756 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_26.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 18032 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_26.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_195
timestamp 1586364061
transform 1 0 19044 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_191
timestamp 1586364061
transform 1 0 18676 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 19228 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 18860 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 18492 0 -1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_26.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_7_207
timestamp 1586364061
transform 1 0 20148 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_203
timestamp 1586364061
transform 1 0 19780 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_206
timestamp 1586364061
transform 1 0 20056 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_6_199
timestamp 1586364061
transform 1 0 19412 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 19964 0 1 5984
box -38 -48 222 592
use scs8hd_buf_2  _064_
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_213
timestamp 1586364061
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_210
timestamp 1586364061
transform 1 0 20424 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 20516 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 20332 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 20516 0 1 5984
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 22908 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 22540 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_234
timestamp 1586364061
transform 1 0 22632 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_7_230
timestamp 1586364061
transform 1 0 22264 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_235
timestamp 1586364061
transform 1 0 22724 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_22.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 24104 0 1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_right_track_22.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 23368 0 -1 5984
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 23920 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 23276 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_239
timestamp 1586364061
transform 1 0 23092 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_243
timestamp 1586364061
transform 1 0 23460 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_6_265
timestamp 1586364061
transform 1 0 25484 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_6_261
timestamp 1586364061
transform 1 0 25116 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_273
timestamp 1586364061
transform 1 0 26220 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_273
timestamp 1586364061
transform 1 0 26220 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 26036 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use scs8hd_buf_2  _061_
timestamp 1586364061
transform 1 0 8004 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_6  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_74
timestamp 1586364061
transform 1 0 7912 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_79
timestamp 1586364061
transform 1 0 8372 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_91
timestamp 1586364061
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 14536 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_141
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_148
timestamp 1586364061
transform 1 0 14720 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_152
timestamp 1586364061
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_right_track_26.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 16008 0 -1 7072
box -38 -48 1786 592
use scs8hd_mux2_2  mux_right_track_26.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18492 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_181
timestamp 1586364061
transform 1 0 17756 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_186
timestamp 1586364061
transform 1 0 18216 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_198
timestamp 1586364061
transform 1 0 19320 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_2  _066_
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 19504 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 19872 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 20516 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_206
timestamp 1586364061
transform 1 0 20056 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_210
timestamp 1586364061
transform 1 0 20424 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_213
timestamp 1586364061
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use scs8hd_buf_4  mux_right_track_18.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22724 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 21436 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_219
timestamp 1586364061
transform 1 0 21252 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_223
timestamp 1586364061
transform 1 0 21620 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_233
timestamp 1586364061
transform 1 0 22540 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_237
timestamp 1586364061
transform 1 0 22908 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_22.mux_l1_in_0_
timestamp 1586364061
transform 1 0 23276 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_22.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 24288 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_22.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 24656 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_250
timestamp 1586364061
transform 1 0 24104 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_254
timestamp 1586364061
transform 1 0 24472 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_20.mux_l1_in_0_
timestamp 1586364061
transform 1 0 24840 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_267
timestamp 1586364061
transform 1 0 25668 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_51
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_59
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_110
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 774 592
use scs8hd_mux2_2  mux_right_track_24.mux_l1_in_0_
timestamp 1586364061
transform 1 0 14536 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 14352 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_143
timestamp 1586364061
transform 1 0 14260 0 1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_155
timestamp 1586364061
transform 1 0 15364 0 1 7072
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_track_26.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_159
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_162
timestamp 1586364061
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_16.mux_l2_in_0_
timestamp 1586364061
transform 1 0 20516 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 19964 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 20332 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_203
timestamp 1586364061
transform 1 0 19780 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_207
timestamp 1586364061
transform 1 0 20148 0 1 7072
box -38 -48 222 592
use scs8hd_buf_4  mux_right_track_20.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22264 0 1 7072
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 21528 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 21896 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_220
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_224
timestamp 1586364061
transform 1 0 21712 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_228
timestamp 1586364061
transform 1 0 22080 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_236
timestamp 1586364061
transform 1 0 22816 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_20.mux_l2_in_0_
timestamp 1586364061
transform 1 0 23920 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_20.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_240
timestamp 1586364061
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _067_
timestamp 1586364061
transform 1 0 25484 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_20.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 24932 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 26036 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 25300 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_261
timestamp 1586364061
transform 1 0 25116 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_273
timestamp 1586364061
transform 1 0 26220 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_56
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_80
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_117
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14536 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_141
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_148
timestamp 1586364061
transform 1 0 14720 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_152
timestamp 1586364061
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use scs8hd_conb_1  _032_
timestamp 1586364061
transform 1 0 16928 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16744 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_168
timestamp 1586364061
transform 1 0 16560 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_175
timestamp 1586364061
transform 1 0 17204 0 -1 8160
box -38 -48 774 592
use scs8hd_mux2_2  mux_right_track_16.mux_l1_in_1_
timestamp 1586364061
transform 1 0 19228 0 -1 8160
box -38 -48 866 592
use scs8hd_buf_4  mux_right_track_26.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 17940 0 -1 8160
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_26.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 18676 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_189
timestamp 1586364061
transform 1 0 18492 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_193
timestamp 1586364061
transform 1 0 18860 0 -1 8160
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_16.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 20516 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_206
timestamp 1586364061
transform 1 0 20056 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_210
timestamp 1586364061
transform 1 0 20424 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_213
timestamp 1586364061
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_18.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 22816 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_234
timestamp 1586364061
transform 1 0 22632 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_238
timestamp 1586364061
transform 1 0 23000 0 -1 8160
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_20.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 23920 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_20.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 23644 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 23276 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_243
timestamp 1586364061
transform 1 0 23460 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_247
timestamp 1586364061
transform 1 0 23828 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_267
timestamp 1586364061
transform 1 0 25668 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_39
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_98
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_110
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_147
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_11_155
timestamp 1586364061
transform 1 0 15364 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_158
timestamp 1586364061
transform 1 0 15640 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 15824 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_162
timestamp 1586364061
transform 1 0 16008 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_175
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_179
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 18308 0 1 8160
box -38 -48 222 592
use scs8hd_conb_1  _054_
timestamp 1586364061
transform 1 0 18492 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_192
timestamp 1586364061
transform 1 0 18768 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_196
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 18952 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 19320 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_18.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 21068 0 1 8160
box -38 -48 1786 592
use scs8hd_mux2_2  mux_right_track_16.mux_l1_in_0_
timestamp 1586364061
transform 1 0 19504 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_18.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 20884 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 20516 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_209
timestamp 1586364061
transform 1 0 20332 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_213
timestamp 1586364061
transform 1 0 20700 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_18.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_236
timestamp 1586364061
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_20.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_20.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_240
timestamp 1586364061
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 25576 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 25944 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 26312 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_264
timestamp 1586364061
transform 1 0 25392 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_268
timestamp 1586364061
transform 1 0 25760 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_272
timestamp 1586364061
transform 1 0 26128 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_276
timestamp 1586364061
transform 1 0 26496 0 1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 13340 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 13708 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_131
timestamp 1586364061
transform 1 0 13156 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_135
timestamp 1586364061
transform 1 0 13524 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_139
timestamp 1586364061
transform 1 0 13892 0 -1 9248
box -38 -48 590 592
use scs8hd_decap_6  FILLER_12_147
timestamp 1586364061
transform 1 0 14628 0 -1 9248
box -38 -48 590 592
use scs8hd_decap_8  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 774 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l3_in_0_
timestamp 1586364061
transform 1 0 16284 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  FILLER_12_162
timestamp 1586364061
transform 1 0 16008 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_174
timestamp 1586364061
transform 1 0 17112 0 -1 9248
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_right_track_16.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18308 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_182
timestamp 1586364061
transform 1 0 17848 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_186
timestamp 1586364061
transform 1 0 18216 0 -1 9248
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_18.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 21068 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_206
timestamp 1586364061
transform 1 0 20056 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_210
timestamp 1586364061
transform 1 0 20424 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_2  _062_
timestamp 1586364061
transform 1 0 21252 0 -1 9248
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_18.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 22356 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_223
timestamp 1586364061
transform 1 0 21620 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_229
timestamp 1586364061
transform 1 0 22172 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 24288 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 24656 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_250
timestamp 1586364061
transform 1 0 24104 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_254
timestamp 1586364061
transform 1 0 24472 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_20.mux_l1_in_1_
timestamp 1586364061
transform 1 0 24840 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_267
timestamp 1586364061
transform 1 0 25668 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_74
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_98
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 10856 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_110
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_105
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_108
timestamp 1586364061
transform 1 0 11040 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_14_128
timestamp 1586364061
transform 1 0 12880 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_120
timestamp 1586364061
transform 1 0 12144 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 12696 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l2_in_1_
timestamp 1586364061
transform 1 0 12880 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_138
timestamp 1586364061
transform 1 0 13800 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_137
timestamp 1586364061
transform 1 0 13708 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l3_in_0_
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_8  FILLER_14_142
timestamp 1586364061
transform 1 0 14168 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_141
timestamp 1586364061
transform 1 0 14076 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 13892 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 13984 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_158
timestamp 1586364061
transform 1 0 15640 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_3  FILLER_14_150
timestamp 1586364061
transform 1 0 14904 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 14444 0 1 9248
box -38 -48 1786 592
use scs8hd_conb_1  _049_
timestamp 1586364061
transform 1 0 16928 0 1 9248
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15916 0 -1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 16376 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 16744 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 15732 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_164
timestamp 1586364061
transform 1 0 16192 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_168
timestamp 1586364061
transform 1 0 16560 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1786 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l1_in_2_
timestamp 1586364061
transform 1 0 18400 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 18216 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_180
timestamp 1586364061
transform 1 0 17664 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_197
timestamp 1586364061
transform 1 0 19228 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_201
timestamp 1586364061
transform 1 0 19596 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_13_207
timestamp 1586364061
transform 1 0 20148 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_203
timestamp 1586364061
transform 1 0 19780 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 19412 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 19964 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_209
timestamp 1586364061
transform 1 0 20332 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_212
timestamp 1586364061
transform 1 0 20608 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 20424 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 20792 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_17.mux_l3_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use scs8hd_conb_1  _029_
timestamp 1586364061
transform 1 0 20976 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_228
timestamp 1586364061
transform 1 0 22080 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_224
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_223
timestamp 1586364061
transform 1 0 21620 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_219
timestamp 1586364061
transform 1 0 21252 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 21896 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 21436 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 21804 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_18.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21988 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_236
timestamp 1586364061
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 22264 0 -1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_18.mux_l1_in_1_
timestamp 1586364061
transform 1 0 22448 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_247
timestamp 1586364061
transform 1 0 23828 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_241
timestamp 1586364061
transform 1 0 23276 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_240
timestamp 1586364061
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 23644 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_18.mux_l1_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_254
timestamp 1586364061
transform 1 0 24472 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 24656 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_33.mux_l2_in_0_
timestamp 1586364061
transform 1 0 24012 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_8  FILLER_14_264
timestamp 1586364061
transform 1 0 25392 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_4  FILLER_14_258
timestamp 1586364061
transform 1 0 24840 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_266
timestamp 1586364061
transform 1 0 25576 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_258
timestamp 1586364061
transform 1 0 24840 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 25208 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 25024 0 1 9248
box -38 -48 222 592
use scs8hd_buf_2  _065_
timestamp 1586364061
transform 1 0 25208 0 1 9248
box -38 -48 406 592
use scs8hd_decap_3  FILLER_14_272
timestamp 1586364061
transform 1 0 26128 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_6  FILLER_13_270
timestamp 1586364061
transform 1 0 25944 0 1 9248
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 25760 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_276
timestamp 1586364061
transform 1 0 26496 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 406 592
use scs8hd_conb_1  _048_
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10856 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10488 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_104
timestamp 1586364061
transform 1 0 10672 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_108
timestamp 1586364061
transform 1 0 11040 0 1 10336
box -38 -48 314 592
use scs8hd_decap_6  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 13064 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12604 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_127
timestamp 1586364061
transform 1 0 12788 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_151
timestamp 1586364061
transform 1 0 14996 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_155
timestamp 1586364061
transform 1 0 15364 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_158
timestamp 1586364061
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l2_in_1_
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_162
timestamp 1586364061
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_17.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18952 0 1 10336
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 18216 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 18584 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_188
timestamp 1586364061
transform 1 0 18400 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_192
timestamp 1586364061
transform 1 0 18768 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 20884 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_213
timestamp 1586364061
transform 1 0 20700 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_217
timestamp 1586364061
transform 1 0 21068 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_17.mux_l1_in_0_
timestamp 1586364061
transform 1 0 21436 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 21252 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_230
timestamp 1586364061
transform 1 0 22264 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_234
timestamp 1586364061
transform 1 0 22632 0 1 10336
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_track_33.mux_l1_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 24656 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_240
timestamp 1586364061
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_254
timestamp 1586364061
transform 1 0 24472 0 1 10336
box -38 -48 222 592
use scs8hd_buf_2  _063_
timestamp 1586364061
transform 1 0 25208 0 1 10336
box -38 -48 406 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 25760 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_258
timestamp 1586364061
transform 1 0 24840 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_266
timestamp 1586364061
transform 1 0 25576 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_270
timestamp 1586364061
transform 1 0 25944 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_276
timestamp 1586364061
transform 1 0 26496 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10856 0 -1 11424
box -38 -48 866 592
use scs8hd_fill_1  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_115
timestamp 1586364061
transform 1 0 11684 0 -1 11424
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12420 0 -1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 12236 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 15456 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 14812 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_142
timestamp 1586364061
transform 1 0 14168 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_148
timestamp 1586364061
transform 1 0 14720 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_151
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_158
timestamp 1586364061
transform 1 0 15640 0 -1 11424
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l2_in_0_
timestamp 1586364061
transform 1 0 16468 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 16284 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 15916 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_163
timestamp 1586364061
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_176
timestamp 1586364061
transform 1 0 17296 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l1_in_1_
timestamp 1586364061
transform 1 0 18032 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 19044 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17848 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_180
timestamp 1586364061
transform 1 0 17664 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_193
timestamp 1586364061
transform 1 0 18860 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_197
timestamp 1586364061
transform 1 0 19228 0 -1 11424
box -38 -48 590 592
use scs8hd_conb_1  _055_
timestamp 1586364061
transform 1 0 19780 0 -1 11424
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_track_17.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_206
timestamp 1586364061
transform 1 0 20056 0 -1 11424
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 22816 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_234
timestamp 1586364061
transform 1 0 22632 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_238
timestamp 1586364061
transform 1 0 23000 0 -1 11424
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_bottom_track_33.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 23920 0 -1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 23644 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_244
timestamp 1586364061
transform 1 0 23552 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_247
timestamp 1586364061
transform 1 0 23828 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_267
timestamp 1586364061
transform 1 0 25668 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_98
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 12052 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 11316 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_110
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_113
timestamp 1586364061
transform 1 0 11500 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_117
timestamp 1586364061
transform 1 0 11868 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12880 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 12696 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_121
timestamp 1586364061
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_137
timestamp 1586364061
transform 1 0 13708 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l3_in_0_
timestamp 1586364061
transform 1 0 14812 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 13892 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_141
timestamp 1586364061
transform 1 0 14076 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_145
timestamp 1586364061
transform 1 0 14444 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_158
timestamp 1586364061
transform 1 0 15640 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l2_in_1_
timestamp 1586364061
transform 1 0 16376 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_162
timestamp 1586364061
transform 1 0 16008 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_175
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l1_in_2_
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_179
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_193
timestamp 1586364061
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_197
timestamp 1586364061
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _044_
timestamp 1586364061
transform 1 0 20056 0 1 11424
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_track_17.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 21068 0 1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 20516 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 19412 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_201
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_205
timestamp 1586364061
transform 1 0 19964 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_209
timestamp 1586364061
transform 1 0 20332 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_213
timestamp 1586364061
transform 1 0 20700 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_236
timestamp 1586364061
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_33.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 24104 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23920 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_240
timestamp 1586364061
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l1_in_1_
timestamp 1586364061
transform 1 0 11684 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_18_105
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_113
timestamp 1586364061
transform 1 0 11500 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l1_in_2_
timestamp 1586364061
transform 1 0 13248 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 12880 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_124
timestamp 1586364061
transform 1 0 12512 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_130
timestamp 1586364061
transform 1 0 13064 0 -1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 15364 0 -1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14260 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_149
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17296 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_174
timestamp 1586364061
transform 1 0 17112 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_178
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 17848 0 -1 12512
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 17664 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_17.mux_l1_in_1_
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_201
timestamp 1586364061
transform 1 0 19596 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_205
timestamp 1586364061
transform 1 0 19964 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_208
timestamp 1586364061
transform 1 0 20240 0 -1 12512
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 22448 0 -1 12512
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 21896 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_224
timestamp 1586364061
transform 1 0 21712 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_228
timestamp 1586364061
transform 1 0 22080 0 -1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 24748 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 24380 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_255
timestamp 1586364061
transform 1 0 24564 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_2  _056_
timestamp 1586364061
transform 1 0 24932 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_68
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_80
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_105
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_106
timestamp 1586364061
transform 1 0 10856 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11040 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_111
timestamp 1586364061
transform 1 0 11316 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 11408 0 -1 13600
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13800 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_131
timestamp 1586364061
transform 1 0 13156 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_20_137
timestamp 1586364061
transform 1 0 13708 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_20_148
timestamp 1586364061
transform 1 0 14720 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_144
timestamp 1586364061
transform 1 0 14352 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_140
timestamp 1586364061
transform 1 0 13984 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_148
timestamp 1586364061
transform 1 0 14720 0 1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_19_142
timestamp 1586364061
transform 1 0 14168 0 1 12512
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14536 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14168 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_158
timestamp 1586364061
transform 1 0 15640 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 14812 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 14996 0 1 12512
box -38 -48 1786 592
use scs8hd_conb_1  _043_
timestamp 1586364061
transform 1 0 15732 0 -1 13600
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 16744 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 16376 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 16928 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_170
timestamp 1586364061
transform 1 0 16744 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_174
timestamp 1586364061
transform 1 0 17112 0 1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_162
timestamp 1586364061
transform 1 0 16008 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_168
timestamp 1586364061
transform 1 0 16560 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_186
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_183
timestamp 1586364061
transform 1 0 17940 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_179
timestamp 1586364061
transform 1 0 17572 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 18032 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l1_in_1_
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_196
timestamp 1586364061
transform 1 0 19136 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_197
timestamp 1586364061
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_193
timestamp 1586364061
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 19320 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 19780 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 19688 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_201
timestamp 1586364061
transform 1 0 19596 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_200
timestamp 1586364061
transform 1 0 19504 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_205
timestamp 1586364061
transform 1 0 19964 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_204
timestamp 1586364061
transform 1 0 19872 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_208
timestamp 1586364061
transform 1 0 20240 0 -1 13600
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_17.mux_l2_in_0_
timestamp 1586364061
transform 1 0 20056 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_212
timestamp 1586364061
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_215
timestamp 1586364061
transform 1 0 20884 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 20424 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 21068 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_17.mux_l2_in_1_
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_219
timestamp 1586364061
transform 1 0 21252 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 21436 0 1 12512
box -38 -48 222 592
use scs8hd_conb_1  _036_
timestamp 1586364061
transform 1 0 21620 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_224
timestamp 1586364061
transform 1 0 21712 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_226
timestamp 1586364061
transform 1 0 21896 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 21988 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_229
timestamp 1586364061
transform 1 0 22172 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_230
timestamp 1586364061
transform 1 0 22264 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 22356 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 22080 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_237
timestamp 1586364061
transform 1 0 22908 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_233
timestamp 1586364061
transform 1 0 22540 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_236
timestamp 1586364061
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 22632 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 23000 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_240
timestamp 1586364061
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_33.mux_l1_in_1_
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l1_in_0_
timestamp 1586364061
transform 1 0 23184 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_253
timestamp 1586364061
transform 1 0 24380 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_249
timestamp 1586364061
transform 1 0 24012 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_254
timestamp 1586364061
transform 1 0 24472 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 24564 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 24196 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l2_in_1_
timestamp 1586364061
transform 1 0 24748 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_8  FILLER_20_266
timestamp 1586364061
transform 1 0 25576 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_265
timestamp 1586364061
transform 1 0 25484 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_259
timestamp 1586364061
transform 1 0 24932 0 1 12512
box -38 -48 314 592
use scs8hd_conb_1  _047_
timestamp 1586364061
transform 1 0 25208 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_274
timestamp 1586364061
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 25668 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_39
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_21_59
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_74
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_86
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_98
timestamp 1586364061
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 12052 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 11684 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_110
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_117
timestamp 1586364061
transform 1 0 11868 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_121
timestamp 1586364061
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 12604 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_conb_1  _046_
timestamp 1586364061
transform 1 0 12788 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_134
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_130
timestamp 1586364061
transform 1 0 13064 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 13800 0 1 13600
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_21_157
timestamp 1586364061
transform 1 0 15548 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_2.mux_l1_in_1_
timestamp 1586364061
transform 1 0 16376 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 16192 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_161
timestamp 1586364061
transform 1 0 15916 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_175
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 18860 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 18676 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 18308 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_179
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_189
timestamp 1586364061
transform 1 0 18492 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 20424 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 19872 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_202
timestamp 1586364061
transform 1 0 19688 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_206
timestamp 1586364061
transform 1 0 20056 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l3_in_0_
timestamp 1586364061
transform 1 0 21988 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 21436 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 21804 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_219
timestamp 1586364061
transform 1 0 21252 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_223
timestamp 1586364061
transform 1 0 21620 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_236
timestamp 1586364061
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 24104 0 1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 23920 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_240
timestamp 1586364061
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_44
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_56
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_68
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_80
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l3_in_0_
timestamp 1586364061
transform 1 0 12052 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_12  FILLER_22_105
timestamp 1586364061
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_22_117
timestamp 1586364061
transform 1 0 11868 0 -1 14688
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 13340 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_128
timestamp 1586364061
transform 1 0 12880 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_132
timestamp 1586364061
transform 1 0 13248 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_135
timestamp 1586364061
transform 1 0 13524 0 -1 14688
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l1_in_1_
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_145
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_163
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_168
timestamp 1586364061
transform 1 0 16560 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  FILLER_22_176
timestamp 1586364061
transform 1 0 17296 0 -1 14688
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 17756 0 -1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 17572 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 20424 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 19688 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_200
timestamp 1586364061
transform 1 0 19504 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_204
timestamp 1586364061
transform 1 0 19872 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_208
timestamp 1586364061
transform 1 0 20240 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_212
timestamp 1586364061
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 22816 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_234
timestamp 1586364061
transform 1 0 22632 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_238
timestamp 1586364061
transform 1 0 23000 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 23736 0 -1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 23552 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 23184 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_242
timestamp 1586364061
transform 1 0 23368 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_265
timestamp 1586364061
transform 1 0 25484 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_273
timestamp 1586364061
transform 1 0 26220 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_59
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_74
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_86
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_98
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_110
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 13340 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 12972 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 12604 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_127
timestamp 1586364061
transform 1 0 12788 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_131
timestamp 1586364061
transform 1 0 13156 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_2.mux_l2_in_1_
timestamp 1586364061
transform 1 0 15272 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 15088 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 14720 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_144
timestamp 1586364061
transform 1 0 14352 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_150
timestamp 1586364061
transform 1 0 14904 0 1 14688
box -38 -48 222 592
use scs8hd_conb_1  _038_
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 16284 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 16652 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_163
timestamp 1586364061
transform 1 0 16100 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_167
timestamp 1586364061
transform 1 0 16468 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_174
timestamp 1586364061
transform 1 0 17112 0 1 14688
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 18676 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 18492 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_188
timestamp 1586364061
transform 1 0 18400 0 1 14688
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 20056 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 19688 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_200
timestamp 1586364061
transform 1 0 19504 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_204
timestamp 1586364061
transform 1 0 19872 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 22448 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_227
timestamp 1586364061
transform 1 0 21988 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_231
timestamp 1586364061
transform 1 0 22356 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_234
timestamp 1586364061
transform 1 0 22632 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_238
timestamp 1586364061
transform 1 0 23000 0 1 14688
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l2_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 24656 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_254
timestamp 1586364061
transform 1 0 24472 0 1 14688
box -38 -48 222 592
use scs8hd_conb_1  _045_
timestamp 1586364061
transform 1 0 25208 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 25024 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_258
timestamp 1586364061
transform 1 0 24840 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_265
timestamp 1586364061
transform 1 0 25484 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_56
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9844 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_97
timestamp 1586364061
transform 1 0 10028 0 -1 15776
box -38 -48 774 592
use scs8hd_mux2_2  mux_top_track_4.mux_l1_in_0_
timestamp 1586364061
transform 1 0 11776 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_107
timestamp 1586364061
transform 1 0 10948 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_1  FILLER_24_115
timestamp 1586364061
transform 1 0 11684 0 -1 15776
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l2_in_1_
timestamp 1586364061
transform 1 0 13340 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 13156 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_125
timestamp 1586364061
transform 1 0 12604 0 -1 15776
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14352 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_142
timestamp 1586364061
transform 1 0 14168 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_146
timestamp 1586364061
transform 1 0 14536 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_150
timestamp 1586364061
transform 1 0 14904 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17204 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_173
timestamp 1586364061
transform 1 0 17020 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_177
timestamp 1586364061
transform 1 0 17388 0 -1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 17756 0 -1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 17572 0 -1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 19872 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 20240 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_200
timestamp 1586364061
transform 1 0 19504 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_206
timestamp 1586364061
transform 1 0 20056 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_210
timestamp 1586364061
transform 1 0 20424 0 -1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_24.mux_l2_in_1_
timestamp 1586364061
transform 1 0 22448 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 21896 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 22264 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_224
timestamp 1586364061
transform 1 0 21712 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_228
timestamp 1586364061
transform 1 0 22080 0 -1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l1_in_1_
timestamp 1586364061
transform 1 0 24288 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 24012 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 23644 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_241
timestamp 1586364061
transform 1 0 23276 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_247
timestamp 1586364061
transform 1 0 23828 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_251
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 25300 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_261
timestamp 1586364061
transform 1 0 25116 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_265
timestamp 1586364061
transform 1 0 25484 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_273
timestamp 1586364061
transform 1 0 26220 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_74
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 10212 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9844 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9476 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_86
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_90
timestamp 1586364061
transform 1 0 9384 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_93
timestamp 1586364061
transform 1 0 9660 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_97
timestamp 1586364061
transform 1 0 10028 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_4.mux_l1_in_2_
timestamp 1586364061
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_101
timestamp 1586364061
transform 1 0 10396 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 13616 0 1 15776
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 13064 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 12604 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_127
timestamp 1586364061
transform 1 0 12788 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_132
timestamp 1586364061
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 15548 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_155
timestamp 1586364061
transform 1 0 15364 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_2.mux_l2_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 16192 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_159
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_163
timestamp 1586364061
transform 1 0 16100 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_175
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_24.mux_l1_in_0_
timestamp 1586364061
transform 1 0 18308 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 19320 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_179
timestamp 1586364061
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_196
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 19872 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 19688 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_200
timestamp 1586364061
transform 1 0 19504 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_213
timestamp 1586364061
transform 1 0 20700 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_217
timestamp 1586364061
transform 1 0 21068 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 21436 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 21252 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_230
timestamp 1586364061
transform 1 0 22264 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_234
timestamp 1586364061
transform 1 0 22632 0 1 15776
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_top_track_32.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 24012 0 1 15776
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 23828 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 25944 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_268
timestamp 1586364061
transform 1 0 25760 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_272
timestamp 1586364061
transform 1 0 26128 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_276
timestamp 1586364061
transform 1 0 26496 0 1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_27_86
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_96
timestamp 1586364061
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_92
timestamp 1586364061
transform 1 0 9568 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 9384 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9844 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_12  FILLER_26_80
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_27_100
timestamp 1586364061
transform 1 0 10304 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_108
timestamp 1586364061
transform 1 0 11040 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_104
timestamp 1586364061
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 10856 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_4.mux_l2_in_1_
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11224 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11408 0 -1 16864
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_4.mux_l3_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_136
timestamp 1586364061
transform 1 0 13616 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_138
timestamp 1586364061
transform 1 0 13800 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_135
timestamp 1586364061
transform 1 0 13524 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_131
timestamp 1586364061
transform 1 0 13156 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 13432 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 13616 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_145
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14628 0 -1 16864
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_4.mux_l1_in_1_
timestamp 1586364061
transform 1 0 13984 0 1 16864
box -38 -48 866 592
use scs8hd_buf_4  mux_top_track_2.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 13892 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_156
timestamp 1586364061
transform 1 0 15456 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_153
timestamp 1586364061
transform 1 0 15180 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_149
timestamp 1586364061
transform 1 0 14812 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_149
timestamp 1586364061
transform 1 0 14812 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 15640 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 15272 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_2.mux_l3_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_4  FILLER_27_160
timestamp 1586364061
transform 1 0 15824 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_168
timestamp 1586364061
transform 1 0 16560 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_163
timestamp 1586364061
transform 1 0 16100 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16376 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16192 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_2.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_175
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_172
timestamp 1586364061
transform 1 0 16928 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 16744 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use scs8hd_buf_4  mux_top_track_0.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 17020 0 -1 16864
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 17756 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_179
timestamp 1586364061
transform 1 0 17572 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_183
timestamp 1586364061
transform 1 0 17940 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_179
timestamp 1586364061
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 18308 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 18124 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_16.mux_l1_in_1_
timestamp 1586364061
transform 1 0 18308 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_198
timestamp 1586364061
transform 1 0 19320 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_196
timestamp 1586364061
transform 1 0 19136 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 19320 0 -1 16864
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_16.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18492 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_202
timestamp 1586364061
transform 1 0 19688 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_208
timestamp 1586364061
transform 1 0 20240 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_204
timestamp 1586364061
transform 1 0 19872 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_200
timestamp 1586364061
transform 1 0 19504 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 19504 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 20056 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 19872 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_16.mux_l1_in_0_
timestamp 1586364061
transform 1 0 20056 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_215
timestamp 1586364061
transform 1 0 20884 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_212
timestamp 1586364061
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 21068 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 21068 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_27_223
timestamp 1586364061
transform 1 0 21620 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_219
timestamp 1586364061
transform 1 0 21252 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_223
timestamp 1586364061
transform 1 0 21620 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_219
timestamp 1586364061
transform 1 0 21252 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 21712 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 21436 0 -1 16864
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_24.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21896 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_235
timestamp 1586364061
transform 1 0 22724 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 22908 0 1 16864
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 21804 0 -1 16864
box -38 -48 1786 592
use scs8hd_decap_3  FILLER_27_239
timestamp 1586364061
transform 1 0 23092 0 1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_26_244
timestamp 1586364061
transform 1 0 23552 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_254
timestamp 1586364061
transform 1 0 24472 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_250
timestamp 1586364061
transform 1 0 24104 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 24288 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23920 0 -1 16864
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_32.mux_l1_in_0_
timestamp 1586364061
transform 1 0 24564 0 -1 16864
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 1786 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_264
timestamp 1586364061
transform 1 0 25392 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_26_272
timestamp 1586364061
transform 1 0 26128 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_264
timestamp 1586364061
transform 1 0 25392 0 1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_27_276
timestamp 1586364061
transform 1 0 26496 0 1 16864
box -38 -48 130 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use scs8hd_mux2_2  mux_top_track_8.mux_l1_in_2_
timestamp 1586364061
transform 1 0 9752 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_88
timestamp 1586364061
transform 1 0 9200 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 11316 0 -1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 11132 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_103
timestamp 1586364061
transform 1 0 10580 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_107
timestamp 1586364061
transform 1 0 10948 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 13248 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13616 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_130
timestamp 1586364061
transform 1 0 13064 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_134
timestamp 1586364061
transform 1 0 13432 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_138
timestamp 1586364061
transform 1 0 13800 0 -1 17952
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_8.mux_l3_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 13984 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14352 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_142
timestamp 1586364061
transform 1 0 14168 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_146
timestamp 1586364061
transform 1 0 14536 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_150
timestamp 1586364061
transform 1 0 14904 0 -1 17952
box -38 -48 130 592
use scs8hd_conb_1  _037_
timestamp 1586364061
transform 1 0 17296 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17112 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_163
timestamp 1586364061
transform 1 0 16100 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_6  FILLER_28_168
timestamp 1586364061
transform 1 0 16560 0 -1 17952
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_top_track_16.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18308 0 -1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 18032 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_179
timestamp 1586364061
transform 1 0 17572 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_183
timestamp 1586364061
transform 1 0 17940 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_186
timestamp 1586364061
transform 1 0 18216 0 -1 17952
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 20240 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_206
timestamp 1586364061
transform 1 0 20056 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_210
timestamp 1586364061
transform 1 0 20424 0 -1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 22816 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_234
timestamp 1586364061
transform 1 0 22632 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_238
timestamp 1586364061
transform 1 0 23000 0 -1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_32.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 23920 0 -1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 23644 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 23184 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_242
timestamp 1586364061
transform 1 0 23368 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_28_247
timestamp 1586364061
transform 1 0 23828 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_267
timestamp 1586364061
transform 1 0 25668 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_39
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 590 592
use scs8hd_mux2_2  mux_right_track_10.mux_l2_in_1_
timestamp 1586364061
transform 1 0 9476 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 9292 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 8924 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 8556 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_80
timestamp 1586364061
transform 1 0 8464 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_83
timestamp 1586364061
transform 1 0 8740 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_87
timestamp 1586364061
transform 1 0 9108 0 1 17952
box -38 -48 222 592
use scs8hd_conb_1  _041_
timestamp 1586364061
transform 1 0 11316 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 12052 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 11132 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10488 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_100
timestamp 1586364061
transform 1 0 10304 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_104
timestamp 1586364061
transform 1 0 10672 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_108
timestamp 1586364061
transform 1 0 11040 0 1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_29_121
timestamp 1586364061
transform 1 0 12236 0 1 17952
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 15456 0 1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 15272 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 14904 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 14536 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_142
timestamp 1586364061
transform 1 0 14168 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_148
timestamp 1586364061
transform 1 0 14720 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_152
timestamp 1586364061
transform 1 0 15088 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_175
timestamp 1586364061
transform 1 0 17204 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_16.mux_l2_in_1_
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_179
timestamp 1586364061
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_193
timestamp 1586364061
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_197
timestamp 1586364061
transform 1 0 19228 0 1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_16.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 19596 0 1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 19412 0 1 17952
box -38 -48 222 592
use scs8hd_buf_4  mux_top_track_24.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22080 0 1 17952
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 23000 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 21804 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_220
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_224
timestamp 1586364061
transform 1 0 21712 0 1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_29_227
timestamp 1586364061
transform 1 0 21988 0 1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_234
timestamp 1586364061
transform 1 0 22632 0 1 17952
box -38 -48 406 592
use scs8hd_mux2_2  mux_top_track_32.mux_l2_in_0_
timestamp 1586364061
transform 1 0 24288 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 24104 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_240
timestamp 1586364061
transform 1 0 23184 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_249
timestamp 1586364061
transform 1 0 24012 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 25300 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 25668 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_261
timestamp 1586364061
transform 1 0 25116 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_265
timestamp 1586364061
transform 1 0 25484 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 8004 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_30_74
timestamp 1586364061
transform 1 0 7912 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_77
timestamp 1586364061
transform 1 0 8188 0 -1 19040
box -38 -48 1142 592
use scs8hd_mux2_2  mux_right_track_10.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_89
timestamp 1586364061
transform 1 0 9292 0 -1 19040
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_track_8.mux_l1_in_1_
timestamp 1586364061
transform 1 0 12052 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 10672 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_106
timestamp 1586364061
transform 1 0 10856 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_30_114
timestamp 1586364061
transform 1 0 11592 0 -1 19040
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13064 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 13432 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_128
timestamp 1586364061
transform 1 0 12880 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_132
timestamp 1586364061
transform 1 0 13248 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_8.mux_l2_in_1_
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14628 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_145
timestamp 1586364061
transform 1 0 14444 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_149
timestamp 1586364061
transform 1 0 14812 0 -1 19040
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_16.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 17112 0 -1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 16284 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 16652 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_163
timestamp 1586364061
transform 1 0 16100 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_167
timestamp 1586364061
transform 1 0 16468 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_171
timestamp 1586364061
transform 1 0 16836 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 19044 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_193
timestamp 1586364061
transform 1 0 18860 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_197
timestamp 1586364061
transform 1 0 19228 0 -1 19040
box -38 -48 406 592
use scs8hd_conb_1  _039_
timestamp 1586364061
transform 1 0 19780 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 21160 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 19596 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 20240 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_206
timestamp 1586364061
transform 1 0 20056 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_210
timestamp 1586364061
transform 1 0 20424 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_24.mux_l3_in_0_
timestamp 1586364061
transform 1 0 21804 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 21528 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 22816 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_220
timestamp 1586364061
transform 1 0 21344 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_224
timestamp 1586364061
transform 1 0 21712 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_234
timestamp 1586364061
transform 1 0 22632 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_238
timestamp 1586364061
transform 1 0 23000 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_32.mux_l2_in_1_
timestamp 1586364061
transform 1 0 23828 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 23184 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23552 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_242
timestamp 1586364061
transform 1 0 23368 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_246
timestamp 1586364061
transform 1 0 23736 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_256
timestamp 1586364061
transform 1 0 24656 0 -1 19040
box -38 -48 222 592
use scs8hd_conb_1  _040_
timestamp 1586364061
transform 1 0 25392 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 24840 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 25208 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_260
timestamp 1586364061
transform 1 0 25024 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_267
timestamp 1586364061
transform 1 0 25668 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_10.mux_l3_in_0_
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_31_70
timestamp 1586364061
transform 1 0 7544 0 1 19040
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_10.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 9568 0 1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 9384 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_84
timestamp 1586364061
transform 1 0 8832 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_88
timestamp 1586364061
transform 1 0 9200 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11500 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_111
timestamp 1586364061
transform 1 0 11316 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_115
timestamp 1586364061
transform 1 0 11684 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_119
timestamp 1586364061
transform 1 0 12052 0 1 19040
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 13800 0 1 19040
box -38 -48 1786 592
use scs8hd_buf_4  mux_top_track_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 13156 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13616 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_129
timestamp 1586364061
transform 1 0 12972 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_133
timestamp 1586364061
transform 1 0 13340 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_157
timestamp 1586364061
transform 1 0 15548 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_8.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16284 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16100 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 17296 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_161
timestamp 1586364061
transform 1 0 15916 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_174
timestamp 1586364061
transform 1 0 17112 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_178
timestamp 1586364061
transform 1 0 17480 0 1 19040
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_track_14.mux_l3_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 19044 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_193
timestamp 1586364061
transform 1 0 18860 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_197
timestamp 1586364061
transform 1 0 19228 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_16.mux_l3_in_0_
timestamp 1586364061
transform 1 0 19596 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 21160 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 20792 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 19412 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_210
timestamp 1586364061
transform 1 0 20424 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_216
timestamp 1586364061
transform 1 0 20976 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 22724 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 22356 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_229
timestamp 1586364061
transform 1 0 22172 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_233
timestamp 1586364061
transform 1 0 22540 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_237
timestamp 1586364061
transform 1 0 22908 0 1 19040
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_32.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 24104 0 1 19040
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 23920 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_241
timestamp 1586364061
transform 1 0 23276 0 1 19040
box -38 -48 130 592
use scs8hd_decap_3  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 26036 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_273
timestamp 1586364061
transform 1 0 26220 0 1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 8004 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_32_74
timestamp 1586364061
transform 1 0 7912 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_6  FILLER_32_77
timestamp 1586364061
transform 1 0 8188 0 -1 20128
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 8740 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_85
timestamp 1586364061
transform 1 0 8924 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_32_91
timestamp 1586364061
transform 1 0 9476 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_right_track_12.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10488 0 -1 20128
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_32_101
timestamp 1586364061
transform 1 0 10396 0 -1 20128
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_12.mux_l2_in_1_
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 12420 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_121
timestamp 1586364061
transform 1 0 12236 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_125
timestamp 1586364061
transform 1 0 12604 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_138
timestamp 1586364061
transform 1 0 13800 0 -1 20128
box -38 -48 222 592
use scs8hd_conb_1  _042_
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 13984 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_142
timestamp 1586364061
transform 1 0 14168 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_3  FILLER_32_150
timestamp 1586364061
transform 1 0 14904 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_157
timestamp 1586364061
transform 1 0 15548 0 -1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_14.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 16284 0 -1 20128
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 15732 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 16100 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_161
timestamp 1586364061
transform 1 0 15916 0 -1 20128
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_14.mux_l2_in_1_
timestamp 1586364061
transform 1 0 18768 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 18216 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_184
timestamp 1586364061
transform 1 0 18032 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_188
timestamp 1586364061
transform 1 0 18400 0 -1 20128
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 21160 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 19780 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 20148 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_201
timestamp 1586364061
transform 1 0 19596 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_205
timestamp 1586364061
transform 1 0 19964 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_209
timestamp 1586364061
transform 1 0 20332 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_track_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 22724 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 22172 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_231
timestamp 1586364061
transform 1 0 22356 0 -1 20128
box -38 -48 406 592
use scs8hd_mux2_2  mux_top_track_32.mux_l3_in_0_
timestamp 1586364061
transform 1 0 24288 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 24104 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 23736 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_244
timestamp 1586364061
transform 1 0 23552 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_248
timestamp 1586364061
transform 1 0 23920 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_261
timestamp 1586364061
transform 1 0 25116 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_32_273
timestamp 1586364061
transform 1 0 26220 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_34_69
timestamp 1586364061
transform 1 0 7452 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_64
timestamp 1586364061
transform 1 0 6992 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 7268 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_73
timestamp 1586364061
transform 1 0 7820 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_77
timestamp 1586364061
transform 1 0 8188 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_73
timestamp 1586364061
transform 1 0 7820 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_70
timestamp 1586364061
transform 1 0 7544 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 7636 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 7636 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 8372 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 8004 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_10.mux_l1_in_0_
timestamp 1586364061
transform 1 0 8004 0 -1 21216
box -38 -48 866 592
use scs8hd_conb_1  _051_
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_10.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 8740 0 1 20128
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9016 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_81
timestamp 1586364061
transform 1 0 8556 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_84
timestamp 1586364061
transform 1 0 8832 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_88
timestamp 1586364061
transform 1 0 9200 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_8  FILLER_34_96
timestamp 1586364061
transform 1 0 9936 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  FILLER_34_106
timestamp 1586364061
transform 1 0 10856 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 11132 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10672 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_111
timestamp 1586364061
transform 1 0 11316 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_117
timestamp 1586364061
transform 1 0 11868 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_114
timestamp 1586364061
transform 1 0 11592 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 11500 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12052 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11684 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_102
timestamp 1586364061
transform 1 0 10488 0 1 20128
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_track_12.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11684 0 -1 21216
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_right_track_12.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 12880 0 1 20128
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 12696 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 13616 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_121
timestamp 1586364061
transform 1 0 12236 0 1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_134
timestamp 1586364061
transform 1 0 13432 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_138
timestamp 1586364061
transform 1 0 13800 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_145
timestamp 1586364061
transform 1 0 14444 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_2  FILLER_33_147
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 13984 0 -1 21216
box -38 -48 222 592
use scs8hd_conb_1  _052_
timestamp 1586364061
transform 1 0 14168 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_151
timestamp 1586364061
transform 1 0 14996 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 14812 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 15180 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_12.mux_l3_in_0_
timestamp 1586364061
transform 1 0 15364 0 1 20128
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_14.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1786 592
use scs8hd_conb_1  _053_
timestamp 1586364061
transform 1 0 16928 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 17204 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 16376 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_164
timestamp 1586364061
transform 1 0 16192 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_168
timestamp 1586364061
transform 1 0 16560 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_175
timestamp 1586364061
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_173
timestamp 1586364061
transform 1 0 17020 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_177
timestamp 1586364061
transform 1 0 17388 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_179
timestamp 1586364061
transform 1 0 17572 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17572 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_14.mux_l2_in_0_
timestamp 1586364061
transform 1 0 17756 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_194
timestamp 1586364061
transform 1 0 18952 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 19136 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 18768 0 -1 21216
box -38 -48 222 592
use scs8hd_buf_4  mux_top_track_16.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 19320 0 -1 21216
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_right_track_14.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_34_208
timestamp 1586364061
transform 1 0 20240 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_204
timestamp 1586364061
transform 1 0 19872 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_203
timestamp 1586364061
transform 1 0 19780 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 20056 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 20148 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_213
timestamp 1586364061
transform 1 0 20700 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_209
timestamp 1586364061
transform 1 0 20332 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 20516 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 20884 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 21068 0 1 20128
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 22540 0 -1 21216
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 23000 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 21896 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 22264 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_236
timestamp 1586364061
transform 1 0 22816 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_224
timestamp 1586364061
transform 1 0 21712 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_228
timestamp 1586364061
transform 1 0 22080 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_232
timestamp 1586364061
transform 1 0 22448 0 -1 21216
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 24104 0 1 20128
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23920 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_240
timestamp 1586364061
transform 1 0 23184 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_34_252
timestamp 1586364061
transform 1 0 24288 0 -1 21216
box -38 -48 774 592
use scs8hd_conb_1  _050_
timestamp 1586364061
transform 1 0 25024 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_10.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 8096 0 1 21216
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 7544 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 7176 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_68
timestamp 1586364061
transform 1 0 7360 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_72
timestamp 1586364061
transform 1 0 7728 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_95
timestamp 1586364061
transform 1 0 9844 0 1 21216
box -38 -48 590 592
use scs8hd_mux2_2  mux_right_track_12.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10672 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 11684 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10488 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_101
timestamp 1586364061
transform 1 0 10396 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_113
timestamp 1586364061
transform 1 0 11500 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_117
timestamp 1586364061
transform 1 0 11868 0 1 21216
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_track_12.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12696 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 13708 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_14.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15088 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 14904 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 14536 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 14076 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_139
timestamp 1586364061
transform 1 0 13892 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_143
timestamp 1586364061
transform 1 0 14260 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_148
timestamp 1586364061
transform 1 0 14720 0 1 21216
box -38 -48 222 592
use scs8hd_buf_4  mux_top_track_8.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16652 0 1 21216
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 16100 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 16468 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_161
timestamp 1586364061
transform 1 0 15916 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_165
timestamp 1586364061
transform 1 0 16284 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_175
timestamp 1586364061
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use scs8hd_conb_1  _028_
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_track_2.mux_l1_in_2_
timestamp 1586364061
transform 1 0 19228 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 19044 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 18676 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_179
timestamp 1586364061
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_187
timestamp 1586364061
transform 1 0 18308 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_193
timestamp 1586364061
transform 1 0 18860 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 21160 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 20792 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_206
timestamp 1586364061
transform 1 0 20056 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_210
timestamp 1586364061
transform 1 0 20424 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_216
timestamp 1586364061
transform 1 0 20976 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 21712 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 21528 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 22816 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_233
timestamp 1586364061
transform 1 0 22540 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_238
timestamp 1586364061
transform 1 0 23000 0 1 21216
box -38 -48 222 592
use scs8hd_buf_4  mux_top_track_32.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23920 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23184 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24656 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_242
timestamp 1586364061
transform 1 0 23368 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_254
timestamp 1586364061
transform 1 0 24472 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_258
timestamp 1586364061
transform 1 0 24840 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_270
timestamp 1586364061
transform 1 0 25944 0 1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_35_276
timestamp 1586364061
transform 1 0 26496 0 1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 406 592
use scs8hd_conb_1  _035_
timestamp 1586364061
transform 1 0 6624 0 -1 22304
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_track_8.mux_l3_in_0_
timestamp 1586364061
transform 1 0 7636 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 7452 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_63
timestamp 1586364061
transform 1 0 6900 0 -1 22304
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 10212 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 590 592
use scs8hd_mux2_2  mux_right_track_6.mux_l1_in_3_
timestamp 1586364061
transform 1 0 11132 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 10672 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_101
timestamp 1586364061
transform 1 0 10396 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_36_106
timestamp 1586364061
transform 1 0 10856 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_4  FILLER_36_118
timestamp 1586364061
transform 1 0 11960 0 -1 22304
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_track_4.mux_l1_in_1_
timestamp 1586364061
transform 1 0 13432 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12696 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 13064 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 12328 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_124
timestamp 1586364061
transform 1 0 12512 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_128
timestamp 1586364061
transform 1 0 12880 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_132
timestamp 1586364061
transform 1 0 13248 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_4.mux_l1_in_3_
timestamp 1586364061
transform 1 0 15640 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 15456 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 14996 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_143
timestamp 1586364061
transform 1 0 14260 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_2.mux_l1_in_3_
timestamp 1586364061
transform 1 0 17204 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 16652 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_167
timestamp 1586364061
transform 1 0 16468 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_171
timestamp 1586364061
transform 1 0 16836 0 -1 22304
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_track_2.mux_l2_in_1_
timestamp 1586364061
transform 1 0 18768 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 18492 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_184
timestamp 1586364061
transform 1 0 18032 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_188
timestamp 1586364061
transform 1 0 18400 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_191
timestamp 1586364061
transform 1 0 18676 0 -1 22304
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 21068 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 19780 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20148 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_201
timestamp 1586364061
transform 1 0 19596 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_205
timestamp 1586364061
transform 1 0 19964 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_209
timestamp 1586364061
transform 1 0 20332 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_213
timestamp 1586364061
transform 1 0 20700 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 21620 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 21436 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_219
timestamp 1586364061
transform 1 0 21252 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_232
timestamp 1586364061
transform 1 0 22448 0 -1 22304
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 23184 0 -1 22304
box -38 -48 1786 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_259
timestamp 1586364061
transform 1 0 24932 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_36_271
timestamp 1586364061
transform 1 0 26036 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 7728 0 1 22304
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 7544 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6992 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_66
timestamp 1586364061
transform 1 0 7176 0 1 22304
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_track_8.mux_l2_in_1_
timestamp 1586364061
transform 1 0 10212 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 10028 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 9660 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_91
timestamp 1586364061
transform 1 0 9476 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_95
timestamp 1586364061
transform 1 0 9844 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_108
timestamp 1586364061
transform 1 0 11040 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_112
timestamp 1586364061
transform 1 0 11408 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_118
timestamp 1586364061
transform 1 0 11960 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_6.mux_l1_in_1_
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 13432 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_132
timestamp 1586364061
transform 1 0 13248 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_136
timestamp 1586364061
transform 1 0 13616 0 1 22304
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_track_4.mux_l3_in_0_
timestamp 1586364061
transform 1 0 14996 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 14812 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 14444 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14076 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_140
timestamp 1586364061
transform 1 0 13984 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_143
timestamp 1586364061
transform 1 0 14260 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_147
timestamp 1586364061
transform 1 0 14628 0 1 22304
box -38 -48 222 592
use scs8hd_buf_2  _109_
timestamp 1586364061
transform 1 0 16744 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 17296 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 16008 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_160
timestamp 1586364061
transform 1 0 15824 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_164
timestamp 1586364061
transform 1 0 16192 0 1 22304
box -38 -48 590 592
use scs8hd_fill_2  FILLER_37_174
timestamp 1586364061
transform 1 0 17112 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_178
timestamp 1586364061
transform 1 0 17480 0 1 22304
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18492 0 1 22304
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 18308 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_track_2.mux_l3_in_0_
timestamp 1586364061
transform 1 0 20976 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 20792 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 20424 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_208
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_212
timestamp 1586364061
transform 1 0 20608 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 21988 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 22356 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_225
timestamp 1586364061
transform 1 0 21804 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_229
timestamp 1586364061
transform 1 0 22172 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_233
timestamp 1586364061
transform 1 0 22540 0 1 22304
box -38 -48 774 592
use scs8hd_buf_2  _099_
timestamp 1586364061
transform 1 0 24564 0 1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 24380 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_241
timestamp 1586364061
transform 1 0 23276 0 1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 25116 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_259
timestamp 1586364061
transform 1 0 24932 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_263
timestamp 1586364061
transform 1 0 25300 0 1 22304
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_37_275
timestamp 1586364061
transform 1 0 26404 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6992 0 -1 23392
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_right_track_6.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 10120 0 -1 23392
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 9936 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_83
timestamp 1586364061
transform 1 0 8740 0 -1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_38_91
timestamp 1586364061
transform 1 0 9476 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 12052 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_6.mux_l2_in_1_
timestamp 1586364061
transform 1 0 12604 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 12420 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13616 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_121
timestamp 1586364061
transform 1 0 12236 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_134
timestamp 1586364061
transform 1 0 13432 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_138
timestamp 1586364061
transform 1 0 13800 0 -1 23392
box -38 -48 222 592
use scs8hd_conb_1  _034_
timestamp 1586364061
transform 1 0 14168 0 -1 23392
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 13984 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 14996 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_145
timestamp 1586364061
transform 1 0 14444 0 -1 23392
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 17204 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_173
timestamp 1586364061
transform 1 0 17020 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_177
timestamp 1586364061
transform 1 0 17388 0 -1 23392
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_6.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 17756 0 -1 23392
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17572 0 -1 23392
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 20976 0 -1 23392
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 19872 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 20608 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 20240 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_200
timestamp 1586364061
transform 1 0 19504 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_38_206
timestamp 1586364061
transform 1 0 20056 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_210
timestamp 1586364061
transform 1 0 20424 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 22908 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_235
timestamp 1586364061
transform 1 0 22724 0 -1 23392
box -38 -48 222 592
use scs8hd_buf_2  _098_
timestamp 1586364061
transform 1 0 24564 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_259
timestamp 1586364061
transform 1 0 24932 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_38_271
timestamp 1586364061
transform 1 0 26036 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_15
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_27
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_39
timestamp 1586364061
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_51
timestamp 1586364061
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_2  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_64
timestamp 1586364061
transform 1 0 6992 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_66
timestamp 1586364061
transform 1 0 7176 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 7176 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6992 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 7360 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 6808 0 -1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 7544 0 -1 24480
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 7728 0 -1 24480
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7544 0 1 23392
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_40_81
timestamp 1586364061
transform 1 0 8556 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_6  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 590 592
use scs8hd_decap_3  FILLER_40_89
timestamp 1586364061
transform 1 0 9292 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_96
timestamp 1586364061
transform 1 0 9936 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_93
timestamp 1586364061
transform 1 0 9660 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_89
timestamp 1586364061
transform 1 0 9292 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9752 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_40_99
timestamp 1586364061
transform 1 0 10212 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_6.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 10488 0 -1 24480
box -38 -48 1786 592
use scs8hd_mux2_2  mux_right_track_6.mux_l3_in_0_
timestamp 1586364061
transform 1 0 10304 0 1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11316 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 10304 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 11684 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_109
timestamp 1586364061
transform 1 0 11132 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_113
timestamp 1586364061
transform 1 0 11500 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_117
timestamp 1586364061
transform 1 0 11868 0 1 23392
box -38 -48 314 592
use scs8hd_decap_4  FILLER_40_125
timestamp 1586364061
transform 1 0 12604 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_121
timestamp 1586364061
transform 1 0 12236 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_127
timestamp 1586364061
transform 1 0 12788 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 12420 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_buf_2  _114_
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_131
timestamp 1586364061
transform 1 0 13156 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_131
timestamp 1586364061
transform 1 0 13156 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12972 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13340 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13340 0 -1 24480
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 1786 592
use scs8hd_mux2_2  mux_right_track_4.mux_l2_in_1_
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 15456 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 14996 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_154
timestamp 1586364061
transform 1 0 15272 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_158
timestamp 1586364061
transform 1 0 15640 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_142
timestamp 1586364061
transform 1 0 14168 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_1  FILLER_40_150
timestamp 1586364061
transform 1 0 14904 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_40_168
timestamp 1586364061
transform 1 0 16560 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_40_163
timestamp 1586364061
transform 1 0 16100 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_162
timestamp 1586364061
transform 1 0 16008 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 15824 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16192 0 1 23392
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_2.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 23392
box -38 -48 866 592
use scs8hd_decap_8  FILLER_40_175
timestamp 1586364061
transform 1 0 17204 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_175
timestamp 1586364061
transform 1 0 17204 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _111_
timestamp 1586364061
transform 1 0 16836 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_187
timestamp 1586364061
transform 1 0 18308 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_179
timestamp 1586364061
transform 1 0 17572 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_6.mux_l1_in_2_
timestamp 1586364061
transform 1 0 18216 0 1 23392
box -38 -48 866 592
use scs8hd_buf_2  _108_
timestamp 1586364061
transform 1 0 17940 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_191
timestamp 1586364061
transform 1 0 18676 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_195
timestamp 1586364061
transform 1 0 19044 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 18860 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 19228 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 18492 0 -1 24480
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_2.mux_l2_in_0_
timestamp 1586364061
transform 1 0 19044 0 -1 24480
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 19872 0 1 23392
box -38 -48 1786 592
use scs8hd_mux2_2  mux_right_track_4.mux_l1_in_2_
timestamp 1586364061
transform 1 0 20976 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 19688 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 20056 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_199
timestamp 1586364061
transform 1 0 19412 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_40_204
timestamp 1586364061
transform 1 0 19872 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_40_208
timestamp 1586364061
transform 1 0 20240 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_40_225
timestamp 1586364061
transform 1 0 21804 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_227
timestamp 1586364061
transform 1 0 21988 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_223
timestamp 1586364061
transform 1 0 21620 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 21804 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_235
timestamp 1586364061
transform 1 0 22724 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 22172 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _104_
timestamp 1586364061
transform 1 0 22356 0 1 23392
box -38 -48 406 592
use scs8hd_buf_2  _103_
timestamp 1586364061
transform 1 0 22540 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_8  FILLER_40_237
timestamp 1586364061
transform 1 0 22908 0 -1 24480
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 22908 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_239
timestamp 1586364061
transform 1 0 23092 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 23368 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_buf_2  _101_
timestamp 1586364061
transform 1 0 23644 0 -1 24480
box -38 -48 406 592
use scs8hd_buf_2  _100_
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 406 592
use scs8hd_decap_8  FILLER_40_249
timestamp 1586364061
transform 1 0 24012 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_253
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_249
timestamp 1586364061
transform 1 0 24012 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 24564 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 24196 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _097_
timestamp 1586364061
transform 1 0 24748 0 -1 24480
box -38 -48 406 592
use scs8hd_buf_2  _096_
timestamp 1586364061
transform 1 0 24748 0 1 23392
box -38 -48 406 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 25300 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_261
timestamp 1586364061
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_265
timestamp 1586364061
transform 1 0 25484 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_261
timestamp 1586364061
transform 1 0 25116 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_40_273
timestamp 1586364061
transform 1 0 26220 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_57
timestamp 1586364061
transform 1 0 6348 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_8.mux_l1_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 7820 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_71
timestamp 1586364061
transform 1 0 7636 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_75
timestamp 1586364061
transform 1 0 8004 0 1 24480
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9936 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 9568 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_87
timestamp 1586364061
transform 1 0 9108 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_91
timestamp 1586364061
transform 1 0 9476 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_94
timestamp 1586364061
transform 1 0 9752 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_6.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10488 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10304 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 11500 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_111
timestamp 1586364061
transform 1 0 11316 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_115
timestamp 1586364061
transform 1 0 11684 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_119
timestamp 1586364061
transform 1 0 12052 0 1 24480
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_4.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12972 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12788 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_138
timestamp 1586364061
transform 1 0 13800 0 1 24480
box -38 -48 222 592
use scs8hd_buf_2  _112_
timestamp 1586364061
transform 1 0 15640 0 1 24480
box -38 -48 406 592
use scs8hd_buf_2  _115_
timestamp 1586364061
transform 1 0 14536 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 15088 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 13984 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_142
timestamp 1586364061
transform 1 0 14168 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_150
timestamp 1586364061
transform 1 0 14904 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_154
timestamp 1586364061
transform 1 0 15272 0 1 24480
box -38 -48 406 592
use scs8hd_buf_2  _110_
timestamp 1586364061
transform 1 0 16744 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 16192 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 17296 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_162
timestamp 1586364061
transform 1 0 16008 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_166
timestamp 1586364061
transform 1 0 16376 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_174
timestamp 1586364061
transform 1 0 17112 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_178
timestamp 1586364061
transform 1 0 17480 0 1 24480
box -38 -48 406 592
use scs8hd_buf_2  _106_
timestamp 1586364061
transform 1 0 18400 0 1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 18952 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 19320 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 18216 0 1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_182
timestamp 1586364061
transform 1 0 17848 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_192
timestamp 1586364061
transform 1 0 18768 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 222 592
use scs8hd_buf_2  _105_
timestamp 1586364061
transform 1 0 21068 0 1 24480
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_track_2.mux_l1_in_1_
timestamp 1586364061
transform 1 0 19504 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 20516 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_209
timestamp 1586364061
transform 1 0 20332 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_213
timestamp 1586364061
transform 1 0 20700 0 1 24480
box -38 -48 406 592
use scs8hd_buf_2  _102_
timestamp 1586364061
transform 1 0 22172 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 22724 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 21620 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_221
timestamp 1586364061
transform 1 0 21436 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_225
timestamp 1586364061
transform 1 0 21804 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_233
timestamp 1586364061
transform 1 0 22540 0 1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_41_237
timestamp 1586364061
transform 1 0 22908 0 1 24480
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_41_243
timestamp 1586364061
transform 1 0 23460 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_mux2_2  mux_right_track_6.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9936 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_fill_2  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10948 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 11316 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_105
timestamp 1586364061
transform 1 0 10764 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_109
timestamp 1586364061
transform 1 0 11132 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_113
timestamp 1586364061
transform 1 0 11500 0 -1 25568
box -38 -48 774 592
use scs8hd_buf_2  _113_
timestamp 1586364061
transform 1 0 12972 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_3  FILLER_42_121
timestamp 1586364061
transform 1 0 12236 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_133
timestamp 1586364061
transform 1 0 13340 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_145
timestamp 1586364061
transform 1 0 14444 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_2  FILLER_42_153
timestamp 1586364061
transform 1 0 15180 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 406 592
use scs8hd_conb_1  _033_
timestamp 1586364061
transform 1 0 15916 0 -1 25568
box -38 -48 314 592
use scs8hd_fill_1  FILLER_42_160
timestamp 1586364061
transform 1 0 15824 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_164
timestamp 1586364061
transform 1 0 16192 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_42_176
timestamp 1586364061
transform 1 0 17296 0 -1 25568
box -38 -48 774 592
use scs8hd_buf_2  _107_
timestamp 1586364061
transform 1 0 19136 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_42_184
timestamp 1586364061
transform 1 0 18032 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_1  FILLER_42_195
timestamp 1586364061
transform 1 0 19044 0 -1 25568
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 19688 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_200
timestamp 1586364061
transform 1 0 19504 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_42_204
timestamp 1586364061
transform 1 0 19872 0 -1 25568
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_42_216
timestamp 1586364061
transform 1 0 20976 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 294 0 350 480 6 bottom_left_grid_pin_1_
port 0 nsew default input
rlabel metal2 s 27526 0 27582 480 6 ccff_head
port 1 nsew default input
rlabel metal3 s 0 6944 480 7064 6 ccff_tail
port 2 nsew default tristate
rlabel metal3 s 27520 11840 28000 11960 6 chanx_right_in[0]
port 3 nsew default input
rlabel metal3 s 27520 17688 28000 17808 6 chanx_right_in[10]
port 4 nsew default input
rlabel metal3 s 27520 18368 28000 18488 6 chanx_right_in[11]
port 5 nsew default input
rlabel metal3 s 27520 18912 28000 19032 6 chanx_right_in[12]
port 6 nsew default input
rlabel metal3 s 27520 19456 28000 19576 6 chanx_right_in[13]
port 7 nsew default input
rlabel metal3 s 27520 20000 28000 20120 6 chanx_right_in[14]
port 8 nsew default input
rlabel metal3 s 27520 20680 28000 20800 6 chanx_right_in[15]
port 9 nsew default input
rlabel metal3 s 27520 21224 28000 21344 6 chanx_right_in[16]
port 10 nsew default input
rlabel metal3 s 27520 21768 28000 21888 6 chanx_right_in[17]
port 11 nsew default input
rlabel metal3 s 27520 22448 28000 22568 6 chanx_right_in[18]
port 12 nsew default input
rlabel metal3 s 27520 22992 28000 23112 6 chanx_right_in[19]
port 13 nsew default input
rlabel metal3 s 27520 12520 28000 12640 6 chanx_right_in[1]
port 14 nsew default input
rlabel metal3 s 27520 13064 28000 13184 6 chanx_right_in[2]
port 15 nsew default input
rlabel metal3 s 27520 13608 28000 13728 6 chanx_right_in[3]
port 16 nsew default input
rlabel metal3 s 27520 14288 28000 14408 6 chanx_right_in[4]
port 17 nsew default input
rlabel metal3 s 27520 14832 28000 14952 6 chanx_right_in[5]
port 18 nsew default input
rlabel metal3 s 27520 15376 28000 15496 6 chanx_right_in[6]
port 19 nsew default input
rlabel metal3 s 27520 15920 28000 16040 6 chanx_right_in[7]
port 20 nsew default input
rlabel metal3 s 27520 16600 28000 16720 6 chanx_right_in[8]
port 21 nsew default input
rlabel metal3 s 27520 17144 28000 17264 6 chanx_right_in[9]
port 22 nsew default input
rlabel metal3 s 27520 280 28000 400 6 chanx_right_out[0]
port 23 nsew default tristate
rlabel metal3 s 27520 5992 28000 6112 6 chanx_right_out[10]
port 24 nsew default tristate
rlabel metal3 s 27520 6672 28000 6792 6 chanx_right_out[11]
port 25 nsew default tristate
rlabel metal3 s 27520 7216 28000 7336 6 chanx_right_out[12]
port 26 nsew default tristate
rlabel metal3 s 27520 7760 28000 7880 6 chanx_right_out[13]
port 27 nsew default tristate
rlabel metal3 s 27520 8440 28000 8560 6 chanx_right_out[14]
port 28 nsew default tristate
rlabel metal3 s 27520 8984 28000 9104 6 chanx_right_out[15]
port 29 nsew default tristate
rlabel metal3 s 27520 9528 28000 9648 6 chanx_right_out[16]
port 30 nsew default tristate
rlabel metal3 s 27520 10072 28000 10192 6 chanx_right_out[17]
port 31 nsew default tristate
rlabel metal3 s 27520 10752 28000 10872 6 chanx_right_out[18]
port 32 nsew default tristate
rlabel metal3 s 27520 11296 28000 11416 6 chanx_right_out[19]
port 33 nsew default tristate
rlabel metal3 s 27520 824 28000 944 6 chanx_right_out[1]
port 34 nsew default tristate
rlabel metal3 s 27520 1368 28000 1488 6 chanx_right_out[2]
port 35 nsew default tristate
rlabel metal3 s 27520 1912 28000 2032 6 chanx_right_out[3]
port 36 nsew default tristate
rlabel metal3 s 27520 2592 28000 2712 6 chanx_right_out[4]
port 37 nsew default tristate
rlabel metal3 s 27520 3136 28000 3256 6 chanx_right_out[5]
port 38 nsew default tristate
rlabel metal3 s 27520 3680 28000 3800 6 chanx_right_out[6]
port 39 nsew default tristate
rlabel metal3 s 27520 4360 28000 4480 6 chanx_right_out[7]
port 40 nsew default tristate
rlabel metal3 s 27520 4904 28000 5024 6 chanx_right_out[8]
port 41 nsew default tristate
rlabel metal3 s 27520 5448 28000 5568 6 chanx_right_out[9]
port 42 nsew default tristate
rlabel metal2 s 938 0 994 480 6 chany_bottom_in[0]
port 43 nsew default input
rlabel metal2 s 7562 0 7618 480 6 chany_bottom_in[10]
port 44 nsew default input
rlabel metal2 s 8206 0 8262 480 6 chany_bottom_in[11]
port 45 nsew default input
rlabel metal2 s 8942 0 8998 480 6 chany_bottom_in[12]
port 46 nsew default input
rlabel metal2 s 9586 0 9642 480 6 chany_bottom_in[13]
port 47 nsew default input
rlabel metal2 s 10230 0 10286 480 6 chany_bottom_in[14]
port 48 nsew default input
rlabel metal2 s 10874 0 10930 480 6 chany_bottom_in[15]
port 49 nsew default input
rlabel metal2 s 11610 0 11666 480 6 chany_bottom_in[16]
port 50 nsew default input
rlabel metal2 s 12254 0 12310 480 6 chany_bottom_in[17]
port 51 nsew default input
rlabel metal2 s 12898 0 12954 480 6 chany_bottom_in[18]
port 52 nsew default input
rlabel metal2 s 13542 0 13598 480 6 chany_bottom_in[19]
port 53 nsew default input
rlabel metal2 s 1582 0 1638 480 6 chany_bottom_in[1]
port 54 nsew default input
rlabel metal2 s 2226 0 2282 480 6 chany_bottom_in[2]
port 55 nsew default input
rlabel metal2 s 2870 0 2926 480 6 chany_bottom_in[3]
port 56 nsew default input
rlabel metal2 s 3606 0 3662 480 6 chany_bottom_in[4]
port 57 nsew default input
rlabel metal2 s 4250 0 4306 480 6 chany_bottom_in[5]
port 58 nsew default input
rlabel metal2 s 4894 0 4950 480 6 chany_bottom_in[6]
port 59 nsew default input
rlabel metal2 s 5538 0 5594 480 6 chany_bottom_in[7]
port 60 nsew default input
rlabel metal2 s 6274 0 6330 480 6 chany_bottom_in[8]
port 61 nsew default input
rlabel metal2 s 6918 0 6974 480 6 chany_bottom_in[9]
port 62 nsew default input
rlabel metal2 s 14278 0 14334 480 6 chany_bottom_out[0]
port 63 nsew default tristate
rlabel metal2 s 20902 0 20958 480 6 chany_bottom_out[10]
port 64 nsew default tristate
rlabel metal2 s 21546 0 21602 480 6 chany_bottom_out[11]
port 65 nsew default tristate
rlabel metal2 s 22190 0 22246 480 6 chany_bottom_out[12]
port 66 nsew default tristate
rlabel metal2 s 22926 0 22982 480 6 chany_bottom_out[13]
port 67 nsew default tristate
rlabel metal2 s 23570 0 23626 480 6 chany_bottom_out[14]
port 68 nsew default tristate
rlabel metal2 s 24214 0 24270 480 6 chany_bottom_out[15]
port 69 nsew default tristate
rlabel metal2 s 24858 0 24914 480 6 chany_bottom_out[16]
port 70 nsew default tristate
rlabel metal2 s 25594 0 25650 480 6 chany_bottom_out[17]
port 71 nsew default tristate
rlabel metal2 s 26238 0 26294 480 6 chany_bottom_out[18]
port 72 nsew default tristate
rlabel metal2 s 26882 0 26938 480 6 chany_bottom_out[19]
port 73 nsew default tristate
rlabel metal2 s 14922 0 14978 480 6 chany_bottom_out[1]
port 74 nsew default tristate
rlabel metal2 s 15566 0 15622 480 6 chany_bottom_out[2]
port 75 nsew default tristate
rlabel metal2 s 16210 0 16266 480 6 chany_bottom_out[3]
port 76 nsew default tristate
rlabel metal2 s 16854 0 16910 480 6 chany_bottom_out[4]
port 77 nsew default tristate
rlabel metal2 s 17590 0 17646 480 6 chany_bottom_out[5]
port 78 nsew default tristate
rlabel metal2 s 18234 0 18290 480 6 chany_bottom_out[6]
port 79 nsew default tristate
rlabel metal2 s 18878 0 18934 480 6 chany_bottom_out[7]
port 80 nsew default tristate
rlabel metal2 s 19522 0 19578 480 6 chany_bottom_out[8]
port 81 nsew default tristate
rlabel metal2 s 20258 0 20314 480 6 chany_bottom_out[9]
port 82 nsew default tristate
rlabel metal2 s 938 27520 994 28000 6 chany_top_in[0]
port 83 nsew default input
rlabel metal2 s 7746 27520 7802 28000 6 chany_top_in[10]
port 84 nsew default input
rlabel metal2 s 8390 27520 8446 28000 6 chany_top_in[11]
port 85 nsew default input
rlabel metal2 s 9126 27520 9182 28000 6 chany_top_in[12]
port 86 nsew default input
rlabel metal2 s 9770 27520 9826 28000 6 chany_top_in[13]
port 87 nsew default input
rlabel metal2 s 10506 27520 10562 28000 6 chany_top_in[14]
port 88 nsew default input
rlabel metal2 s 11150 27520 11206 28000 6 chany_top_in[15]
port 89 nsew default input
rlabel metal2 s 11886 27520 11942 28000 6 chany_top_in[16]
port 90 nsew default input
rlabel metal2 s 12530 27520 12586 28000 6 chany_top_in[17]
port 91 nsew default input
rlabel metal2 s 13174 27520 13230 28000 6 chany_top_in[18]
port 92 nsew default input
rlabel metal2 s 13910 27520 13966 28000 6 chany_top_in[19]
port 93 nsew default input
rlabel metal2 s 1582 27520 1638 28000 6 chany_top_in[1]
port 94 nsew default input
rlabel metal2 s 2318 27520 2374 28000 6 chany_top_in[2]
port 95 nsew default input
rlabel metal2 s 2962 27520 3018 28000 6 chany_top_in[3]
port 96 nsew default input
rlabel metal2 s 3698 27520 3754 28000 6 chany_top_in[4]
port 97 nsew default input
rlabel metal2 s 4342 27520 4398 28000 6 chany_top_in[5]
port 98 nsew default input
rlabel metal2 s 4986 27520 5042 28000 6 chany_top_in[6]
port 99 nsew default input
rlabel metal2 s 5722 27520 5778 28000 6 chany_top_in[7]
port 100 nsew default input
rlabel metal2 s 6366 27520 6422 28000 6 chany_top_in[8]
port 101 nsew default input
rlabel metal2 s 7102 27520 7158 28000 6 chany_top_in[9]
port 102 nsew default input
rlabel metal2 s 14554 27520 14610 28000 6 chany_top_out[0]
port 103 nsew default tristate
rlabel metal2 s 21362 27520 21418 28000 6 chany_top_out[10]
port 104 nsew default tristate
rlabel metal2 s 22098 27520 22154 28000 6 chany_top_out[11]
port 105 nsew default tristate
rlabel metal2 s 22742 27520 22798 28000 6 chany_top_out[12]
port 106 nsew default tristate
rlabel metal2 s 23478 27520 23534 28000 6 chany_top_out[13]
port 107 nsew default tristate
rlabel metal2 s 24122 27520 24178 28000 6 chany_top_out[14]
port 108 nsew default tristate
rlabel metal2 s 24766 27520 24822 28000 6 chany_top_out[15]
port 109 nsew default tristate
rlabel metal2 s 25502 27520 25558 28000 6 chany_top_out[16]
port 110 nsew default tristate
rlabel metal2 s 26146 27520 26202 28000 6 chany_top_out[17]
port 111 nsew default tristate
rlabel metal2 s 26882 27520 26938 28000 6 chany_top_out[18]
port 112 nsew default tristate
rlabel metal2 s 27526 27520 27582 28000 6 chany_top_out[19]
port 113 nsew default tristate
rlabel metal2 s 15290 27520 15346 28000 6 chany_top_out[1]
port 114 nsew default tristate
rlabel metal2 s 15934 27520 15990 28000 6 chany_top_out[2]
port 115 nsew default tristate
rlabel metal2 s 16578 27520 16634 28000 6 chany_top_out[3]
port 116 nsew default tristate
rlabel metal2 s 17314 27520 17370 28000 6 chany_top_out[4]
port 117 nsew default tristate
rlabel metal2 s 17958 27520 18014 28000 6 chany_top_out[5]
port 118 nsew default tristate
rlabel metal2 s 18694 27520 18750 28000 6 chany_top_out[6]
port 119 nsew default tristate
rlabel metal2 s 19338 27520 19394 28000 6 chany_top_out[7]
port 120 nsew default tristate
rlabel metal2 s 20074 27520 20130 28000 6 chany_top_out[8]
port 121 nsew default tristate
rlabel metal2 s 20718 27520 20774 28000 6 chany_top_out[9]
port 122 nsew default tristate
rlabel metal3 s 0 20952 480 21072 6 prog_clk
port 123 nsew default input
rlabel metal3 s 27520 23536 28000 23656 6 right_top_grid_pin_42_
port 124 nsew default input
rlabel metal3 s 27520 24080 28000 24200 6 right_top_grid_pin_43_
port 125 nsew default input
rlabel metal3 s 27520 24760 28000 24880 6 right_top_grid_pin_44_
port 126 nsew default input
rlabel metal3 s 27520 25304 28000 25424 6 right_top_grid_pin_45_
port 127 nsew default input
rlabel metal3 s 27520 25848 28000 25968 6 right_top_grid_pin_46_
port 128 nsew default input
rlabel metal3 s 27520 26528 28000 26648 6 right_top_grid_pin_47_
port 129 nsew default input
rlabel metal3 s 27520 27072 28000 27192 6 right_top_grid_pin_48_
port 130 nsew default input
rlabel metal3 s 27520 27616 28000 27736 6 right_top_grid_pin_49_
port 131 nsew default input
rlabel metal2 s 294 27520 350 28000 6 top_left_grid_pin_1_
port 132 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 133 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 134 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
