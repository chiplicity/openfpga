* NGSPICE file created from cby_3__1_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand2_4 abstract view
.subckt scs8hd_nand2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor3_4 abstract view
.subckt scs8hd_nor3_4 A B C Y vgnd vpwr
.ends

.subckt cby_3__1_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] chany_bottom_in[0] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_out[0] chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3]
+ chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7]
+ chany_bottom_out[8] chany_top_in[0] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_out[0] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4]
+ chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8] data_in enable
+ left_grid_pin_1_ left_grid_pin_5_ left_grid_pin_9_ right_grid_pin_0_ right_grid_pin_10_
+ right_grid_pin_12_ right_grid_pin_14_ right_grid_pin_2_ right_grid_pin_4_ right_grid_pin_6_
+ right_grid_pin_8_ vpwr vgnd
XFILLER_13_100 vpwr vgnd scs8hd_fill_2
XFILLER_26_96 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_5.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_29 vpwr vgnd scs8hd_fill_2
XFILLER_47_18 vpwr vgnd scs8hd_fill_2
XFILLER_63_39 vgnd vpwr scs8hd_decap_12
XFILLER_10_125 vgnd vpwr scs8hd_decap_12
XFILLER_12_32 vgnd vpwr scs8hd_decap_3
XFILLER_12_65 vgnd vpwr scs8hd_decap_3
XFILLER_12_87 vgnd vpwr scs8hd_decap_4
XFILLER_37_40 vpwr vgnd scs8hd_fill_2
XFILLER_37_73 vgnd vpwr scs8hd_decap_3
XANTENNA__124__A _132_/A vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_2_.latch/Q mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_left_ipin_6.LATCH_4_.latch/Q mux_left_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_0.LATCH_1_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
X_200_ chany_top_in[0] chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _159_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__209__A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
X_131_ _139_/A _131_/B _131_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_42 vpwr vgnd scs8hd_fill_2
XFILLER_23_75 vpwr vgnd scs8hd_fill_2
XFILLER_48_83 vpwr vgnd scs8hd_fill_2
XANTENNA__110__C address[3] vgnd vpwr scs8hd_diode_2
XFILLER_9_77 vpwr vgnd scs8hd_fill_2
XANTENNA__119__A _110_/A vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_4.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_left_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_47_139 vgnd vpwr scs8hd_decap_6
XFILLER_47_106 vgnd vpwr scs8hd_decap_4
XFILLER_18_42 vpwr vgnd scs8hd_fill_2
XFILLER_34_41 vgnd vpwr scs8hd_decap_3
XFILLER_50_84 vgnd vpwr scs8hd_decap_8
XFILLER_50_73 vpwr vgnd scs8hd_fill_2
X_114_ _132_/A _118_/B _114_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__121__B _120_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_5.INVTX1_5_.scs8hd_inv_1 chany_top_in[5] mux_left_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_right_ipin_2.LATCH_1_.latch data_in _161_/A _157_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_32 vpwr vgnd scs8hd_fill_2
XFILLER_20_43 vpwr vgnd scs8hd_fill_2
XFILLER_29_74 vpwr vgnd scs8hd_fill_2
XFILLER_45_62 vgnd vpwr scs8hd_decap_3
Xmux_left_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_ipin_2.LATCH_1_.latch/Q mux_left_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_109 vgnd vpwr scs8hd_fill_1
XFILLER_61_94 vpwr vgnd scs8hd_fill_2
XFILLER_61_83 vgnd vpwr scs8hd_decap_8
XFILLER_6_23 vpwr vgnd scs8hd_fill_2
XANTENNA__116__B _118_/B vgnd vpwr scs8hd_diode_2
XANTENNA__132__A _132_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_89 vgnd vpwr scs8hd_decap_3
XFILLER_6_56 vpwr vgnd scs8hd_fill_2
XFILLER_6_45 vpwr vgnd scs8hd_fill_2
XFILLER_13_3 vpwr vgnd scs8hd_fill_2
XFILLER_15_10 vgnd vpwr scs8hd_decap_4
XFILLER_25_120 vpwr vgnd scs8hd_fill_2
XFILLER_40_145 vgnd vpwr scs8hd_fill_1
XFILLER_31_53 vpwr vgnd scs8hd_fill_2
XFILLER_56_83 vpwr vgnd scs8hd_fill_2
XFILLER_56_72 vgnd vpwr scs8hd_decap_8
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_101 vgnd vpwr scs8hd_decap_3
XFILLER_31_123 vgnd vpwr scs8hd_decap_12
XANTENNA__127__A _135_/A vgnd vpwr scs8hd_diode_2
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_145 vgnd vpwr scs8hd_fill_1
XFILLER_13_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_85 vgnd vpwr scs8hd_decap_6
XFILLER_3_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_7.LATCH_0_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_ipin_6.LATCH_2_.latch/Q mux_left_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _186_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_108 vgnd vpwr scs8hd_decap_12
XFILLER_10_137 vgnd vpwr scs8hd_decap_8
XFILLER_12_44 vpwr vgnd scs8hd_fill_2
XFILLER_53_84 vpwr vgnd scs8hd_fill_2
XFILLER_53_51 vgnd vpwr scs8hd_decap_4
XANTENNA__124__B _124_/B vgnd vpwr scs8hd_diode_2
XANTENNA__140__A _132_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_1.LATCH_5_.latch data_in mem_left_ipin_1.LATCH_5_.latch/Q _173_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_left_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_ipin_4.LATCH_0_.latch/Q mux_left_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
X_130_ _130_/A _131_/B vgnd vpwr scs8hd_buf_1
XFILLER_23_54 vgnd vpwr scs8hd_decap_4
XFILLER_48_51 vgnd vpwr scs8hd_decap_4
XANTENNA__110__D _110_/D vgnd vpwr scs8hd_diode_2
XFILLER_64_94 vgnd vpwr scs8hd_decap_12
XFILLER_0_25 vgnd vpwr scs8hd_decap_4
XFILLER_0_36 vgnd vpwr scs8hd_fill_1
XANTENNA__119__B address[4] vgnd vpwr scs8hd_diode_2
XANTENNA__135__A _135_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_34 vpwr vgnd scs8hd_fill_2
XFILLER_43_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_1.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_ipin_1.LATCH_3_.latch/Q mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_18_32 vgnd vpwr scs8hd_fill_1
X_113_ _100_/B _132_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mem_right_ipin_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_107 vgnd vpwr scs8hd_decap_12
XFILLER_61_143 vgnd vpwr scs8hd_decap_3
XFILLER_61_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_5.INVTX1_5_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_2.INVTX1_1_.scs8hd_inv_1 chany_top_in[1] mux_left_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_ipin_5.LATCH_1_.latch_SLEEPB _127_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_20_66 vpwr vgnd scs8hd_fill_2
XFILLER_45_52 vgnd vpwr scs8hd_decap_3
XFILLER_43_121 vgnd vpwr scs8hd_fill_1
XANTENNA__132__B _131_/B vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_3.INVTX1_5_.scs8hd_inv_1 chany_top_in[7] mux_left_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_40_113 vgnd vpwr scs8hd_decap_12
XFILLER_40_102 vpwr vgnd scs8hd_fill_2
XFILLER_15_44 vpwr vgnd scs8hd_fill_2
XFILLER_25_143 vgnd vpwr scs8hd_decap_3
XFILLER_15_99 vgnd vpwr scs8hd_decap_12
XFILLER_31_21 vpwr vgnd scs8hd_fill_2
XFILLER_56_40 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_left_ipin_5.LATCH_4_.latch/Q mux_left_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_135 vgnd vpwr scs8hd_decap_8
XANTENNA__127__B _124_/B vgnd vpwr scs8hd_diode_2
XANTENNA__143__A _135_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_9 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_ipin_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_26_32 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_ipin_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_135 vgnd vpwr scs8hd_decap_8
XFILLER_42_64 vpwr vgnd scs8hd_fill_2
XFILLER_3_36 vpwr vgnd scs8hd_fill_2
XANTENNA__138__A _137_/X vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_2.LATCH_1_.latch data_in mem_left_ipin_2.LATCH_1_.latch/Q _085_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_ipin_4.tap_buf4_0_.scs8hd_inv_1_A mux_left_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_3.LATCH_2_.latch_SLEEPB _103_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_53 vpwr vgnd scs8hd_fill_2
XFILLER_37_86 vgnd vpwr scs8hd_fill_1
XFILLER_5_120 vpwr vgnd scs8hd_fill_2
Xmem_left_ipin_4.LATCH_4_.latch data_in mem_left_ipin_4.LATCH_4_.latch/Q _114_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__140__B _139_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_ipin_1.LATCH_1_.latch/Q mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_3 vgnd vpwr scs8hd_decap_6
XANTENNA__119__C _095_/C vgnd vpwr scs8hd_diode_2
X_189_ _189_/HI _189_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_6.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__135__B _131_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_3.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA__151__A _151_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_4.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_ipin_5.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_7.INVTX1_3_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_11 vgnd vpwr scs8hd_decap_3
XFILLER_18_66 vgnd vpwr scs8hd_decap_4
X_112_ _139_/A _118_/B _112_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_59_95 vgnd vpwr scs8hd_decap_3
XFILLER_59_73 vpwr vgnd scs8hd_fill_2
XFILLER_59_51 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_0.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[7] mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_38_119 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1 mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ right_grid_pin_2_ vgnd vpwr scs8hd_inv_1
XANTENNA__146__A _145_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_108 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_23 vgnd vpwr scs8hd_decap_4
XFILLER_20_89 vgnd vpwr scs8hd_fill_1
XFILLER_45_31 vgnd vpwr scs8hd_decap_4
XFILLER_45_97 vpwr vgnd scs8hd_fill_2
XFILLER_43_111 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_ipin_5.LATCH_2_.latch/Q mux_left_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_left_ipin_1.LATCH_3_.latch_SLEEPB _175_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_125 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_1.LATCH_0_.latch_SLEEPB _156_/Y vgnd vpwr scs8hd_diode_2
XFILLER_25_100 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_5.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_77 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_0.INVTX1_1_.scs8hd_inv_1 chany_top_in[0] mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__B _139_/B vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_ipin_3.LATCH_0_.latch/Q mux_left_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_left_ipin_5.LATCH_0_.latch data_in mem_left_ipin_5.LATCH_0_.latch/Q _128_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_55 vgnd vpwr scs8hd_decap_8
XFILLER_26_66 vgnd vpwr scs8hd_decap_4
XFILLER_42_32 vgnd vpwr scs8hd_decap_4
XFILLER_26_88 vgnd vpwr scs8hd_decap_4
Xmem_right_ipin_0.LATCH_4_.latch data_in mem_right_ipin_0.LATCH_4_.latch/Q _150_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_1.INVTX1_5_.scs8hd_inv_1 chany_top_in[5] mux_left_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_15 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__154__A _144_/A vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_ipin_0.LATCH_3_.latch/Q mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmem_left_ipin_7.LATCH_3_.latch data_in mem_left_ipin_7.LATCH_3_.latch/Q _141_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_106 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _187_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_21 vgnd vpwr scs8hd_decap_4
XFILLER_37_98 vgnd vpwr scs8hd_decap_6
XFILLER_53_75 vgnd vpwr scs8hd_decap_4
XFILLER_5_143 vgnd vpwr scs8hd_decap_3
XANTENNA__149__A _139_/A vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_7.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[6] mux_left_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_59_128 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_ipin_7.LATCH_1_.latch/Q mux_left_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_5.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_23_12 vpwr vgnd scs8hd_fill_2
XFILLER_23_23 vpwr vgnd scs8hd_fill_2
XFILLER_2_102 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_63 vgnd vpwr scs8hd_decap_12
X_188_ _188_/HI _188_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__151__B _149_/B vgnd vpwr scs8hd_diode_2
XFILLER_29_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_7.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_23 vgnd vpwr scs8hd_decap_4
Xmux_left_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_ipin_4.LATCH_4_.latch/Q mux_left_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_34_88 vpwr vgnd scs8hd_fill_2
XFILLER_50_32 vgnd vpwr scs8hd_decap_6
X_111_ _110_/X _118_/B vgnd vpwr scs8hd_buf_1
XFILLER_61_123 vgnd vpwr scs8hd_decap_12
XANTENNA__162__A _162_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_145 vgnd vpwr scs8hd_fill_1
XFILLER_1_81 vpwr vgnd scs8hd_fill_2
XANTENNA__072__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_29_44 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_55 vgnd vpwr scs8hd_decap_4
XFILLER_45_76 vpwr vgnd scs8hd_fill_2
XFILLER_6_15 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_7 vgnd vpwr scs8hd_decap_12
XFILLER_19_120 vpwr vgnd scs8hd_fill_2
XANTENNA__157__A _077_/B vgnd vpwr scs8hd_diode_2
XFILLER_34_145 vgnd vpwr scs8hd_fill_1
Xmem_right_ipin_1.LATCH_0_.latch data_in _160_/A _156_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_25_112 vgnd vpwr scs8hd_decap_8
XFILLER_25_123 vgnd vpwr scs8hd_decap_12
XFILLER_40_137 vgnd vpwr scs8hd_decap_8
XANTENNA__067__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_15_57 vpwr vgnd scs8hd_fill_2
XFILLER_31_34 vpwr vgnd scs8hd_fill_2
XFILLER_56_53 vgnd vpwr scs8hd_decap_6
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_3 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_1_.latch/Q mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_104 vpwr vgnd scs8hd_fill_2
XFILLER_22_115 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_5.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_104 vpwr vgnd scs8hd_fill_2
XFILLER_26_23 vgnd vpwr scs8hd_decap_4
XFILLER_42_77 vpwr vgnd scs8hd_fill_2
XFILLER_59_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_ipin_6.LATCH_3_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__154__B _149_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_130 vgnd vpwr scs8hd_decap_12
XANTENNA__170__A _088_/B vgnd vpwr scs8hd_diode_2
XANTENNA__080__A _069_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__149__B _149_/B vgnd vpwr scs8hd_diode_2
XANTENNA__165__A _179_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_70 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_ipin_4.LATCH_2_.latch/Q mux_left_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__075__A _093_/A vgnd vpwr scs8hd_diode_2
XFILLER_48_32 vgnd vpwr scs8hd_decap_6
XFILLER_48_87 vgnd vpwr scs8hd_decap_3
XFILLER_64_75 vgnd vpwr scs8hd_decap_12
X_187_ _187_/HI _187_/LO vgnd vpwr scs8hd_conb_1
XFILLER_50_7 vgnd vpwr scs8hd_decap_12
Xmem_left_ipin_0.LATCH_4_.latch data_in mem_left_ipin_0.LATCH_4_.latch/Q _166_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_left_ipin_5.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[4] mux_left_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_55_132 vgnd vpwr scs8hd_decap_12
XFILLER_18_46 vpwr vgnd scs8hd_fill_2
X_110_ _110_/A address[4] address[3] _110_/D _110_/X vgnd vpwr scs8hd_or4_4
XFILLER_34_67 vpwr vgnd scs8hd_fill_2
XFILLER_50_77 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_ipin_2.LATCH_0_.latch/Q mux_left_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_61_135 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_121 vgnd vpwr scs8hd_fill_1
XFILLER_37_143 vgnd vpwr scs8hd_decap_3
XFILLER_52_113 vgnd vpwr scs8hd_decap_12
XFILLER_52_102 vgnd vpwr scs8hd_decap_8
XANTENNA__072__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_20_47 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_4.LATCH_4_.latch_SLEEPB _114_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_12 vpwr vgnd scs8hd_fill_2
XFILLER_29_23 vpwr vgnd scs8hd_fill_2
XFILLER_29_78 vpwr vgnd scs8hd_fill_2
XFILLER_61_98 vgnd vpwr scs8hd_decap_12
XFILLER_61_65 vpwr vgnd scs8hd_fill_2
XFILLER_6_27 vpwr vgnd scs8hd_fill_2
XFILLER_13_7 vgnd vpwr scs8hd_decap_12
XFILLER_19_143 vgnd vpwr scs8hd_decap_3
XANTENNA__157__B _147_/D vgnd vpwr scs8hd_diode_2
XFILLER_34_102 vpwr vgnd scs8hd_fill_2
XFILLER_34_113 vgnd vpwr scs8hd_decap_12
XANTENNA__173__A _179_/B vgnd vpwr scs8hd_diode_2
XFILLER_25_135 vgnd vpwr scs8hd_decap_8
XANTENNA__083__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_31_57 vpwr vgnd scs8hd_fill_2
XFILLER_56_32 vpwr vgnd scs8hd_fill_2
XFILLER_56_87 vgnd vpwr scs8hd_decap_3
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_102 vgnd vpwr scs8hd_decap_12
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_ipin_6.LATCH_1_.latch/Q mux_left_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__168__A _102_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_127 vgnd vpwr scs8hd_decap_12
XFILLER_7_92 vgnd vpwr scs8hd_fill_1
XANTENNA__078__A _078_/A vgnd vpwr scs8hd_diode_2
XFILLER_42_45 vpwr vgnd scs8hd_fill_2
XFILLER_9_109 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_142 vgnd vpwr scs8hd_decap_4
XANTENNA__170__B _168_/B vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_left_ipin_3.LATCH_4_.latch/Q mux_left_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_15 vgnd vpwr scs8hd_decap_4
XFILLER_12_48 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _188_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__080__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_37_78 vgnd vpwr scs8hd_decap_8
XFILLER_53_88 vgnd vpwr scs8hd_decap_3
XFILLER_53_22 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_ipin_2.LATCH_5_.latch_SLEEPB _179_/Y vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_1.LATCH_0_.latch data_in mem_left_ipin_1.LATCH_0_.latch/Q _178_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_123 vgnd vpwr scs8hd_decap_12
XFILLER_5_112 vgnd vpwr scs8hd_decap_8
XFILLER_5_101 vgnd vpwr scs8hd_decap_4
XANTENNA__165__B _168_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__075__B _095_/B vgnd vpwr scs8hd_diode_2
XANTENNA__091__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_58 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_48_66 vpwr vgnd scs8hd_fill_2
XFILLER_64_87 vgnd vpwr scs8hd_decap_6
XFILLER_64_32 vgnd vpwr scs8hd_decap_12
XFILLER_0_18 vgnd vpwr scs8hd_decap_4
Xmem_left_ipin_3.LATCH_3_.latch data_in mem_left_ipin_3.LATCH_3_.latch/Q _101_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_38 vgnd vpwr scs8hd_decap_4
X_186_ _186_/HI _186_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_ipin_4.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA__176__A _102_/A vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _188_/HI mem_left_ipin_7.LATCH_5_.latch/Q
+ mux_left_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_55_144 vpwr vgnd scs8hd_fill_2
XANTENNA__086__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_34_46 vpwr vgnd scs8hd_fill_2
XFILLER_59_32 vpwr vgnd scs8hd_fill_2
XFILLER_1_3 vgnd vpwr scs8hd_decap_12
X_169_ _104_/A _168_/B _169_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XFILLER_52_125 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_61_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_ipin_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_3.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[3] mux_left_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_ipin_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__157__C _069_/C vgnd vpwr scs8hd_diode_2
XFILLER_34_125 vgnd vpwr scs8hd_decap_12
XANTENNA__173__B _177_/B vgnd vpwr scs8hd_diode_2
XFILLER_40_106 vgnd vpwr scs8hd_decap_4
XFILLER_15_48 vpwr vgnd scs8hd_fill_2
XANTENNA__083__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_3.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_0.LATCH_3_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
XFILLER_56_11 vgnd vpwr scs8hd_decap_3
XFILLER_16_114 vgnd vpwr scs8hd_decap_12
XPHY_120 vgnd vpwr scs8hd_decap_3
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_106 vgnd vpwr scs8hd_decap_12
XFILLER_21_91 vpwr vgnd scs8hd_fill_2
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_ipin_3.LATCH_2_.latch/Q mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA__168__B _168_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_139 vgnd vpwr scs8hd_decap_6
XFILLER_7_71 vpwr vgnd scs8hd_fill_2
XANTENNA__094__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_26_36 vpwr vgnd scs8hd_fill_2
XANTENNA__179__A _079_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_5.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_12_27 vpwr vgnd scs8hd_fill_2
XANTENNA__080__C address[0] vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_ipin_1.LATCH_0_.latch/Q mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_left_ipin_6.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__089__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_37_57 vpwr vgnd scs8hd_fill_2
XFILLER_53_34 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_7.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_135 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_ipin_2.INVTX1_1_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_64_3 vgnd vpwr scs8hd_decap_12
Xmem_left_ipin_6.LATCH_2_.latch data_in mem_left_ipin_6.LATCH_2_.latch/Q _134_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_83 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_6.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__075__C address[3] vgnd vpwr scs8hd_diode_2
XFILLER_48_23 vgnd vpwr scs8hd_decap_8
XFILLER_64_44 vgnd vpwr scs8hd_decap_12
XFILLER_9_17 vpwr vgnd scs8hd_fill_2
X_185_ _185_/HI _185_/LO vgnd vpwr scs8hd_conb_1
XFILLER_64_145 vgnd vpwr scs8hd_fill_1
XANTENNA__176__B _177_/B vgnd vpwr scs8hd_diode_2
XANTENNA__192__A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_5.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_112 vpwr vgnd scs8hd_fill_2
XANTENNA__086__B address[2] vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_4.tap_buf4_0_.scs8hd_inv_1 mux_left_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ right_grid_pin_8_ vgnd vpwr scs8hd_inv_1
XFILLER_18_59 vgnd vpwr scs8hd_decap_4
XFILLER_59_77 vpwr vgnd scs8hd_fill_2
XFILLER_59_55 vgnd vpwr scs8hd_decap_4
Xmux_left_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_ipin_5.LATCH_1_.latch/Q mux_left_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_left_ipin_7.LATCH_5_.latch_SLEEPB _139_/Y vgnd vpwr scs8hd_diode_2
X_168_ _102_/A _168_/B _168_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_80 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_099_ _099_/A _100_/B vgnd vpwr scs8hd_buf_1
XFILLER_27_3 vgnd vpwr scs8hd_decap_12
XFILLER_52_137 vgnd vpwr scs8hd_decap_8
XFILLER_1_73 vpwr vgnd scs8hd_fill_2
XFILLER_37_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_ipin_1.LATCH_0_.latch_SLEEPB _178_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_5_ vgnd vpwr scs8hd_inv_1
XFILLER_45_57 vpwr vgnd scs8hd_fill_2
XFILLER_45_35 vgnd vpwr scs8hd_fill_1
XFILLER_43_126 vgnd vpwr scs8hd_decap_12
XFILLER_43_115 vgnd vpwr scs8hd_decap_6
XANTENNA__097__A _139_/A vgnd vpwr scs8hd_diode_2
XFILLER_61_56 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_123 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_left_ipin_2.LATCH_4_.latch/Q mux_left_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_34_137 vgnd vpwr scs8hd_decap_8
XFILLER_15_16 vpwr vgnd scs8hd_fill_2
XFILLER_15_27 vpwr vgnd scs8hd_fill_2
XANTENNA__083__C _069_/C vgnd vpwr scs8hd_diode_2
XFILLER_56_23 vgnd vpwr scs8hd_decap_8
XFILLER_16_126 vgnd vpwr scs8hd_decap_12
XPHY_121 vgnd vpwr scs8hd_decap_3
XPHY_110 vgnd vpwr scs8hd_decap_3
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_118 vgnd vpwr scs8hd_decap_4
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1 vgnd vpwr scs8hd_decap_3
Xmux_left_ipin_1.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[1] mux_left_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_15 vgnd vpwr scs8hd_decap_4
XFILLER_3_19 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _187_/HI mem_left_ipin_6.LATCH_5_.latch/Q
+ mux_left_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__179__B _179_/B vgnd vpwr scs8hd_diode_2
XANTENNA__195__A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_7.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_36 vpwr vgnd scs8hd_fill_2
XFILLER_53_57 vpwr vgnd scs8hd_fill_2
XFILLER_57_3 vgnd vpwr scs8hd_decap_12
XFILLER_23_38 vpwr vgnd scs8hd_fill_2
XFILLER_23_49 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_56 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_184_ _184_/HI _184_/LO vgnd vpwr scs8hd_conb_1
XFILLER_49_121 vgnd vpwr scs8hd_fill_1
XFILLER_29_7 vpwr vgnd scs8hd_fill_2
XFILLER_49_143 vgnd vpwr scs8hd_decap_3
XANTENNA__086__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XFILLER_59_23 vgnd vpwr scs8hd_decap_3
XFILLER_46_102 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_ipin_2.LATCH_2_.latch/Q mux_left_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_40_80 vgnd vpwr scs8hd_decap_4
X_098_ address[1] _098_/B address[0] _099_/A vgnd vpwr scs8hd_or3_4
X_167_ _151_/A _168_/B _167_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_113 vgnd vpwr scs8hd_decap_8
XFILLER_1_85 vpwr vgnd scs8hd_fill_2
XFILLER_37_135 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_14 vpwr vgnd scs8hd_fill_2
XFILLER_28_102 vgnd vpwr scs8hd_decap_12
XANTENNA__097__B _101_/B vgnd vpwr scs8hd_diode_2
XFILLER_43_138 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_135 vgnd vpwr scs8hd_decap_8
Xmux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_0_.latch/Q mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__198__A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_38 vpwr vgnd scs8hd_fill_2
XPHY_100 vgnd vpwr scs8hd_decap_3
XFILLER_16_138 vgnd vpwr scs8hd_decap_8
XPHY_122 vgnd vpwr scs8hd_decap_3
XPHY_111 vgnd vpwr scs8hd_decap_3
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_22_108 vgnd vpwr scs8hd_decap_4
XFILLER_7_95 vgnd vpwr scs8hd_fill_1
XFILLER_7_51 vpwr vgnd scs8hd_fill_2
XFILLER_30_141 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_ipin_6.LATCH_0_.latch_SLEEPB _136_/Y vgnd vpwr scs8hd_diode_2
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XFILLER_13_108 vgnd vpwr scs8hd_decap_12
XFILLER_16_71 vpwr vgnd scs8hd_fill_2
XFILLER_16_82 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_ipin_4.LATCH_1_.latch/Q mux_left_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_37_15 vgnd vpwr scs8hd_decap_4
XFILLER_27_70 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_9 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_ipin_1.INVTX1_5_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_48_47 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_ipin_1.LATCH_4_.latch/Q mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_13_72 vpwr vgnd scs8hd_fill_2
X_183_ _183_/HI _183_/LO vgnd vpwr scs8hd_conb_1
XFILLER_49_111 vgnd vpwr scs8hd_decap_8
XFILLER_64_125 vgnd vpwr scs8hd_decap_12
XFILLER_38_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_2.LATCH_2_.latch data_in mem_left_ipin_2.LATCH_2_.latch/Q _082_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_left_ipin_6.INVTX1_3_.scs8hd_inv_1 chany_top_in[5] mux_left_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_46_114 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_ipin_4.LATCH_1_.latch_SLEEPB _117_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_166_ _132_/A _168_/B _166_/Y vgnd vpwr scs8hd_nor2_4
X_097_ _139_/A _101_/B _097_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_49_90 vpwr vgnd scs8hd_fill_2
XFILLER_1_53 vpwr vgnd scs8hd_fill_2
XFILLER_20_29 vpwr vgnd scs8hd_fill_2
Xmem_left_ipin_4.LATCH_5_.latch data_in mem_left_ipin_4.LATCH_5_.latch/Q _112_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_16 vpwr vgnd scs8hd_fill_2
XFILLER_29_27 vpwr vgnd scs8hd_fill_2
XFILLER_45_48 vpwr vgnd scs8hd_fill_2
XFILLER_28_114 vgnd vpwr scs8hd_decap_12
XFILLER_61_69 vgnd vpwr scs8hd_decap_3
XFILLER_10_73 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _186_/HI mem_left_ipin_5.LATCH_5_.latch/Q
+ mux_left_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_10_84 vgnd vpwr scs8hd_decap_6
XFILLER_19_82 vpwr vgnd scs8hd_fill_2
XFILLER_19_93 vpwr vgnd scs8hd_fill_2
XFILLER_34_106 vgnd vpwr scs8hd_decap_4
XFILLER_35_92 vgnd vpwr scs8hd_fill_1
X_149_ _139_/A _149_/B _149_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_32_3 vgnd vpwr scs8hd_decap_8
XFILLER_31_17 vpwr vgnd scs8hd_fill_2
XFILLER_56_36 vpwr vgnd scs8hd_fill_2
XPHY_123 vgnd vpwr scs8hd_decap_3
XPHY_112 vgnd vpwr scs8hd_decap_3
XPHY_101 vgnd vpwr scs8hd_decap_3
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_ipin_3.tap_buf4_0_.scs8hd_inv_1_A mux_left_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_42_49 vpwr vgnd scs8hd_fill_2
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_8_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_60 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_2.LATCH_2_.latch_SLEEPB _082_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_19 vgnd vpwr scs8hd_fill_1
Xmux_left_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_ipin_1.LATCH_2_.latch/Q mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_53_15 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_ipin_3.INVTX1_3_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_5.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_7.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_48_15 vgnd vpwr scs8hd_decap_4
XFILLER_2_119 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_145 vgnd vpwr scs8hd_fill_1
X_182_ _182_/HI _182_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_40 vpwr vgnd scs8hd_fill_2
XFILLER_13_62 vgnd vpwr scs8hd_decap_3
XFILLER_49_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_1_130 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_5.LATCH_1_.latch data_in mem_left_ipin_5.LATCH_1_.latch/Q _127_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_64_137 vgnd vpwr scs8hd_decap_8
XANTENNA__100__A _101_/B vgnd vpwr scs8hd_diode_2
XFILLER_62_3 vgnd vpwr scs8hd_decap_12
Xmem_right_ipin_0.LATCH_5_.latch data_in mem_right_ipin_0.LATCH_5_.latch/Q _149_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_left_ipin_3.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_50_38 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_36 vpwr vgnd scs8hd_fill_2
XFILLER_46_126 vgnd vpwr scs8hd_decap_12
Xmem_left_ipin_7.LATCH_4_.latch data_in mem_left_ipin_7.LATCH_4_.latch/Q _140_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_165_ _179_/B _168_/B _165_/Y vgnd vpwr scs8hd_nor2_4
X_096_ _095_/X _101_/B vgnd vpwr scs8hd_buf_1
XFILLER_1_32 vpwr vgnd scs8hd_fill_2
XFILLER_1_98 vpwr vgnd scs8hd_fill_2
XFILLER_20_19 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_0.LATCH_3_.latch_SLEEPB _167_/Y vgnd vpwr scs8hd_diode_2
XFILLER_45_38 vgnd vpwr scs8hd_fill_1
XFILLER_28_126 vgnd vpwr scs8hd_decap_12
XFILLER_61_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_41 vgnd vpwr scs8hd_decap_3
XFILLER_10_52 vpwr vgnd scs8hd_fill_2
XFILLER_19_104 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_0.LATCH_0_.latch_SLEEPB _154_/Y vgnd vpwr scs8hd_diode_2
X_148_ _148_/A _149_/B vgnd vpwr scs8hd_buf_1
Xmux_left_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_ipin_3.LATCH_1_.latch/Q mux_left_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_3 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_4.INVTX1_3_.scs8hd_inv_1 chany_top_in[4] mux_left_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_079_ _133_/A _079_/B _079_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_124 vgnd vpwr scs8hd_decap_3
XPHY_113 vgnd vpwr scs8hd_decap_3
XPHY_102 vgnd vpwr scs8hd_decap_3
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_40 vpwr vgnd scs8hd_fill_2
XFILLER_21_62 vgnd vpwr scs8hd_fill_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_left_ipin_7.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_95 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_7.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_81 vpwr vgnd scs8hd_fill_2
XFILLER_62_80 vgnd vpwr scs8hd_decap_12
XFILLER_7_20 vgnd vpwr scs8hd_decap_3
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_7_75 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_ipin_0.LATCH_4_.latch/Q mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_26_29 vpwr vgnd scs8hd_fill_2
XFILLER_42_39 vgnd vpwr scs8hd_decap_4
XFILLER_21_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_32_83 vpwr vgnd scs8hd_fill_2
XANTENNA__103__A _142_/A vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_ipin_7.LATCH_2_.latch/Q mux_left_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_5.INVTX1_1_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_53_38 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_1.LATCH_1_.latch data_in _159_/A _155_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_27_83 vpwr vgnd scs8hd_fill_2
XFILLER_4_32 vpwr vgnd scs8hd_fill_2
XFILLER_4_87 vpwr vgnd scs8hd_fill_2
XFILLER_23_19 vpwr vgnd scs8hd_fill_2
XFILLER_58_113 vgnd vpwr scs8hd_decap_12
XFILLER_58_102 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _185_/HI mem_left_ipin_4.LATCH_5_.latch/Q
+ mux_left_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_64_15 vgnd vpwr scs8hd_decap_12
X_181_ _181_/HI _181_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_85 vpwr vgnd scs8hd_fill_2
XFILLER_13_96 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_5.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_7.tap_buf4_0_.scs8hd_inv_1 mux_left_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ right_grid_pin_14_ vgnd vpwr scs8hd_inv_1
XFILLER_49_135 vgnd vpwr scs8hd_decap_8
XANTENNA__100__B _100_/B vgnd vpwr scs8hd_diode_2
XFILLER_55_3 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_ipin_7.LATCH_2_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
XFILLER_55_116 vgnd vpwr scs8hd_decap_4
XFILLER_34_29 vpwr vgnd scs8hd_fill_2
XFILLER_59_15 vgnd vpwr scs8hd_decap_8
XFILLER_46_138 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_1.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__201__A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
X_164_ _164_/A _168_/B vgnd vpwr scs8hd_buf_1
X_095_ _110_/A _095_/B _095_/C _095_/D _095_/X vgnd vpwr scs8hd_or4_4
XFILLER_1_22 vgnd vpwr scs8hd_fill_1
XFILLER_1_77 vpwr vgnd scs8hd_fill_2
XANTENNA__111__A _110_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_138 vgnd vpwr scs8hd_decap_8
XFILLER_61_27 vgnd vpwr scs8hd_decap_12
XFILLER_19_40 vpwr vgnd scs8hd_fill_2
XFILLER_51_60 vgnd vpwr scs8hd_fill_1
X_147_ _110_/A address[4] address[3] _147_/D _148_/A vgnd vpwr scs8hd_or4_4
X_078_ _078_/A _079_/B vgnd vpwr scs8hd_buf_1
XANTENNA__106__A _088_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_3 vgnd vpwr scs8hd_decap_8
Xmux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_2_.latch/Q mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_108 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_4.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_125 vgnd vpwr scs8hd_decap_3
XPHY_114 vgnd vpwr scs8hd_decap_3
XPHY_103 vgnd vpwr scs8hd_decap_3
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_left_ipin_0.LATCH_5_.latch data_in mem_left_ipin_0.LATCH_5_.latch/Q _165_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_74 vpwr vgnd scs8hd_fill_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_26_19 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_ipin_5.LATCH_3_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_2.INVTX1_3_.scs8hd_inv_1 chany_top_in[2] mux_left_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_7.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_41 vpwr vgnd scs8hd_fill_2
XFILLER_16_52 vgnd vpwr scs8hd_decap_8
XANTENNA__103__B _101_/B vgnd vpwr scs8hd_diode_2
XFILLER_57_81 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__204__A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_27_40 vpwr vgnd scs8hd_fill_2
XFILLER_27_62 vgnd vpwr scs8hd_fill_1
XFILLER_43_94 vpwr vgnd scs8hd_fill_2
XFILLER_4_66 vpwr vgnd scs8hd_fill_2
XANTENNA__114__A _132_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_58_125 vgnd vpwr scs8hd_decap_12
XFILLER_64_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_53 vpwr vgnd scs8hd_fill_2
X_180_ _079_/B _100_/B _180_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_110 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_ipin_2.LATCH_1_.latch/Q mux_left_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_64_106 vgnd vpwr scs8hd_decap_12
XFILLER_38_72 vgnd vpwr scs8hd_decap_4
XFILLER_38_83 vgnd vpwr scs8hd_decap_8
XFILLER_54_82 vpwr vgnd scs8hd_fill_2
XFILLER_54_71 vpwr vgnd scs8hd_fill_2
XANTENNA__109__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_48_3 vgnd vpwr scs8hd_decap_12
XFILLER_24_41 vgnd vpwr scs8hd_decap_3
XFILLER_24_63 vpwr vgnd scs8hd_fill_2
X_163_ _110_/A address[4] address[3] _095_/D _164_/A vgnd vpwr scs8hd_or4_4
X_094_ address[3] _095_/C vgnd vpwr scs8hd_inv_8
XANTENNA_mem_left_ipin_3.LATCH_4_.latch_SLEEPB _100_/Y vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_1.LATCH_1_.latch data_in mem_left_ipin_1.LATCH_1_.latch/Q _177_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_18 vpwr vgnd scs8hd_fill_2
XFILLER_61_39 vpwr vgnd scs8hd_fill_2
XFILLER_51_120 vpwr vgnd scs8hd_fill_2
XFILLER_35_73 vpwr vgnd scs8hd_fill_2
XFILLER_35_95 vgnd vpwr scs8hd_fill_1
Xmux_left_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_ipin_6.LATCH_2_.latch/Q mux_left_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
X_146_ _145_/X _147_/D vgnd vpwr scs8hd_buf_1
XANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _162_/A vgnd vpwr
+ scs8hd_diode_2
X_077_ _095_/D _077_/B _078_/A vgnd vpwr scs8hd_or2_4
XANTENNA__122__A _121_/X vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_3.LATCH_4_.latch data_in mem_left_ipin_3.LATCH_4_.latch/Q _100_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_33_120 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_0_.latch/Q mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_126 vgnd vpwr scs8hd_decap_3
XPHY_115 vgnd vpwr scs8hd_decap_3
XANTENNA__207__A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XPHY_104 vgnd vpwr scs8hd_decap_3
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_131 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_53 vpwr vgnd scs8hd_fill_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_62_93 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_0.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[8] mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_7_88 vgnd vpwr scs8hd_decap_4
XFILLER_7_55 vpwr vgnd scs8hd_fill_2
XANTENNA__117__A _135_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_145 vgnd vpwr scs8hd_fill_1
Xmux_left_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _184_/HI mem_left_ipin_3.LATCH_5_.latch/Q
+ mux_left_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_7_99 vpwr vgnd scs8hd_fill_2
X_129_ _077_/B _110_/D _130_/A vgnd vpwr scs8hd_or2_4
XFILLER_21_123 vgnd vpwr scs8hd_decap_12
XFILLER_16_75 vpwr vgnd scs8hd_fill_2
XFILLER_16_86 vgnd vpwr scs8hd_decap_6
XFILLER_12_145 vgnd vpwr scs8hd_fill_1
XFILLER_32_96 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_1.LATCH_5_.latch_SLEEPB _173_/Y vgnd vpwr scs8hd_diode_2
XFILLER_53_18 vgnd vpwr scs8hd_decap_4
XFILLER_5_108 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_62 vpwr vgnd scs8hd_fill_2
XFILLER_43_51 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_0.INVTX1_3_.scs8hd_inv_1 chany_top_in[4] mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_right_ipin_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__114__B _118_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_4.INVTX1_5_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA__130__A _130_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_23 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_ipin_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_58_137 vgnd vpwr scs8hd_decap_8
XFILLER_13_21 vpwr vgnd scs8hd_fill_2
XFILLER_8_3 vgnd vpwr scs8hd_decap_8
XFILLER_64_118 vgnd vpwr scs8hd_decap_6
XFILLER_54_61 vgnd vpwr scs8hd_fill_1
XANTENNA__109__B _145_/B vgnd vpwr scs8hd_diode_2
XANTENNA__125__A _133_/A vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_6.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[1] mux_left_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_50_19 vgnd vpwr scs8hd_decap_12
Xmem_left_ipin_4.LATCH_0_.latch data_in mem_left_ipin_4.LATCH_0_.latch/Q _118_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_162_ _162_/A _162_/Y vgnd vpwr scs8hd_inv_8
XFILLER_24_86 vgnd vpwr scs8hd_fill_1
X_093_ _093_/A _110_/A vgnd vpwr scs8hd_buf_1
XFILLER_40_52 vpwr vgnd scs8hd_fill_2
XFILLER_49_94 vpwr vgnd scs8hd_fill_2
XFILLER_60_121 vgnd vpwr scs8hd_decap_12
XFILLER_1_57 vpwr vgnd scs8hd_fill_2
XFILLER_60_3 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_7.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[7] mux_left_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_51_143 vgnd vpwr scs8hd_decap_3
Xmem_left_ipin_6.LATCH_3_.latch data_in mem_left_ipin_6.LATCH_3_.latch/Q _133_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_77 vgnd vpwr scs8hd_decap_4
XFILLER_19_53 vpwr vgnd scs8hd_fill_2
XFILLER_42_121 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_ipin_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_86 vpwr vgnd scs8hd_fill_2
XFILLER_19_97 vpwr vgnd scs8hd_fill_2
XFILLER_51_40 vpwr vgnd scs8hd_fill_2
X_145_ address[5] _145_/B _145_/X vgnd vpwr scs8hd_or2_4
X_076_ _075_/X _077_/B vgnd vpwr scs8hd_buf_1
XFILLER_33_143 vgnd vpwr scs8hd_decap_3
XPHY_116 vgnd vpwr scs8hd_decap_3
XPHY_105 vgnd vpwr scs8hd_decap_3
XFILLER_24_143 vgnd vpwr scs8hd_decap_3
XPHY_127 vgnd vpwr scs8hd_decap_3
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_5.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_143 vgnd vpwr scs8hd_decap_3
XANTENNA__133__A _133_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_34 vpwr vgnd scs8hd_fill_2
XFILLER_7_12 vpwr vgnd scs8hd_fill_2
XANTENNA__117__B _118_/B vgnd vpwr scs8hd_diode_2
X_128_ _144_/A _124_/B _128_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_3 vgnd vpwr scs8hd_decap_6
XFILLER_21_135 vgnd vpwr scs8hd_decap_8
Xmux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_ipin_1.LATCH_1_.latch/Q mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_102 vgnd vpwr scs8hd_decap_8
XFILLER_12_113 vgnd vpwr scs8hd_decap_12
XFILLER_16_10 vpwr vgnd scs8hd_fill_2
XFILLER_8_106 vgnd vpwr scs8hd_decap_12
XFILLER_32_64 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_2.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_57_94 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__128__A _144_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_3.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_6.INVTX1_3_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_4.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_27_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_5.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1 mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ right_grid_pin_0_ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_19 vgnd vpwr scs8hd_fill_1
Xmem_right_ipin_0.LATCH_0_.latch data_in mem_right_ipin_0.LATCH_0_.latch/Q _154_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_ipin_5.LATCH_2_.latch/Q mux_left_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_134 vgnd vpwr scs8hd_decap_12
XFILLER_38_96 vpwr vgnd scs8hd_fill_2
XANTENNA__125__B _124_/B vgnd vpwr scs8hd_diode_2
XANTENNA__141__A _133_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_6.LATCH_5_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
X_161_ _161_/A _161_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mem_left_ipin_0.LATCH_0_.latch_SLEEPB _170_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_7.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_86 vgnd vpwr scs8hd_decap_4
X_092_ _179_/B _139_/A vgnd vpwr scs8hd_buf_1
Xmux_left_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _183_/HI mem_left_ipin_2.LATCH_5_.latch/Q
+ mux_left_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_49_73 vpwr vgnd scs8hd_fill_2
XFILLER_49_40 vpwr vgnd scs8hd_fill_2
XFILLER_1_36 vpwr vgnd scs8hd_fill_2
XFILLER_60_133 vgnd vpwr scs8hd_decap_12
XFILLER_53_3 vgnd vpwr scs8hd_decap_12
XANTENNA__136__A _144_/A vgnd vpwr scs8hd_diode_2
XFILLER_51_100 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_12 vpwr vgnd scs8hd_fill_2
XFILLER_10_23 vpwr vgnd scs8hd_fill_2
XFILLER_10_56 vgnd vpwr scs8hd_decap_4
Xmux_left_ipin_4.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[3] mux_left_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_65 vpwr vgnd scs8hd_fill_2
XFILLER_19_108 vgnd vpwr scs8hd_decap_12
XFILLER_42_133 vgnd vpwr scs8hd_decap_12
XFILLER_35_53 vgnd vpwr scs8hd_decap_3
XFILLER_51_96 vpwr vgnd scs8hd_fill_2
XFILLER_51_85 vpwr vgnd scs8hd_fill_2
X_144_ _144_/A _139_/B _144_/Y vgnd vpwr scs8hd_nor2_4
X_075_ _093_/A _095_/B address[3] _075_/X vgnd vpwr scs8hd_or3_4
XANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_128 vgnd vpwr scs8hd_decap_3
XPHY_117 vgnd vpwr scs8hd_decap_3
XPHY_106 vgnd vpwr scs8hd_decap_3
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_ipin_5.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[5] mux_left_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_22 vgnd vpwr scs8hd_decap_3
XFILLER_46_85 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_15_111 vgnd vpwr scs8hd_decap_8
XANTENNA__133__B _131_/B vgnd vpwr scs8hd_diode_2
X_127_ _135_/A _124_/B _127_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_21_114 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_ipin_4.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_8_118 vgnd vpwr scs8hd_decap_12
XFILLER_12_125 vgnd vpwr scs8hd_decap_12
XFILLER_32_43 vpwr vgnd scs8hd_fill_2
XFILLER_32_87 vgnd vpwr scs8hd_decap_3
XFILLER_57_51 vgnd vpwr scs8hd_decap_4
XFILLER_57_73 vpwr vgnd scs8hd_fill_2
XANTENNA__144__A _144_/A vgnd vpwr scs8hd_diode_2
XANTENNA__128__B _124_/B vgnd vpwr scs8hd_diode_2
XFILLER_27_87 vpwr vgnd scs8hd_fill_2
XFILLER_43_75 vpwr vgnd scs8hd_fill_2
XFILLER_4_36 vpwr vgnd scs8hd_fill_2
XANTENNA__139__A _139_/A vgnd vpwr scs8hd_diode_2
XFILLER_58_106 vgnd vpwr scs8hd_decap_4
XFILLER_1_102 vgnd vpwr scs8hd_decap_4
XFILLER_13_89 vgnd vpwr scs8hd_decap_4
XFILLER_38_53 vpwr vgnd scs8hd_fill_2
XANTENNA__141__B _139_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_4.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_11 vgnd vpwr scs8hd_decap_3
X_160_ _160_/A _160_/Y vgnd vpwr scs8hd_inv_8
X_091_ _091_/A _179_/B vgnd vpwr scs8hd_buf_1
XFILLER_40_32 vgnd vpwr scs8hd_decap_6
XFILLER_45_120 vpwr vgnd scs8hd_fill_2
XFILLER_1_15 vgnd vpwr scs8hd_fill_1
XFILLER_37_109 vpwr vgnd scs8hd_fill_2
XFILLER_60_145 vgnd vpwr scs8hd_fill_1
XANTENNA__136__B _131_/B vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_2.INVTX1_1_.scs8hd_inv_1 chany_top_in[1] mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__152__A _142_/A vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_1_.latch/Q mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_46_3 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _161_/A mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_51_123 vgnd vpwr scs8hd_decap_12
XFILLER_51_112 vgnd vpwr scs8hd_decap_8
XFILLER_10_46 vgnd vpwr scs8hd_decap_3
XFILLER_19_22 vgnd vpwr scs8hd_decap_3
XFILLER_42_145 vgnd vpwr scs8hd_fill_1
XFILLER_35_65 vpwr vgnd scs8hd_fill_2
XFILLER_51_53 vgnd vpwr scs8hd_decap_4
X_143_ _135_/A _139_/B _143_/Y vgnd vpwr scs8hd_nor2_4
X_074_ address[4] _095_/B vgnd vpwr scs8hd_inv_8
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_0.LATCH_0_.latch data_in mem_left_ipin_0.LATCH_0_.latch/Q _170_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_112 vgnd vpwr scs8hd_decap_8
XFILLER_33_123 vgnd vpwr scs8hd_decap_12
XANTENNA__147__A _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_91 vgnd vpwr scs8hd_fill_1
XPHY_129 vgnd vpwr scs8hd_decap_3
XPHY_118 vgnd vpwr scs8hd_decap_3
XPHY_107 vgnd vpwr scs8hd_decap_3
XFILLER_21_78 vpwr vgnd scs8hd_fill_2
XFILLER_46_64 vgnd vpwr scs8hd_decap_6
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_123 vgnd vpwr scs8hd_decap_12
Xmem_left_ipin_2.LATCH_3_.latch data_in mem_left_ipin_2.LATCH_3_.latch/Q _079_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_left_ipin_2.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[1] mux_left_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_ipin_5.LATCH_0_.latch_SLEEPB _128_/Y vgnd vpwr scs8hd_diode_2
X_126_ _142_/A _124_/B _126_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_30_6 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_ipin_4.LATCH_2_.latch/Q mux_left_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_23 vpwr vgnd scs8hd_fill_2
XFILLER_12_137 vgnd vpwr scs8hd_decap_8
XFILLER_16_45 vpwr vgnd scs8hd_fill_2
XFILLER_32_11 vgnd vpwr scs8hd_decap_3
XFILLER_32_77 vgnd vpwr scs8hd_decap_4
Xmux_left_ipin_3.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[7] mux_left_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__144__B _139_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_109_ address[5] _145_/B _110_/D vgnd vpwr scs8hd_nand2_4
XANTENNA__160__A _160_/A vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _182_/HI mem_left_ipin_1.LATCH_5_.latch/Q
+ mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__070__A _069_/X vgnd vpwr scs8hd_diode_2
XFILLER_27_66 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_0.LATCH_5_.latch_SLEEPB _149_/Y vgnd vpwr scs8hd_diode_2
XFILLER_43_98 vpwr vgnd scs8hd_fill_2
XFILLER_4_15 vgnd vpwr scs8hd_fill_1
XANTENNA__139__B _139_/B vgnd vpwr scs8hd_diode_2
XANTENNA__155__A _120_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_13_57 vpwr vgnd scs8hd_fill_2
XFILLER_13_68 vpwr vgnd scs8hd_fill_2
XFILLER_1_114 vpwr vgnd scs8hd_fill_2
XFILLER_49_107 vpwr vgnd scs8hd_fill_2
XFILLER_38_32 vgnd vpwr scs8hd_decap_4
XFILLER_54_86 vgnd vpwr scs8hd_decap_4
XFILLER_54_75 vgnd vpwr scs8hd_decap_4
XFILLER_54_53 vgnd vpwr scs8hd_decap_8
XFILLER_54_20 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _161_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_63_143 vgnd vpwr scs8hd_decap_3
XFILLER_63_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_ipin_3.LATCH_1_.latch_SLEEPB _105_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_23 vgnd vpwr scs8hd_decap_4
XFILLER_24_67 vpwr vgnd scs8hd_fill_2
X_090_ address[1] _098_/B _069_/C _091_/A vgnd vpwr scs8hd_or3_4
XFILLER_24_89 vgnd vpwr scs8hd_decap_3
XFILLER_49_53 vpwr vgnd scs8hd_fill_2
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
XFILLER_45_143 vgnd vpwr scs8hd_decap_3
XANTENNA__152__B _149_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_2.tap_buf4_0_.scs8hd_inv_1_A mux_left_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_3 vgnd vpwr scs8hd_decap_8
XFILLER_51_135 vgnd vpwr scs8hd_decap_8
XFILLER_27_121 vgnd vpwr scs8hd_fill_1
XFILLER_27_143 vgnd vpwr scs8hd_decap_3
XFILLER_35_33 vgnd vpwr scs8hd_decap_3
X_142_ _142_/A _139_/B _142_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_35_88 vgnd vpwr scs8hd_decap_4
XFILLER_51_65 vpwr vgnd scs8hd_fill_2
X_073_ enable _093_/A vgnd vpwr scs8hd_inv_8
XANTENNA__147__B address[4] vgnd vpwr scs8hd_diode_2
XFILLER_33_135 vgnd vpwr scs8hd_decap_8
XANTENNA__163__A _110_/A vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_5.LATCH_2_.latch data_in mem_left_ipin_5.LATCH_2_.latch/Q _126_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_ipin_0.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_119 vgnd vpwr scs8hd_decap_3
XPHY_108 vgnd vpwr scs8hd_decap_3
XANTENNA__073__A enable vgnd vpwr scs8hd_diode_2
XFILLER_21_57 vpwr vgnd scs8hd_fill_2
XFILLER_46_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_135 vgnd vpwr scs8hd_decap_8
X_125_ _133_/A _124_/B _125_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_59 vpwr vgnd scs8hd_fill_2
XFILLER_30_105 vgnd vpwr scs8hd_decap_12
XFILLER_11_90 vpwr vgnd scs8hd_fill_2
Xmem_left_ipin_7.LATCH_5_.latch data_in mem_left_ipin_7.LATCH_5_.latch/Q _139_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__158__A _077_/B vgnd vpwr scs8hd_diode_2
XANTENNA__068__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_1.LATCH_2_.latch_SLEEPB _176_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_3.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
X_108_ address[6] _145_/B vgnd vpwr scs8hd_inv_8
XFILLER_21_3 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_0.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_ipin_7.INVTX1_5_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_27_23 vpwr vgnd scs8hd_fill_2
XFILLER_43_55 vgnd vpwr scs8hd_decap_6
XFILLER_43_22 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _159_/A mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_4_145 vgnd vpwr scs8hd_fill_1
XFILLER_4_49 vpwr vgnd scs8hd_fill_2
XANTENNA__155__B _147_/D vgnd vpwr scs8hd_diode_2
XANTENNA__171__A _095_/D vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_1.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[5] mux_left_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_7.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_25 vpwr vgnd scs8hd_fill_2
XFILLER_13_36 vpwr vgnd scs8hd_fill_2
XANTENNA__081__A _080_/X vgnd vpwr scs8hd_diode_2
XFILLER_1_126 vpwr vgnd scs8hd_fill_2
XFILLER_54_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__166__A _132_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_70 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_7.INVTX1_1_.scs8hd_inv_1 chany_top_in[2] mux_left_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__076__A _075_/X vgnd vpwr scs8hd_diode_2
XFILLER_24_46 vgnd vpwr scs8hd_decap_6
XFILLER_40_23 vpwr vgnd scs8hd_fill_2
XFILLER_40_56 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_ipin_3.LATCH_2_.latch/Q mux_left_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_57 vpwr vgnd scs8hd_fill_2
XFILLER_27_100 vpwr vgnd scs8hd_fill_2
XFILLER_27_111 vpwr vgnd scs8hd_fill_2
XFILLER_35_23 vgnd vpwr scs8hd_decap_3
X_141_ _133_/A _139_/B _141_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_51_33 vgnd vpwr scs8hd_fill_1
X_072_ address[5] address[6] _095_/D vgnd vpwr scs8hd_or2_4
XANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__147__C address[3] vgnd vpwr scs8hd_diode_2
XANTENNA__163__B address[4] vgnd vpwr scs8hd_diode_2
XFILLER_51_3 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _181_/HI mem_left_ipin_0.LATCH_5_.latch/Q
+ mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_5.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_109 vgnd vpwr scs8hd_decap_3
XFILLER_21_36 vpwr vgnd scs8hd_fill_2
XFILLER_46_11 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_ipin_5.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_62_32 vgnd vpwr scs8hd_decap_12
XFILLER_30_117 vgnd vpwr scs8hd_decap_12
X_124_ _132_/A _124_/B _124_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_38 vpwr vgnd scs8hd_fill_2
XFILLER_7_16 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_6.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__158__B _147_/D vgnd vpwr scs8hd_diode_2
XFILLER_16_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_7.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__174__A _100_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_5.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__084__A _083_/X vgnd vpwr scs8hd_diode_2
XFILLER_57_98 vpwr vgnd scs8hd_fill_2
XFILLER_57_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_143 vgnd vpwr scs8hd_decap_3
XFILLER_7_121 vgnd vpwr scs8hd_fill_1
X_107_ _144_/A _101_/B _107_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__169__A _104_/A vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_3.tap_buf4_0_.scs8hd_inv_1 mux_left_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ right_grid_pin_6_ vgnd vpwr scs8hd_inv_1
XFILLER_27_57 vpwr vgnd scs8hd_fill_2
XANTENNA__079__A _133_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_113 vgnd vpwr scs8hd_decap_12
XFILLER_4_102 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_4.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__155__C _069_/C vgnd vpwr scs8hd_diode_2
XANTENNA__171__B _120_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_1_ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_ipin_6.LATCH_2_.latch_SLEEPB _134_/Y vgnd vpwr scs8hd_diode_2
XFILLER_38_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_123 vgnd vpwr scs8hd_decap_12
XANTENNA__166__B _168_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_7.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_60 vgnd vpwr scs8hd_fill_1
XFILLER_54_145 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__092__A _179_/B vgnd vpwr scs8hd_diode_2
XFILLER_49_77 vpwr vgnd scs8hd_fill_2
XFILLER_1_18 vpwr vgnd scs8hd_fill_2
XFILLER_45_123 vgnd vpwr scs8hd_decap_12
XANTENNA__177__A _104_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_145 vgnd vpwr scs8hd_fill_1
XFILLER_51_104 vgnd vpwr scs8hd_decap_6
XFILLER_10_16 vpwr vgnd scs8hd_fill_2
XFILLER_10_27 vpwr vgnd scs8hd_fill_2
XFILLER_19_36 vpwr vgnd scs8hd_fill_2
XFILLER_19_69 vpwr vgnd scs8hd_fill_2
XFILLER_42_104 vpwr vgnd scs8hd_fill_2
XANTENNA__087__A _086_/X vgnd vpwr scs8hd_diode_2
XFILLER_27_123 vgnd vpwr scs8hd_decap_12
X_140_ _132_/A _139_/B _140_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_51_89 vpwr vgnd scs8hd_fill_2
X_071_ _151_/A _133_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_5.INVTX1_1_.scs8hd_inv_1 chany_top_in[0] mux_left_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_ipin_7.tap_buf4_0_.scs8hd_inv_1_A mux_left_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XPHY_90 vgnd vpwr scs8hd_decap_3
XANTENNA__147__D _147_/D vgnd vpwr scs8hd_diode_2
XANTENNA__163__C address[3] vgnd vpwr scs8hd_diode_2
XFILLER_44_3 vgnd vpwr scs8hd_decap_8
XFILLER_21_15 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_ipin_0.LATCH_3_.latch/Q mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_46_23 vgnd vpwr scs8hd_decap_8
XFILLER_62_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_6.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_7.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_46_89 vgnd vpwr scs8hd_fill_1
XFILLER_30_129 vgnd vpwr scs8hd_decap_12
X_123_ _139_/A _124_/B _123_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_left_ipin_4.LATCH_3_.latch_SLEEPB _115_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_6.INVTX1_5_.scs8hd_inv_1 chany_top_in[6] mux_left_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__158__C address[0] vgnd vpwr scs8hd_diode_2
XANTENNA__174__B _177_/B vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_1.LATCH_2_.latch data_in mem_left_ipin_1.LATCH_2_.latch/Q _176_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_47 vgnd vpwr scs8hd_decap_4
XFILLER_57_77 vpwr vgnd scs8hd_fill_2
X_106_ _088_/B _144_/A vgnd vpwr scs8hd_buf_1
XANTENNA__169__B _168_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_3.LATCH_5_.latch data_in mem_left_ipin_3.LATCH_5_.latch/Q _097_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _162_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_36 vpwr vgnd scs8hd_fill_2
XANTENNA__079__B _079_/B vgnd vpwr scs8hd_diode_2
XFILLER_43_79 vpwr vgnd scs8hd_fill_2
XFILLER_43_46 vgnd vpwr scs8hd_decap_3
XFILLER_43_35 vpwr vgnd scs8hd_fill_2
XANTENNA__095__A _110_/A vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_ipin_2.LATCH_2_.latch/Q mux_left_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_125 vgnd vpwr scs8hd_decap_12
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_90 vgnd vpwr scs8hd_decap_3
XFILLER_57_143 vgnd vpwr scs8hd_decap_3
XFILLER_57_121 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_4.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_68 vpwr vgnd scs8hd_fill_2
XFILLER_38_79 vpwr vgnd scs8hd_fill_2
XFILLER_54_45 vpwr vgnd scs8hd_fill_2
XFILLER_63_135 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_ipin_2.LATCH_4_.latch_SLEEPB _180_/Y vgnd vpwr scs8hd_diode_2
XFILLER_39_143 vgnd vpwr scs8hd_decap_3
XFILLER_39_121 vgnd vpwr scs8hd_fill_1
XFILLER_5_83 vpwr vgnd scs8hd_fill_2
XFILLER_54_102 vpwr vgnd scs8hd_fill_2
XFILLER_40_69 vgnd vpwr scs8hd_decap_8
XFILLER_45_135 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_ipin_2.LATCH_1_.latch_SLEEPB _157_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_91 vgnd vpwr scs8hd_fill_1
XANTENNA__177__B _177_/B vgnd vpwr scs8hd_diode_2
XFILLER_36_102 vpwr vgnd scs8hd_fill_2
XFILLER_36_113 vgnd vpwr scs8hd_decap_12
XANTENNA__193__A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_1_.latch/Q mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_15 vgnd vpwr scs8hd_fill_1
XFILLER_27_135 vgnd vpwr scs8hd_decap_8
XFILLER_35_58 vgnd vpwr scs8hd_decap_3
XFILLER_35_69 vpwr vgnd scs8hd_fill_2
XFILLER_51_57 vgnd vpwr scs8hd_fill_1
X_070_ _069_/X _151_/A vgnd vpwr scs8hd_buf_1
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
XFILLER_18_102 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_91 vgnd vpwr scs8hd_decap_3
XPHY_80 vgnd vpwr scs8hd_decap_3
X_199_ chany_top_in[1] chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA__163__D _095_/D vgnd vpwr scs8hd_diode_2
XFILLER_2_84 vgnd vpwr scs8hd_decap_4
XFILLER_2_73 vpwr vgnd scs8hd_fill_2
XFILLER_37_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__098__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_62_56 vgnd vpwr scs8hd_decap_12
X_122_ _121_/X _124_/B vgnd vpwr scs8hd_buf_1
XFILLER_23_9 vgnd vpwr scs8hd_fill_1
Xmem_left_ipin_4.LATCH_1_.latch data_in mem_left_ipin_4.LATCH_1_.latch/Q _117_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_21_108 vgnd vpwr scs8hd_decap_4
Xmux_left_ipin_3.INVTX1_1_.scs8hd_inv_1 chany_top_in[2] mux_left_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_16_27 vpwr vgnd scs8hd_fill_2
XFILLER_20_130 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_ipin_0.LATCH_5_.latch_SLEEPB _165_/Y vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_6.LATCH_4_.latch data_in mem_left_ipin_6.LATCH_4_.latch/Q _132_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_123 vgnd vpwr scs8hd_decap_12
X_105_ _135_/A _101_/B _105_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_right_ipin_0.LATCH_2_.latch_SLEEPB _152_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_83 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_4.INVTX1_5_.scs8hd_inv_1 chany_top_in[8] mux_left_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_15 vgnd vpwr scs8hd_fill_1
XANTENNA__095__B _095_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_137 vgnd vpwr scs8hd_decap_8
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_81 vgnd vpwr scs8hd_fill_1
Xmux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ _162_/A mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_ipin_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__196__A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_118 vgnd vpwr scs8hd_decap_4
XFILLER_57_111 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _190_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_48_144 vpwr vgnd scs8hd_fill_2
XFILLER_28_91 vgnd vpwr scs8hd_fill_1
XFILLER_54_125 vgnd vpwr scs8hd_decap_12
XFILLER_40_15 vgnd vpwr scs8hd_decap_4
XFILLER_49_57 vpwr vgnd scs8hd_fill_2
XFILLER_14_60 vpwr vgnd scs8hd_fill_2
XFILLER_36_125 vgnd vpwr scs8hd_decap_12
XFILLER_35_15 vgnd vpwr scs8hd_decap_8
XFILLER_51_36 vpwr vgnd scs8hd_fill_2
XFILLER_51_69 vgnd vpwr scs8hd_decap_3
Xmem_right_ipin_0.LATCH_1_.latch data_in mem_right_ipin_0.LATCH_1_.latch/Q _153_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_18_114 vgnd vpwr scs8hd_decap_12
XPHY_92 vgnd vpwr scs8hd_decap_3
XPHY_81 vgnd vpwr scs8hd_decap_3
XFILLER_25_81 vgnd vpwr scs8hd_decap_4
XPHY_70 vgnd vpwr scs8hd_decap_3
X_198_ chany_top_in[2] chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_left_ipin_7.LATCH_4_.latch_SLEEPB _140_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_ipin_1.LATCH_2_.latch/Q mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_106 vgnd vpwr scs8hd_decap_4
Xmem_left_ipin_7.LATCH_0_.latch data_in mem_left_ipin_7.LATCH_0_.latch/Q _144_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_47 vgnd vpwr scs8hd_decap_8
XANTENNA__098__B _098_/B vgnd vpwr scs8hd_diode_2
XFILLER_62_68 vgnd vpwr scs8hd_decap_12
X_121_ _110_/D _120_/X _121_/X vgnd vpwr scs8hd_or2_4
XFILLER_11_94 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_2.INVTX1_3_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_36_91 vgnd vpwr scs8hd_fill_1
XANTENNA__199__A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_7.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_6.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_20_142 vgnd vpwr scs8hd_decap_4
XFILLER_32_27 vpwr vgnd scs8hd_fill_2
XFILLER_57_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_7_135 vgnd vpwr scs8hd_decap_8
XFILLER_11_120 vpwr vgnd scs8hd_fill_2
X_104_ _104_/A _135_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mem_left_ipin_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_43_15 vgnd vpwr scs8hd_decap_4
XANTENNA__095__C _095_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[0] mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_60 vgnd vpwr scs8hd_fill_1
XFILLER_12_3 vgnd vpwr scs8hd_decap_12
XFILLER_57_123 vgnd vpwr scs8hd_decap_12
XFILLER_38_15 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_ipin_5.LATCH_5_.latch_SLEEPB _123_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_2.INVTX1_5_.scs8hd_inv_1 chany_top_in[6] mux_left_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_28_81 vpwr vgnd scs8hd_fill_2
XFILLER_5_52 vpwr vgnd scs8hd_fill_2
XFILLER_39_123 vgnd vpwr scs8hd_decap_12
XFILLER_54_137 vgnd vpwr scs8hd_decap_8
XFILLER_40_27 vgnd vpwr scs8hd_decap_4
XFILLER_40_38 vgnd vpwr scs8hd_fill_1
XFILLER_49_36 vpwr vgnd scs8hd_fill_2
XFILLER_49_25 vpwr vgnd scs8hd_fill_2
XFILLER_45_104 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_6.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_30_93 vgnd vpwr scs8hd_decap_12
XFILLER_36_137 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_ipin_7.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_27_104 vpwr vgnd scs8hd_fill_2
XFILLER_27_115 vgnd vpwr scs8hd_decap_6
XFILLER_35_38 vgnd vpwr scs8hd_decap_4
XFILLER_51_15 vgnd vpwr scs8hd_decap_12
XPHY_82 vgnd vpwr scs8hd_decap_3
XFILLER_18_126 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_33_107 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_93 vgnd vpwr scs8hd_decap_3
X_197_ chany_top_in[3] chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_4.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_21_18 vpwr vgnd scs8hd_fill_2
XANTENNA__098__C address[0] vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ _160_/A mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
X_120_ _119_/X _120_/X vgnd vpwr scs8hd_buf_1
XANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_4.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_40 vpwr vgnd scs8hd_fill_2
XFILLER_11_73 vpwr vgnd scs8hd_fill_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XFILLER_57_36 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_6.tap_buf4_0_.scs8hd_inv_1 mux_left_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ right_grid_pin_12_ vgnd vpwr scs8hd_inv_1
XFILLER_7_103 vgnd vpwr scs8hd_decap_12
XFILLER_11_143 vgnd vpwr scs8hd_decap_3
XFILLER_22_72 vpwr vgnd scs8hd_fill_2
X_103_ _142_/A _101_/B _103_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_47_91 vpwr vgnd scs8hd_fill_2
XFILLER_14_7 vgnd vpwr scs8hd_decap_6
XFILLER_8_41 vgnd vpwr scs8hd_decap_3
Xmem_left_ipin_0.LATCH_1_.latch data_in mem_left_ipin_0.LATCH_1_.latch/Q _169_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__095__D _095_/D vgnd vpwr scs8hd_diode_2
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_71 vpwr vgnd scs8hd_fill_2
Xmem_left_ipin_2.LATCH_4_.latch data_in mem_left_ipin_2.LATCH_4_.latch/Q _180_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_27 vgnd vpwr scs8hd_decap_4
XFILLER_57_135 vgnd vpwr scs8hd_decap_8
XFILLER_54_15 vgnd vpwr scs8hd_fill_1
XFILLER_38_49 vpwr vgnd scs8hd_fill_2
XFILLER_48_124 vgnd vpwr scs8hd_decap_12
XFILLER_48_113 vgnd vpwr scs8hd_decap_8
XFILLER_48_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _191_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _191_/HI _161_/Y mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_2_.latch/Q mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_97 vpwr vgnd scs8hd_fill_2
XFILLER_39_135 vgnd vpwr scs8hd_decap_8
XFILLER_39_113 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_6.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_84 vgnd vpwr scs8hd_decap_8
XFILLER_30_61 vgnd vpwr scs8hd_fill_1
XFILLER_30_83 vgnd vpwr scs8hd_decap_8
XFILLER_39_92 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_0.INVTX1_5_.scs8hd_inv_1 chany_top_in[8] mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__101__A _133_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_18 vpwr vgnd scs8hd_fill_2
XFILLER_42_108 vgnd vpwr scs8hd_decap_4
XFILLER_51_27 vgnd vpwr scs8hd_decap_6
Xmux_left_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_ipin_7.LATCH_0_.latch/Q mux_left_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_138 vgnd vpwr scs8hd_decap_8
XPHY_94 vgnd vpwr scs8hd_decap_3
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_50 vgnd vpwr scs8hd_decap_3
XFILLER_25_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XFILLER_41_71 vpwr vgnd scs8hd_fill_2
X_196_ chany_top_in[4] chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_32 vgnd vpwr scs8hd_decap_3
XFILLER_2_54 vpwr vgnd scs8hd_fill_2
XFILLER_24_119 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_6.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[5] mux_left_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_ipin_4.LATCH_0_.latch_SLEEPB _118_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _161_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_15 vgnd vpwr scs8hd_decap_12
XFILLER_15_119 vgnd vpwr scs8hd_decap_3
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
X_179_ _079_/B _179_/B _179_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
XFILLER_57_15 vgnd vpwr scs8hd_decap_6
Xmem_left_ipin_3.LATCH_0_.latch data_in mem_left_ipin_3.LATCH_0_.latch/Q _107_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_115 vgnd vpwr scs8hd_decap_6
XFILLER_22_40 vgnd vpwr scs8hd_decap_4
XFILLER_22_84 vpwr vgnd scs8hd_fill_2
X_102_ _102_/A _142_/A vgnd vpwr scs8hd_buf_1
XFILLER_8_64 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_43_39 vpwr vgnd scs8hd_fill_2
Xmem_left_ipin_5.LATCH_3_.latch data_in mem_left_ipin_5.LATCH_3_.latch/Q _125_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_62 vpwr vgnd scs8hd_fill_2
XFILLER_17_73 vpwr vgnd scs8hd_fill_2
XFILLER_17_95 vpwr vgnd scs8hd_fill_2
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__104__A _104_/A vgnd vpwr scs8hd_diode_2
XFILLER_58_91 vgnd vpwr scs8hd_fill_1
XFILLER_54_49 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_2.LATCH_1_.latch_SLEEPB _085_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1_A mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_136 vgnd vpwr scs8hd_decap_8
XFILLER_28_61 vgnd vpwr scs8hd_decap_4
XFILLER_44_82 vpwr vgnd scs8hd_fill_2
XFILLER_5_87 vgnd vpwr scs8hd_decap_4
XFILLER_54_106 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_0_.latch/Q mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_60_109 vgnd vpwr scs8hd_decap_12
XFILLER_14_96 vgnd vpwr scs8hd_decap_8
XFILLER_30_51 vpwr vgnd scs8hd_fill_2
XFILLER_39_71 vpwr vgnd scs8hd_fill_2
XFILLER_36_106 vgnd vpwr scs8hd_decap_4
XANTENNA__101__B _101_/B vgnd vpwr scs8hd_diode_2
XFILLER_35_29 vpwr vgnd scs8hd_fill_2
XANTENNA__202__A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XPHY_95 vgnd vpwr scs8hd_decap_3
XPHY_84 vgnd vpwr scs8hd_decap_3
XFILLER_41_120 vpwr vgnd scs8hd_fill_2
XPHY_40 vgnd vpwr scs8hd_decap_3
XFILLER_25_62 vgnd vpwr scs8hd_fill_1
XPHY_51 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
X_195_ chany_top_in[5] chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_2_77 vgnd vpwr scs8hd_decap_4
XANTENNA__112__A _139_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_88 vgnd vpwr scs8hd_fill_1
XFILLER_32_131 vgnd vpwr scs8hd_decap_12
XFILLER_62_27 vgnd vpwr scs8hd_decap_4
XFILLER_11_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_3.INVTX1_5_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_14_120 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_ipin_0.LATCH_2_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
XFILLER_52_71 vgnd vpwr scs8hd_decap_4
XANTENNA__107__A _144_/A vgnd vpwr scs8hd_diode_2
X_178_ _088_/B _177_/B _178_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_right_ipin_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_3 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_ipin_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_4.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[4] mux_left_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _190_/HI _159_/Y mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_112 vgnd vpwr scs8hd_decap_8
XFILLER_11_123 vgnd vpwr scs8hd_decap_12
X_101_ _133_/A _101_/B _101_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_8_87 vgnd vpwr scs8hd_decap_3
XFILLER_27_19 vpwr vgnd scs8hd_fill_2
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_52 vpwr vgnd scs8hd_fill_2
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_40 vpwr vgnd scs8hd_fill_2
XFILLER_33_95 vgnd vpwr scs8hd_decap_3
XANTENNA__120__A _119_/X vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_ipin_6.LATCH_0_.latch/Q mux_left_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_57_115 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_54_28 vgnd vpwr scs8hd_decap_3
XANTENNA__205__A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_0_133 vgnd vpwr scs8hd_decap_12
XFILLER_60_60 vgnd vpwr scs8hd_fill_1
XFILLER_5_22 vpwr vgnd scs8hd_fill_2
XANTENNA__115__A _133_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_66 vpwr vgnd scs8hd_fill_2
XFILLER_10_3 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_left_ipin_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_19 vgnd vpwr scs8hd_fill_1
XFILLER_14_64 vpwr vgnd scs8hd_fill_2
XFILLER_14_75 vpwr vgnd scs8hd_fill_2
XFILLER_55_93 vpwr vgnd scs8hd_fill_2
XFILLER_58_3 vgnd vpwr scs8hd_decap_12
XFILLER_50_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_4.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_7.LATCH_1_.latch_SLEEPB _143_/Y vgnd vpwr scs8hd_diode_2
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_143 vgnd vpwr scs8hd_decap_3
XFILLER_41_40 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_1.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_25_41 vpwr vgnd scs8hd_fill_2
XFILLER_25_52 vgnd vpwr scs8hd_decap_3
XFILLER_25_96 vpwr vgnd scs8hd_fill_2
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_74 vgnd vpwr scs8hd_decap_3
XFILLER_41_95 vpwr vgnd scs8hd_fill_2
X_194_ chany_top_in[6] chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_2_23 vgnd vpwr scs8hd_decap_8
XANTENNA__112__B _118_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_ipin_5.INVTX1_3_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_23_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_ipin_3.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_11_21 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_7.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_4.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_132 vgnd vpwr scs8hd_decap_12
XFILLER_36_84 vgnd vpwr scs8hd_decap_4
XFILLER_52_50 vgnd vpwr scs8hd_decap_8
X_177_ _104_/A _177_/B _177_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__107__B _101_/B vgnd vpwr scs8hd_diode_2
XANTENNA__123__A _139_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_5.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_102 vpwr vgnd scs8hd_fill_2
XANTENNA__208__A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_11_135 vgnd vpwr scs8hd_decap_8
XFILLER_22_53 vpwr vgnd scs8hd_fill_2
X_100_ _101_/B _100_/B _100_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_8_11 vgnd vpwr scs8hd_decap_3
XANTENNA__118__A _144_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_77 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XFILLER_43_19 vgnd vpwr scs8hd_fill_1
XFILLER_17_31 vpwr vgnd scs8hd_fill_2
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_120 vpwr vgnd scs8hd_fill_2
XFILLER_58_71 vgnd vpwr scs8hd_decap_8
Xmux_left_ipin_2.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[2] mux_left_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_ipin_5.LATCH_2_.latch_SLEEPB _126_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_6.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_123 vgnd vpwr scs8hd_fill_1
XFILLER_0_145 vgnd vpwr scs8hd_fill_1
XFILLER_28_41 vgnd vpwr scs8hd_decap_3
XFILLER_28_85 vgnd vpwr scs8hd_decap_6
Xmem_left_ipin_1.LATCH_3_.latch data_in mem_left_ipin_1.LATCH_3_.latch/Q _175_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_60_72 vpwr vgnd scs8hd_fill_2
XFILLER_5_56 vpwr vgnd scs8hd_fill_2
XANTENNA__115__B _118_/B vgnd vpwr scs8hd_diode_2
XANTENNA__131__A _139_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_105 vpwr vgnd scs8hd_fill_2
XFILLER_62_141 vgnd vpwr scs8hd_decap_4
XFILLER_54_119 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_6.tap_buf4_0_.scs8hd_inv_1_A mux_left_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_49_29 vpwr vgnd scs8hd_fill_2
XFILLER_45_108 vgnd vpwr scs8hd_decap_12
XFILLER_14_32 vpwr vgnd scs8hd_fill_2
XFILLER_14_43 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_64 vpwr vgnd scs8hd_fill_2
XFILLER_55_50 vgnd vpwr scs8hd_fill_1
XANTENNA__126__A _142_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_3.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_right_ipin_0.LATCH_4_.latch/Q mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_7.INVTX1_1_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XPHY_64 vgnd vpwr scs8hd_decap_3
X_193_ chany_top_in[7] chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
XPHY_97 vgnd vpwr scs8hd_decap_3
XPHY_86 vgnd vpwr scs8hd_decap_3
XPHY_75 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_4.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_100 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_3.LATCH_3_.latch_SLEEPB _101_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_77 vpwr vgnd scs8hd_fill_2
XFILLER_14_144 vpwr vgnd scs8hd_fill_2
XFILLER_52_84 vpwr vgnd scs8hd_fill_2
X_176_ _102_/A _177_/B _176_/Y vgnd vpwr scs8hd_nor2_4
Xmux_left_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_ipin_5.LATCH_0_.latch/Q mux_left_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__123__B _124_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_32 vgnd vpwr scs8hd_fill_1
XFILLER_22_76 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_3 vgnd vpwr scs8hd_decap_4
XFILLER_47_73 vgnd vpwr scs8hd_fill_1
XFILLER_8_23 vpwr vgnd scs8hd_fill_2
XANTENNA__118__B _118_/B vgnd vpwr scs8hd_diode_2
XANTENNA__134__A _142_/A vgnd vpwr scs8hd_diode_2
X_159_ _159_/A _159_/Y vgnd vpwr scs8hd_inv_8
XFILLER_33_3 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_0.INVTX1_3_.scs8hd_inv_1 chany_top_in[7] mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_10 vpwr vgnd scs8hd_fill_2
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_53 vpwr vgnd scs8hd_fill_2
XFILLER_33_75 vpwr vgnd scs8hd_fill_2
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_143 vgnd vpwr scs8hd_decap_3
XFILLER_58_83 vpwr vgnd scs8hd_fill_2
XANTENNA__129__A _077_/B vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_4.LATCH_2_.latch data_in mem_left_ipin_4.LATCH_2_.latch/Q _116_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_1.LATCH_4_.latch_SLEEPB _174_/Y vgnd vpwr scs8hd_diode_2
XFILLER_48_106 vgnd vpwr scs8hd_decap_4
XFILLER_44_41 vpwr vgnd scs8hd_fill_2
XFILLER_60_84 vpwr vgnd scs8hd_fill_2
XANTENNA__131__B _131_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_6.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_35 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_1.LATCH_1_.latch_SLEEPB _155_/Y vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_6.LATCH_5_.latch data_in mem_left_ipin_6.LATCH_5_.latch/Q _131_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_2_.latch/Q mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_ipin_0.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[4] mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_49_19 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_10 vgnd vpwr scs8hd_decap_4
XFILLER_30_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_62 vgnd vpwr scs8hd_decap_3
XANTENNA__126__B _124_/B vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _142_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_120 vpwr vgnd scs8hd_fill_2
XFILLER_50_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_98 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_decap_3
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XFILLER_41_112 vpwr vgnd scs8hd_fill_2
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_26_131 vgnd vpwr scs8hd_decap_12
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_76 vgnd vpwr scs8hd_decap_3
XFILLER_41_75 vpwr vgnd scs8hd_fill_2
XFILLER_41_53 vpwr vgnd scs8hd_fill_2
X_192_ chany_top_in[8] chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_2_58 vpwr vgnd scs8hd_fill_2
XFILLER_17_131 vgnd vpwr scs8hd_decap_3
XANTENNA__137__A _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_63_3 vgnd vpwr scs8hd_decap_12
XFILLER_23_112 vpwr vgnd scs8hd_fill_2
XFILLER_23_123 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_7.INVTX1_3_.scs8hd_inv_1 chany_top_in[6] mux_left_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_175_ _151_/A _177_/B _175_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_3_90 vpwr vgnd scs8hd_fill_2
XFILLER_22_88 vpwr vgnd scs8hd_fill_2
XFILLER_63_51 vgnd vpwr scs8hd_decap_8
XFILLER_47_52 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ _162_/Y mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_63_62 vgnd vpwr scs8hd_decap_12
XFILLER_8_46 vgnd vpwr scs8hd_decap_3
Xmem_right_ipin_0.LATCH_2_.latch data_in mem_right_ipin_0.LATCH_2_.latch/Q _152_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__134__B _131_/B vgnd vpwr scs8hd_diode_2
X_089_ address[2] _098_/B vgnd vpwr scs8hd_inv_8
X_158_ _077_/B _147_/D address[0] _158_/Y vgnd vpwr scs8hd_nor3_4
XANTENNA__150__A _132_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _160_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_44 vpwr vgnd scs8hd_fill_2
XFILLER_17_77 vgnd vpwr scs8hd_decap_4
XFILLER_17_99 vpwr vgnd scs8hd_fill_2
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_left_ipin_7.LATCH_1_.latch data_in mem_left_ipin_7.LATCH_1_.latch/Q _143_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_58_51 vgnd vpwr scs8hd_decap_6
XANTENNA__129__B _110_/D vgnd vpwr scs8hd_diode_2
XANTENNA__145__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_0_103 vgnd vpwr scs8hd_decap_8
XFILLER_44_86 vgnd vpwr scs8hd_decap_6
XFILLER_60_52 vgnd vpwr scs8hd_decap_8
XFILLER_53_143 vgnd vpwr scs8hd_decap_3
XFILLER_14_23 vgnd vpwr scs8hd_decap_6
Xmux_left_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_ipin_4.LATCH_0_.latch/Q mux_left_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_55 vgnd vpwr scs8hd_decap_6
XFILLER_39_75 vpwr vgnd scs8hd_fill_2
XFILLER_39_53 vpwr vgnd scs8hd_fill_2
XFILLER_55_74 vpwr vgnd scs8hd_fill_2
XANTENNA__142__B _139_/B vgnd vpwr scs8hd_diode_2
XFILLER_50_102 vgnd vpwr scs8hd_decap_12
XFILLER_35_143 vgnd vpwr scs8hd_decap_3
XFILLER_50_135 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_ipin_6.LATCH_4_.latch_SLEEPB _132_/Y vgnd vpwr scs8hd_diode_2
XPHY_99 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_decap_3
XFILLER_41_135 vgnd vpwr scs8hd_decap_8
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XFILLER_25_22 vpwr vgnd scs8hd_fill_2
XFILLER_25_77 vpwr vgnd scs8hd_fill_2
XFILLER_26_143 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_77 vgnd vpwr scs8hd_decap_3
XFILLER_41_21 vgnd vpwr scs8hd_fill_1
X_191_ _191_/HI _191_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_ipin_2.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_2_37 vpwr vgnd scs8hd_fill_2
XFILLER_2_15 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__137__B _095_/B vgnd vpwr scs8hd_diode_2
XFILLER_56_3 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_ipin_6.INVTX1_5_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__153__A _135_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_135 vgnd vpwr scs8hd_decap_8
XFILLER_11_57 vpwr vgnd scs8hd_fill_2
XFILLER_36_32 vpwr vgnd scs8hd_fill_2
XFILLER_36_65 vpwr vgnd scs8hd_fill_2
X_174_ _100_/B _177_/B _174_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__148__A _148_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _181_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_23 vgnd vpwr scs8hd_decap_4
XFILLER_63_74 vgnd vpwr scs8hd_decap_12
XFILLER_8_58 vgnd vpwr scs8hd_decap_4
XFILLER_6_120 vgnd vpwr scs8hd_decap_12
X_157_ _077_/B _147_/D _069_/C _157_/Y vgnd vpwr scs8hd_nor3_4
Xmux_left_ipin_5.INVTX1_3_.scs8hd_inv_1 chany_top_in[4] mux_left_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__150__B _149_/B vgnd vpwr scs8hd_diode_2
X_088_ _079_/B _088_/B _088_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_left_ipin_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_56 vpwr vgnd scs8hd_fill_2
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_123 vgnd vpwr scs8hd_decap_12
XFILLER_3_112 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_ipin_4.LATCH_5_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__145__B _145_/B vgnd vpwr scs8hd_diode_2
XANTENNA__161__A _161_/A vgnd vpwr scs8hd_diode_2
X_209_ chany_bottom_in[0] chany_top_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_4.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__071__A _151_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_115 vpwr vgnd scs8hd_fill_2
XFILLER_28_11 vgnd vpwr scs8hd_decap_3
XFILLER_60_97 vgnd vpwr scs8hd_decap_12
XFILLER_60_42 vgnd vpwr scs8hd_fill_1
XANTENNA__156__A _120_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_13 vgnd vpwr scs8hd_fill_1
XFILLER_14_79 vgnd vpwr scs8hd_decap_3
Xmem_left_ipin_0.LATCH_2_.latch data_in mem_left_ipin_0.LATCH_2_.latch/Q _168_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_30_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_55_53 vpwr vgnd scs8hd_fill_2
XFILLER_55_31 vpwr vgnd scs8hd_fill_2
XFILLER_55_20 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_4.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_55_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_5.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_50_114 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_ipin_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_4.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XPHY_12 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ _160_/Y mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
Xmem_left_ipin_2.LATCH_5_.latch data_in mem_left_ipin_2.LATCH_5_.latch/Q _179_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_100 vgnd vpwr scs8hd_decap_4
Xmux_left_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_left_ipin_7.LATCH_3_.latch/Q mux_left_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XPHY_89 vgnd vpwr scs8hd_decap_3
X_190_ _190_/HI _190_/LO vgnd vpwr scs8hd_conb_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_78 vgnd vpwr scs8hd_decap_3
XFILLER_41_99 vpwr vgnd scs8hd_fill_2
XFILLER_17_144 vpwr vgnd scs8hd_fill_2
XANTENNA__153__B _149_/B vgnd vpwr scs8hd_diode_2
XANTENNA__137__C _095_/C vgnd vpwr scs8hd_diode_2
XFILLER_49_3 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_2.tap_buf4_0_.scs8hd_inv_1 mux_left_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ right_grid_pin_4_ vgnd vpwr scs8hd_inv_1
Xmux_right_ipin_2.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[1] mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_25 vpwr vgnd scs8hd_fill_2
XFILLER_11_36 vpwr vgnd scs8hd_fill_2
XFILLER_36_55 vgnd vpwr scs8hd_fill_1
XFILLER_36_88 vgnd vpwr scs8hd_fill_1
XFILLER_52_32 vgnd vpwr scs8hd_decap_3
X_173_ _179_/B _177_/B _173_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_6.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_106 vgnd vpwr scs8hd_decap_12
XANTENNA__164__A _164_/A vgnd vpwr scs8hd_diode_2
XANTENNA__074__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_22_57 vgnd vpwr scs8hd_decap_4
XFILLER_47_87 vpwr vgnd scs8hd_fill_2
XFILLER_47_65 vpwr vgnd scs8hd_fill_2
XFILLER_63_86 vgnd vpwr scs8hd_decap_12
XFILLER_6_132 vgnd vpwr scs8hd_decap_12
X_156_ _120_/X _147_/D address[0] _156_/Y vgnd vpwr scs8hd_nor3_4
X_087_ _086_/X _088_/B vgnd vpwr scs8hd_buf_1
XANTENNA__159__A _159_/A vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_ipin_3.LATCH_0_.latch/Q mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__069__A _069_/A vgnd vpwr scs8hd_diode_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_23 vpwr vgnd scs8hd_fill_2
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_135 vgnd vpwr scs8hd_decap_8
X_139_ _139_/A _139_/B _139_/Y vgnd vpwr scs8hd_nor2_4
X_208_ chany_bottom_in[1] chany_top_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_31_3 vgnd vpwr scs8hd_decap_3
Xmux_left_ipin_3.INVTX1_3_.scs8hd_inv_1 chany_top_in[3] mux_left_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_56_131 vgnd vpwr scs8hd_decap_12
XFILLER_56_120 vgnd vpwr scs8hd_decap_8
XFILLER_28_23 vgnd vpwr scs8hd_decap_8
XFILLER_28_67 vgnd vpwr scs8hd_decap_3
XFILLER_44_66 vgnd vpwr scs8hd_fill_1
XFILLER_44_11 vgnd vpwr scs8hd_decap_3
XFILLER_60_76 vgnd vpwr scs8hd_decap_4
XFILLER_47_120 vpwr vgnd scs8hd_fill_2
XFILLER_39_109 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_145 vgnd vpwr scs8hd_fill_1
Xmem_left_ipin_3.LATCH_1_.latch data_in mem_left_ipin_3.LATCH_1_.latch/Q _105_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_ipin_0.LATCH_4_.latch_SLEEPB _150_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__156__B _147_/D vgnd vpwr scs8hd_diode_2
XANTENNA__172__A _172_/A vgnd vpwr scs8hd_diode_2
XFILLER_53_123 vgnd vpwr scs8hd_decap_12
XFILLER_53_112 vpwr vgnd scs8hd_fill_2
XFILLER_38_131 vgnd vpwr scs8hd_decap_12
XFILLER_14_47 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_ipin_7.LATCH_1_.latch/Q mux_left_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__082__A _079_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_79 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_6.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_39_88 vpwr vgnd scs8hd_fill_2
XFILLER_29_120 vpwr vgnd scs8hd_fill_2
XFILLER_39_11 vgnd vpwr scs8hd_fill_1
XFILLER_39_22 vgnd vpwr scs8hd_decap_3
XFILLER_44_145 vgnd vpwr scs8hd_fill_1
Xmem_left_ipin_5.LATCH_4_.latch data_in mem_left_ipin_5.LATCH_4_.latch/Q _124_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_35_112 vgnd vpwr scs8hd_decap_8
XANTENNA__167__A _151_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_123 vgnd vpwr scs8hd_decap_12
XFILLER_6_81 vpwr vgnd scs8hd_fill_2
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XANTENNA__077__A _095_/D vgnd vpwr scs8hd_diode_2
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_79 vgnd vpwr scs8hd_decap_3
XFILLER_25_57 vpwr vgnd scs8hd_fill_2
XPHY_57 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_ipin_3.LATCH_0_.latch_SLEEPB _107_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_123 vgnd vpwr scs8hd_decap_8
XANTENNA__137__D _110_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_15 vgnd vpwr scs8hd_fill_1
XFILLER_14_104 vgnd vpwr scs8hd_fill_1
XFILLER_36_45 vpwr vgnd scs8hd_fill_2
XFILLER_52_88 vpwr vgnd scs8hd_fill_2
X_172_ _172_/A _177_/B vgnd vpwr scs8hd_buf_1
XFILLER_20_118 vgnd vpwr scs8hd_decap_12
XFILLER_61_3 vgnd vpwr scs8hd_decap_12
XANTENNA__180__A _079_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _182_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_107 vgnd vpwr scs8hd_decap_3
XFILLER_22_36 vpwr vgnd scs8hd_fill_2
XANTENNA__090__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_47_44 vpwr vgnd scs8hd_fill_2
XFILLER_63_98 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_0.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[3] mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_27 vpwr vgnd scs8hd_fill_2
X_086_ address[1] address[2] address[0] _086_/X vgnd vpwr scs8hd_or3_4
XFILLER_6_144 vpwr vgnd scs8hd_fill_2
X_155_ _120_/X _147_/D _069_/C _155_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_12_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1_A mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__175__A _151_/A vgnd vpwr scs8hd_diode_2
XANTENNA__069__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_17_14 vpwr vgnd scs8hd_fill_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__085__A _079_/B vgnd vpwr scs8hd_diode_2
XFILLER_33_57 vpwr vgnd scs8hd_fill_2
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_58_87 vpwr vgnd scs8hd_fill_2
XFILLER_58_32 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_left_ipin_1.LATCH_1_.latch_SLEEPB _177_/Y vgnd vpwr scs8hd_diode_2
X_207_ chany_bottom_in[2] chany_top_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_23_90 vgnd vpwr scs8hd_decap_3
X_138_ _137_/X _139_/B vgnd vpwr scs8hd_buf_1
X_069_ _069_/A address[2] _069_/C _069_/X vgnd vpwr scs8hd_or3_4
XFILLER_24_3 vgnd vpwr scs8hd_decap_8
Xmux_left_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_left_ipin_6.LATCH_3_.latch/Q mux_left_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_1_.latch/Q mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_92 vpwr vgnd scs8hd_fill_2
Xmem_left_ipin_6.LATCH_0_.latch data_in mem_left_ipin_6.LATCH_0_.latch/Q _136_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_56_143 vgnd vpwr scs8hd_decap_3
XFILLER_44_23 vpwr vgnd scs8hd_fill_2
XFILLER_28_46 vgnd vpwr scs8hd_decap_6
XFILLER_44_45 vpwr vgnd scs8hd_fill_2
XFILLER_60_88 vgnd vpwr scs8hd_decap_4
XFILLER_5_39 vpwr vgnd scs8hd_fill_2
XANTENNA__156__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_53_135 vgnd vpwr scs8hd_decap_8
XFILLER_53_102 vpwr vgnd scs8hd_fill_2
XFILLER_38_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__082__B _102_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_36 vpwr vgnd scs8hd_fill_2
XFILLER_55_11 vgnd vpwr scs8hd_decap_3
Xmux_left_ipin_1.INVTX1_3_.scs8hd_inv_1 chany_top_in[1] mux_left_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_143 vgnd vpwr scs8hd_decap_3
XFILLER_39_34 vpwr vgnd scs8hd_fill_2
XFILLER_44_113 vgnd vpwr scs8hd_decap_12
XFILLER_44_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_135 vgnd vpwr scs8hd_decap_8
XANTENNA__167__B _168_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_60 vpwr vgnd scs8hd_fill_2
XFILLER_41_116 vpwr vgnd scs8hd_fill_2
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XANTENNA__077__B _077_/B vgnd vpwr scs8hd_diode_2
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XPHY_69 vgnd vpwr scs8hd_decap_3
XFILLER_41_79 vgnd vpwr scs8hd_decap_3
XFILLER_41_57 vpwr vgnd scs8hd_fill_2
XANTENNA__093__A _093_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_18 vpwr vgnd scs8hd_fill_2
XFILLER_15_91 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_ipin_2.LATCH_0_.latch/Q mux_left_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_ipin_7.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[2] mux_left_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_31_90 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _159_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__178__A _088_/B vgnd vpwr scs8hd_diode_2
XFILLER_23_116 vgnd vpwr scs8hd_decap_6
XANTENNA__088__A _079_/B vgnd vpwr scs8hd_diode_2
XFILLER_52_23 vpwr vgnd scs8hd_fill_2
XFILLER_52_67 vpwr vgnd scs8hd_fill_2
X_171_ _095_/D _120_/X _172_/A vgnd vpwr scs8hd_or2_4
XFILLER_54_3 vgnd vpwr scs8hd_decap_12
XANTENNA__180__B _100_/B vgnd vpwr scs8hd_diode_2
XFILLER_3_94 vpwr vgnd scs8hd_fill_2
XFILLER_22_15 vgnd vpwr scs8hd_decap_4
XANTENNA__090__B _098_/B vgnd vpwr scs8hd_diode_2
X_154_ _144_/A _149_/B _154_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_12_70 vgnd vpwr scs8hd_decap_4
X_085_ _079_/B _104_/A _085_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__175__B _177_/B vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_ipin_6.LATCH_1_.latch/Q mux_left_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_right_ipin_2.LATCH_0_.latch data_in _162_/A _158_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__069__C _069_/C vgnd vpwr scs8hd_diode_2
XFILLER_17_48 vpwr vgnd scs8hd_fill_2
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__085__B _104_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_36 vpwr vgnd scs8hd_fill_2
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_206_ chany_bottom_in[3] chany_top_out[3] vgnd vpwr scs8hd_buf_2
X_137_ _110_/A _095_/B _095_/C _110_/D _137_/X vgnd vpwr scs8hd_or4_4
X_068_ address[0] _069_/C vgnd vpwr scs8hd_inv_8
XFILLER_17_3 vpwr vgnd scs8hd_fill_2
XFILLER_0_129 vpwr vgnd scs8hd_fill_2
XANTENNA__096__A _095_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_91 vgnd vpwr scs8hd_fill_1
XFILLER_38_100 vgnd vpwr scs8hd_decap_4
XFILLER_14_16 vpwr vgnd scs8hd_fill_2
XFILLER_39_57 vpwr vgnd scs8hd_fill_2
XFILLER_55_78 vpwr vgnd scs8hd_fill_2
XFILLER_44_125 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_1.INVTX1_3_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_20_81 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_6.LATCH_1_.latch_SLEEPB _135_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_5.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XFILLER_25_15 vgnd vpwr scs8hd_fill_1
XFILLER_25_37 vpwr vgnd scs8hd_fill_2
XFILLER_25_48 vpwr vgnd scs8hd_fill_2
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_41_36 vpwr vgnd scs8hd_fill_2
XFILLER_41_25 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_6.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_136 vgnd vpwr scs8hd_decap_8
Xmem_left_ipin_1.LATCH_4_.latch data_in mem_left_ipin_1.LATCH_4_.latch/Q _174_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__194__A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__178__B _177_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__088__B _088_/B vgnd vpwr scs8hd_diode_2
XFILLER_36_69 vgnd vpwr scs8hd_decap_4
X_170_ _088_/B _168_/B _170_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_left_ipin_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_left_ipin_5.LATCH_3_.latch/Q mux_left_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_9_121 vgnd vpwr scs8hd_fill_1
XFILLER_9_143 vgnd vpwr scs8hd_decap_3
XFILLER_47_3 vgnd vpwr scs8hd_decap_8
XFILLER_3_73 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _183_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_left_ipin_5.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_left_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__090__C _069_/C vgnd vpwr scs8hd_diode_2
XANTENNA__099__A _099_/A vgnd vpwr scs8hd_diode_2
XFILLER_47_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _189_/HI vgnd vpwr
+ scs8hd_diode_2
X_153_ _135_/A _149_/B _153_/Y vgnd vpwr scs8hd_nor2_4
X_084_ _083_/X _104_/A vgnd vpwr scs8hd_buf_1
XFILLER_19_7 vgnd vpwr scs8hd_decap_8
Xmux_left_ipin_6.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[6] mux_left_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_ipin_4.LATCH_2_.latch_SLEEPB _116_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_27 vpwr vgnd scs8hd_fill_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_15 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_4.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_5.tap_buf4_0_.scs8hd_inv_1_A mux_left_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_136_ _144_/A _131_/B _136_/Y vgnd vpwr scs8hd_nor2_4
X_205_ chany_bottom_in[4] chany_top_out[4] vgnd vpwr scs8hd_buf_2
X_067_ address[1] _069_/A vgnd vpwr scs8hd_inv_8
XFILLER_0_52 vpwr vgnd scs8hd_fill_2
XFILLER_0_74 vpwr vgnd scs8hd_fill_2
XFILLER_0_85 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_6.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_7.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_119 vgnd vpwr scs8hd_decap_4
XFILLER_44_69 vpwr vgnd scs8hd_fill_2
XFILLER_44_58 vgnd vpwr scs8hd_decap_8
XFILLER_60_35 vgnd vpwr scs8hd_decap_4
Xmux_left_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_ipin_1.LATCH_0_.latch/Q mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_47_145 vgnd vpwr scs8hd_fill_1
XFILLER_47_123 vpwr vgnd scs8hd_fill_2
XFILLER_47_112 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_81 vpwr vgnd scs8hd_fill_2
X_119_ _110_/A address[4] _095_/C _119_/X vgnd vpwr scs8hd_or3_4
XANTENNA_mux_left_ipin_3.INVTX1_1_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _189_/HI mem_right_ipin_0.LATCH_5_.latch/Q
+ mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__197__A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_30_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_7.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_55_57 vpwr vgnd scs8hd_fill_2
XFILLER_55_46 vgnd vpwr scs8hd_decap_4
XFILLER_44_137 vgnd vpwr scs8hd_decap_8
XFILLER_29_123 vgnd vpwr scs8hd_decap_12
Xmem_left_ipin_2.LATCH_0_.latch data_in mem_left_ipin_2.LATCH_0_.latch/Q _088_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_50_118 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_49 vgnd vpwr scs8hd_decap_3
XFILLER_41_15 vgnd vpwr scs8hd_decap_6
Xmux_left_ipin_5.tap_buf4_0_.scs8hd_inv_1 mux_left_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ right_grid_pin_10_ vgnd vpwr scs8hd_inv_1
XFILLER_9_6 vpwr vgnd scs8hd_fill_2
Xmem_left_ipin_4.LATCH_3_.latch data_in mem_left_ipin_4.LATCH_3_.latch/Q _115_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_left_ipin_2.LATCH_3_.latch_SLEEPB _079_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_107 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_ipin_5.LATCH_1_.latch/Q mux_left_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_49_7 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_2.LATCH_0_.latch_SLEEPB _158_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_107 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_6.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XFILLER_7_3 vgnd vpwr scs8hd_decap_6
Xmux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_9_ vgnd vpwr scs8hd_inv_1
XFILLER_42_91 vgnd vpwr scs8hd_fill_1
XFILLER_47_69 vgnd vpwr scs8hd_decap_4
XFILLER_47_25 vpwr vgnd scs8hd_fill_2
XFILLER_47_14 vpwr vgnd scs8hd_fill_2
X_152_ _142_/A _149_/B _152_/Y vgnd vpwr scs8hd_nor2_4
X_083_ address[1] address[2] _069_/C _083_/X vgnd vpwr scs8hd_or3_4
XFILLER_12_61 vpwr vgnd scs8hd_fill_2
XFILLER_12_83 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_59_121 vgnd vpwr scs8hd_fill_1
XFILLER_59_132 vgnd vpwr scs8hd_decap_12
XFILLER_58_57 vgnd vpwr scs8hd_fill_1
Xmux_left_ipin_3.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[2] mux_left_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_204_ chany_bottom_in[5] chany_top_out[5] vgnd vpwr scs8hd_buf_2
X_135_ _135_/A _131_/B _135_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_left_ipin_0.LATCH_4_.latch_SLEEPB _166_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_5.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_73 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_ipin_7.LATCH_0_.latch/Q mux_left_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_16 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_ipin_0.LATCH_1_.latch_SLEEPB _153_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_4.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[8] mux_left_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_62_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_118_ _144_/A _118_/B _118_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_22_3 vgnd vpwr scs8hd_decap_12
XFILLER_53_116 vgnd vpwr scs8hd_decap_6
Xmem_right_ipin_0.LATCH_3_.latch data_in mem_right_ipin_0.LATCH_3_.latch/Q _151_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_135 vgnd vpwr scs8hd_decap_8
Xmux_left_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_left_ipin_4.LATCH_3_.latch/Q mux_left_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _160_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_45_80 vpwr vgnd scs8hd_fill_2
XFILLER_35_105 vgnd vpwr scs8hd_decap_4
Xmem_left_ipin_7.LATCH_2_.latch data_in mem_left_ipin_7.LATCH_2_.latch/Q _142_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_6_41 vpwr vgnd scs8hd_fill_2
XFILLER_6_96 vgnd vpwr scs8hd_decap_12
XFILLER_6_85 vpwr vgnd scs8hd_fill_2
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_32_119 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_15 vgnd vpwr scs8hd_decap_8
XFILLER_14_108 vgnd vpwr scs8hd_decap_12
XFILLER_36_49 vgnd vpwr scs8hd_decap_6
XFILLER_52_37 vpwr vgnd scs8hd_fill_2
XFILLER_9_123 vgnd vpwr scs8hd_decap_12
XFILLER_42_81 vpwr vgnd scs8hd_fill_2
XFILLER_3_53 vpwr vgnd scs8hd_fill_2
XFILLER_22_29 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_0_.latch/Q mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _184_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_47_48 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_7.LATCH_3_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
X_151_ _151_/A _149_/B _151_/Y vgnd vpwr scs8hd_nor2_4
X_082_ _079_/B _102_/A _082_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_52_3 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[0] mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_107 vgnd vpwr scs8hd_decap_3
XFILLER_59_144 vpwr vgnd scs8hd_fill_2
XFILLER_58_47 vpwr vgnd scs8hd_fill_2
XFILLER_58_25 vgnd vpwr scs8hd_decap_6
X_203_ chany_bottom_in[6] chany_top_out[6] vgnd vpwr scs8hd_buf_2
X_134_ _142_/A _131_/B _134_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_0_32 vgnd vpwr scs8hd_decap_4
XFILLER_9_96 vpwr vgnd scs8hd_fill_2
XFILLER_56_103 vgnd vpwr scs8hd_decap_6
XFILLER_44_16 vgnd vpwr scs8hd_decap_4
XFILLER_60_15 vgnd vpwr scs8hd_decap_12
XFILLER_44_27 vgnd vpwr scs8hd_decap_4
Xmux_left_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_ipin_4.LATCH_1_.latch/Q mux_left_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_62_117 vgnd vpwr scs8hd_decap_12
X_117_ _135_/A _118_/B _117_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_34_71 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_1.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_59_90 vgnd vpwr scs8hd_decap_3
XFILLER_53_106 vgnd vpwr scs8hd_decap_4
XFILLER_15_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_38 vpwr vgnd scs8hd_fill_2
XFILLER_44_106 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_2.INVTX1_5_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_20_62 vpwr vgnd scs8hd_fill_2
XFILLER_29_93 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_ipin_5.LATCH_4_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_2.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[6] mux_left_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_64 vgnd vpwr scs8hd_fill_1
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_25_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_17_106 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_62 vgnd vpwr scs8hd_fill_1
XFILLER_15_95 vpwr vgnd scs8hd_fill_2
XFILLER_31_94 vpwr vgnd scs8hd_fill_2
XANTENNA__102__A _102_/A vgnd vpwr scs8hd_diode_2
XFILLER_52_27 vgnd vpwr scs8hd_decap_4
XFILLER_42_60 vpwr vgnd scs8hd_fill_2
XFILLER_9_113 vgnd vpwr scs8hd_decap_8
XFILLER_9_135 vgnd vpwr scs8hd_decap_8
XFILLER_13_120 vpwr vgnd scs8hd_fill_2
Xmem_left_ipin_0.LATCH_3_.latch data_in mem_left_ipin_0.LATCH_3_.latch/Q _167_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_72 vgnd vpwr scs8hd_decap_3
Xmux_left_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_ipin_6.LATCH_0_.latch/Q mux_left_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_32 vpwr vgnd scs8hd_fill_2
XFILLER_22_19 vgnd vpwr scs8hd_fill_1
XFILLER_63_15 vgnd vpwr scs8hd_decap_12
XFILLER_63_59 vpwr vgnd scs8hd_fill_2
X_150_ _132_/A _149_/B _150_/Y vgnd vpwr scs8hd_nor2_4
X_081_ _080_/X _102_/A vgnd vpwr scs8hd_buf_1
XFILLER_10_145 vgnd vpwr scs8hd_fill_1
XFILLER_45_3 vgnd vpwr scs8hd_decap_6
Xmux_left_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_ipin_3.LATCH_3_.latch/Q mux_left_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mem_left_ipin_3.LATCH_5_.latch_SLEEPB _097_/Y vgnd vpwr scs8hd_diode_2
XFILLER_59_123 vgnd vpwr scs8hd_fill_1
XFILLER_59_101 vgnd vpwr scs8hd_decap_12
XFILLER_58_15 vgnd vpwr scs8hd_decap_8
XANTENNA__200__A chany_top_in[0] vgnd vpwr scs8hd_diode_2
X_202_ chany_bottom_in[7] chany_top_out[7] vgnd vpwr scs8hd_buf_2
X_133_ _133_/A _131_/B _133_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_95 vgnd vpwr scs8hd_decap_3
XFILLER_2_130 vgnd vpwr scs8hd_decap_12
XFILLER_48_70 vpwr vgnd scs8hd_fill_2
XFILLER_0_22 vgnd vpwr scs8hd_fill_1
XANTENNA__110__A _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_53 vpwr vgnd scs8hd_fill_2
XFILLER_60_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_6.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_62_129 vgnd vpwr scs8hd_decap_12
XFILLER_34_50 vgnd vpwr scs8hd_decap_6
XFILLER_50_60 vpwr vgnd scs8hd_fill_2
X_116_ _142_/A _118_/B _116_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__105__A _135_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_4.INVTX1_3_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_55_16 vpwr vgnd scs8hd_fill_2
XFILLER_29_104 vpwr vgnd scs8hd_fill_2
XFILLER_39_17 vgnd vpwr scs8hd_decap_3
Xmux_left_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_ipin_7.LATCH_4_.latch/Q mux_left_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_right_ipin_0.INVTX1_5_.scs8hd_inv_1 chany_top_in[8] mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_ipin_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_85 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_ipin_3.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_45_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_76 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_ipin_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_26_107 vgnd vpwr scs8hd_decap_12
XFILLER_41_29 vpwr vgnd scs8hd_fill_2
XFILLER_17_118 vgnd vpwr scs8hd_decap_4
XFILLER_15_52 vgnd vpwr scs8hd_decap_3
XFILLER_15_74 vgnd vpwr scs8hd_decap_6
XFILLER_31_73 vpwr vgnd scs8hd_fill_2
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_143 vgnd vpwr scs8hd_decap_3
Xmux_left_ipin_0.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[8] mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_36_29 vpwr vgnd scs8hd_fill_2
Xmem_left_ipin_3.LATCH_2_.latch data_in mem_left_ipin_3.LATCH_2_.latch/Q _103_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__203__A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_26_40 vgnd vpwr scs8hd_decap_4
XFILLER_26_84 vpwr vgnd scs8hd_fill_2
XFILLER_13_143 vgnd vpwr scs8hd_decap_3
XANTENNA__113__A _100_/B vgnd vpwr scs8hd_diode_2
XFILLER_3_77 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_ipin_3.LATCH_1_.latch/Q mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_left_ipin_5.LATCH_5_.latch data_in mem_left_ipin_5.LATCH_5_.latch/Q _123_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _185_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_63_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_ipin_7.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_080_ _069_/A address[2] address[0] _080_/X vgnd vpwr scs8hd_or3_4
XFILLER_10_102 vpwr vgnd scs8hd_fill_2
XFILLER_10_113 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_6.INVTX1_1_.scs8hd_inv_1 chany_top_in[1] mux_left_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
XFILLER_53_71 vpwr vgnd scs8hd_fill_2
XANTENNA__108__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_38_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_19 vpwr vgnd scs8hd_fill_2
XFILLER_59_113 vgnd vpwr scs8hd_decap_8
Xmux_left_ipin_7.INVTX1_5_.scs8hd_inv_1 chany_top_in[7] mux_left_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_132_ _132_/A _131_/B _132_/Y vgnd vpwr scs8hd_nor2_4
X_201_ chany_bottom_in[8] chany_top_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_2_142 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_3.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_56 vgnd vpwr scs8hd_decap_4
XFILLER_0_78 vgnd vpwr scs8hd_decap_4
XANTENNA__110__B address[4] vgnd vpwr scs8hd_diode_2
XFILLER_9_21 vpwr vgnd scs8hd_fill_2
XFILLER_9_10 vpwr vgnd scs8hd_fill_2
XFILLER_0_89 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_2.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_ipin_7.LATCH_2_.latch/Q mux_left_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_60_39 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_ipin_6.INVTX1_1_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_47_127 vgnd vpwr scs8hd_decap_12
XFILLER_18_63 vgnd vpwr scs8hd_fill_1
XFILLER_18_85 vgnd vpwr scs8hd_decap_6
XFILLER_34_84 vpwr vgnd scs8hd_fill_2
XFILLER_50_50 vgnd vpwr scs8hd_decap_8
X_115_ _133_/A _118_/B _115_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__105__B _101_/B vgnd vpwr scs8hd_diode_2
XANTENNA__121__A _110_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_28 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__206__A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_29_40 vpwr vgnd scs8hd_fill_2
XFILLER_29_51 vpwr vgnd scs8hd_fill_2
XFILLER_29_62 vgnd vpwr scs8hd_decap_3
Xmux_left_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_ipin_5.LATCH_0_.latch/Q mux_left_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_61_60 vgnd vpwr scs8hd_fill_1
XANTENNA__116__A _142_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_2.LATCH_0_.latch_SLEEPB _088_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_119 vgnd vpwr scs8hd_decap_12
XFILLER_15_31 vpwr vgnd scs8hd_fill_2
Xmem_left_ipin_6.LATCH_1_.latch data_in mem_left_ipin_6.LATCH_1_.latch/Q _135_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_56_93 vgnd vpwr scs8hd_fill_1
Xmux_left_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_left_ipin_2.LATCH_3_.latch/Q mux_left_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
.ends

