VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cbx_1__0_
  CLASS BLOCK ;
  FOREIGN cbx_1__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 90.000 BY 83.600 ;
  PIN bottom_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 2.400 ;
    END
  END bottom_grid_pin_0_
  PIN bottom_grid_pin_10_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 2.400 ;
    END
  END bottom_grid_pin_10_
  PIN bottom_grid_pin_12_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 2.400 ;
    END
  END bottom_grid_pin_12_
  PIN bottom_grid_pin_14_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 2.400 ;
    END
  END bottom_grid_pin_14_
  PIN bottom_grid_pin_16_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 2.400 ;
    END
  END bottom_grid_pin_16_
  PIN bottom_grid_pin_2_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 2.400 ;
    END
  END bottom_grid_pin_2_
  PIN bottom_grid_pin_4_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 2.400 ;
    END
  END bottom_grid_pin_4_
  PIN bottom_grid_pin_6_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 2.400 ;
    END
  END bottom_grid_pin_6_
  PIN bottom_grid_pin_8_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 2.400 ;
    END
  END bottom_grid_pin_8_
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 2.400 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 2.400 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 2.400 43.480 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 2.400 64.560 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 2.400 66.600 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 2.400 69.320 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 2.400 71.360 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 2.400 73.400 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 2.400 75.440 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 2.400 77.480 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 2.400 79.520 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 2.400 81.560 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 2.400 83.600 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 2.400 45.520 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 2.400 47.560 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 2.400 49.600 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 2.400 52.320 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 2.400 54.360 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 2.400 56.400 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 2.400 58.440 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 2.400 60.480 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 2.400 62.520 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 2.400 1.320 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 2.400 22.400 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 2.400 24.440 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 2.400 26.480 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 2.400 28.520 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 2.400 30.560 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.000 2.400 32.600 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 2.400 35.320 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 2.400 37.360 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 2.400 39.400 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 2.400 41.440 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 2.400 3.360 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 2.400 5.400 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 2.400 7.440 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 2.400 9.480 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 2.400 11.520 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 2.400 13.560 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 2.400 15.600 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 2.400 18.320 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 2.400 20.360 ;
    END
  END chanx_left_out[9]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 87.600 42.880 90.000 43.480 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 87.600 63.960 90.000 64.560 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 87.600 66.000 90.000 66.600 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 87.600 68.720 90.000 69.320 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 87.600 70.760 90.000 71.360 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 87.600 72.800 90.000 73.400 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 87.600 74.840 90.000 75.440 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 87.600 76.880 90.000 77.480 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 87.600 78.920 90.000 79.520 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 87.600 80.960 90.000 81.560 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 87.600 83.000 90.000 83.600 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 87.600 44.920 90.000 45.520 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 87.600 46.960 90.000 47.560 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 87.600 49.000 90.000 49.600 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 87.600 51.720 90.000 52.320 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 87.600 53.760 90.000 54.360 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 87.600 55.800 90.000 56.400 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 87.600 57.840 90.000 58.440 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 87.600 59.880 90.000 60.480 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 87.600 61.920 90.000 62.520 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 87.600 0.720 90.000 1.320 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 87.600 21.800 90.000 22.400 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 87.600 23.840 90.000 24.440 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 87.600 25.880 90.000 26.480 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 87.600 27.920 90.000 28.520 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 87.600 29.960 90.000 30.560 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 87.600 32.000 90.000 32.600 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 87.600 34.720 90.000 35.320 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 87.600 36.760 90.000 37.360 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 87.600 38.800 90.000 39.400 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 87.600 40.840 90.000 41.440 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 87.600 2.760 90.000 3.360 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 87.600 4.800 90.000 5.400 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 87.600 6.840 90.000 7.440 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 87.600 8.880 90.000 9.480 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 87.600 10.920 90.000 11.520 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 87.600 12.960 90.000 13.560 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 87.600 15.000 90.000 15.600 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 87.600 17.720 90.000 18.320 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 87.600 19.760 90.000 20.360 ;
    END
  END chanx_right_out[9]
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 2.400 ;
    END
  END prog_clk
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 17.880 10.640 19.480 73.680 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 31.040 10.640 32.640 73.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 84.180 73.525 ;
      LAYER met1 ;
        RECT 3.750 10.640 86.410 76.460 ;
      LAYER met2 ;
        RECT 3.780 2.680 86.380 83.485 ;
        RECT 4.330 0.835 10.850 2.680 ;
        RECT 11.690 0.835 18.210 2.680 ;
        RECT 19.050 0.835 26.030 2.680 ;
        RECT 26.870 0.835 33.390 2.680 ;
        RECT 34.230 0.835 40.750 2.680 ;
        RECT 41.590 0.835 48.570 2.680 ;
        RECT 49.410 0.835 55.930 2.680 ;
        RECT 56.770 0.835 63.290 2.680 ;
        RECT 64.130 0.835 71.110 2.680 ;
        RECT 71.950 0.835 78.470 2.680 ;
        RECT 79.310 0.835 85.830 2.680 ;
      LAYER met3 ;
        RECT 2.800 82.600 87.200 83.465 ;
        RECT 2.400 81.960 87.600 82.600 ;
        RECT 2.800 80.560 87.200 81.960 ;
        RECT 2.400 79.920 87.600 80.560 ;
        RECT 2.800 78.520 87.200 79.920 ;
        RECT 2.400 77.880 87.600 78.520 ;
        RECT 2.800 76.480 87.200 77.880 ;
        RECT 2.400 75.840 87.600 76.480 ;
        RECT 2.800 74.440 87.200 75.840 ;
        RECT 2.400 73.800 87.600 74.440 ;
        RECT 2.800 72.400 87.200 73.800 ;
        RECT 2.400 71.760 87.600 72.400 ;
        RECT 2.800 70.360 87.200 71.760 ;
        RECT 2.400 69.720 87.600 70.360 ;
        RECT 2.800 68.320 87.200 69.720 ;
        RECT 2.400 67.000 87.600 68.320 ;
        RECT 2.800 65.600 87.200 67.000 ;
        RECT 2.400 64.960 87.600 65.600 ;
        RECT 2.800 63.560 87.200 64.960 ;
        RECT 2.400 62.920 87.600 63.560 ;
        RECT 2.800 61.520 87.200 62.920 ;
        RECT 2.400 60.880 87.600 61.520 ;
        RECT 2.800 59.480 87.200 60.880 ;
        RECT 2.400 58.840 87.600 59.480 ;
        RECT 2.800 57.440 87.200 58.840 ;
        RECT 2.400 56.800 87.600 57.440 ;
        RECT 2.800 55.400 87.200 56.800 ;
        RECT 2.400 54.760 87.600 55.400 ;
        RECT 2.800 53.360 87.200 54.760 ;
        RECT 2.400 52.720 87.600 53.360 ;
        RECT 2.800 51.320 87.200 52.720 ;
        RECT 2.400 50.000 87.600 51.320 ;
        RECT 2.800 48.600 87.200 50.000 ;
        RECT 2.400 47.960 87.600 48.600 ;
        RECT 2.800 46.560 87.200 47.960 ;
        RECT 2.400 45.920 87.600 46.560 ;
        RECT 2.800 44.520 87.200 45.920 ;
        RECT 2.400 43.880 87.600 44.520 ;
        RECT 2.800 42.480 87.200 43.880 ;
        RECT 2.400 41.840 87.600 42.480 ;
        RECT 2.800 40.440 87.200 41.840 ;
        RECT 2.400 39.800 87.600 40.440 ;
        RECT 2.800 38.400 87.200 39.800 ;
        RECT 2.400 37.760 87.600 38.400 ;
        RECT 2.800 36.360 87.200 37.760 ;
        RECT 2.400 35.720 87.600 36.360 ;
        RECT 2.800 34.320 87.200 35.720 ;
        RECT 2.400 33.000 87.600 34.320 ;
        RECT 2.800 31.600 87.200 33.000 ;
        RECT 2.400 30.960 87.600 31.600 ;
        RECT 2.800 29.560 87.200 30.960 ;
        RECT 2.400 28.920 87.600 29.560 ;
        RECT 2.800 27.520 87.200 28.920 ;
        RECT 2.400 26.880 87.600 27.520 ;
        RECT 2.800 25.480 87.200 26.880 ;
        RECT 2.400 24.840 87.600 25.480 ;
        RECT 2.800 23.440 87.200 24.840 ;
        RECT 2.400 22.800 87.600 23.440 ;
        RECT 2.800 21.400 87.200 22.800 ;
        RECT 2.400 20.760 87.600 21.400 ;
        RECT 2.800 19.360 87.200 20.760 ;
        RECT 2.400 18.720 87.600 19.360 ;
        RECT 2.800 17.320 87.200 18.720 ;
        RECT 2.400 16.000 87.600 17.320 ;
        RECT 2.800 14.600 87.200 16.000 ;
        RECT 2.400 13.960 87.600 14.600 ;
        RECT 2.800 12.560 87.200 13.960 ;
        RECT 2.400 11.920 87.600 12.560 ;
        RECT 2.800 10.520 87.200 11.920 ;
        RECT 2.400 9.880 87.600 10.520 ;
        RECT 2.800 8.480 87.200 9.880 ;
        RECT 2.400 7.840 87.600 8.480 ;
        RECT 2.800 6.440 87.200 7.840 ;
        RECT 2.400 5.800 87.600 6.440 ;
        RECT 2.800 4.400 87.200 5.800 ;
        RECT 2.400 3.760 87.600 4.400 ;
        RECT 2.800 2.360 87.200 3.760 ;
        RECT 2.400 1.720 87.600 2.360 ;
        RECT 2.800 0.855 87.200 1.720 ;
      LAYER met4 ;
        RECT 44.200 10.640 74.225 73.680 ;
  END
END cbx_1__0_
END LIBRARY

