magic
tech EFS8A
magscale 1 2
timestamp 1602531303
<< locali >>
rect 11471 24225 11598 24259
rect 1443 22049 1478 22083
rect 3007 22049 3042 22083
rect 5359 18921 5365 18955
rect 7567 18921 7573 18955
rect 11431 18921 11437 18955
rect 5359 18853 5393 18921
rect 7567 18853 7601 18921
rect 11431 18853 11465 18921
rect 1443 18785 1478 18819
rect 3801 18207 3835 18309
rect 5359 18071 5393 18139
rect 5359 18037 5365 18071
rect 15243 17697 15370 17731
rect 10051 14569 10057 14603
rect 3617 14331 3651 14569
rect 10051 14501 10085 14569
rect 8493 12631 8527 12801
rect 17233 12257 17394 12291
rect 17233 12087 17267 12257
rect 4813 10455 4847 10625
rect 7757 8823 7791 8925
rect 10333 8279 10367 8381
rect 5273 7735 5307 7837
rect 8211 6953 8217 6987
rect 8211 6885 8245 6953
rect 15347 5253 15485 5287
rect 11483 2601 11621 2635
<< viali >>
rect 6260 24225 6294 24259
rect 7364 24225 7398 24259
rect 11437 24225 11471 24259
rect 23556 24225 23590 24259
rect 24660 24225 24694 24259
rect 24731 24089 24765 24123
rect 6331 24021 6365 24055
rect 7435 24021 7469 24055
rect 10241 24021 10275 24055
rect 11667 24021 11701 24055
rect 23627 24021 23661 24055
rect 2513 23817 2547 23851
rect 6285 23817 6319 23851
rect 7849 23817 7883 23851
rect 11621 23817 11655 23851
rect 14381 23817 14415 23851
rect 17417 23817 17451 23851
rect 22385 23817 22419 23851
rect 23949 23817 23983 23851
rect 25145 23817 25179 23851
rect 25513 23817 25547 23851
rect 2191 23749 2225 23783
rect 8217 23681 8251 23715
rect 8907 23681 8941 23715
rect 10241 23681 10275 23715
rect 2120 23613 2154 23647
rect 7364 23613 7398 23647
rect 8804 23613 8838 23647
rect 9229 23613 9263 23647
rect 13896 23613 13930 23647
rect 16932 23613 16966 23647
rect 21900 23613 21934 23647
rect 24660 23613 24694 23647
rect 10333 23545 10367 23579
rect 10885 23545 10919 23579
rect 7435 23477 7469 23511
rect 10057 23477 10091 23511
rect 13967 23477 14001 23511
rect 17003 23477 17037 23511
rect 21971 23477 22005 23511
rect 24731 23477 24765 23511
rect 1593 23273 1627 23307
rect 3065 23273 3099 23307
rect 6929 23205 6963 23239
rect 9873 23205 9907 23239
rect 11437 23205 11471 23239
rect 1409 23137 1443 23171
rect 2881 23137 2915 23171
rect 6837 23069 6871 23103
rect 9781 23069 9815 23103
rect 10241 23069 10275 23103
rect 11345 23069 11379 23103
rect 11621 23069 11655 23103
rect 7389 23001 7423 23035
rect 5917 22729 5951 22763
rect 6653 22729 6687 22763
rect 11713 22729 11747 22763
rect 7849 22661 7883 22695
rect 6929 22593 6963 22627
rect 7389 22593 7423 22627
rect 8861 22593 8895 22627
rect 9505 22593 9539 22627
rect 11069 22593 11103 22627
rect 11345 22593 11379 22627
rect 3065 22525 3099 22559
rect 10149 22525 10183 22559
rect 10793 22525 10827 22559
rect 15368 22525 15402 22559
rect 1685 22457 1719 22491
rect 7021 22457 7055 22491
rect 8953 22457 8987 22491
rect 2513 22389 2547 22423
rect 2789 22389 2823 22423
rect 3249 22389 3283 22423
rect 6285 22389 6319 22423
rect 8677 22389 8711 22423
rect 9781 22389 9815 22423
rect 15439 22389 15473 22423
rect 15853 22389 15887 22423
rect 3111 22185 3145 22219
rect 4215 22185 4249 22219
rect 6837 22185 6871 22219
rect 8861 22185 8895 22219
rect 9873 22185 9907 22219
rect 1409 22049 1443 22083
rect 2973 22049 3007 22083
rect 4144 22049 4178 22083
rect 6745 22049 6779 22083
rect 9689 22049 9723 22083
rect 5089 21981 5123 22015
rect 10333 21981 10367 22015
rect 1547 21913 1581 21947
rect 1869 21845 1903 21879
rect 2237 21845 2271 21879
rect 1593 21641 1627 21675
rect 3249 21641 3283 21675
rect 4445 21641 4479 21675
rect 9689 21641 9723 21675
rect 10609 21641 10643 21675
rect 1961 21505 1995 21539
rect 3801 21505 3835 21539
rect 8677 21505 8711 21539
rect 5089 21437 5123 21471
rect 8585 21437 8619 21471
rect 9137 21437 9171 21471
rect 10425 21437 10459 21471
rect 2053 21369 2087 21403
rect 2605 21369 2639 21403
rect 3525 21369 3559 21403
rect 3617 21369 3651 21403
rect 4997 21369 5031 21403
rect 2973 21301 3007 21335
rect 4905 21301 4939 21335
rect 6469 21301 6503 21335
rect 11069 21301 11103 21335
rect 3525 21097 3559 21131
rect 4077 21097 4111 21131
rect 9827 21097 9861 21131
rect 2145 21029 2179 21063
rect 2697 21029 2731 21063
rect 5365 21029 5399 21063
rect 7573 20961 7607 20995
rect 9724 20961 9758 20995
rect 2053 20893 2087 20927
rect 5273 20893 5307 20927
rect 5549 20893 5583 20927
rect 7297 20893 7331 20927
rect 11437 20893 11471 20927
rect 1547 20553 1581 20587
rect 6009 20553 6043 20587
rect 9229 20553 9263 20587
rect 11391 20553 11425 20587
rect 12633 20553 12667 20587
rect 14105 20553 14139 20587
rect 25145 20553 25179 20587
rect 5181 20485 5215 20519
rect 8769 20485 8803 20519
rect 2973 20417 3007 20451
rect 3249 20417 3283 20451
rect 4629 20417 4663 20451
rect 1444 20349 1478 20383
rect 1869 20349 1903 20383
rect 9597 20349 9631 20383
rect 9781 20349 9815 20383
rect 11320 20349 11354 20383
rect 12449 20349 12483 20383
rect 13001 20349 13035 20383
rect 13620 20349 13654 20383
rect 24660 20349 24694 20383
rect 2789 20281 2823 20315
rect 3065 20281 3099 20315
rect 4721 20281 4755 20315
rect 5641 20281 5675 20315
rect 7113 20281 7147 20315
rect 7665 20281 7699 20315
rect 8217 20281 8251 20315
rect 8309 20281 8343 20315
rect 9689 20281 9723 20315
rect 2329 20213 2363 20247
rect 4445 20213 4479 20247
rect 8033 20213 8067 20247
rect 11805 20213 11839 20247
rect 13691 20213 13725 20247
rect 24731 20213 24765 20247
rect 1869 20009 1903 20043
rect 2973 20009 3007 20043
rect 4629 20009 4663 20043
rect 7573 20009 7607 20043
rect 1961 19941 1995 19975
rect 4997 19941 5031 19975
rect 5549 19941 5583 19975
rect 6653 19941 6687 19975
rect 8217 19941 8251 19975
rect 8769 19941 8803 19975
rect 9873 19941 9907 19975
rect 11713 19941 11747 19975
rect 11805 19941 11839 19975
rect 13185 19941 13219 19975
rect 2329 19873 2363 19907
rect 13461 19873 13495 19907
rect 4905 19805 4939 19839
rect 6561 19805 6595 19839
rect 7205 19805 7239 19839
rect 8125 19805 8159 19839
rect 9781 19805 9815 19839
rect 12357 19805 12391 19839
rect 10333 19737 10367 19771
rect 7849 19669 7883 19703
rect 12633 19669 12667 19703
rect 5641 19465 5675 19499
rect 6561 19465 6595 19499
rect 8401 19465 8435 19499
rect 8769 19465 8803 19499
rect 12173 19465 12207 19499
rect 13461 19465 13495 19499
rect 4905 19397 4939 19431
rect 11897 19397 11931 19431
rect 7481 19329 7515 19363
rect 10885 19329 10919 19363
rect 11483 19329 11517 19363
rect 12541 19329 12575 19363
rect 12817 19329 12851 19363
rect 2605 19261 2639 19295
rect 3341 19261 3375 19295
rect 3433 19261 3467 19295
rect 4077 19261 4111 19295
rect 9321 19261 9355 19295
rect 9873 19261 9907 19295
rect 11161 19261 11195 19295
rect 11380 19261 11414 19295
rect 4353 19193 4387 19227
rect 4445 19193 4479 19227
rect 7297 19193 7331 19227
rect 7802 19193 7836 19227
rect 12633 19193 12667 19227
rect 2053 19125 2087 19159
rect 5365 19125 5399 19159
rect 6101 19125 6135 19159
rect 9597 19125 9631 19159
rect 10057 19125 10091 19159
rect 4353 18921 4387 18955
rect 5365 18921 5399 18955
rect 5917 18921 5951 18955
rect 7573 18921 7607 18955
rect 8125 18921 8159 18955
rect 8493 18921 8527 18955
rect 11437 18921 11471 18955
rect 11989 18921 12023 18955
rect 12541 18921 12575 18955
rect 12909 18853 12943 18887
rect 13001 18853 13035 18887
rect 1409 18785 1443 18819
rect 2697 18785 2731 18819
rect 2881 18785 2915 18819
rect 3157 18717 3191 18751
rect 4997 18717 5031 18751
rect 7205 18717 7239 18751
rect 9965 18717 9999 18751
rect 11069 18717 11103 18751
rect 13185 18717 13219 18751
rect 1547 18581 1581 18615
rect 7021 18581 7055 18615
rect 8861 18581 8895 18615
rect 1593 18377 1627 18411
rect 3525 18377 3559 18411
rect 5917 18377 5951 18411
rect 7941 18377 7975 18411
rect 9965 18377 9999 18411
rect 11161 18377 11195 18411
rect 13461 18377 13495 18411
rect 3249 18309 3283 18343
rect 3801 18309 3835 18343
rect 7665 18241 7699 18275
rect 8585 18241 8619 18275
rect 8861 18241 8895 18275
rect 9597 18241 9631 18275
rect 10149 18241 10183 18275
rect 12817 18241 12851 18275
rect 2329 18173 2363 18207
rect 3801 18173 3835 18207
rect 3893 18173 3927 18207
rect 4997 18173 5031 18207
rect 6653 18173 6687 18207
rect 6929 18173 6963 18207
rect 7389 18173 7423 18207
rect 2237 18105 2271 18139
rect 2691 18105 2725 18139
rect 4445 18105 4479 18139
rect 4813 18105 4847 18139
rect 8401 18105 8435 18139
rect 8677 18105 8711 18139
rect 10241 18105 10275 18139
rect 10793 18105 10827 18139
rect 12541 18105 12575 18139
rect 12633 18105 12667 18139
rect 5365 18037 5399 18071
rect 11437 18037 11471 18071
rect 11805 18037 11839 18071
rect 12265 18037 12299 18071
rect 4997 17833 5031 17867
rect 5273 17833 5307 17867
rect 5641 17833 5675 17867
rect 13185 17833 13219 17867
rect 4398 17765 4432 17799
rect 7205 17765 7239 17799
rect 7481 17765 7515 17799
rect 8217 17765 8251 17799
rect 8769 17765 8803 17799
rect 9873 17765 9907 17799
rect 9965 17765 9999 17799
rect 10517 17765 10551 17799
rect 11666 17765 11700 17799
rect 12909 17765 12943 17799
rect 1444 17697 1478 17731
rect 2697 17697 2731 17731
rect 2881 17697 2915 17731
rect 3157 17697 3191 17731
rect 6469 17697 6503 17731
rect 7021 17697 7055 17731
rect 12265 17697 12299 17731
rect 13093 17697 13127 17731
rect 13553 17697 13587 17731
rect 15209 17697 15243 17731
rect 4077 17629 4111 17663
rect 8125 17629 8159 17663
rect 11345 17629 11379 17663
rect 1547 17493 1581 17527
rect 1961 17493 1995 17527
rect 2329 17493 2363 17527
rect 7849 17493 7883 17527
rect 15439 17493 15473 17527
rect 1593 17289 1627 17323
rect 2881 17289 2915 17323
rect 7021 17289 7055 17323
rect 9505 17289 9539 17323
rect 10885 17289 10919 17323
rect 11345 17289 11379 17323
rect 11805 17289 11839 17323
rect 12265 17289 12299 17323
rect 12725 17289 12759 17323
rect 13461 17289 13495 17323
rect 9137 17221 9171 17255
rect 13829 17153 13863 17187
rect 15393 17153 15427 17187
rect 1844 17085 1878 17119
rect 3525 17085 3559 17119
rect 4537 17085 4571 17119
rect 4629 17085 4663 17119
rect 5089 17085 5123 17119
rect 5641 17085 5675 17119
rect 6561 17085 6595 17119
rect 8217 17085 8251 17119
rect 9965 17085 9999 17119
rect 12541 17085 12575 17119
rect 3801 17017 3835 17051
rect 8538 17017 8572 17051
rect 9873 17017 9907 17051
rect 10327 17017 10361 17051
rect 1915 16949 1949 16983
rect 2513 16949 2547 16983
rect 4169 16949 4203 16983
rect 4721 16949 4755 16983
rect 7757 16949 7791 16983
rect 8125 16949 8159 16983
rect 3893 16745 3927 16779
rect 6745 16745 6779 16779
rect 9413 16745 9447 16779
rect 2513 16677 2547 16711
rect 2605 16677 2639 16711
rect 4261 16677 4295 16711
rect 6146 16677 6180 16711
rect 8401 16677 8435 16711
rect 9965 16677 9999 16711
rect 11069 16677 11103 16711
rect 1476 16609 1510 16643
rect 7665 16609 7699 16643
rect 8125 16609 8159 16643
rect 10609 16609 10643 16643
rect 10885 16609 10919 16643
rect 11989 16609 12023 16643
rect 4169 16541 4203 16575
rect 4445 16541 4479 16575
rect 5825 16541 5859 16575
rect 11897 16541 11931 16575
rect 3065 16473 3099 16507
rect 1547 16405 1581 16439
rect 1869 16405 1903 16439
rect 2329 16405 2363 16439
rect 3525 16405 3559 16439
rect 5089 16405 5123 16439
rect 8677 16405 8711 16439
rect 2513 16201 2547 16235
rect 4077 16201 4111 16235
rect 7665 16201 7699 16235
rect 9137 16201 9171 16235
rect 9505 16201 9539 16235
rect 11989 16201 12023 16235
rect 1501 16065 1535 16099
rect 2145 16065 2179 16099
rect 3341 16065 3375 16099
rect 10057 16065 10091 16099
rect 4537 15997 4571 16031
rect 5089 15997 5123 16031
rect 6193 15997 6227 16031
rect 8217 15997 8251 16031
rect 10701 15997 10735 16031
rect 11621 15997 11655 16031
rect 12541 15997 12575 16031
rect 1593 15929 1627 15963
rect 3065 15929 3099 15963
rect 3157 15929 3191 15963
rect 6837 15929 6871 15963
rect 7389 15929 7423 15963
rect 8538 15929 8572 15963
rect 10149 15929 10183 15963
rect 12449 15929 12483 15963
rect 2881 15861 2915 15895
rect 4629 15861 4663 15895
rect 5917 15861 5951 15895
rect 8033 15861 8067 15895
rect 9781 15861 9815 15895
rect 11069 15861 11103 15895
rect 1409 15657 1443 15691
rect 2237 15657 2271 15691
rect 3433 15657 3467 15691
rect 4997 15657 5031 15691
rect 10057 15657 10091 15691
rect 3893 15589 3927 15623
rect 4398 15589 4432 15623
rect 6193 15589 6227 15623
rect 8309 15589 8343 15623
rect 10425 15589 10459 15623
rect 11897 15589 11931 15623
rect 11989 15589 12023 15623
rect 1961 15521 1995 15555
rect 2421 15521 2455 15555
rect 2973 15521 3007 15555
rect 7573 15521 7607 15555
rect 8033 15521 8067 15555
rect 4077 15453 4111 15487
rect 6101 15453 6135 15487
rect 6377 15453 6411 15487
rect 10333 15453 10367 15487
rect 10977 15453 11011 15487
rect 12541 15453 12575 15487
rect 13369 15453 13403 15487
rect 8953 15385 8987 15419
rect 5273 15317 5307 15351
rect 5641 15317 5675 15351
rect 7205 15317 7239 15351
rect 8585 15317 8619 15351
rect 12817 15317 12851 15351
rect 1593 15113 1627 15147
rect 2513 15113 2547 15147
rect 3985 15113 4019 15147
rect 6653 15113 6687 15147
rect 8493 15113 8527 15147
rect 9965 15113 9999 15147
rect 11713 15113 11747 15147
rect 25145 15113 25179 15147
rect 9597 15045 9631 15079
rect 5917 14977 5951 15011
rect 7849 14977 7883 15011
rect 10241 14977 10275 15011
rect 1409 14909 1443 14943
rect 1961 14909 1995 14943
rect 3065 14909 3099 14943
rect 7113 14909 7147 14943
rect 7573 14909 7607 14943
rect 8677 14909 8711 14943
rect 10425 14909 10459 14943
rect 11345 14909 11379 14943
rect 12081 14909 12115 14943
rect 12817 14909 12851 14943
rect 19016 14909 19050 14943
rect 19441 14909 19475 14943
rect 24660 14909 24694 14943
rect 3386 14841 3420 14875
rect 4721 14841 4755 14875
rect 5273 14841 5307 14875
rect 5365 14841 5399 14875
rect 8217 14841 8251 14875
rect 8998 14841 9032 14875
rect 10746 14841 10780 14875
rect 12449 14841 12483 14875
rect 2973 14773 3007 14807
rect 4261 14773 4295 14807
rect 5089 14773 5123 14807
rect 6285 14773 6319 14807
rect 14013 14773 14047 14807
rect 19119 14773 19153 14807
rect 24731 14773 24765 14807
rect 3433 14569 3467 14603
rect 3617 14569 3651 14603
rect 6745 14569 6779 14603
rect 10057 14569 10091 14603
rect 10609 14569 10643 14603
rect 11253 14569 11287 14603
rect 11805 14569 11839 14603
rect 3157 14501 3191 14535
rect 1476 14433 1510 14467
rect 2697 14433 2731 14467
rect 2973 14433 3007 14467
rect 5819 14501 5853 14535
rect 8401 14501 8435 14535
rect 12173 14501 12207 14535
rect 12265 14501 12299 14535
rect 4445 14433 4479 14467
rect 4997 14433 5031 14467
rect 7665 14433 7699 14467
rect 8125 14433 8159 14467
rect 13737 14433 13771 14467
rect 15336 14433 15370 14467
rect 5457 14365 5491 14399
rect 9689 14365 9723 14399
rect 12541 14365 12575 14399
rect 13645 14365 13679 14399
rect 1547 14297 1581 14331
rect 3617 14297 3651 14331
rect 7113 14297 7147 14331
rect 1869 14229 1903 14263
rect 2329 14229 2363 14263
rect 3801 14229 3835 14263
rect 4353 14229 4387 14263
rect 4629 14229 4663 14263
rect 5365 14229 5399 14263
rect 6377 14229 6411 14263
rect 7573 14229 7607 14263
rect 8769 14229 8803 14263
rect 9045 14229 9079 14263
rect 9505 14229 9539 14263
rect 10885 14229 10919 14263
rect 15439 14229 15473 14263
rect 1593 14025 1627 14059
rect 4169 14025 4203 14059
rect 9505 14025 9539 14059
rect 12173 14025 12207 14059
rect 13185 14025 13219 14059
rect 13553 14025 13587 14059
rect 15669 14025 15703 14059
rect 11253 13957 11287 13991
rect 12633 13957 12667 13991
rect 2513 13889 2547 13923
rect 6653 13889 6687 13923
rect 9321 13889 9355 13923
rect 11805 13889 11839 13923
rect 13737 13889 13771 13923
rect 14657 13889 14691 13923
rect 1409 13821 1443 13855
rect 2973 13821 3007 13855
rect 3341 13821 3375 13855
rect 3525 13821 3559 13855
rect 4537 13821 4571 13855
rect 4629 13821 4663 13855
rect 5457 13821 5491 13855
rect 5641 13821 5675 13855
rect 6837 13821 6871 13855
rect 6929 13821 6963 13855
rect 8217 13821 8251 13855
rect 8585 13821 8619 13855
rect 9229 13821 9263 13855
rect 10333 13821 10367 13855
rect 10885 13821 10919 13855
rect 11161 13821 11195 13855
rect 12449 13821 12483 13855
rect 2145 13753 2179 13787
rect 3801 13753 3835 13787
rect 10149 13753 10183 13787
rect 13829 13753 13863 13787
rect 14381 13753 14415 13787
rect 4721 13685 4755 13719
rect 6009 13685 6043 13719
rect 7941 13685 7975 13719
rect 9873 13685 9907 13719
rect 15209 13685 15243 13719
rect 1961 13481 1995 13515
rect 4721 13481 4755 13515
rect 6009 13481 6043 13515
rect 8585 13481 8619 13515
rect 9413 13481 9447 13515
rect 12633 13481 12667 13515
rect 24731 13481 24765 13515
rect 6561 13413 6595 13447
rect 7205 13413 7239 13447
rect 7297 13413 7331 13447
rect 11621 13413 11655 13447
rect 11713 13413 11747 13447
rect 12909 13413 12943 13447
rect 13829 13413 13863 13447
rect 14381 13413 14415 13447
rect 1409 13345 1443 13379
rect 3065 13345 3099 13379
rect 4629 13345 4663 13379
rect 5273 13345 5307 13379
rect 5457 13345 5491 13379
rect 9781 13345 9815 13379
rect 10241 13345 10275 13379
rect 12265 13345 12299 13379
rect 15301 13345 15335 13379
rect 24660 13345 24694 13379
rect 3157 13277 3191 13311
rect 7573 13277 7607 13311
rect 10517 13277 10551 13311
rect 13737 13277 13771 13311
rect 3801 13209 3835 13243
rect 1593 13141 1627 13175
rect 2329 13141 2363 13175
rect 3525 13141 3559 13175
rect 4537 13141 4571 13175
rect 6929 13141 6963 13175
rect 8125 13141 8159 13175
rect 8861 13141 8895 13175
rect 10793 13141 10827 13175
rect 11161 13141 11195 13175
rect 15485 13141 15519 13175
rect 1593 12937 1627 12971
rect 1961 12937 1995 12971
rect 2513 12937 2547 12971
rect 7113 12937 7147 12971
rect 9321 12937 9355 12971
rect 13369 12937 13403 12971
rect 13645 12937 13679 12971
rect 15301 12937 15335 12971
rect 24685 12937 24719 12971
rect 4353 12869 4387 12903
rect 9137 12869 9171 12903
rect 3065 12801 3099 12835
rect 7665 12801 7699 12835
rect 8493 12801 8527 12835
rect 9229 12801 9263 12835
rect 10425 12801 10459 12835
rect 12449 12801 12483 12835
rect 1409 12733 1443 12767
rect 4905 12733 4939 12767
rect 5457 12733 5491 12767
rect 5917 12733 5951 12767
rect 2881 12665 2915 12699
rect 3157 12665 3191 12699
rect 3709 12665 3743 12699
rect 7389 12665 7423 12699
rect 7481 12665 7515 12699
rect 8861 12733 8895 12767
rect 9008 12733 9042 12767
rect 14105 12733 14139 12767
rect 14289 12733 14323 12767
rect 10333 12665 10367 12699
rect 10787 12665 10821 12699
rect 12770 12665 12804 12699
rect 14197 12665 14231 12699
rect 4629 12597 4663 12631
rect 4997 12597 5031 12631
rect 6561 12597 6595 12631
rect 8309 12597 8343 12631
rect 8493 12597 8527 12631
rect 8677 12597 8711 12631
rect 9873 12597 9907 12631
rect 11345 12597 11379 12631
rect 11713 12597 11747 12631
rect 12265 12597 12299 12631
rect 15761 12597 15795 12631
rect 1593 12393 1627 12427
rect 3525 12393 3559 12427
rect 4353 12393 4387 12427
rect 6745 12393 6779 12427
rect 8861 12393 8895 12427
rect 10793 12393 10827 12427
rect 11069 12393 11103 12427
rect 12449 12393 12483 12427
rect 2605 12325 2639 12359
rect 3157 12325 3191 12359
rect 6146 12325 6180 12359
rect 8309 12325 8343 12359
rect 10425 12325 10459 12359
rect 11437 12325 11471 12359
rect 15485 12325 15519 12359
rect 1409 12257 1443 12291
rect 4261 12257 4295 12291
rect 4629 12257 4663 12291
rect 5825 12257 5859 12291
rect 7573 12257 7607 12291
rect 9689 12257 9723 12291
rect 10241 12257 10275 12291
rect 13461 12257 13495 12291
rect 2513 12189 2547 12223
rect 3893 12189 3927 12223
rect 7941 12189 7975 12223
rect 11345 12189 11379 12223
rect 12817 12189 12851 12223
rect 15393 12189 15427 12223
rect 16037 12189 16071 12223
rect 7849 12121 7883 12155
rect 9229 12121 9263 12155
rect 11897 12121 11931 12155
rect 13921 12121 13955 12155
rect 17463 12121 17497 12155
rect 1961 12053 1995 12087
rect 2237 12053 2271 12087
rect 5089 12053 5123 12087
rect 5457 12053 5491 12087
rect 7297 12053 7331 12087
rect 7711 12053 7745 12087
rect 17233 12053 17267 12087
rect 4261 11849 4295 11883
rect 4997 11849 5031 11883
rect 7849 11849 7883 11883
rect 9229 11849 9263 11883
rect 10149 11849 10183 11883
rect 10701 11849 10735 11883
rect 11897 11849 11931 11883
rect 13553 11849 13587 11883
rect 14289 11849 14323 11883
rect 4886 11781 4920 11815
rect 5181 11781 5215 11815
rect 7343 11781 7377 11815
rect 7481 11781 7515 11815
rect 8907 11781 8941 11815
rect 9045 11781 9079 11815
rect 13829 11781 13863 11815
rect 2973 11713 3007 11747
rect 5089 11713 5123 11747
rect 7573 11713 7607 11747
rect 8585 11713 8619 11747
rect 9137 11713 9171 11747
rect 14473 11713 14507 11747
rect 15117 11713 15151 11747
rect 16957 11713 16991 11747
rect 1409 11645 1443 11679
rect 4629 11645 4663 11679
rect 10793 11645 10827 11679
rect 11345 11645 11379 11679
rect 12633 11645 12667 11679
rect 16037 11645 16071 11679
rect 2881 11577 2915 11611
rect 3294 11577 3328 11611
rect 4721 11577 4755 11611
rect 6561 11577 6595 11611
rect 7205 11577 7239 11611
rect 8769 11577 8803 11611
rect 11529 11577 11563 11611
rect 12995 11577 13029 11611
rect 14565 11577 14599 11611
rect 15945 11577 15979 11611
rect 1593 11509 1627 11543
rect 2053 11509 2087 11543
rect 2421 11509 2455 11543
rect 3893 11509 3927 11543
rect 5825 11509 5859 11543
rect 6193 11509 6227 11543
rect 7021 11509 7055 11543
rect 8217 11509 8251 11543
rect 9873 11509 9907 11543
rect 12265 11509 12299 11543
rect 15393 11509 15427 11543
rect 15761 11509 15795 11543
rect 17417 11509 17451 11543
rect 1409 11305 1443 11339
rect 4721 11305 4755 11339
rect 5549 11305 5583 11339
rect 7941 11305 7975 11339
rect 9137 11305 9171 11339
rect 11253 11305 11287 11339
rect 13829 11305 13863 11339
rect 2421 11237 2455 11271
rect 7113 11237 7147 11271
rect 8309 11237 8343 11271
rect 12081 11237 12115 11271
rect 12357 11237 12391 11271
rect 13271 11237 13305 11271
rect 14473 11237 14507 11271
rect 15393 11237 15427 11271
rect 15485 11237 15519 11271
rect 16037 11237 16071 11271
rect 3065 11169 3099 11203
rect 4905 11169 4939 11203
rect 7297 11169 7331 11203
rect 9689 11169 9723 11203
rect 11437 11169 11471 11203
rect 11897 11169 11931 11203
rect 12909 11169 12943 11203
rect 16900 11169 16934 11203
rect 5273 11101 5307 11135
rect 6377 11101 6411 11135
rect 7665 11101 7699 11135
rect 9836 11101 9870 11135
rect 10057 11101 10091 11135
rect 10425 11101 10459 11135
rect 10885 11101 10919 11135
rect 3709 11033 3743 11067
rect 6837 11033 6871 11067
rect 7573 11033 7607 11067
rect 9965 11033 9999 11067
rect 2145 10965 2179 10999
rect 4353 10965 4387 10999
rect 5043 10965 5077 10999
rect 5181 10965 5215 10999
rect 6009 10965 6043 10999
rect 7435 10965 7469 10999
rect 8769 10965 8803 10999
rect 12817 10965 12851 10999
rect 17003 10965 17037 10999
rect 2513 10761 2547 10795
rect 3893 10761 3927 10795
rect 6561 10761 6595 10795
rect 9045 10761 9079 10795
rect 9413 10761 9447 10795
rect 12173 10761 12207 10795
rect 14197 10761 14231 10795
rect 15669 10761 15703 10795
rect 15991 10761 16025 10795
rect 16865 10761 16899 10795
rect 24777 10761 24811 10795
rect 2218 10693 2252 10727
rect 2329 10693 2363 10727
rect 3755 10693 3789 10727
rect 4997 10693 5031 10727
rect 6285 10693 6319 10727
rect 7343 10693 7377 10727
rect 7481 10693 7515 10727
rect 8309 10693 8343 10727
rect 8907 10693 8941 10727
rect 10149 10693 10183 10727
rect 14933 10693 14967 10727
rect 15301 10693 15335 10727
rect 2421 10625 2455 10659
rect 3157 10625 3191 10659
rect 3985 10625 4019 10659
rect 4813 10625 4847 10659
rect 7573 10625 7607 10659
rect 8585 10625 8619 10659
rect 9137 10625 9171 10659
rect 9781 10625 9815 10659
rect 13277 10625 13311 10659
rect 1961 10557 1995 10591
rect 2053 10489 2087 10523
rect 3617 10489 3651 10523
rect 4353 10489 4387 10523
rect 5273 10557 5307 10591
rect 7205 10557 7239 10591
rect 8769 10557 8803 10591
rect 10793 10557 10827 10591
rect 11345 10557 11379 10591
rect 15888 10557 15922 10591
rect 16313 10557 16347 10591
rect 24593 10557 24627 10591
rect 25145 10557 25179 10591
rect 11529 10489 11563 10523
rect 12817 10489 12851 10523
rect 12909 10489 12943 10523
rect 14381 10489 14415 10523
rect 14473 10489 14507 10523
rect 3433 10421 3467 10455
rect 4813 10421 4847 10455
rect 5641 10421 5675 10455
rect 7021 10421 7055 10455
rect 7849 10421 7883 10455
rect 10701 10421 10735 10455
rect 11805 10421 11839 10455
rect 13737 10421 13771 10455
rect 1593 10217 1627 10251
rect 2881 10217 2915 10251
rect 5181 10217 5215 10251
rect 6837 10217 6871 10251
rect 8769 10217 8803 10251
rect 12357 10217 12391 10251
rect 14381 10217 14415 10251
rect 7389 10149 7423 10183
rect 8493 10149 8527 10183
rect 9413 10149 9447 10183
rect 9873 10149 9907 10183
rect 13179 10149 13213 10183
rect 15485 10149 15519 10183
rect 24317 10149 24351 10183
rect 1409 10081 1443 10115
rect 2145 10081 2179 10115
rect 2605 10081 2639 10115
rect 2789 10081 2823 10115
rect 4169 10081 4203 10115
rect 4537 10081 4571 10115
rect 4721 10081 4755 10115
rect 5733 10081 5767 10115
rect 5880 10081 5914 10115
rect 11253 10081 11287 10115
rect 11713 10081 11747 10115
rect 12817 10081 12851 10115
rect 6101 10013 6135 10047
rect 7757 10013 7791 10047
rect 9781 10013 9815 10047
rect 10057 10013 10091 10047
rect 11989 10013 12023 10047
rect 15393 10013 15427 10047
rect 15669 10013 15703 10047
rect 24225 10013 24259 10047
rect 2421 9945 2455 9979
rect 6009 9945 6043 9979
rect 7205 9945 7239 9979
rect 7665 9945 7699 9979
rect 13737 9945 13771 9979
rect 24777 9945 24811 9979
rect 3709 9877 3743 9911
rect 5549 9877 5583 9911
rect 6377 9877 6411 9911
rect 7527 9877 7561 9911
rect 8033 9877 8067 9911
rect 10793 9877 10827 9911
rect 12725 9877 12759 9911
rect 3893 9673 3927 9707
rect 4629 9673 4663 9707
rect 7481 9673 7515 9707
rect 7849 9673 7883 9707
rect 11713 9673 11747 9707
rect 15025 9673 15059 9707
rect 16221 9673 16255 9707
rect 25053 9673 25087 9707
rect 6653 9605 6687 9639
rect 7370 9605 7404 9639
rect 14013 9605 14047 9639
rect 1777 9537 1811 9571
rect 7573 9537 7607 9571
rect 14197 9537 14231 9571
rect 16589 9537 16623 9571
rect 24409 9537 24443 9571
rect 24685 9537 24719 9571
rect 1593 9469 1627 9503
rect 2145 9469 2179 9503
rect 3525 9469 3559 9503
rect 3709 9469 3743 9503
rect 5089 9469 5123 9503
rect 5825 9469 5859 9503
rect 8769 9469 8803 9503
rect 10517 9469 10551 9503
rect 12449 9469 12483 9503
rect 23765 9469 23799 9503
rect 4353 9401 4387 9435
rect 6193 9401 6227 9435
rect 7205 9401 7239 9435
rect 9090 9401 9124 9435
rect 10333 9401 10367 9435
rect 10838 9401 10872 9435
rect 12173 9401 12207 9435
rect 12770 9401 12804 9435
rect 13645 9401 13679 9435
rect 14749 9401 14783 9435
rect 15301 9401 15335 9435
rect 15393 9401 15427 9435
rect 15945 9401 15979 9435
rect 2421 9333 2455 9367
rect 2789 9333 2823 9367
rect 5457 9333 5491 9367
rect 7021 9333 7055 9367
rect 8217 9333 8251 9367
rect 8585 9333 8619 9367
rect 9689 9333 9723 9367
rect 9965 9333 9999 9367
rect 11437 9333 11471 9367
rect 13369 9333 13403 9367
rect 16773 9333 16807 9367
rect 23489 9333 23523 9367
rect 3157 9129 3191 9163
rect 3433 9129 3467 9163
rect 4353 9129 4387 9163
rect 6285 9129 6319 9163
rect 7481 9129 7515 9163
rect 12265 9129 12299 9163
rect 13921 9129 13955 9163
rect 6469 9061 6503 9095
rect 7849 9061 7883 9095
rect 9873 9061 9907 9095
rect 11069 9061 11103 9095
rect 11989 9061 12023 9095
rect 12633 9061 12667 9095
rect 13363 9061 13397 9095
rect 15669 9061 15703 9095
rect 16221 9061 16255 9095
rect 24225 9061 24259 9095
rect 1593 8993 1627 9027
rect 2973 8993 3007 9027
rect 4997 8993 5031 9027
rect 8033 8993 8067 9027
rect 8493 8993 8527 9027
rect 8769 8993 8803 9027
rect 11529 8993 11563 9027
rect 11805 8993 11839 9027
rect 13001 8993 13035 9027
rect 17116 8993 17150 9027
rect 24777 8993 24811 9027
rect 3801 8925 3835 8959
rect 4905 8925 4939 8959
rect 6837 8925 6871 8959
rect 7757 8925 7791 8959
rect 9781 8925 9815 8959
rect 15577 8925 15611 8959
rect 24133 8925 24167 8959
rect 2697 8857 2731 8891
rect 5917 8857 5951 8891
rect 9413 8857 9447 8891
rect 10333 8857 10367 8891
rect 1685 8789 1719 8823
rect 4813 8789 4847 8823
rect 6607 8789 6641 8823
rect 6745 8789 6779 8823
rect 7113 8789 7147 8823
rect 7757 8789 7791 8823
rect 9045 8789 9079 8823
rect 10701 8789 10735 8823
rect 14289 8789 14323 8823
rect 14565 8789 14599 8823
rect 17187 8789 17221 8823
rect 4353 8585 4387 8619
rect 5457 8585 5491 8619
rect 10057 8585 10091 8619
rect 11713 8585 11747 8619
rect 13645 8585 13679 8619
rect 16773 8585 16807 8619
rect 17141 8585 17175 8619
rect 3341 8517 3375 8551
rect 5641 8517 5675 8551
rect 7021 8517 7055 8551
rect 11989 8517 12023 8551
rect 13277 8517 13311 8551
rect 24777 8517 24811 8551
rect 3709 8449 3743 8483
rect 5549 8449 5583 8483
rect 8309 8449 8343 8483
rect 9781 8449 9815 8483
rect 14933 8449 14967 8483
rect 15577 8449 15611 8483
rect 15761 8449 15795 8483
rect 1593 8381 1627 8415
rect 1777 8381 1811 8415
rect 2421 8381 2455 8415
rect 3157 8381 3191 8415
rect 4169 8381 4203 8415
rect 5328 8381 5362 8415
rect 7297 8381 7331 8415
rect 7849 8381 7883 8415
rect 8677 8381 8711 8415
rect 9137 8381 9171 8415
rect 9505 8381 9539 8415
rect 10333 8381 10367 8415
rect 10609 8381 10643 8415
rect 11069 8381 11103 8415
rect 16313 8381 16347 8415
rect 24593 8381 24627 8415
rect 25145 8381 25179 8415
rect 2145 8313 2179 8347
rect 5181 8313 5215 8347
rect 8033 8313 8067 8347
rect 11345 8313 11379 8347
rect 12725 8313 12759 8347
rect 12817 8313 12851 8347
rect 14289 8313 14323 8347
rect 14381 8313 14415 8347
rect 2973 8245 3007 8279
rect 3985 8245 4019 8279
rect 4997 8245 5031 8279
rect 6561 8245 6595 8279
rect 10333 8245 10367 8279
rect 10425 8245 10459 8279
rect 14105 8245 14139 8279
rect 24041 8245 24075 8279
rect 24501 8245 24535 8279
rect 2237 8041 2271 8075
rect 3157 8041 3191 8075
rect 4537 8041 4571 8075
rect 5825 8041 5859 8075
rect 6561 8041 6595 8075
rect 9045 8041 9079 8075
rect 10793 8041 10827 8075
rect 11253 8041 11287 8075
rect 14105 8041 14139 8075
rect 14565 8041 14599 8075
rect 16313 8041 16347 8075
rect 1547 7973 1581 8007
rect 9413 7973 9447 8007
rect 11707 7973 11741 8007
rect 13093 7973 13127 8007
rect 15301 7973 15335 8007
rect 1444 7905 1478 7939
rect 2973 7905 3007 7939
rect 4997 7905 5031 7939
rect 5549 7905 5583 7939
rect 7021 7905 7055 7939
rect 7389 7905 7423 7939
rect 7573 7905 7607 7939
rect 8033 7905 8067 7939
rect 9781 7905 9815 7939
rect 10241 7905 10275 7939
rect 11345 7905 11379 7939
rect 12725 7905 12759 7939
rect 13369 7905 13403 7939
rect 15393 7905 15427 7939
rect 5273 7837 5307 7871
rect 8309 7837 8343 7871
rect 10517 7837 10551 7871
rect 4905 7769 4939 7803
rect 8585 7769 8619 7803
rect 1869 7701 1903 7735
rect 5181 7701 5215 7735
rect 5273 7701 5307 7735
rect 6377 7701 6411 7735
rect 12265 7701 12299 7735
rect 1823 7497 1857 7531
rect 2145 7497 2179 7531
rect 2973 7497 3007 7531
rect 4077 7497 4111 7531
rect 5089 7497 5123 7531
rect 5733 7497 5767 7531
rect 8493 7497 8527 7531
rect 9781 7497 9815 7531
rect 10149 7497 10183 7531
rect 11897 7497 11931 7531
rect 12173 7497 12207 7531
rect 13645 7497 13679 7531
rect 15393 7497 15427 7531
rect 24731 7497 24765 7531
rect 2605 7361 2639 7395
rect 12449 7361 12483 7395
rect 14289 7361 14323 7395
rect 14565 7361 14599 7395
rect 1752 7293 1786 7327
rect 3893 7293 3927 7327
rect 4353 7293 4387 7327
rect 4905 7293 4939 7327
rect 7113 7293 7147 7327
rect 7573 7293 7607 7327
rect 10793 7293 10827 7327
rect 11253 7293 11287 7327
rect 24660 7293 24694 7327
rect 5365 7225 5399 7259
rect 8125 7225 8159 7259
rect 8769 7225 8803 7259
rect 8861 7225 8895 7259
rect 9413 7225 9447 7259
rect 11529 7225 11563 7259
rect 12770 7225 12804 7259
rect 14381 7225 14415 7259
rect 6561 7157 6595 7191
rect 7389 7157 7423 7191
rect 10609 7157 10643 7191
rect 13369 7157 13403 7191
rect 14105 7157 14139 7191
rect 25145 7157 25179 7191
rect 1915 6953 1949 6987
rect 4813 6953 4847 6987
rect 7113 6953 7147 6987
rect 7665 6953 7699 6987
rect 8217 6953 8251 6987
rect 9413 6953 9447 6987
rect 9965 6953 9999 6987
rect 10885 6953 10919 6987
rect 12449 6953 12483 6987
rect 12817 6953 12851 6987
rect 13829 6885 13863 6919
rect 14381 6885 14415 6919
rect 15301 6885 15335 6919
rect 1844 6817 1878 6851
rect 4629 6817 4663 6851
rect 6101 6817 6135 6851
rect 9873 6817 9907 6851
rect 11345 6817 11379 6851
rect 15945 6817 15979 6851
rect 7849 6749 7883 6783
rect 11253 6749 11287 6783
rect 13737 6749 13771 6783
rect 6285 6681 6319 6715
rect 13461 6681 13495 6715
rect 8769 6613 8803 6647
rect 9045 6613 9079 6647
rect 2329 6409 2363 6443
rect 6193 6409 6227 6443
rect 9413 6409 9447 6443
rect 11345 6409 11379 6443
rect 13185 6409 13219 6443
rect 14473 6409 14507 6443
rect 15945 6409 15979 6443
rect 1547 6341 1581 6375
rect 5365 6341 5399 6375
rect 10885 6341 10919 6375
rect 7665 6273 7699 6307
rect 10057 6273 10091 6307
rect 10333 6273 10367 6307
rect 13461 6273 13495 6307
rect 14105 6273 14139 6307
rect 15301 6273 15335 6307
rect 1444 6205 1478 6239
rect 5181 6205 5215 6239
rect 5641 6205 5675 6239
rect 6653 6205 6687 6239
rect 7021 6205 7055 6239
rect 8493 6205 8527 6239
rect 9781 6205 9815 6239
rect 1869 6137 1903 6171
rect 8814 6137 8848 6171
rect 10425 6137 10459 6171
rect 13553 6137 13587 6171
rect 15025 6137 15059 6171
rect 15117 6137 15151 6171
rect 4629 6069 4663 6103
rect 8033 6069 8067 6103
rect 8309 6069 8343 6103
rect 14841 6069 14875 6103
rect 6193 5865 6227 5899
rect 8861 5865 8895 5899
rect 13737 5865 13771 5899
rect 9873 5797 9907 5831
rect 11253 5797 11287 5831
rect 12586 5797 12620 5831
rect 15301 5797 15335 5831
rect 6009 5729 6043 5763
rect 7481 5729 7515 5763
rect 7941 5729 7975 5763
rect 8493 5729 8527 5763
rect 12265 5729 12299 5763
rect 14080 5729 14114 5763
rect 15393 5729 15427 5763
rect 8217 5661 8251 5695
rect 9781 5661 9815 5695
rect 10425 5661 10459 5695
rect 14933 5661 14967 5695
rect 10793 5525 10827 5559
rect 13185 5525 13219 5559
rect 14151 5525 14185 5559
rect 14565 5525 14599 5559
rect 6009 5321 6043 5355
rect 7297 5321 7331 5355
rect 9689 5321 9723 5355
rect 11161 5321 11195 5355
rect 12265 5321 12299 5355
rect 13001 5321 13035 5355
rect 13461 5321 13495 5355
rect 22247 5321 22281 5355
rect 14289 5253 14323 5287
rect 14657 5253 14691 5287
rect 15485 5253 15519 5287
rect 16037 5253 16071 5287
rect 8401 5185 8435 5219
rect 10241 5185 10275 5219
rect 10517 5185 10551 5219
rect 12541 5185 12575 5219
rect 7113 5117 7147 5151
rect 15276 5117 15310 5151
rect 22176 5117 22210 5151
rect 8722 5049 8756 5083
rect 10057 5049 10091 5083
rect 10333 5049 10367 5083
rect 13737 5049 13771 5083
rect 13829 5049 13863 5083
rect 15761 5049 15795 5083
rect 7665 4981 7699 5015
rect 8309 4981 8343 5015
rect 9321 4981 9355 5015
rect 22661 4981 22695 5015
rect 7481 4777 7515 4811
rect 7941 4777 7975 4811
rect 8401 4777 8435 4811
rect 10149 4777 10183 4811
rect 23811 4777 23845 4811
rect 13829 4709 13863 4743
rect 10460 4641 10494 4675
rect 10563 4641 10597 4675
rect 11437 4641 11471 4675
rect 15301 4641 15335 4675
rect 23740 4641 23774 4675
rect 13737 4573 13771 4607
rect 14013 4573 14047 4607
rect 11621 4437 11655 4471
rect 15485 4437 15519 4471
rect 7573 4233 7607 4267
rect 10885 4233 10919 4267
rect 11437 4233 11471 4267
rect 13185 4233 13219 4267
rect 15301 4233 15335 4267
rect 8125 4097 8159 4131
rect 9965 4029 9999 4063
rect 13461 4029 13495 4063
rect 24660 4029 24694 4063
rect 8446 3961 8480 3995
rect 9873 3961 9907 3995
rect 14105 3961 14139 3995
rect 14381 3961 14415 3995
rect 7941 3893 7975 3927
rect 9045 3893 9079 3927
rect 9781 3893 9815 3927
rect 23949 3893 23983 3927
rect 24731 3893 24765 3927
rect 25145 3893 25179 3927
rect 13737 3689 13771 3723
rect 9965 3621 9999 3655
rect 8677 3553 8711 3587
rect 8033 3485 8067 3519
rect 9873 3485 9907 3519
rect 11345 3485 11379 3519
rect 10425 3417 10459 3451
rect 8033 3145 8067 3179
rect 9229 3145 9263 3179
rect 9597 3145 9631 3179
rect 10701 3077 10735 3111
rect 7665 3009 7699 3043
rect 10425 3009 10459 3043
rect 11288 2941 11322 2975
rect 11713 2941 11747 2975
rect 7297 2873 7331 2907
rect 8217 2873 8251 2907
rect 8309 2873 8343 2907
rect 8861 2873 8895 2907
rect 9781 2873 9815 2907
rect 9873 2873 9907 2907
rect 11069 2873 11103 2907
rect 11391 2873 11425 2907
rect 5687 2601 5721 2635
rect 7067 2601 7101 2635
rect 8079 2601 8113 2635
rect 11621 2601 11655 2635
rect 13047 2601 13081 2635
rect 9597 2533 9631 2567
rect 9965 2533 9999 2567
rect 20545 2533 20579 2567
rect 5584 2465 5618 2499
rect 6996 2465 7030 2499
rect 7389 2465 7423 2499
rect 8008 2465 8042 2499
rect 11412 2465 11446 2499
rect 12944 2465 12978 2499
rect 18797 2465 18831 2499
rect 19349 2465 19383 2499
rect 19993 2465 20027 2499
rect 24660 2465 24694 2499
rect 9229 2397 9263 2431
rect 9873 2397 9907 2431
rect 10149 2397 10183 2431
rect 13369 2397 13403 2431
rect 20177 2329 20211 2363
rect 6009 2261 6043 2295
rect 8493 2261 8527 2295
rect 11805 2261 11839 2295
rect 18981 2261 19015 2295
rect 24731 2261 24765 2295
rect 25145 2261 25179 2295
<< metal1 >>
rect 14 27072 20 27124
rect 72 27112 78 27124
rect 750 27112 756 27124
rect 72 27084 756 27112
rect 72 27072 78 27084
rect 750 27072 756 27084
rect 808 27072 814 27124
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 23934 24324 23940 24336
rect 23559 24296 23940 24324
rect 6270 24265 6276 24268
rect 6248 24259 6276 24265
rect 6248 24256 6260 24259
rect 6183 24228 6260 24256
rect 6248 24225 6260 24228
rect 6328 24256 6334 24268
rect 7006 24256 7012 24268
rect 6328 24228 7012 24256
rect 6248 24219 6276 24225
rect 6270 24216 6276 24219
rect 6328 24216 6334 24228
rect 7006 24216 7012 24228
rect 7064 24216 7070 24268
rect 7352 24259 7410 24265
rect 7352 24225 7364 24259
rect 7398 24256 7410 24259
rect 8202 24256 8208 24268
rect 7398 24228 8208 24256
rect 7398 24225 7410 24228
rect 7352 24219 7410 24225
rect 8202 24216 8208 24228
rect 8260 24216 8266 24268
rect 11425 24259 11483 24265
rect 11425 24225 11437 24259
rect 11471 24256 11483 24259
rect 11606 24256 11612 24268
rect 11471 24228 11612 24256
rect 11471 24225 11483 24228
rect 11425 24219 11483 24225
rect 11606 24216 11612 24228
rect 11664 24216 11670 24268
rect 23559 24265 23587 24296
rect 23934 24284 23940 24296
rect 23992 24324 23998 24336
rect 25406 24324 25412 24336
rect 23992 24296 25412 24324
rect 23992 24284 23998 24296
rect 25406 24284 25412 24296
rect 25464 24284 25470 24336
rect 23544 24259 23602 24265
rect 23544 24225 23556 24259
rect 23590 24225 23602 24259
rect 23544 24219 23602 24225
rect 24648 24259 24706 24265
rect 24648 24225 24660 24259
rect 24694 24256 24706 24259
rect 25130 24256 25136 24268
rect 24694 24228 25136 24256
rect 24694 24225 24706 24228
rect 24648 24219 24706 24225
rect 25130 24216 25136 24228
rect 25188 24216 25194 24268
rect 22186 24080 22192 24132
rect 22244 24120 22250 24132
rect 24719 24123 24777 24129
rect 24719 24120 24731 24123
rect 22244 24092 24731 24120
rect 22244 24080 22250 24092
rect 24719 24089 24731 24092
rect 24765 24089 24777 24123
rect 24719 24083 24777 24089
rect 6319 24055 6377 24061
rect 6319 24021 6331 24055
rect 6365 24052 6377 24055
rect 6730 24052 6736 24064
rect 6365 24024 6736 24052
rect 6365 24021 6377 24024
rect 6319 24015 6377 24021
rect 6730 24012 6736 24024
rect 6788 24012 6794 24064
rect 6822 24012 6828 24064
rect 6880 24052 6886 24064
rect 7423 24055 7481 24061
rect 7423 24052 7435 24055
rect 6880 24024 7435 24052
rect 6880 24012 6886 24024
rect 7423 24021 7435 24024
rect 7469 24021 7481 24055
rect 10226 24052 10232 24064
rect 10187 24024 10232 24052
rect 7423 24015 7481 24021
rect 10226 24012 10232 24024
rect 10284 24012 10290 24064
rect 11330 24012 11336 24064
rect 11388 24052 11394 24064
rect 11655 24055 11713 24061
rect 11655 24052 11667 24055
rect 11388 24024 11667 24052
rect 11388 24012 11394 24024
rect 11655 24021 11667 24024
rect 11701 24021 11713 24055
rect 11655 24015 11713 24021
rect 20622 24012 20628 24064
rect 20680 24052 20686 24064
rect 23615 24055 23673 24061
rect 23615 24052 23627 24055
rect 20680 24024 23627 24052
rect 20680 24012 20686 24024
rect 23615 24021 23627 24024
rect 23661 24021 23673 24055
rect 23615 24015 23673 24021
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 2498 23848 2504 23860
rect 2459 23820 2504 23848
rect 2498 23808 2504 23820
rect 2556 23808 2562 23860
rect 6270 23848 6276 23860
rect 6231 23820 6276 23848
rect 6270 23808 6276 23820
rect 6328 23808 6334 23860
rect 7837 23851 7895 23857
rect 7837 23817 7849 23851
rect 7883 23848 7895 23851
rect 8938 23848 8944 23860
rect 7883 23820 8944 23848
rect 7883 23817 7895 23820
rect 7837 23811 7895 23817
rect 2179 23783 2237 23789
rect 2179 23749 2191 23783
rect 2225 23780 2237 23783
rect 7742 23780 7748 23792
rect 2225 23752 7748 23780
rect 2225 23749 2237 23752
rect 2179 23743 2237 23749
rect 7742 23740 7748 23752
rect 7800 23740 7806 23792
rect 2108 23647 2166 23653
rect 2108 23613 2120 23647
rect 2154 23644 2166 23647
rect 2498 23644 2504 23656
rect 2154 23616 2504 23644
rect 2154 23613 2166 23616
rect 2108 23607 2166 23613
rect 2498 23604 2504 23616
rect 2556 23604 2562 23656
rect 7352 23647 7410 23653
rect 7352 23613 7364 23647
rect 7398 23644 7410 23647
rect 7852 23644 7880 23811
rect 8938 23808 8944 23820
rect 8996 23808 9002 23860
rect 11606 23848 11612 23860
rect 11567 23820 11612 23848
rect 11606 23808 11612 23820
rect 11664 23808 11670 23860
rect 14369 23851 14427 23857
rect 14369 23817 14381 23851
rect 14415 23848 14427 23851
rect 15470 23848 15476 23860
rect 14415 23820 15476 23848
rect 14415 23817 14427 23820
rect 14369 23811 14427 23817
rect 8202 23712 8208 23724
rect 8163 23684 8208 23712
rect 8202 23672 8208 23684
rect 8260 23672 8266 23724
rect 8895 23715 8953 23721
rect 8895 23681 8907 23715
rect 8941 23712 8953 23715
rect 10226 23712 10232 23724
rect 8941 23684 10232 23712
rect 8941 23681 8953 23684
rect 8895 23675 8953 23681
rect 10226 23672 10232 23684
rect 10284 23672 10290 23724
rect 7398 23616 7880 23644
rect 8792 23647 8850 23653
rect 7398 23613 7410 23616
rect 7352 23607 7410 23613
rect 8792 23613 8804 23647
rect 8838 23644 8850 23647
rect 9217 23647 9275 23653
rect 9217 23644 9229 23647
rect 8838 23616 9229 23644
rect 8838 23613 8850 23616
rect 8792 23607 8850 23613
rect 9217 23613 9229 23616
rect 9263 23613 9275 23647
rect 9217 23607 9275 23613
rect 13884 23647 13942 23653
rect 13884 23613 13896 23647
rect 13930 23644 13942 23647
rect 14384 23644 14412 23811
rect 15470 23808 15476 23820
rect 15528 23808 15534 23860
rect 17405 23851 17463 23857
rect 17405 23817 17417 23851
rect 17451 23848 17463 23851
rect 18782 23848 18788 23860
rect 17451 23820 18788 23848
rect 17451 23817 17463 23820
rect 17405 23811 17463 23817
rect 13930 23616 14412 23644
rect 16920 23647 16978 23653
rect 13930 23613 13942 23616
rect 13884 23607 13942 23613
rect 16920 23613 16932 23647
rect 16966 23644 16978 23647
rect 17420 23644 17448 23811
rect 18782 23808 18788 23820
rect 18840 23808 18846 23860
rect 22373 23851 22431 23857
rect 22373 23817 22385 23851
rect 22419 23848 22431 23851
rect 23750 23848 23756 23860
rect 22419 23820 23756 23848
rect 22419 23817 22431 23820
rect 22373 23811 22431 23817
rect 16966 23616 17448 23644
rect 21888 23647 21946 23653
rect 16966 23613 16978 23616
rect 16920 23607 16978 23613
rect 21888 23613 21900 23647
rect 21934 23644 21946 23647
rect 22388 23644 22416 23811
rect 23750 23808 23756 23820
rect 23808 23808 23814 23860
rect 23934 23848 23940 23860
rect 23895 23820 23940 23848
rect 23934 23808 23940 23820
rect 23992 23808 23998 23860
rect 25130 23848 25136 23860
rect 25091 23820 25136 23848
rect 25130 23808 25136 23820
rect 25188 23808 25194 23860
rect 25501 23851 25559 23857
rect 25501 23817 25513 23851
rect 25547 23848 25559 23851
rect 27062 23848 27068 23860
rect 25547 23820 27068 23848
rect 25547 23817 25559 23820
rect 25501 23811 25559 23817
rect 21934 23616 22416 23644
rect 24648 23647 24706 23653
rect 21934 23613 21946 23616
rect 21888 23607 21946 23613
rect 24648 23613 24660 23647
rect 24694 23644 24706 23647
rect 25516 23644 25544 23811
rect 27062 23808 27068 23820
rect 27120 23808 27126 23860
rect 24694 23616 25544 23644
rect 24694 23613 24706 23616
rect 24648 23607 24706 23613
rect 5994 23536 6000 23588
rect 6052 23576 6058 23588
rect 8807 23576 8835 23607
rect 6052 23548 8835 23576
rect 10321 23579 10379 23585
rect 6052 23536 6058 23548
rect 10321 23545 10333 23579
rect 10367 23545 10379 23579
rect 10321 23539 10379 23545
rect 10873 23579 10931 23585
rect 10873 23545 10885 23579
rect 10919 23576 10931 23579
rect 11606 23576 11612 23588
rect 10919 23548 11612 23576
rect 10919 23545 10931 23548
rect 10873 23539 10931 23545
rect 6638 23468 6644 23520
rect 6696 23508 6702 23520
rect 7423 23511 7481 23517
rect 7423 23508 7435 23511
rect 6696 23480 7435 23508
rect 6696 23468 6702 23480
rect 7423 23477 7435 23480
rect 7469 23477 7481 23511
rect 7423 23471 7481 23477
rect 9950 23468 9956 23520
rect 10008 23508 10014 23520
rect 10045 23511 10103 23517
rect 10045 23508 10057 23511
rect 10008 23480 10057 23508
rect 10008 23468 10014 23480
rect 10045 23477 10057 23480
rect 10091 23508 10103 23511
rect 10336 23508 10364 23539
rect 11606 23536 11612 23548
rect 11664 23536 11670 23588
rect 10091 23480 10364 23508
rect 10091 23477 10103 23480
rect 10045 23471 10103 23477
rect 13722 23468 13728 23520
rect 13780 23508 13786 23520
rect 13955 23511 14013 23517
rect 13955 23508 13967 23511
rect 13780 23480 13967 23508
rect 13780 23468 13786 23480
rect 13955 23477 13967 23480
rect 14001 23477 14013 23511
rect 13955 23471 14013 23477
rect 15746 23468 15752 23520
rect 15804 23508 15810 23520
rect 16991 23511 17049 23517
rect 16991 23508 17003 23511
rect 15804 23480 17003 23508
rect 15804 23468 15810 23480
rect 16991 23477 17003 23480
rect 17037 23477 17049 23511
rect 16991 23471 17049 23477
rect 19978 23468 19984 23520
rect 20036 23508 20042 23520
rect 21959 23511 22017 23517
rect 21959 23508 21971 23511
rect 20036 23480 21971 23508
rect 20036 23468 20042 23480
rect 21959 23477 21971 23480
rect 22005 23477 22017 23511
rect 21959 23471 22017 23477
rect 23934 23468 23940 23520
rect 23992 23508 23998 23520
rect 24719 23511 24777 23517
rect 24719 23508 24731 23511
rect 23992 23480 24731 23508
rect 23992 23468 23998 23480
rect 24719 23477 24731 23480
rect 24765 23477 24777 23511
rect 24719 23471 24777 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 1578 23304 1584 23316
rect 1539 23276 1584 23304
rect 1578 23264 1584 23276
rect 1636 23264 1642 23316
rect 3053 23307 3111 23313
rect 3053 23273 3065 23307
rect 3099 23304 3111 23307
rect 3970 23304 3976 23316
rect 3099 23276 3976 23304
rect 3099 23273 3111 23276
rect 3053 23267 3111 23273
rect 3970 23264 3976 23276
rect 4028 23264 4034 23316
rect 6914 23236 6920 23248
rect 6875 23208 6920 23236
rect 6914 23196 6920 23208
rect 6972 23196 6978 23248
rect 9766 23196 9772 23248
rect 9824 23236 9830 23248
rect 9861 23239 9919 23245
rect 9861 23236 9873 23239
rect 9824 23208 9873 23236
rect 9824 23196 9830 23208
rect 9861 23205 9873 23208
rect 9907 23205 9919 23239
rect 11422 23236 11428 23248
rect 11383 23208 11428 23236
rect 9861 23199 9919 23205
rect 11422 23196 11428 23208
rect 11480 23196 11486 23248
rect 1394 23168 1400 23180
rect 1355 23140 1400 23168
rect 1394 23128 1400 23140
rect 1452 23128 1458 23180
rect 2498 23128 2504 23180
rect 2556 23168 2562 23180
rect 2869 23171 2927 23177
rect 2869 23168 2881 23171
rect 2556 23140 2881 23168
rect 2556 23128 2562 23140
rect 2869 23137 2881 23140
rect 2915 23137 2927 23171
rect 2869 23131 2927 23137
rect 6546 23060 6552 23112
rect 6604 23100 6610 23112
rect 6822 23100 6828 23112
rect 6604 23072 6828 23100
rect 6604 23060 6610 23072
rect 6822 23060 6828 23072
rect 6880 23060 6886 23112
rect 9769 23103 9827 23109
rect 9769 23069 9781 23103
rect 9815 23100 9827 23103
rect 10134 23100 10140 23112
rect 9815 23072 10140 23100
rect 9815 23069 9827 23072
rect 9769 23063 9827 23069
rect 10134 23060 10140 23072
rect 10192 23060 10198 23112
rect 10226 23060 10232 23112
rect 10284 23100 10290 23112
rect 11330 23100 11336 23112
rect 10284 23072 10329 23100
rect 11291 23072 11336 23100
rect 10284 23060 10290 23072
rect 11330 23060 11336 23072
rect 11388 23060 11394 23112
rect 11606 23100 11612 23112
rect 11567 23072 11612 23100
rect 11606 23060 11612 23072
rect 11664 23060 11670 23112
rect 7374 23032 7380 23044
rect 7335 23004 7380 23032
rect 7374 22992 7380 23004
rect 7432 22992 7438 23044
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 5905 22763 5963 22769
rect 5905 22729 5917 22763
rect 5951 22760 5963 22763
rect 6546 22760 6552 22772
rect 5951 22732 6552 22760
rect 5951 22729 5963 22732
rect 5905 22723 5963 22729
rect 6546 22720 6552 22732
rect 6604 22720 6610 22772
rect 6641 22763 6699 22769
rect 6641 22729 6653 22763
rect 6687 22760 6699 22763
rect 6914 22760 6920 22772
rect 6687 22732 6920 22760
rect 6687 22729 6699 22732
rect 6641 22723 6699 22729
rect 6914 22720 6920 22732
rect 6972 22720 6978 22772
rect 11330 22720 11336 22772
rect 11388 22760 11394 22772
rect 11701 22763 11759 22769
rect 11701 22760 11713 22763
rect 11388 22732 11713 22760
rect 11388 22720 11394 22732
rect 11701 22729 11713 22732
rect 11747 22729 11759 22763
rect 11701 22723 11759 22729
rect 7837 22695 7895 22701
rect 7837 22692 7849 22695
rect 6932 22664 7849 22692
rect 6730 22584 6736 22636
rect 6788 22624 6794 22636
rect 6932 22633 6960 22664
rect 7837 22661 7849 22664
rect 7883 22661 7895 22695
rect 7837 22655 7895 22661
rect 6917 22627 6975 22633
rect 6917 22624 6929 22627
rect 6788 22596 6929 22624
rect 6788 22584 6794 22596
rect 6917 22593 6929 22596
rect 6963 22593 6975 22627
rect 7374 22624 7380 22636
rect 7335 22596 7380 22624
rect 6917 22587 6975 22593
rect 7374 22584 7380 22596
rect 7432 22584 7438 22636
rect 7742 22584 7748 22636
rect 7800 22624 7806 22636
rect 8846 22624 8852 22636
rect 7800 22596 8852 22624
rect 7800 22584 7806 22596
rect 8846 22584 8852 22596
rect 8904 22584 8910 22636
rect 9490 22624 9496 22636
rect 9403 22596 9496 22624
rect 9490 22584 9496 22596
rect 9548 22624 9554 22636
rect 10226 22624 10232 22636
rect 9548 22596 10232 22624
rect 9548 22584 9554 22596
rect 10226 22584 10232 22596
rect 10284 22584 10290 22636
rect 11057 22627 11115 22633
rect 11057 22593 11069 22627
rect 11103 22624 11115 22627
rect 11333 22627 11391 22633
rect 11333 22624 11345 22627
rect 11103 22596 11345 22624
rect 11103 22593 11115 22596
rect 11057 22587 11115 22593
rect 11333 22593 11345 22596
rect 11379 22624 11391 22627
rect 11422 22624 11428 22636
rect 11379 22596 11428 22624
rect 11379 22593 11391 22596
rect 11333 22587 11391 22593
rect 11422 22584 11428 22596
rect 11480 22584 11486 22636
rect 2774 22516 2780 22568
rect 2832 22556 2838 22568
rect 3053 22559 3111 22565
rect 3053 22556 3065 22559
rect 2832 22528 3065 22556
rect 2832 22516 2838 22528
rect 3053 22525 3065 22528
rect 3099 22525 3111 22559
rect 3053 22519 3111 22525
rect 9950 22516 9956 22568
rect 10008 22556 10014 22568
rect 10137 22559 10195 22565
rect 10137 22556 10149 22559
rect 10008 22528 10149 22556
rect 10008 22516 10014 22528
rect 10137 22525 10149 22528
rect 10183 22556 10195 22559
rect 10778 22556 10784 22568
rect 10183 22528 10784 22556
rect 10183 22525 10195 22528
rect 10137 22519 10195 22525
rect 10778 22516 10784 22528
rect 10836 22516 10842 22568
rect 15356 22559 15414 22565
rect 15356 22525 15368 22559
rect 15402 22556 15414 22559
rect 15838 22556 15844 22568
rect 15402 22528 15844 22556
rect 15402 22525 15414 22528
rect 15356 22519 15414 22525
rect 15838 22516 15844 22528
rect 15896 22516 15902 22568
rect 1394 22448 1400 22500
rect 1452 22488 1458 22500
rect 1673 22491 1731 22497
rect 1673 22488 1685 22491
rect 1452 22460 1685 22488
rect 1452 22448 1458 22460
rect 1673 22457 1685 22460
rect 1719 22488 1731 22491
rect 3326 22488 3332 22500
rect 1719 22460 3332 22488
rect 1719 22457 1731 22460
rect 1673 22451 1731 22457
rect 3326 22448 3332 22460
rect 3384 22448 3390 22500
rect 7009 22491 7067 22497
rect 7009 22457 7021 22491
rect 7055 22457 7067 22491
rect 7009 22451 7067 22457
rect 8941 22491 8999 22497
rect 8941 22457 8953 22491
rect 8987 22457 8999 22491
rect 8941 22451 8999 22457
rect 2498 22420 2504 22432
rect 2459 22392 2504 22420
rect 2498 22380 2504 22392
rect 2556 22380 2562 22432
rect 2774 22420 2780 22432
rect 2735 22392 2780 22420
rect 2774 22380 2780 22392
rect 2832 22380 2838 22432
rect 3234 22420 3240 22432
rect 3195 22392 3240 22420
rect 3234 22380 3240 22392
rect 3292 22380 3298 22432
rect 6273 22423 6331 22429
rect 6273 22389 6285 22423
rect 6319 22420 6331 22423
rect 6730 22420 6736 22432
rect 6319 22392 6736 22420
rect 6319 22389 6331 22392
rect 6273 22383 6331 22389
rect 6730 22380 6736 22392
rect 6788 22420 6794 22432
rect 7024 22420 7052 22451
rect 8662 22420 8668 22432
rect 6788 22392 7052 22420
rect 8623 22392 8668 22420
rect 6788 22380 6794 22392
rect 8662 22380 8668 22392
rect 8720 22420 8726 22432
rect 8956 22420 8984 22451
rect 8720 22392 8984 22420
rect 8720 22380 8726 22392
rect 9122 22380 9128 22432
rect 9180 22420 9186 22432
rect 9766 22420 9772 22432
rect 9180 22392 9772 22420
rect 9180 22380 9186 22392
rect 9766 22380 9772 22392
rect 9824 22380 9830 22432
rect 15427 22423 15485 22429
rect 15427 22389 15439 22423
rect 15473 22420 15485 22423
rect 15562 22420 15568 22432
rect 15473 22392 15568 22420
rect 15473 22389 15485 22392
rect 15427 22383 15485 22389
rect 15562 22380 15568 22392
rect 15620 22380 15626 22432
rect 15838 22420 15844 22432
rect 15799 22392 15844 22420
rect 15838 22380 15844 22392
rect 15896 22380 15902 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 2498 22176 2504 22228
rect 2556 22216 2562 22228
rect 3099 22219 3157 22225
rect 3099 22216 3111 22219
rect 2556 22188 3111 22216
rect 2556 22176 2562 22188
rect 3099 22185 3111 22188
rect 3145 22185 3157 22219
rect 3099 22179 3157 22185
rect 3326 22176 3332 22228
rect 3384 22216 3390 22228
rect 4203 22219 4261 22225
rect 4203 22216 4215 22219
rect 3384 22188 4215 22216
rect 3384 22176 3390 22188
rect 4203 22185 4215 22188
rect 4249 22185 4261 22219
rect 4203 22179 4261 22185
rect 6825 22219 6883 22225
rect 6825 22185 6837 22219
rect 6871 22216 6883 22219
rect 6914 22216 6920 22228
rect 6871 22188 6920 22216
rect 6871 22185 6883 22188
rect 6825 22179 6883 22185
rect 6914 22176 6920 22188
rect 6972 22176 6978 22228
rect 8846 22216 8852 22228
rect 8807 22188 8852 22216
rect 8846 22176 8852 22188
rect 8904 22176 8910 22228
rect 9861 22219 9919 22225
rect 9861 22185 9873 22219
rect 9907 22216 9919 22219
rect 10686 22216 10692 22228
rect 9907 22188 10692 22216
rect 9907 22185 9919 22188
rect 9861 22179 9919 22185
rect 10686 22176 10692 22188
rect 10744 22176 10750 22228
rect 1397 22083 1455 22089
rect 1397 22049 1409 22083
rect 1443 22080 1455 22083
rect 1486 22080 1492 22092
rect 1443 22052 1492 22080
rect 1443 22049 1455 22052
rect 1397 22043 1455 22049
rect 1486 22040 1492 22052
rect 1544 22040 1550 22092
rect 2961 22083 3019 22089
rect 2961 22049 2973 22083
rect 3007 22080 3019 22083
rect 3050 22080 3056 22092
rect 3007 22052 3056 22080
rect 3007 22049 3019 22052
rect 2961 22043 3019 22049
rect 3050 22040 3056 22052
rect 3108 22040 3114 22092
rect 4132 22083 4190 22089
rect 4132 22049 4144 22083
rect 4178 22080 4190 22083
rect 4430 22080 4436 22092
rect 4178 22052 4436 22080
rect 4178 22049 4190 22052
rect 4132 22043 4190 22049
rect 4430 22040 4436 22052
rect 4488 22040 4494 22092
rect 6730 22080 6736 22092
rect 6691 22052 6736 22080
rect 6730 22040 6736 22052
rect 6788 22040 6794 22092
rect 9674 22080 9680 22092
rect 9635 22052 9680 22080
rect 9674 22040 9680 22052
rect 9732 22040 9738 22092
rect 5074 22012 5080 22024
rect 5035 21984 5080 22012
rect 5074 21972 5080 21984
rect 5132 21972 5138 22024
rect 10318 22012 10324 22024
rect 10279 21984 10324 22012
rect 10318 21972 10324 21984
rect 10376 21972 10382 22024
rect 1535 21947 1593 21953
rect 1535 21913 1547 21947
rect 1581 21944 1593 21947
rect 1581 21916 1992 21944
rect 1581 21913 1593 21916
rect 1535 21907 1593 21913
rect 1964 21888 1992 21916
rect 1854 21876 1860 21888
rect 1815 21848 1860 21876
rect 1854 21836 1860 21848
rect 1912 21836 1918 21888
rect 1946 21836 1952 21888
rect 2004 21876 2010 21888
rect 2225 21879 2283 21885
rect 2225 21876 2237 21879
rect 2004 21848 2237 21876
rect 2004 21836 2010 21848
rect 2225 21845 2237 21848
rect 2271 21845 2283 21879
rect 2225 21839 2283 21845
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1486 21632 1492 21684
rect 1544 21672 1550 21684
rect 1581 21675 1639 21681
rect 1581 21672 1593 21675
rect 1544 21644 1593 21672
rect 1544 21632 1550 21644
rect 1581 21641 1593 21644
rect 1627 21641 1639 21675
rect 3234 21672 3240 21684
rect 3195 21644 3240 21672
rect 1581 21635 1639 21641
rect 3234 21632 3240 21644
rect 3292 21632 3298 21684
rect 4430 21672 4436 21684
rect 4391 21644 4436 21672
rect 4430 21632 4436 21644
rect 4488 21632 4494 21684
rect 9674 21672 9680 21684
rect 9635 21644 9680 21672
rect 9674 21632 9680 21644
rect 9732 21632 9738 21684
rect 9858 21632 9864 21684
rect 9916 21672 9922 21684
rect 10597 21675 10655 21681
rect 10597 21672 10609 21675
rect 9916 21644 10609 21672
rect 9916 21632 9922 21644
rect 10597 21641 10609 21644
rect 10643 21641 10655 21675
rect 10597 21635 10655 21641
rect 1946 21536 1952 21548
rect 1907 21508 1952 21536
rect 1946 21496 1952 21508
rect 2004 21496 2010 21548
rect 3050 21496 3056 21548
rect 3108 21536 3114 21548
rect 3789 21539 3847 21545
rect 3789 21536 3801 21539
rect 3108 21508 3801 21536
rect 3108 21496 3114 21508
rect 3789 21505 3801 21508
rect 3835 21505 3847 21539
rect 8662 21536 8668 21548
rect 8623 21508 8668 21536
rect 3789 21499 3847 21505
rect 8662 21496 8668 21508
rect 8720 21496 8726 21548
rect 5077 21471 5135 21477
rect 5077 21437 5089 21471
rect 5123 21437 5135 21471
rect 5077 21431 5135 21437
rect 8573 21471 8631 21477
rect 8573 21437 8585 21471
rect 8619 21468 8631 21471
rect 9122 21468 9128 21480
rect 8619 21440 9128 21468
rect 8619 21437 8631 21440
rect 8573 21431 8631 21437
rect 1946 21360 1952 21412
rect 2004 21400 2010 21412
rect 2041 21403 2099 21409
rect 2041 21400 2053 21403
rect 2004 21372 2053 21400
rect 2004 21360 2010 21372
rect 2041 21369 2053 21372
rect 2087 21369 2099 21403
rect 2041 21363 2099 21369
rect 2593 21403 2651 21409
rect 2593 21369 2605 21403
rect 2639 21400 2651 21403
rect 2682 21400 2688 21412
rect 2639 21372 2688 21400
rect 2639 21369 2651 21372
rect 2593 21363 2651 21369
rect 2682 21360 2688 21372
rect 2740 21360 2746 21412
rect 3510 21400 3516 21412
rect 3471 21372 3516 21400
rect 3510 21360 3516 21372
rect 3568 21360 3574 21412
rect 3605 21403 3663 21409
rect 3605 21369 3617 21403
rect 3651 21369 3663 21403
rect 4982 21400 4988 21412
rect 4943 21372 4988 21400
rect 3605 21363 3663 21369
rect 2961 21335 3019 21341
rect 2961 21301 2973 21335
rect 3007 21332 3019 21335
rect 3050 21332 3056 21344
rect 3007 21304 3056 21332
rect 3007 21301 3019 21304
rect 2961 21295 3019 21301
rect 3050 21292 3056 21304
rect 3108 21292 3114 21344
rect 3234 21292 3240 21344
rect 3292 21332 3298 21344
rect 3620 21332 3648 21363
rect 4982 21360 4988 21372
rect 5040 21360 5046 21412
rect 4890 21332 4896 21344
rect 3292 21304 3648 21332
rect 4851 21304 4896 21332
rect 3292 21292 3298 21304
rect 4890 21292 4896 21304
rect 4948 21332 4954 21344
rect 5092 21332 5120 21431
rect 9122 21428 9128 21440
rect 9180 21428 9186 21480
rect 10413 21471 10471 21477
rect 10413 21437 10425 21471
rect 10459 21468 10471 21471
rect 10459 21440 11100 21468
rect 10459 21437 10471 21440
rect 10413 21431 10471 21437
rect 11072 21344 11100 21440
rect 4948 21304 5120 21332
rect 6457 21335 6515 21341
rect 4948 21292 4954 21304
rect 6457 21301 6469 21335
rect 6503 21332 6515 21335
rect 6730 21332 6736 21344
rect 6503 21304 6736 21332
rect 6503 21301 6515 21304
rect 6457 21295 6515 21301
rect 6730 21292 6736 21304
rect 6788 21292 6794 21344
rect 11054 21332 11060 21344
rect 11015 21304 11060 21332
rect 11054 21292 11060 21304
rect 11112 21292 11118 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 3510 21128 3516 21140
rect 3471 21100 3516 21128
rect 3510 21088 3516 21100
rect 3568 21128 3574 21140
rect 4065 21131 4123 21137
rect 4065 21128 4077 21131
rect 3568 21100 4077 21128
rect 3568 21088 3574 21100
rect 4065 21097 4077 21100
rect 4111 21097 4123 21131
rect 4065 21091 4123 21097
rect 9674 21088 9680 21140
rect 9732 21128 9738 21140
rect 9815 21131 9873 21137
rect 9815 21128 9827 21131
rect 9732 21100 9827 21128
rect 9732 21088 9738 21100
rect 9815 21097 9827 21100
rect 9861 21097 9873 21131
rect 9815 21091 9873 21097
rect 2133 21063 2191 21069
rect 2133 21029 2145 21063
rect 2179 21060 2191 21063
rect 2314 21060 2320 21072
rect 2179 21032 2320 21060
rect 2179 21029 2191 21032
rect 2133 21023 2191 21029
rect 2314 21020 2320 21032
rect 2372 21020 2378 21072
rect 2682 21060 2688 21072
rect 2643 21032 2688 21060
rect 2682 21020 2688 21032
rect 2740 21020 2746 21072
rect 5350 21060 5356 21072
rect 5311 21032 5356 21060
rect 5350 21020 5356 21032
rect 5408 21020 5414 21072
rect 7558 20992 7564 21004
rect 7519 20964 7564 20992
rect 7558 20952 7564 20964
rect 7616 20952 7622 21004
rect 9214 20952 9220 21004
rect 9272 20992 9278 21004
rect 9712 20995 9770 21001
rect 9712 20992 9724 20995
rect 9272 20964 9724 20992
rect 9272 20952 9278 20964
rect 9712 20961 9724 20964
rect 9758 20961 9770 20995
rect 9712 20955 9770 20961
rect 2038 20924 2044 20936
rect 1999 20896 2044 20924
rect 2038 20884 2044 20896
rect 2096 20884 2102 20936
rect 5261 20927 5319 20933
rect 5261 20893 5273 20927
rect 5307 20893 5319 20927
rect 5534 20924 5540 20936
rect 5495 20896 5540 20924
rect 5261 20887 5319 20893
rect 5276 20856 5304 20887
rect 5534 20884 5540 20896
rect 5592 20884 5598 20936
rect 7282 20924 7288 20936
rect 7243 20896 7288 20924
rect 7282 20884 7288 20896
rect 7340 20884 7346 20936
rect 11422 20924 11428 20936
rect 11383 20896 11428 20924
rect 11422 20884 11428 20896
rect 11480 20884 11486 20936
rect 5994 20856 6000 20868
rect 5276 20828 6000 20856
rect 5994 20816 6000 20828
rect 6052 20816 6058 20868
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1535 20587 1593 20593
rect 1535 20553 1547 20587
rect 1581 20584 1593 20587
rect 2038 20584 2044 20596
rect 1581 20556 2044 20584
rect 1581 20553 1593 20556
rect 1535 20547 1593 20553
rect 2038 20544 2044 20556
rect 2096 20544 2102 20596
rect 5994 20584 6000 20596
rect 5955 20556 6000 20584
rect 5994 20544 6000 20556
rect 6052 20544 6058 20596
rect 9214 20584 9220 20596
rect 8772 20556 9220 20584
rect 8772 20528 8800 20556
rect 9214 20544 9220 20556
rect 9272 20544 9278 20596
rect 11054 20544 11060 20596
rect 11112 20584 11118 20596
rect 11379 20587 11437 20593
rect 11379 20584 11391 20587
rect 11112 20556 11391 20584
rect 11112 20544 11118 20556
rect 11379 20553 11391 20556
rect 11425 20553 11437 20587
rect 11379 20547 11437 20553
rect 12621 20587 12679 20593
rect 12621 20553 12633 20587
rect 12667 20584 12679 20587
rect 13906 20584 13912 20596
rect 12667 20556 13912 20584
rect 12667 20553 12679 20556
rect 12621 20547 12679 20553
rect 13906 20544 13912 20556
rect 13964 20544 13970 20596
rect 14093 20587 14151 20593
rect 14093 20553 14105 20587
rect 14139 20584 14151 20587
rect 22094 20584 22100 20596
rect 14139 20556 22100 20584
rect 14139 20553 14151 20556
rect 14093 20547 14151 20553
rect 4430 20476 4436 20528
rect 4488 20516 4494 20528
rect 5166 20516 5172 20528
rect 4488 20488 5172 20516
rect 4488 20476 4494 20488
rect 5166 20476 5172 20488
rect 5224 20476 5230 20528
rect 8754 20516 8760 20528
rect 8667 20488 8760 20516
rect 8754 20476 8760 20488
rect 8812 20476 8818 20528
rect 2682 20408 2688 20460
rect 2740 20448 2746 20460
rect 2961 20451 3019 20457
rect 2961 20448 2973 20451
rect 2740 20420 2973 20448
rect 2740 20408 2746 20420
rect 2961 20417 2973 20420
rect 3007 20417 3019 20451
rect 2961 20411 3019 20417
rect 3050 20408 3056 20460
rect 3108 20448 3114 20460
rect 3237 20451 3295 20457
rect 3237 20448 3249 20451
rect 3108 20420 3249 20448
rect 3108 20408 3114 20420
rect 3237 20417 3249 20420
rect 3283 20417 3295 20451
rect 4614 20448 4620 20460
rect 4527 20420 4620 20448
rect 3237 20411 3295 20417
rect 4614 20408 4620 20420
rect 4672 20448 4678 20460
rect 5074 20448 5080 20460
rect 4672 20420 5080 20448
rect 4672 20408 4678 20420
rect 5074 20408 5080 20420
rect 5132 20408 5138 20460
rect 1118 20340 1124 20392
rect 1176 20380 1182 20392
rect 1432 20383 1490 20389
rect 1432 20380 1444 20383
rect 1176 20352 1444 20380
rect 1176 20340 1182 20352
rect 1432 20349 1444 20352
rect 1478 20380 1490 20383
rect 1857 20383 1915 20389
rect 1857 20380 1869 20383
rect 1478 20352 1869 20380
rect 1478 20349 1490 20352
rect 1432 20343 1490 20349
rect 1857 20349 1869 20352
rect 1903 20349 1915 20383
rect 9582 20380 9588 20392
rect 9495 20352 9588 20380
rect 1857 20343 1915 20349
rect 9582 20340 9588 20352
rect 9640 20380 9646 20392
rect 9769 20383 9827 20389
rect 9769 20380 9781 20383
rect 9640 20352 9781 20380
rect 9640 20340 9646 20352
rect 9769 20349 9781 20352
rect 9815 20349 9827 20383
rect 9769 20343 9827 20349
rect 11308 20383 11366 20389
rect 11308 20349 11320 20383
rect 11354 20380 11366 20383
rect 11354 20352 11836 20380
rect 11354 20349 11366 20352
rect 11308 20343 11366 20349
rect 2774 20312 2780 20324
rect 2687 20284 2780 20312
rect 2774 20272 2780 20284
rect 2832 20312 2838 20324
rect 3050 20312 3056 20324
rect 2832 20284 3056 20312
rect 2832 20272 2838 20284
rect 3050 20272 3056 20284
rect 3108 20272 3114 20324
rect 4709 20315 4767 20321
rect 4709 20281 4721 20315
rect 4755 20312 4767 20315
rect 4982 20312 4988 20324
rect 4755 20284 4988 20312
rect 4755 20281 4767 20284
rect 4709 20275 4767 20281
rect 2314 20244 2320 20256
rect 2275 20216 2320 20244
rect 2314 20204 2320 20216
rect 2372 20204 2378 20256
rect 4433 20247 4491 20253
rect 4433 20213 4445 20247
rect 4479 20244 4491 20247
rect 4724 20244 4752 20275
rect 4982 20272 4988 20284
rect 5040 20272 5046 20324
rect 5350 20272 5356 20324
rect 5408 20312 5414 20324
rect 5629 20315 5687 20321
rect 5629 20312 5641 20315
rect 5408 20284 5641 20312
rect 5408 20272 5414 20284
rect 5629 20281 5641 20284
rect 5675 20312 5687 20315
rect 5994 20312 6000 20324
rect 5675 20284 6000 20312
rect 5675 20281 5687 20284
rect 5629 20275 5687 20281
rect 5994 20272 6000 20284
rect 6052 20272 6058 20324
rect 7101 20315 7159 20321
rect 7101 20281 7113 20315
rect 7147 20312 7159 20315
rect 7653 20315 7711 20321
rect 7653 20312 7665 20315
rect 7147 20284 7665 20312
rect 7147 20281 7159 20284
rect 7101 20275 7159 20281
rect 7653 20281 7665 20284
rect 7699 20312 7711 20315
rect 8205 20315 8263 20321
rect 8205 20312 8217 20315
rect 7699 20284 8217 20312
rect 7699 20281 7711 20284
rect 7653 20275 7711 20281
rect 8205 20281 8217 20284
rect 8251 20281 8263 20315
rect 8205 20275 8263 20281
rect 8297 20315 8355 20321
rect 8297 20281 8309 20315
rect 8343 20312 8355 20315
rect 9677 20315 9735 20321
rect 9677 20312 9689 20315
rect 8343 20284 9689 20312
rect 8343 20281 8355 20284
rect 8297 20275 8355 20281
rect 9677 20281 9689 20284
rect 9723 20281 9735 20315
rect 9677 20275 9735 20281
rect 4479 20216 4752 20244
rect 8021 20247 8079 20253
rect 4479 20213 4491 20216
rect 4433 20207 4491 20213
rect 8021 20213 8033 20247
rect 8067 20244 8079 20247
rect 8312 20244 8340 20275
rect 11808 20256 11836 20352
rect 12342 20340 12348 20392
rect 12400 20380 12406 20392
rect 12437 20383 12495 20389
rect 12437 20380 12449 20383
rect 12400 20352 12449 20380
rect 12400 20340 12406 20352
rect 12437 20349 12449 20352
rect 12483 20380 12495 20383
rect 12989 20383 13047 20389
rect 12989 20380 13001 20383
rect 12483 20352 13001 20380
rect 12483 20349 12495 20352
rect 12437 20343 12495 20349
rect 12989 20349 13001 20352
rect 13035 20349 13047 20383
rect 12989 20343 13047 20349
rect 13608 20383 13666 20389
rect 13608 20349 13620 20383
rect 13654 20380 13666 20383
rect 14108 20380 14136 20547
rect 22094 20544 22100 20556
rect 22152 20544 22158 20596
rect 25130 20584 25136 20596
rect 25091 20556 25136 20584
rect 25130 20544 25136 20556
rect 25188 20544 25194 20596
rect 13654 20352 14136 20380
rect 24648 20383 24706 20389
rect 13654 20349 13666 20352
rect 13608 20343 13666 20349
rect 24648 20349 24660 20383
rect 24694 20380 24706 20383
rect 25130 20380 25136 20392
rect 24694 20352 25136 20380
rect 24694 20349 24706 20352
rect 24648 20343 24706 20349
rect 25130 20340 25136 20352
rect 25188 20340 25194 20392
rect 11790 20244 11796 20256
rect 8067 20216 8340 20244
rect 11751 20216 11796 20244
rect 8067 20213 8079 20216
rect 8021 20207 8079 20213
rect 11790 20204 11796 20216
rect 11848 20204 11854 20256
rect 12894 20204 12900 20256
rect 12952 20244 12958 20256
rect 13679 20247 13737 20253
rect 13679 20244 13691 20247
rect 12952 20216 13691 20244
rect 12952 20204 12958 20216
rect 13679 20213 13691 20216
rect 13725 20213 13737 20247
rect 13679 20207 13737 20213
rect 17126 20204 17132 20256
rect 17184 20244 17190 20256
rect 24719 20247 24777 20253
rect 24719 20244 24731 20247
rect 17184 20216 24731 20244
rect 17184 20204 17190 20216
rect 24719 20213 24731 20216
rect 24765 20213 24777 20247
rect 24719 20207 24777 20213
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 1857 20043 1915 20049
rect 1857 20009 1869 20043
rect 1903 20040 1915 20043
rect 2038 20040 2044 20052
rect 1903 20012 2044 20040
rect 1903 20009 1915 20012
rect 1857 20003 1915 20009
rect 2038 20000 2044 20012
rect 2096 20000 2102 20052
rect 2682 20000 2688 20052
rect 2740 20040 2746 20052
rect 2961 20043 3019 20049
rect 2961 20040 2973 20043
rect 2740 20012 2973 20040
rect 2740 20000 2746 20012
rect 2961 20009 2973 20012
rect 3007 20009 3019 20043
rect 4614 20040 4620 20052
rect 4575 20012 4620 20040
rect 2961 20003 3019 20009
rect 4614 20000 4620 20012
rect 4672 20000 4678 20052
rect 7558 20040 7564 20052
rect 7519 20012 7564 20040
rect 7558 20000 7564 20012
rect 7616 20000 7622 20052
rect 1946 19972 1952 19984
rect 1907 19944 1952 19972
rect 1946 19932 1952 19944
rect 2004 19932 2010 19984
rect 4982 19972 4988 19984
rect 4943 19944 4988 19972
rect 4982 19932 4988 19944
rect 5040 19932 5046 19984
rect 5166 19932 5172 19984
rect 5224 19972 5230 19984
rect 5537 19975 5595 19981
rect 5537 19972 5549 19975
rect 5224 19944 5549 19972
rect 5224 19932 5230 19944
rect 5537 19941 5549 19944
rect 5583 19941 5595 19975
rect 5537 19935 5595 19941
rect 6546 19932 6552 19984
rect 6604 19972 6610 19984
rect 6641 19975 6699 19981
rect 6641 19972 6653 19975
rect 6604 19944 6653 19972
rect 6604 19932 6610 19944
rect 6641 19941 6653 19944
rect 6687 19972 6699 19975
rect 7282 19972 7288 19984
rect 6687 19944 7288 19972
rect 6687 19941 6699 19944
rect 6641 19935 6699 19941
rect 7282 19932 7288 19944
rect 7340 19932 7346 19984
rect 8202 19972 8208 19984
rect 8163 19944 8208 19972
rect 8202 19932 8208 19944
rect 8260 19932 8266 19984
rect 8754 19972 8760 19984
rect 8715 19944 8760 19972
rect 8754 19932 8760 19944
rect 8812 19932 8818 19984
rect 9766 19932 9772 19984
rect 9824 19972 9830 19984
rect 9861 19975 9919 19981
rect 9861 19972 9873 19975
rect 9824 19944 9873 19972
rect 9824 19932 9830 19944
rect 9861 19941 9873 19944
rect 9907 19941 9919 19975
rect 9861 19935 9919 19941
rect 11422 19932 11428 19984
rect 11480 19972 11486 19984
rect 11701 19975 11759 19981
rect 11701 19972 11713 19975
rect 11480 19944 11713 19972
rect 11480 19932 11486 19944
rect 11701 19941 11713 19944
rect 11747 19941 11759 19975
rect 11701 19935 11759 19941
rect 11793 19975 11851 19981
rect 11793 19941 11805 19975
rect 11839 19972 11851 19975
rect 11882 19972 11888 19984
rect 11839 19944 11888 19972
rect 11839 19941 11851 19944
rect 11793 19935 11851 19941
rect 11882 19932 11888 19944
rect 11940 19972 11946 19984
rect 13173 19975 13231 19981
rect 13173 19972 13185 19975
rect 11940 19944 13185 19972
rect 11940 19932 11946 19944
rect 13173 19941 13185 19944
rect 13219 19941 13231 19975
rect 13173 19935 13231 19941
rect 2314 19904 2320 19916
rect 2275 19876 2320 19904
rect 2314 19864 2320 19876
rect 2372 19864 2378 19916
rect 13446 19904 13452 19916
rect 13407 19876 13452 19904
rect 13446 19864 13452 19876
rect 13504 19864 13510 19916
rect 4893 19839 4951 19845
rect 4893 19805 4905 19839
rect 4939 19836 4951 19839
rect 5534 19836 5540 19848
rect 4939 19808 5540 19836
rect 4939 19805 4951 19808
rect 4893 19799 4951 19805
rect 5534 19796 5540 19808
rect 5592 19796 5598 19848
rect 6086 19796 6092 19848
rect 6144 19836 6150 19848
rect 6549 19839 6607 19845
rect 6549 19836 6561 19839
rect 6144 19808 6561 19836
rect 6144 19796 6150 19808
rect 6549 19805 6561 19808
rect 6595 19805 6607 19839
rect 6549 19799 6607 19805
rect 7193 19839 7251 19845
rect 7193 19805 7205 19839
rect 7239 19836 7251 19839
rect 8113 19839 8171 19845
rect 8113 19836 8125 19839
rect 7239 19808 8125 19836
rect 7239 19805 7251 19808
rect 7193 19799 7251 19805
rect 8113 19805 8125 19808
rect 8159 19805 8171 19839
rect 8113 19799 8171 19805
rect 9769 19839 9827 19845
rect 9769 19805 9781 19839
rect 9815 19836 9827 19839
rect 10870 19836 10876 19848
rect 9815 19808 10876 19836
rect 9815 19805 9827 19808
rect 9769 19799 9827 19805
rect 8128 19768 8156 19799
rect 10870 19796 10876 19808
rect 10928 19796 10934 19848
rect 11790 19796 11796 19848
rect 11848 19836 11854 19848
rect 12345 19839 12403 19845
rect 12345 19836 12357 19839
rect 11848 19808 12357 19836
rect 11848 19796 11854 19808
rect 12345 19805 12357 19808
rect 12391 19836 12403 19839
rect 12802 19836 12808 19848
rect 12391 19808 12808 19836
rect 12391 19805 12403 19808
rect 12345 19799 12403 19805
rect 12802 19796 12808 19808
rect 12860 19796 12866 19848
rect 8478 19768 8484 19780
rect 8128 19740 8484 19768
rect 8478 19728 8484 19740
rect 8536 19768 8542 19780
rect 10321 19771 10379 19777
rect 10321 19768 10333 19771
rect 8536 19740 10333 19768
rect 8536 19728 8542 19740
rect 10321 19737 10333 19740
rect 10367 19737 10379 19771
rect 10321 19731 10379 19737
rect 7834 19700 7840 19712
rect 7795 19672 7840 19700
rect 7834 19660 7840 19672
rect 7892 19660 7898 19712
rect 12618 19700 12624 19712
rect 12579 19672 12624 19700
rect 12618 19660 12624 19672
rect 12676 19660 12682 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 5534 19456 5540 19508
rect 5592 19496 5598 19508
rect 5629 19499 5687 19505
rect 5629 19496 5641 19499
rect 5592 19468 5641 19496
rect 5592 19456 5598 19468
rect 5629 19465 5641 19468
rect 5675 19465 5687 19499
rect 6546 19496 6552 19508
rect 6507 19468 6552 19496
rect 5629 19459 5687 19465
rect 6546 19456 6552 19468
rect 6604 19456 6610 19508
rect 8202 19456 8208 19508
rect 8260 19496 8266 19508
rect 8389 19499 8447 19505
rect 8389 19496 8401 19499
rect 8260 19468 8401 19496
rect 8260 19456 8266 19468
rect 8389 19465 8401 19468
rect 8435 19496 8447 19499
rect 8757 19499 8815 19505
rect 8757 19496 8769 19499
rect 8435 19468 8769 19496
rect 8435 19465 8447 19468
rect 8389 19459 8447 19465
rect 8757 19465 8769 19468
rect 8803 19496 8815 19499
rect 9582 19496 9588 19508
rect 8803 19468 9588 19496
rect 8803 19465 8815 19468
rect 8757 19459 8815 19465
rect 9582 19456 9588 19468
rect 9640 19456 9646 19508
rect 11422 19456 11428 19508
rect 11480 19496 11486 19508
rect 12161 19499 12219 19505
rect 12161 19496 12173 19499
rect 11480 19468 12173 19496
rect 11480 19456 11486 19468
rect 12161 19465 12173 19468
rect 12207 19465 12219 19499
rect 13446 19496 13452 19508
rect 13407 19468 13452 19496
rect 12161 19459 12219 19465
rect 13446 19456 13452 19468
rect 13504 19456 13510 19508
rect 4893 19431 4951 19437
rect 4893 19397 4905 19431
rect 4939 19428 4951 19431
rect 5552 19428 5580 19456
rect 11882 19428 11888 19440
rect 4939 19400 5580 19428
rect 11843 19400 11888 19428
rect 4939 19397 4951 19400
rect 4893 19391 4951 19397
rect 11882 19388 11888 19400
rect 11940 19388 11946 19440
rect 7469 19363 7527 19369
rect 7469 19329 7481 19363
rect 7515 19360 7527 19363
rect 7834 19360 7840 19372
rect 7515 19332 7840 19360
rect 7515 19329 7527 19332
rect 7469 19323 7527 19329
rect 7834 19320 7840 19332
rect 7892 19320 7898 19372
rect 10870 19360 10876 19372
rect 10831 19332 10876 19360
rect 10870 19320 10876 19332
rect 10928 19320 10934 19372
rect 11471 19363 11529 19369
rect 11471 19329 11483 19363
rect 11517 19360 11529 19363
rect 12342 19360 12348 19372
rect 11517 19332 12348 19360
rect 11517 19329 11529 19332
rect 11471 19323 11529 19329
rect 12342 19320 12348 19332
rect 12400 19320 12406 19372
rect 12529 19363 12587 19369
rect 12529 19329 12541 19363
rect 12575 19360 12587 19363
rect 12618 19360 12624 19372
rect 12575 19332 12624 19360
rect 12575 19329 12587 19332
rect 12529 19323 12587 19329
rect 12618 19320 12624 19332
rect 12676 19320 12682 19372
rect 12802 19360 12808 19372
rect 12763 19332 12808 19360
rect 12802 19320 12808 19332
rect 12860 19320 12866 19372
rect 2593 19295 2651 19301
rect 2593 19261 2605 19295
rect 2639 19292 2651 19295
rect 3326 19292 3332 19304
rect 2639 19264 3332 19292
rect 2639 19261 2651 19264
rect 2593 19255 2651 19261
rect 3326 19252 3332 19264
rect 3384 19252 3390 19304
rect 3421 19295 3479 19301
rect 3421 19261 3433 19295
rect 3467 19292 3479 19295
rect 4065 19295 4123 19301
rect 4065 19292 4077 19295
rect 3467 19264 4077 19292
rect 3467 19261 3479 19264
rect 3421 19255 3479 19261
rect 4065 19261 4077 19264
rect 4111 19292 4123 19295
rect 9309 19295 9367 19301
rect 4111 19264 4200 19292
rect 4111 19261 4123 19264
rect 4065 19255 4123 19261
rect 2041 19159 2099 19165
rect 2041 19125 2053 19159
rect 2087 19156 2099 19159
rect 2314 19156 2320 19168
rect 2087 19128 2320 19156
rect 2087 19125 2099 19128
rect 2041 19119 2099 19125
rect 2314 19116 2320 19128
rect 2372 19156 2378 19168
rect 3234 19156 3240 19168
rect 2372 19128 3240 19156
rect 2372 19116 2378 19128
rect 3234 19116 3240 19128
rect 3292 19116 3298 19168
rect 4172 19156 4200 19264
rect 9309 19261 9321 19295
rect 9355 19292 9367 19295
rect 9858 19292 9864 19304
rect 9355 19264 9864 19292
rect 9355 19261 9367 19264
rect 9309 19255 9367 19261
rect 9858 19252 9864 19264
rect 9916 19252 9922 19304
rect 10778 19252 10784 19304
rect 10836 19292 10842 19304
rect 11149 19295 11207 19301
rect 11149 19292 11161 19295
rect 10836 19264 11161 19292
rect 10836 19252 10842 19264
rect 11149 19261 11161 19264
rect 11195 19292 11207 19295
rect 11368 19295 11426 19301
rect 11368 19292 11380 19295
rect 11195 19264 11380 19292
rect 11195 19261 11207 19264
rect 11149 19255 11207 19261
rect 11368 19261 11380 19264
rect 11414 19261 11426 19295
rect 11368 19255 11426 19261
rect 4338 19224 4344 19236
rect 4299 19196 4344 19224
rect 4338 19184 4344 19196
rect 4396 19184 4402 19236
rect 4433 19227 4491 19233
rect 4433 19193 4445 19227
rect 4479 19193 4491 19227
rect 4433 19187 4491 19193
rect 4448 19156 4476 19187
rect 5258 19184 5264 19236
rect 5316 19224 5322 19236
rect 7285 19227 7343 19233
rect 7285 19224 7297 19227
rect 5316 19196 7297 19224
rect 5316 19184 5322 19196
rect 7285 19193 7297 19196
rect 7331 19224 7343 19227
rect 7466 19224 7472 19236
rect 7331 19196 7472 19224
rect 7331 19193 7343 19196
rect 7285 19187 7343 19193
rect 7466 19184 7472 19196
rect 7524 19224 7530 19236
rect 7790 19227 7848 19233
rect 7790 19224 7802 19227
rect 7524 19196 7802 19224
rect 7524 19184 7530 19196
rect 7790 19193 7802 19196
rect 7836 19193 7848 19227
rect 7790 19187 7848 19193
rect 12621 19227 12679 19233
rect 12621 19193 12633 19227
rect 12667 19193 12679 19227
rect 12621 19187 12679 19193
rect 4172 19128 4476 19156
rect 4982 19116 4988 19168
rect 5040 19156 5046 19168
rect 5353 19159 5411 19165
rect 5353 19156 5365 19159
rect 5040 19128 5365 19156
rect 5040 19116 5046 19128
rect 5353 19125 5365 19128
rect 5399 19156 5411 19159
rect 5902 19156 5908 19168
rect 5399 19128 5908 19156
rect 5399 19125 5411 19128
rect 5353 19119 5411 19125
rect 5902 19116 5908 19128
rect 5960 19116 5966 19168
rect 6086 19156 6092 19168
rect 6047 19128 6092 19156
rect 6086 19116 6092 19128
rect 6144 19116 6150 19168
rect 7558 19116 7564 19168
rect 7616 19156 7622 19168
rect 9585 19159 9643 19165
rect 9585 19156 9597 19159
rect 7616 19128 9597 19156
rect 7616 19116 7622 19128
rect 9585 19125 9597 19128
rect 9631 19156 9643 19159
rect 9766 19156 9772 19168
rect 9631 19128 9772 19156
rect 9631 19125 9643 19128
rect 9585 19119 9643 19125
rect 9766 19116 9772 19128
rect 9824 19116 9830 19168
rect 10042 19156 10048 19168
rect 10003 19128 10048 19156
rect 10042 19116 10048 19128
rect 10100 19116 10106 19168
rect 12526 19116 12532 19168
rect 12584 19156 12590 19168
rect 12636 19156 12664 19187
rect 13446 19156 13452 19168
rect 12584 19128 13452 19156
rect 12584 19116 12590 19128
rect 13446 19116 13452 19128
rect 13504 19116 13510 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 4338 18952 4344 18964
rect 4299 18924 4344 18952
rect 4338 18912 4344 18924
rect 4396 18912 4402 18964
rect 5258 18912 5264 18964
rect 5316 18952 5322 18964
rect 5353 18955 5411 18961
rect 5353 18952 5365 18955
rect 5316 18924 5365 18952
rect 5316 18912 5322 18924
rect 5353 18921 5365 18924
rect 5399 18921 5411 18955
rect 5902 18952 5908 18964
rect 5863 18924 5908 18952
rect 5353 18915 5411 18921
rect 5902 18912 5908 18924
rect 5960 18912 5966 18964
rect 7466 18912 7472 18964
rect 7524 18952 7530 18964
rect 7561 18955 7619 18961
rect 7561 18952 7573 18955
rect 7524 18924 7573 18952
rect 7524 18912 7530 18924
rect 7561 18921 7573 18924
rect 7607 18921 7619 18955
rect 7561 18915 7619 18921
rect 7650 18912 7656 18964
rect 7708 18952 7714 18964
rect 8113 18955 8171 18961
rect 8113 18952 8125 18955
rect 7708 18924 8125 18952
rect 7708 18912 7714 18924
rect 8113 18921 8125 18924
rect 8159 18921 8171 18955
rect 8478 18952 8484 18964
rect 8439 18924 8484 18952
rect 8113 18915 8171 18921
rect 8478 18912 8484 18924
rect 8536 18912 8542 18964
rect 11146 18912 11152 18964
rect 11204 18952 11210 18964
rect 11425 18955 11483 18961
rect 11425 18952 11437 18955
rect 11204 18924 11437 18952
rect 11204 18912 11210 18924
rect 11425 18921 11437 18924
rect 11471 18921 11483 18955
rect 11425 18915 11483 18921
rect 11977 18955 12035 18961
rect 11977 18921 11989 18955
rect 12023 18952 12035 18955
rect 12526 18952 12532 18964
rect 12023 18924 12532 18952
rect 12023 18921 12035 18924
rect 11977 18915 12035 18921
rect 12526 18912 12532 18924
rect 12584 18912 12590 18964
rect 12894 18884 12900 18896
rect 12855 18856 12900 18884
rect 12894 18844 12900 18856
rect 12952 18844 12958 18896
rect 12986 18844 12992 18896
rect 13044 18884 13050 18896
rect 13044 18856 13089 18884
rect 13044 18844 13050 18856
rect 1394 18816 1400 18828
rect 1355 18788 1400 18816
rect 1394 18776 1400 18788
rect 1452 18776 1458 18828
rect 2682 18816 2688 18828
rect 2643 18788 2688 18816
rect 2682 18776 2688 18788
rect 2740 18776 2746 18828
rect 2866 18816 2872 18828
rect 2827 18788 2872 18816
rect 2866 18776 2872 18788
rect 2924 18776 2930 18828
rect 3326 18776 3332 18828
rect 3384 18816 3390 18828
rect 5994 18816 6000 18828
rect 3384 18788 6000 18816
rect 3384 18776 3390 18788
rect 5994 18776 6000 18788
rect 6052 18776 6058 18828
rect 3142 18748 3148 18760
rect 3103 18720 3148 18748
rect 3142 18708 3148 18720
rect 3200 18708 3206 18760
rect 4985 18751 5043 18757
rect 4985 18717 4997 18751
rect 5031 18748 5043 18751
rect 5350 18748 5356 18760
rect 5031 18720 5356 18748
rect 5031 18717 5043 18720
rect 4985 18711 5043 18717
rect 5350 18708 5356 18720
rect 5408 18708 5414 18760
rect 7190 18748 7196 18760
rect 7151 18720 7196 18748
rect 7190 18708 7196 18720
rect 7248 18708 7254 18760
rect 9950 18748 9956 18760
rect 9911 18720 9956 18748
rect 9950 18708 9956 18720
rect 10008 18708 10014 18760
rect 11057 18751 11115 18757
rect 11057 18717 11069 18751
rect 11103 18748 11115 18751
rect 11422 18748 11428 18760
rect 11103 18720 11428 18748
rect 11103 18717 11115 18720
rect 11057 18711 11115 18717
rect 11422 18708 11428 18720
rect 11480 18708 11486 18760
rect 13173 18751 13231 18757
rect 13173 18717 13185 18751
rect 13219 18717 13231 18751
rect 13173 18711 13231 18717
rect 12618 18640 12624 18692
rect 12676 18680 12682 18692
rect 13188 18680 13216 18711
rect 12676 18652 13216 18680
rect 12676 18640 12682 18652
rect 1535 18615 1593 18621
rect 1535 18581 1547 18615
rect 1581 18612 1593 18615
rect 2130 18612 2136 18624
rect 1581 18584 2136 18612
rect 1581 18581 1593 18584
rect 1535 18575 1593 18581
rect 2130 18572 2136 18584
rect 2188 18572 2194 18624
rect 3326 18572 3332 18624
rect 3384 18612 3390 18624
rect 4338 18612 4344 18624
rect 3384 18584 4344 18612
rect 3384 18572 3390 18584
rect 4338 18572 4344 18584
rect 4396 18572 4402 18624
rect 7006 18612 7012 18624
rect 6967 18584 7012 18612
rect 7006 18572 7012 18584
rect 7064 18572 7070 18624
rect 8846 18612 8852 18624
rect 8807 18584 8852 18612
rect 8846 18572 8852 18584
rect 8904 18572 8910 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 106 18368 112 18420
rect 164 18408 170 18420
rect 1394 18408 1400 18420
rect 164 18380 1400 18408
rect 164 18368 170 18380
rect 1394 18368 1400 18380
rect 1452 18408 1458 18420
rect 1581 18411 1639 18417
rect 1581 18408 1593 18411
rect 1452 18380 1593 18408
rect 1452 18368 1458 18380
rect 1581 18377 1593 18380
rect 1627 18377 1639 18411
rect 1581 18371 1639 18377
rect 2682 18368 2688 18420
rect 2740 18408 2746 18420
rect 3513 18411 3571 18417
rect 3513 18408 3525 18411
rect 2740 18380 3525 18408
rect 2740 18368 2746 18380
rect 3513 18377 3525 18380
rect 3559 18408 3571 18411
rect 3970 18408 3976 18420
rect 3559 18380 3976 18408
rect 3559 18377 3571 18380
rect 3513 18371 3571 18377
rect 3970 18368 3976 18380
rect 4028 18368 4034 18420
rect 5905 18411 5963 18417
rect 5905 18377 5917 18411
rect 5951 18408 5963 18411
rect 5994 18408 6000 18420
rect 5951 18380 6000 18408
rect 5951 18377 5963 18380
rect 5905 18371 5963 18377
rect 5994 18368 6000 18380
rect 6052 18368 6058 18420
rect 7466 18368 7472 18420
rect 7524 18408 7530 18420
rect 7929 18411 7987 18417
rect 7929 18408 7941 18411
rect 7524 18380 7941 18408
rect 7524 18368 7530 18380
rect 7929 18377 7941 18380
rect 7975 18377 7987 18411
rect 8846 18408 8852 18420
rect 7929 18371 7987 18377
rect 8680 18380 8852 18408
rect 3234 18340 3240 18352
rect 3195 18312 3240 18340
rect 3234 18300 3240 18312
rect 3292 18300 3298 18352
rect 3789 18343 3847 18349
rect 3789 18309 3801 18343
rect 3835 18340 3847 18343
rect 3835 18312 8248 18340
rect 3835 18309 3847 18312
rect 3789 18303 3847 18309
rect 3142 18232 3148 18284
rect 3200 18272 3206 18284
rect 7653 18275 7711 18281
rect 3200 18244 5028 18272
rect 3200 18232 3206 18244
rect 2314 18204 2320 18216
rect 2275 18176 2320 18204
rect 2314 18164 2320 18176
rect 2372 18164 2378 18216
rect 2866 18164 2872 18216
rect 2924 18204 2930 18216
rect 3789 18207 3847 18213
rect 3789 18204 3801 18207
rect 2924 18176 3801 18204
rect 2924 18164 2930 18176
rect 3789 18173 3801 18176
rect 3835 18204 3847 18207
rect 3881 18207 3939 18213
rect 3881 18204 3893 18207
rect 3835 18176 3893 18204
rect 3835 18173 3847 18176
rect 3789 18167 3847 18173
rect 3881 18173 3893 18176
rect 3927 18173 3939 18207
rect 3881 18167 3939 18173
rect 4062 18164 4068 18216
rect 4120 18204 4126 18216
rect 5000 18213 5028 18244
rect 7653 18241 7665 18275
rect 7699 18272 7711 18275
rect 7834 18272 7840 18284
rect 7699 18244 7840 18272
rect 7699 18241 7711 18244
rect 7653 18235 7711 18241
rect 7834 18232 7840 18244
rect 7892 18232 7898 18284
rect 4985 18207 5043 18213
rect 4120 18176 4936 18204
rect 4120 18164 4126 18176
rect 2225 18139 2283 18145
rect 2225 18105 2237 18139
rect 2271 18136 2283 18139
rect 2679 18139 2737 18145
rect 2679 18136 2691 18139
rect 2271 18108 2691 18136
rect 2271 18105 2283 18108
rect 2225 18099 2283 18105
rect 2679 18105 2691 18108
rect 2725 18136 2737 18139
rect 4246 18136 4252 18148
rect 2725 18108 4252 18136
rect 2725 18105 2737 18108
rect 2679 18099 2737 18105
rect 4246 18096 4252 18108
rect 4304 18136 4310 18148
rect 4433 18139 4491 18145
rect 4433 18136 4445 18139
rect 4304 18108 4445 18136
rect 4304 18096 4310 18108
rect 4433 18105 4445 18108
rect 4479 18136 4491 18139
rect 4801 18139 4859 18145
rect 4801 18136 4813 18139
rect 4479 18108 4813 18136
rect 4479 18105 4491 18108
rect 4433 18099 4491 18105
rect 4801 18105 4813 18108
rect 4847 18105 4859 18139
rect 4908 18136 4936 18176
rect 4985 18173 4997 18207
rect 5031 18204 5043 18207
rect 5074 18204 5080 18216
rect 5031 18176 5080 18204
rect 5031 18173 5043 18176
rect 4985 18167 5043 18173
rect 5074 18164 5080 18176
rect 5132 18164 5138 18216
rect 6641 18207 6699 18213
rect 6641 18204 6653 18207
rect 5184 18176 6653 18204
rect 5184 18136 5212 18176
rect 6641 18173 6653 18176
rect 6687 18204 6699 18207
rect 6914 18204 6920 18216
rect 6687 18176 6920 18204
rect 6687 18173 6699 18176
rect 6641 18167 6699 18173
rect 6914 18164 6920 18176
rect 6972 18164 6978 18216
rect 7006 18164 7012 18216
rect 7064 18204 7070 18216
rect 7377 18207 7435 18213
rect 7377 18204 7389 18207
rect 7064 18176 7389 18204
rect 7064 18164 7070 18176
rect 7377 18173 7389 18176
rect 7423 18173 7435 18207
rect 7377 18167 7435 18173
rect 4908 18108 5212 18136
rect 4801 18099 4859 18105
rect 3970 18028 3976 18080
rect 4028 18068 4034 18080
rect 4338 18068 4344 18080
rect 4028 18040 4344 18068
rect 4028 18028 4034 18040
rect 4338 18028 4344 18040
rect 4396 18028 4402 18080
rect 4816 18068 4844 18099
rect 5258 18068 5264 18080
rect 4816 18040 5264 18068
rect 5258 18028 5264 18040
rect 5316 18068 5322 18080
rect 5353 18071 5411 18077
rect 5353 18068 5365 18071
rect 5316 18040 5365 18068
rect 5316 18028 5322 18040
rect 5353 18037 5365 18040
rect 5399 18037 5411 18071
rect 8220 18068 8248 18312
rect 8573 18275 8631 18281
rect 8573 18241 8585 18275
rect 8619 18272 8631 18275
rect 8680 18272 8708 18380
rect 8846 18368 8852 18380
rect 8904 18368 8910 18420
rect 9953 18411 10011 18417
rect 9953 18377 9965 18411
rect 9999 18408 10011 18411
rect 10042 18408 10048 18420
rect 9999 18380 10048 18408
rect 9999 18377 10011 18380
rect 9953 18371 10011 18377
rect 10042 18368 10048 18380
rect 10100 18368 10106 18420
rect 11146 18408 11152 18420
rect 11107 18380 11152 18408
rect 11146 18368 11152 18380
rect 11204 18368 11210 18420
rect 12986 18368 12992 18420
rect 13044 18408 13050 18420
rect 13449 18411 13507 18417
rect 13449 18408 13461 18411
rect 13044 18380 13461 18408
rect 13044 18368 13050 18380
rect 13449 18377 13461 18380
rect 13495 18377 13507 18411
rect 13449 18371 13507 18377
rect 8846 18272 8852 18284
rect 8619 18244 8708 18272
rect 8807 18244 8852 18272
rect 8619 18241 8631 18244
rect 8573 18235 8631 18241
rect 8846 18232 8852 18244
rect 8904 18232 8910 18284
rect 9585 18275 9643 18281
rect 9585 18241 9597 18275
rect 9631 18272 9643 18275
rect 9950 18272 9956 18284
rect 9631 18244 9956 18272
rect 9631 18241 9643 18244
rect 9585 18235 9643 18241
rect 9950 18232 9956 18244
rect 10008 18272 10014 18284
rect 10137 18275 10195 18281
rect 10137 18272 10149 18275
rect 10008 18244 10149 18272
rect 10008 18232 10014 18244
rect 10137 18241 10149 18244
rect 10183 18241 10195 18275
rect 10137 18235 10195 18241
rect 12618 18232 12624 18284
rect 12676 18272 12682 18284
rect 12805 18275 12863 18281
rect 12805 18272 12817 18275
rect 12676 18244 12817 18272
rect 12676 18232 12682 18244
rect 12805 18241 12817 18244
rect 12851 18241 12863 18275
rect 12805 18235 12863 18241
rect 8389 18139 8447 18145
rect 8389 18105 8401 18139
rect 8435 18136 8447 18139
rect 8662 18136 8668 18148
rect 8435 18108 8668 18136
rect 8435 18105 8447 18108
rect 8389 18099 8447 18105
rect 8662 18096 8668 18108
rect 8720 18096 8726 18148
rect 10134 18096 10140 18148
rect 10192 18136 10198 18148
rect 10229 18139 10287 18145
rect 10229 18136 10241 18139
rect 10192 18108 10241 18136
rect 10192 18096 10198 18108
rect 10229 18105 10241 18108
rect 10275 18105 10287 18139
rect 10778 18136 10784 18148
rect 10739 18108 10784 18136
rect 10229 18099 10287 18105
rect 10778 18096 10784 18108
rect 10836 18096 10842 18148
rect 12529 18139 12587 18145
rect 12529 18136 12541 18139
rect 11808 18108 12541 18136
rect 9306 18068 9312 18080
rect 8220 18040 9312 18068
rect 5353 18031 5411 18037
rect 9306 18028 9312 18040
rect 9364 18028 9370 18080
rect 11422 18068 11428 18080
rect 11383 18040 11428 18068
rect 11422 18028 11428 18040
rect 11480 18028 11486 18080
rect 11514 18028 11520 18080
rect 11572 18068 11578 18080
rect 11808 18077 11836 18108
rect 12529 18105 12541 18108
rect 12575 18105 12587 18139
rect 12529 18099 12587 18105
rect 12618 18096 12624 18148
rect 12676 18136 12682 18148
rect 12676 18108 12721 18136
rect 12676 18096 12682 18108
rect 11793 18071 11851 18077
rect 11793 18068 11805 18071
rect 11572 18040 11805 18068
rect 11572 18028 11578 18040
rect 11793 18037 11805 18040
rect 11839 18037 11851 18071
rect 11793 18031 11851 18037
rect 12253 18071 12311 18077
rect 12253 18037 12265 18071
rect 12299 18068 12311 18071
rect 12636 18068 12664 18096
rect 12299 18040 12664 18068
rect 12299 18037 12311 18040
rect 12253 18031 12311 18037
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 3050 17824 3056 17876
rect 3108 17864 3114 17876
rect 4985 17867 5043 17873
rect 4985 17864 4997 17867
rect 3108 17836 4997 17864
rect 3108 17824 3114 17836
rect 4985 17833 4997 17836
rect 5031 17833 5043 17867
rect 4985 17827 5043 17833
rect 5074 17824 5080 17876
rect 5132 17864 5138 17876
rect 5261 17867 5319 17873
rect 5261 17864 5273 17867
rect 5132 17836 5273 17864
rect 5132 17824 5138 17836
rect 5261 17833 5273 17836
rect 5307 17833 5319 17867
rect 5261 17827 5319 17833
rect 5350 17824 5356 17876
rect 5408 17864 5414 17876
rect 5629 17867 5687 17873
rect 5629 17864 5641 17867
rect 5408 17836 5641 17864
rect 5408 17824 5414 17836
rect 5629 17833 5641 17836
rect 5675 17833 5687 17867
rect 5629 17827 5687 17833
rect 11790 17824 11796 17876
rect 11848 17864 11854 17876
rect 13173 17867 13231 17873
rect 13173 17864 13185 17867
rect 11848 17836 13185 17864
rect 11848 17824 11854 17836
rect 13173 17833 13185 17836
rect 13219 17833 13231 17867
rect 13173 17827 13231 17833
rect 4062 17796 4068 17808
rect 2700 17768 4068 17796
rect 2700 17740 2728 17768
rect 4062 17756 4068 17768
rect 4120 17756 4126 17808
rect 4246 17756 4252 17808
rect 4304 17796 4310 17808
rect 4386 17799 4444 17805
rect 4386 17796 4398 17799
rect 4304 17768 4398 17796
rect 4304 17756 4310 17768
rect 4386 17765 4398 17768
rect 4432 17765 4444 17799
rect 4386 17759 4444 17765
rect 1302 17688 1308 17740
rect 1360 17728 1366 17740
rect 1432 17731 1490 17737
rect 1432 17728 1444 17731
rect 1360 17700 1444 17728
rect 1360 17688 1366 17700
rect 1432 17697 1444 17700
rect 1478 17697 1490 17731
rect 2682 17728 2688 17740
rect 2643 17700 2688 17728
rect 1432 17691 1490 17697
rect 2682 17688 2688 17700
rect 2740 17688 2746 17740
rect 2866 17728 2872 17740
rect 2827 17700 2872 17728
rect 2866 17688 2872 17700
rect 2924 17688 2930 17740
rect 3145 17731 3203 17737
rect 3145 17697 3157 17731
rect 3191 17728 3203 17731
rect 5368 17728 5396 17824
rect 7190 17796 7196 17808
rect 7151 17768 7196 17796
rect 7190 17756 7196 17768
rect 7248 17796 7254 17808
rect 7469 17799 7527 17805
rect 7469 17796 7481 17799
rect 7248 17768 7481 17796
rect 7248 17756 7254 17768
rect 7469 17765 7481 17768
rect 7515 17765 7527 17799
rect 7469 17759 7527 17765
rect 7742 17756 7748 17808
rect 7800 17796 7806 17808
rect 8205 17799 8263 17805
rect 8205 17796 8217 17799
rect 7800 17768 8217 17796
rect 7800 17756 7806 17768
rect 8205 17765 8217 17768
rect 8251 17765 8263 17799
rect 8205 17759 8263 17765
rect 8757 17799 8815 17805
rect 8757 17765 8769 17799
rect 8803 17796 8815 17799
rect 8846 17796 8852 17808
rect 8803 17768 8852 17796
rect 8803 17765 8815 17768
rect 8757 17759 8815 17765
rect 8846 17756 8852 17768
rect 8904 17796 8910 17808
rect 9398 17796 9404 17808
rect 8904 17768 9404 17796
rect 8904 17756 8910 17768
rect 9398 17756 9404 17768
rect 9456 17796 9462 17808
rect 9861 17799 9919 17805
rect 9861 17796 9873 17799
rect 9456 17768 9873 17796
rect 9456 17756 9462 17768
rect 9861 17765 9873 17768
rect 9907 17765 9919 17799
rect 9861 17759 9919 17765
rect 9950 17756 9956 17808
rect 10008 17796 10014 17808
rect 10505 17799 10563 17805
rect 10008 17768 10053 17796
rect 10008 17756 10014 17768
rect 10505 17765 10517 17799
rect 10551 17796 10563 17799
rect 10778 17796 10784 17808
rect 10551 17768 10784 17796
rect 10551 17765 10563 17768
rect 10505 17759 10563 17765
rect 10778 17756 10784 17768
rect 10836 17756 10842 17808
rect 11146 17756 11152 17808
rect 11204 17796 11210 17808
rect 11330 17796 11336 17808
rect 11204 17768 11336 17796
rect 11204 17756 11210 17768
rect 11330 17756 11336 17768
rect 11388 17796 11394 17808
rect 11654 17799 11712 17805
rect 11654 17796 11666 17799
rect 11388 17768 11666 17796
rect 11388 17756 11394 17768
rect 11654 17765 11666 17768
rect 11700 17765 11712 17799
rect 12894 17796 12900 17808
rect 12855 17768 12900 17796
rect 11654 17759 11712 17765
rect 12894 17756 12900 17768
rect 12952 17756 12958 17808
rect 3191 17700 5396 17728
rect 6457 17731 6515 17737
rect 3191 17697 3203 17700
rect 3145 17691 3203 17697
rect 6457 17697 6469 17731
rect 6503 17697 6515 17731
rect 7006 17728 7012 17740
rect 6967 17700 7012 17728
rect 6457 17691 6515 17697
rect 4062 17660 4068 17672
rect 4023 17632 4068 17660
rect 4062 17620 4068 17632
rect 4120 17620 4126 17672
rect 4338 17620 4344 17672
rect 4396 17660 4402 17672
rect 6472 17660 6500 17691
rect 7006 17688 7012 17700
rect 7064 17688 7070 17740
rect 12250 17728 12256 17740
rect 12163 17700 12256 17728
rect 12250 17688 12256 17700
rect 12308 17728 12314 17740
rect 12986 17728 12992 17740
rect 12308 17700 12992 17728
rect 12308 17688 12314 17700
rect 12986 17688 12992 17700
rect 13044 17688 13050 17740
rect 13081 17731 13139 17737
rect 13081 17697 13093 17731
rect 13127 17697 13139 17731
rect 13538 17728 13544 17740
rect 13499 17700 13544 17728
rect 13081 17691 13139 17697
rect 6822 17660 6828 17672
rect 4396 17632 6828 17660
rect 4396 17620 4402 17632
rect 6822 17620 6828 17632
rect 6880 17620 6886 17672
rect 8113 17663 8171 17669
rect 8113 17660 8125 17663
rect 7852 17632 8125 17660
rect 1535 17527 1593 17533
rect 1535 17493 1547 17527
rect 1581 17524 1593 17527
rect 1762 17524 1768 17536
rect 1581 17496 1768 17524
rect 1581 17493 1593 17496
rect 1535 17487 1593 17493
rect 1762 17484 1768 17496
rect 1820 17484 1826 17536
rect 1946 17524 1952 17536
rect 1907 17496 1952 17524
rect 1946 17484 1952 17496
rect 2004 17484 2010 17536
rect 2314 17524 2320 17536
rect 2227 17496 2320 17524
rect 2314 17484 2320 17496
rect 2372 17524 2378 17536
rect 4614 17524 4620 17536
rect 2372 17496 4620 17524
rect 2372 17484 2378 17496
rect 4614 17484 4620 17496
rect 4672 17484 4678 17536
rect 7374 17484 7380 17536
rect 7432 17524 7438 17536
rect 7852 17533 7880 17632
rect 8113 17629 8125 17632
rect 8159 17629 8171 17663
rect 8113 17623 8171 17629
rect 11333 17663 11391 17669
rect 11333 17629 11345 17663
rect 11379 17660 11391 17663
rect 11790 17660 11796 17672
rect 11379 17632 11796 17660
rect 11379 17629 11391 17632
rect 11333 17623 11391 17629
rect 11790 17620 11796 17632
rect 11848 17620 11854 17672
rect 13096 17660 13124 17691
rect 13538 17688 13544 17700
rect 13596 17688 13602 17740
rect 15197 17731 15255 17737
rect 15197 17697 15209 17731
rect 15243 17728 15255 17731
rect 15378 17728 15384 17740
rect 15243 17700 15384 17728
rect 15243 17697 15255 17700
rect 15197 17691 15255 17697
rect 15378 17688 15384 17700
rect 15436 17688 15442 17740
rect 13446 17660 13452 17672
rect 12452 17632 13452 17660
rect 9214 17552 9220 17604
rect 9272 17592 9278 17604
rect 11146 17592 11152 17604
rect 9272 17564 11152 17592
rect 9272 17552 9278 17564
rect 11146 17552 11152 17564
rect 11204 17592 11210 17604
rect 12452 17592 12480 17632
rect 13446 17620 13452 17632
rect 13504 17620 13510 17672
rect 11204 17564 12480 17592
rect 11204 17552 11210 17564
rect 7837 17527 7895 17533
rect 7837 17524 7849 17527
rect 7432 17496 7849 17524
rect 7432 17484 7438 17496
rect 7837 17493 7849 17496
rect 7883 17493 7895 17527
rect 7837 17487 7895 17493
rect 14550 17484 14556 17536
rect 14608 17524 14614 17536
rect 15427 17527 15485 17533
rect 15427 17524 15439 17527
rect 14608 17496 15439 17524
rect 14608 17484 14614 17496
rect 15427 17493 15439 17496
rect 15473 17493 15485 17527
rect 15427 17487 15485 17493
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 1302 17280 1308 17332
rect 1360 17320 1366 17332
rect 1581 17323 1639 17329
rect 1581 17320 1593 17323
rect 1360 17292 1593 17320
rect 1360 17280 1366 17292
rect 1581 17289 1593 17292
rect 1627 17289 1639 17323
rect 2866 17320 2872 17332
rect 2827 17292 2872 17320
rect 1581 17283 1639 17289
rect 2866 17280 2872 17292
rect 2924 17280 2930 17332
rect 6822 17280 6828 17332
rect 6880 17320 6886 17332
rect 7009 17323 7067 17329
rect 7009 17320 7021 17323
rect 6880 17292 7021 17320
rect 6880 17280 6886 17292
rect 7009 17289 7021 17292
rect 7055 17320 7067 17323
rect 9214 17320 9220 17332
rect 7055 17292 9220 17320
rect 7055 17289 7067 17292
rect 7009 17283 7067 17289
rect 9214 17280 9220 17292
rect 9272 17280 9278 17332
rect 9493 17323 9551 17329
rect 9493 17289 9505 17323
rect 9539 17320 9551 17323
rect 9858 17320 9864 17332
rect 9539 17292 9864 17320
rect 9539 17289 9551 17292
rect 9493 17283 9551 17289
rect 9858 17280 9864 17292
rect 9916 17320 9922 17332
rect 10873 17323 10931 17329
rect 10873 17320 10885 17323
rect 9916 17292 10885 17320
rect 9916 17280 9922 17292
rect 10873 17289 10885 17292
rect 10919 17289 10931 17323
rect 11330 17320 11336 17332
rect 11291 17292 11336 17320
rect 10873 17283 10931 17289
rect 11330 17280 11336 17292
rect 11388 17280 11394 17332
rect 11790 17320 11796 17332
rect 11751 17292 11796 17320
rect 11790 17280 11796 17292
rect 11848 17280 11854 17332
rect 12250 17320 12256 17332
rect 12211 17292 12256 17320
rect 12250 17280 12256 17292
rect 12308 17280 12314 17332
rect 12618 17280 12624 17332
rect 12676 17320 12682 17332
rect 12713 17323 12771 17329
rect 12713 17320 12725 17323
rect 12676 17292 12725 17320
rect 12676 17280 12682 17292
rect 12713 17289 12725 17292
rect 12759 17289 12771 17323
rect 13446 17320 13452 17332
rect 13407 17292 13452 17320
rect 12713 17283 12771 17289
rect 13446 17280 13452 17292
rect 13504 17280 13510 17332
rect 8662 17212 8668 17264
rect 8720 17252 8726 17264
rect 9125 17255 9183 17261
rect 9125 17252 9137 17255
rect 8720 17224 9137 17252
rect 8720 17212 8726 17224
rect 9125 17221 9137 17224
rect 9171 17252 9183 17255
rect 11974 17252 11980 17264
rect 9171 17224 11980 17252
rect 9171 17221 9183 17224
rect 9125 17215 9183 17221
rect 11974 17212 11980 17224
rect 12032 17212 12038 17264
rect 10870 17144 10876 17196
rect 10928 17184 10934 17196
rect 13538 17184 13544 17196
rect 10928 17156 13544 17184
rect 10928 17144 10934 17156
rect 13538 17144 13544 17156
rect 13596 17184 13602 17196
rect 13817 17187 13875 17193
rect 13817 17184 13829 17187
rect 13596 17156 13829 17184
rect 13596 17144 13602 17156
rect 13817 17153 13829 17156
rect 13863 17153 13875 17187
rect 15378 17184 15384 17196
rect 15339 17156 15384 17184
rect 13817 17147 13875 17153
rect 15378 17144 15384 17156
rect 15436 17144 15442 17196
rect 1832 17119 1890 17125
rect 1832 17085 1844 17119
rect 1878 17116 1890 17119
rect 1946 17116 1952 17128
rect 1878 17088 1952 17116
rect 1878 17085 1890 17088
rect 1832 17079 1890 17085
rect 1946 17076 1952 17088
rect 2004 17076 2010 17128
rect 3510 17116 3516 17128
rect 3471 17088 3516 17116
rect 3510 17076 3516 17088
rect 3568 17076 3574 17128
rect 4525 17119 4583 17125
rect 4525 17085 4537 17119
rect 4571 17116 4583 17119
rect 4617 17119 4675 17125
rect 4617 17116 4629 17119
rect 4571 17088 4629 17116
rect 4571 17085 4583 17088
rect 4525 17079 4583 17085
rect 4617 17085 4629 17088
rect 4663 17116 4675 17119
rect 4982 17116 4988 17128
rect 4663 17088 4988 17116
rect 4663 17085 4675 17088
rect 4617 17079 4675 17085
rect 4982 17076 4988 17088
rect 5040 17076 5046 17128
rect 5074 17076 5080 17128
rect 5132 17116 5138 17128
rect 5629 17119 5687 17125
rect 5629 17116 5641 17119
rect 5132 17088 5641 17116
rect 5132 17076 5138 17088
rect 5629 17085 5641 17088
rect 5675 17085 5687 17119
rect 5629 17079 5687 17085
rect 6549 17119 6607 17125
rect 6549 17085 6561 17119
rect 6595 17116 6607 17119
rect 7006 17116 7012 17128
rect 6595 17088 7012 17116
rect 6595 17085 6607 17088
rect 6549 17079 6607 17085
rect 7006 17076 7012 17088
rect 7064 17116 7070 17128
rect 8018 17116 8024 17128
rect 7064 17088 8024 17116
rect 7064 17076 7070 17088
rect 8018 17076 8024 17088
rect 8076 17076 8082 17128
rect 8205 17119 8263 17125
rect 8205 17085 8217 17119
rect 8251 17116 8263 17119
rect 8294 17116 8300 17128
rect 8251 17088 8300 17116
rect 8251 17085 8263 17088
rect 8205 17079 8263 17085
rect 8294 17076 8300 17088
rect 8352 17076 8358 17128
rect 9950 17116 9956 17128
rect 9911 17088 9956 17116
rect 9950 17076 9956 17088
rect 10008 17076 10014 17128
rect 12250 17076 12256 17128
rect 12308 17116 12314 17128
rect 12529 17119 12587 17125
rect 12529 17116 12541 17119
rect 12308 17088 12541 17116
rect 12308 17076 12314 17088
rect 12529 17085 12541 17088
rect 12575 17085 12587 17119
rect 12529 17079 12587 17085
rect 3786 17048 3792 17060
rect 3747 17020 3792 17048
rect 3786 17008 3792 17020
rect 3844 17008 3850 17060
rect 8526 17051 8584 17057
rect 8526 17048 8538 17051
rect 8128 17020 8538 17048
rect 8128 16992 8156 17020
rect 8526 17017 8538 17020
rect 8572 17048 8584 17051
rect 9861 17051 9919 17057
rect 9861 17048 9873 17051
rect 8572 17020 9873 17048
rect 8572 17017 8584 17020
rect 8526 17011 8584 17017
rect 9861 17017 9873 17020
rect 9907 17048 9919 17051
rect 10315 17051 10373 17057
rect 10315 17048 10327 17051
rect 9907 17020 10327 17048
rect 9907 17017 9919 17020
rect 9861 17011 9919 17017
rect 10315 17017 10327 17020
rect 10361 17048 10373 17051
rect 11330 17048 11336 17060
rect 10361 17020 11336 17048
rect 10361 17017 10373 17020
rect 10315 17011 10373 17017
rect 11330 17008 11336 17020
rect 11388 17008 11394 17060
rect 1670 16940 1676 16992
rect 1728 16980 1734 16992
rect 1903 16983 1961 16989
rect 1903 16980 1915 16983
rect 1728 16952 1915 16980
rect 1728 16940 1734 16952
rect 1903 16949 1915 16952
rect 1949 16949 1961 16983
rect 1903 16943 1961 16949
rect 2501 16983 2559 16989
rect 2501 16949 2513 16983
rect 2547 16980 2559 16983
rect 2682 16980 2688 16992
rect 2547 16952 2688 16980
rect 2547 16949 2559 16952
rect 2501 16943 2559 16949
rect 2682 16940 2688 16952
rect 2740 16980 2746 16992
rect 2866 16980 2872 16992
rect 2740 16952 2872 16980
rect 2740 16940 2746 16952
rect 2866 16940 2872 16952
rect 2924 16940 2930 16992
rect 4157 16983 4215 16989
rect 4157 16949 4169 16983
rect 4203 16980 4215 16983
rect 4246 16980 4252 16992
rect 4203 16952 4252 16980
rect 4203 16949 4215 16952
rect 4157 16943 4215 16949
rect 4246 16940 4252 16952
rect 4304 16940 4310 16992
rect 4706 16980 4712 16992
rect 4667 16952 4712 16980
rect 4706 16940 4712 16952
rect 4764 16940 4770 16992
rect 7742 16980 7748 16992
rect 7703 16952 7748 16980
rect 7742 16940 7748 16952
rect 7800 16940 7806 16992
rect 8110 16980 8116 16992
rect 8071 16952 8116 16980
rect 8110 16940 8116 16952
rect 8168 16940 8174 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 3881 16779 3939 16785
rect 3881 16745 3893 16779
rect 3927 16776 3939 16779
rect 4062 16776 4068 16788
rect 3927 16748 4068 16776
rect 3927 16745 3939 16748
rect 3881 16739 3939 16745
rect 4062 16736 4068 16748
rect 4120 16776 4126 16788
rect 4706 16776 4712 16788
rect 4120 16748 4712 16776
rect 4120 16736 4126 16748
rect 4706 16736 4712 16748
rect 4764 16736 4770 16788
rect 6730 16776 6736 16788
rect 6691 16748 6736 16776
rect 6730 16736 6736 16748
rect 6788 16736 6794 16788
rect 9398 16776 9404 16788
rect 9359 16748 9404 16776
rect 9398 16736 9404 16748
rect 9456 16736 9462 16788
rect 1762 16668 1768 16720
rect 1820 16708 1826 16720
rect 2222 16708 2228 16720
rect 1820 16680 2228 16708
rect 1820 16668 1826 16680
rect 2222 16668 2228 16680
rect 2280 16708 2286 16720
rect 2501 16711 2559 16717
rect 2501 16708 2513 16711
rect 2280 16680 2513 16708
rect 2280 16668 2286 16680
rect 2501 16677 2513 16680
rect 2547 16677 2559 16711
rect 2501 16671 2559 16677
rect 2590 16668 2596 16720
rect 2648 16708 2654 16720
rect 3510 16708 3516 16720
rect 2648 16680 3516 16708
rect 2648 16668 2654 16680
rect 3510 16668 3516 16680
rect 3568 16668 3574 16720
rect 3786 16668 3792 16720
rect 3844 16708 3850 16720
rect 4249 16711 4307 16717
rect 4249 16708 4261 16711
rect 3844 16680 4261 16708
rect 3844 16668 3850 16680
rect 4249 16677 4261 16680
rect 4295 16677 4307 16711
rect 4249 16671 4307 16677
rect 5994 16668 6000 16720
rect 6052 16708 6058 16720
rect 6134 16711 6192 16717
rect 6134 16708 6146 16711
rect 6052 16680 6146 16708
rect 6052 16668 6058 16680
rect 6134 16677 6146 16680
rect 6180 16677 6192 16711
rect 6134 16671 6192 16677
rect 6914 16668 6920 16720
rect 6972 16708 6978 16720
rect 8389 16711 8447 16717
rect 6972 16680 8248 16708
rect 6972 16668 6978 16680
rect 1464 16643 1522 16649
rect 1464 16609 1476 16643
rect 1510 16640 1522 16643
rect 2314 16640 2320 16652
rect 1510 16612 2320 16640
rect 1510 16609 1522 16612
rect 1464 16603 1522 16609
rect 2314 16600 2320 16612
rect 2372 16600 2378 16652
rect 4982 16600 4988 16652
rect 5040 16640 5046 16652
rect 7650 16640 7656 16652
rect 5040 16612 7656 16640
rect 5040 16600 5046 16612
rect 7650 16600 7656 16612
rect 7708 16600 7714 16652
rect 7926 16600 7932 16652
rect 7984 16640 7990 16652
rect 8113 16643 8171 16649
rect 8113 16640 8125 16643
rect 7984 16612 8125 16640
rect 7984 16600 7990 16612
rect 8113 16609 8125 16612
rect 8159 16609 8171 16643
rect 8220 16640 8248 16680
rect 8389 16677 8401 16711
rect 8435 16708 8447 16711
rect 9950 16708 9956 16720
rect 8435 16680 9956 16708
rect 8435 16677 8447 16680
rect 8389 16671 8447 16677
rect 9950 16668 9956 16680
rect 10008 16668 10014 16720
rect 10962 16708 10968 16720
rect 10612 16680 10968 16708
rect 10612 16649 10640 16680
rect 10962 16668 10968 16680
rect 11020 16668 11026 16720
rect 11057 16711 11115 16717
rect 11057 16677 11069 16711
rect 11103 16708 11115 16711
rect 11422 16708 11428 16720
rect 11103 16680 11428 16708
rect 11103 16677 11115 16680
rect 11057 16671 11115 16677
rect 11422 16668 11428 16680
rect 11480 16668 11486 16720
rect 10597 16643 10655 16649
rect 10597 16640 10609 16643
rect 8220 16612 10609 16640
rect 8113 16603 8171 16609
rect 10597 16609 10609 16612
rect 10643 16609 10655 16643
rect 10870 16640 10876 16652
rect 10831 16612 10876 16640
rect 10597 16603 10655 16609
rect 10870 16600 10876 16612
rect 10928 16600 10934 16652
rect 11974 16640 11980 16652
rect 11935 16612 11980 16640
rect 11974 16600 11980 16612
rect 12032 16600 12038 16652
rect 4154 16532 4160 16584
rect 4212 16572 4218 16584
rect 4433 16575 4491 16581
rect 4212 16544 4257 16572
rect 4212 16532 4218 16544
rect 4433 16541 4445 16575
rect 4479 16541 4491 16575
rect 4433 16535 4491 16541
rect 3050 16504 3056 16516
rect 2963 16476 3056 16504
rect 3050 16464 3056 16476
rect 3108 16504 3114 16516
rect 4448 16504 4476 16535
rect 5442 16532 5448 16584
rect 5500 16572 5506 16584
rect 5813 16575 5871 16581
rect 5813 16572 5825 16575
rect 5500 16544 5825 16572
rect 5500 16532 5506 16544
rect 5813 16541 5825 16544
rect 5859 16541 5871 16575
rect 5813 16535 5871 16541
rect 7742 16532 7748 16584
rect 7800 16572 7806 16584
rect 11885 16575 11943 16581
rect 11885 16572 11897 16575
rect 7800 16544 11897 16572
rect 7800 16532 7806 16544
rect 11885 16541 11897 16544
rect 11931 16541 11943 16575
rect 11885 16535 11943 16541
rect 3108 16476 4476 16504
rect 3108 16464 3114 16476
rect 1394 16396 1400 16448
rect 1452 16436 1458 16448
rect 1535 16439 1593 16445
rect 1535 16436 1547 16439
rect 1452 16408 1547 16436
rect 1452 16396 1458 16408
rect 1535 16405 1547 16408
rect 1581 16405 1593 16439
rect 1854 16436 1860 16448
rect 1815 16408 1860 16436
rect 1535 16399 1593 16405
rect 1854 16396 1860 16408
rect 1912 16396 1918 16448
rect 2314 16436 2320 16448
rect 2275 16408 2320 16436
rect 2314 16396 2320 16408
rect 2372 16396 2378 16448
rect 3510 16436 3516 16448
rect 3471 16408 3516 16436
rect 3510 16396 3516 16408
rect 3568 16396 3574 16448
rect 4338 16396 4344 16448
rect 4396 16436 4402 16448
rect 5077 16439 5135 16445
rect 5077 16436 5089 16439
rect 4396 16408 5089 16436
rect 4396 16396 4402 16408
rect 5077 16405 5089 16408
rect 5123 16405 5135 16439
rect 5077 16399 5135 16405
rect 8294 16396 8300 16448
rect 8352 16436 8358 16448
rect 8665 16439 8723 16445
rect 8665 16436 8677 16439
rect 8352 16408 8677 16436
rect 8352 16396 8358 16408
rect 8665 16405 8677 16408
rect 8711 16405 8723 16439
rect 8665 16399 8723 16405
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 2501 16235 2559 16241
rect 2501 16201 2513 16235
rect 2547 16232 2559 16235
rect 2590 16232 2596 16244
rect 2547 16204 2596 16232
rect 2547 16201 2559 16204
rect 2501 16195 2559 16201
rect 2590 16192 2596 16204
rect 2648 16192 2654 16244
rect 3786 16192 3792 16244
rect 3844 16232 3850 16244
rect 4065 16235 4123 16241
rect 4065 16232 4077 16235
rect 3844 16204 4077 16232
rect 3844 16192 3850 16204
rect 4065 16201 4077 16204
rect 4111 16201 4123 16235
rect 7650 16232 7656 16244
rect 7611 16204 7656 16232
rect 4065 16195 4123 16201
rect 7650 16192 7656 16204
rect 7708 16192 7714 16244
rect 9122 16232 9128 16244
rect 9083 16204 9128 16232
rect 9122 16192 9128 16204
rect 9180 16192 9186 16244
rect 9490 16232 9496 16244
rect 9451 16204 9496 16232
rect 9490 16192 9496 16204
rect 9548 16232 9554 16244
rect 11974 16232 11980 16244
rect 9548 16204 10088 16232
rect 11935 16204 11980 16232
rect 9548 16192 9554 16204
rect 1489 16099 1547 16105
rect 1489 16065 1501 16099
rect 1535 16096 1547 16099
rect 1854 16096 1860 16108
rect 1535 16068 1860 16096
rect 1535 16065 1547 16068
rect 1489 16059 1547 16065
rect 1854 16056 1860 16068
rect 1912 16056 1918 16108
rect 2133 16099 2191 16105
rect 2133 16065 2145 16099
rect 2179 16096 2191 16099
rect 2314 16096 2320 16108
rect 2179 16068 2320 16096
rect 2179 16065 2191 16068
rect 2133 16059 2191 16065
rect 2314 16056 2320 16068
rect 2372 16096 2378 16108
rect 10060 16105 10088 16204
rect 11974 16192 11980 16204
rect 12032 16192 12038 16244
rect 3329 16099 3387 16105
rect 3329 16096 3341 16099
rect 2372 16068 3341 16096
rect 2372 16056 2378 16068
rect 3329 16065 3341 16068
rect 3375 16065 3387 16099
rect 3329 16059 3387 16065
rect 10045 16099 10103 16105
rect 10045 16065 10057 16099
rect 10091 16065 10103 16099
rect 10045 16059 10103 16065
rect 10134 16056 10140 16108
rect 10192 16096 10198 16108
rect 10192 16068 11652 16096
rect 10192 16056 10198 16068
rect 4338 15988 4344 16040
rect 4396 16028 4402 16040
rect 4525 16031 4583 16037
rect 4525 16028 4537 16031
rect 4396 16000 4537 16028
rect 4396 15988 4402 16000
rect 4525 15997 4537 16000
rect 4571 15997 4583 16031
rect 5074 16028 5080 16040
rect 5035 16000 5080 16028
rect 4525 15991 4583 15997
rect 5074 15988 5080 16000
rect 5132 15988 5138 16040
rect 5442 15988 5448 16040
rect 5500 16028 5506 16040
rect 6181 16031 6239 16037
rect 6181 16028 6193 16031
rect 5500 16000 6193 16028
rect 5500 15988 5506 16000
rect 6181 15997 6193 16000
rect 6227 15997 6239 16031
rect 8202 16028 8208 16040
rect 8163 16000 8208 16028
rect 6181 15991 6239 15997
rect 8202 15988 8208 16000
rect 8260 15988 8266 16040
rect 10689 16031 10747 16037
rect 10689 15997 10701 16031
rect 10735 16028 10747 16031
rect 10962 16028 10968 16040
rect 10735 16000 10968 16028
rect 10735 15997 10747 16000
rect 10689 15991 10747 15997
rect 10962 15988 10968 16000
rect 11020 15988 11026 16040
rect 11624 16037 11652 16068
rect 11609 16031 11667 16037
rect 11609 15997 11621 16031
rect 11655 16028 11667 16031
rect 12529 16031 12587 16037
rect 12529 16028 12541 16031
rect 11655 16000 12541 16028
rect 11655 15997 11667 16000
rect 11609 15991 11667 15997
rect 12529 15997 12541 16000
rect 12575 15997 12587 16031
rect 12529 15991 12587 15997
rect 1578 15960 1584 15972
rect 1539 15932 1584 15960
rect 1578 15920 1584 15932
rect 1636 15920 1642 15972
rect 3050 15960 3056 15972
rect 3011 15932 3056 15960
rect 3050 15920 3056 15932
rect 3108 15920 3114 15972
rect 3145 15963 3203 15969
rect 3145 15929 3157 15963
rect 3191 15929 3203 15963
rect 3145 15923 3203 15929
rect 2869 15895 2927 15901
rect 2869 15861 2881 15895
rect 2915 15892 2927 15895
rect 2958 15892 2964 15904
rect 2915 15864 2964 15892
rect 2915 15861 2927 15864
rect 2869 15855 2927 15861
rect 2958 15852 2964 15864
rect 3016 15892 3022 15904
rect 3160 15892 3188 15923
rect 5258 15920 5264 15972
rect 5316 15960 5322 15972
rect 6825 15963 6883 15969
rect 6825 15960 6837 15963
rect 5316 15932 6837 15960
rect 5316 15920 5322 15932
rect 6825 15929 6837 15932
rect 6871 15929 6883 15963
rect 6825 15923 6883 15929
rect 7377 15963 7435 15969
rect 7377 15929 7389 15963
rect 7423 15960 7435 15963
rect 7926 15960 7932 15972
rect 7423 15932 7932 15960
rect 7423 15929 7435 15932
rect 7377 15923 7435 15929
rect 7926 15920 7932 15932
rect 7984 15920 7990 15972
rect 8526 15963 8584 15969
rect 8526 15960 8538 15963
rect 8128 15932 8538 15960
rect 8128 15904 8156 15932
rect 8526 15929 8538 15932
rect 8572 15929 8584 15963
rect 8526 15923 8584 15929
rect 10134 15920 10140 15972
rect 10192 15960 10198 15972
rect 10192 15932 10237 15960
rect 10192 15920 10198 15932
rect 10778 15920 10784 15972
rect 10836 15960 10842 15972
rect 12437 15963 12495 15969
rect 12437 15960 12449 15963
rect 10836 15932 12449 15960
rect 10836 15920 10842 15932
rect 12437 15929 12449 15932
rect 12483 15929 12495 15963
rect 12437 15923 12495 15929
rect 4614 15892 4620 15904
rect 3016 15864 3188 15892
rect 4575 15864 4620 15892
rect 3016 15852 3022 15864
rect 4614 15852 4620 15864
rect 4672 15852 4678 15904
rect 5905 15895 5963 15901
rect 5905 15861 5917 15895
rect 5951 15892 5963 15895
rect 5994 15892 6000 15904
rect 5951 15864 6000 15892
rect 5951 15861 5963 15864
rect 5905 15855 5963 15861
rect 5994 15852 6000 15864
rect 6052 15892 6058 15904
rect 8021 15895 8079 15901
rect 8021 15892 8033 15895
rect 6052 15864 8033 15892
rect 6052 15852 6058 15864
rect 8021 15861 8033 15864
rect 8067 15892 8079 15895
rect 8110 15892 8116 15904
rect 8067 15864 8116 15892
rect 8067 15861 8079 15864
rect 8021 15855 8079 15861
rect 8110 15852 8116 15864
rect 8168 15852 8174 15904
rect 9582 15852 9588 15904
rect 9640 15892 9646 15904
rect 9769 15895 9827 15901
rect 9769 15892 9781 15895
rect 9640 15864 9781 15892
rect 9640 15852 9646 15864
rect 9769 15861 9781 15864
rect 9815 15892 9827 15895
rect 10870 15892 10876 15904
rect 9815 15864 10876 15892
rect 9815 15861 9827 15864
rect 9769 15855 9827 15861
rect 10870 15852 10876 15864
rect 10928 15852 10934 15904
rect 11054 15892 11060 15904
rect 11015 15864 11060 15892
rect 11054 15852 11060 15864
rect 11112 15852 11118 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1397 15691 1455 15697
rect 1397 15657 1409 15691
rect 1443 15688 1455 15691
rect 1854 15688 1860 15700
rect 1443 15660 1860 15688
rect 1443 15657 1455 15660
rect 1397 15651 1455 15657
rect 1854 15648 1860 15660
rect 1912 15648 1918 15700
rect 2222 15688 2228 15700
rect 2183 15660 2228 15688
rect 2222 15648 2228 15660
rect 2280 15648 2286 15700
rect 3050 15648 3056 15700
rect 3108 15688 3114 15700
rect 3421 15691 3479 15697
rect 3421 15688 3433 15691
rect 3108 15660 3433 15688
rect 3108 15648 3114 15660
rect 3421 15657 3433 15660
rect 3467 15657 3479 15691
rect 3421 15651 3479 15657
rect 3510 15648 3516 15700
rect 3568 15688 3574 15700
rect 4985 15691 5043 15697
rect 4985 15688 4997 15691
rect 3568 15660 4997 15688
rect 3568 15648 3574 15660
rect 4985 15657 4997 15660
rect 5031 15657 5043 15691
rect 4985 15651 5043 15657
rect 10045 15691 10103 15697
rect 10045 15657 10057 15691
rect 10091 15688 10103 15691
rect 10134 15688 10140 15700
rect 10091 15660 10140 15688
rect 10091 15657 10103 15660
rect 10045 15651 10103 15657
rect 10134 15648 10140 15660
rect 10192 15648 10198 15700
rect 3881 15623 3939 15629
rect 3881 15589 3893 15623
rect 3927 15620 3939 15623
rect 4154 15620 4160 15632
rect 3927 15592 4160 15620
rect 3927 15589 3939 15592
rect 3881 15583 3939 15589
rect 4154 15580 4160 15592
rect 4212 15580 4218 15632
rect 4246 15580 4252 15632
rect 4304 15620 4310 15632
rect 4386 15623 4444 15629
rect 4386 15620 4398 15623
rect 4304 15592 4398 15620
rect 4304 15580 4310 15592
rect 4386 15589 4398 15592
rect 4432 15589 4444 15623
rect 4386 15583 4444 15589
rect 6181 15623 6239 15629
rect 6181 15589 6193 15623
rect 6227 15620 6239 15623
rect 6362 15620 6368 15632
rect 6227 15592 6368 15620
rect 6227 15589 6239 15592
rect 6181 15583 6239 15589
rect 6362 15580 6368 15592
rect 6420 15580 6426 15632
rect 8294 15620 8300 15632
rect 8255 15592 8300 15620
rect 8294 15580 8300 15592
rect 8352 15580 8358 15632
rect 9950 15580 9956 15632
rect 10008 15620 10014 15632
rect 10413 15623 10471 15629
rect 10413 15620 10425 15623
rect 10008 15592 10425 15620
rect 10008 15580 10014 15592
rect 10413 15589 10425 15592
rect 10459 15620 10471 15623
rect 10778 15620 10784 15632
rect 10459 15592 10784 15620
rect 10459 15589 10471 15592
rect 10413 15583 10471 15589
rect 10778 15580 10784 15592
rect 10836 15580 10842 15632
rect 11606 15580 11612 15632
rect 11664 15620 11670 15632
rect 11885 15623 11943 15629
rect 11885 15620 11897 15623
rect 11664 15592 11897 15620
rect 11664 15580 11670 15592
rect 11885 15589 11897 15592
rect 11931 15589 11943 15623
rect 11885 15583 11943 15589
rect 11977 15623 12035 15629
rect 11977 15589 11989 15623
rect 12023 15620 12035 15623
rect 12802 15620 12808 15632
rect 12023 15592 12808 15620
rect 12023 15589 12035 15592
rect 11977 15583 12035 15589
rect 12802 15580 12808 15592
rect 12860 15580 12866 15632
rect 1578 15512 1584 15564
rect 1636 15552 1642 15564
rect 1949 15555 2007 15561
rect 1949 15552 1961 15555
rect 1636 15524 1961 15552
rect 1636 15512 1642 15524
rect 1949 15521 1961 15524
rect 1995 15552 2007 15555
rect 2409 15555 2467 15561
rect 2409 15552 2421 15555
rect 1995 15524 2421 15552
rect 1995 15521 2007 15524
rect 1949 15515 2007 15521
rect 2409 15521 2421 15524
rect 2455 15521 2467 15555
rect 2958 15552 2964 15564
rect 2919 15524 2964 15552
rect 2409 15515 2467 15521
rect 2958 15512 2964 15524
rect 3016 15512 3022 15564
rect 7098 15512 7104 15564
rect 7156 15552 7162 15564
rect 7561 15555 7619 15561
rect 7561 15552 7573 15555
rect 7156 15524 7573 15552
rect 7156 15512 7162 15524
rect 7561 15521 7573 15524
rect 7607 15521 7619 15555
rect 7561 15515 7619 15521
rect 7926 15512 7932 15564
rect 7984 15552 7990 15564
rect 8021 15555 8079 15561
rect 8021 15552 8033 15555
rect 7984 15524 8033 15552
rect 7984 15512 7990 15524
rect 8021 15521 8033 15524
rect 8067 15521 8079 15555
rect 8021 15515 8079 15521
rect 4065 15487 4123 15493
rect 4065 15453 4077 15487
rect 4111 15484 4123 15487
rect 4522 15484 4528 15496
rect 4111 15456 4528 15484
rect 4111 15453 4123 15456
rect 4065 15447 4123 15453
rect 4522 15444 4528 15456
rect 4580 15444 4586 15496
rect 6089 15487 6147 15493
rect 6089 15453 6101 15487
rect 6135 15453 6147 15487
rect 6089 15447 6147 15453
rect 6104 15416 6132 15447
rect 6178 15444 6184 15496
rect 6236 15484 6242 15496
rect 6365 15487 6423 15493
rect 6365 15484 6377 15487
rect 6236 15456 6377 15484
rect 6236 15444 6242 15456
rect 6365 15453 6377 15456
rect 6411 15453 6423 15487
rect 10318 15484 10324 15496
rect 10279 15456 10324 15484
rect 6365 15447 6423 15453
rect 10318 15444 10324 15456
rect 10376 15444 10382 15496
rect 10962 15484 10968 15496
rect 10923 15456 10968 15484
rect 10962 15444 10968 15456
rect 11020 15444 11026 15496
rect 12526 15484 12532 15496
rect 12487 15456 12532 15484
rect 12526 15444 12532 15456
rect 12584 15444 12590 15496
rect 13354 15484 13360 15496
rect 13315 15456 13360 15484
rect 13354 15444 13360 15456
rect 13412 15444 13418 15496
rect 6270 15416 6276 15428
rect 6104 15388 6276 15416
rect 6270 15376 6276 15388
rect 6328 15376 6334 15428
rect 8386 15376 8392 15428
rect 8444 15416 8450 15428
rect 8941 15419 8999 15425
rect 8941 15416 8953 15419
rect 8444 15388 8953 15416
rect 8444 15376 8450 15388
rect 8941 15385 8953 15388
rect 8987 15385 8999 15419
rect 8941 15379 8999 15385
rect 5074 15308 5080 15360
rect 5132 15348 5138 15360
rect 5261 15351 5319 15357
rect 5261 15348 5273 15351
rect 5132 15320 5273 15348
rect 5132 15308 5138 15320
rect 5261 15317 5273 15320
rect 5307 15317 5319 15351
rect 5261 15311 5319 15317
rect 5350 15308 5356 15360
rect 5408 15348 5414 15360
rect 5629 15351 5687 15357
rect 5629 15348 5641 15351
rect 5408 15320 5641 15348
rect 5408 15308 5414 15320
rect 5629 15317 5641 15320
rect 5675 15317 5687 15351
rect 7190 15348 7196 15360
rect 7151 15320 7196 15348
rect 5629 15311 5687 15317
rect 7190 15308 7196 15320
rect 7248 15308 7254 15360
rect 7834 15308 7840 15360
rect 7892 15348 7898 15360
rect 8202 15348 8208 15360
rect 7892 15320 8208 15348
rect 7892 15308 7898 15320
rect 8202 15308 8208 15320
rect 8260 15348 8266 15360
rect 8573 15351 8631 15357
rect 8573 15348 8585 15351
rect 8260 15320 8585 15348
rect 8260 15308 8266 15320
rect 8573 15317 8585 15320
rect 8619 15317 8631 15351
rect 12802 15348 12808 15360
rect 12763 15320 12808 15348
rect 8573 15311 8631 15317
rect 12802 15308 12808 15320
rect 12860 15308 12866 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 1486 15104 1492 15156
rect 1544 15144 1550 15156
rect 1581 15147 1639 15153
rect 1581 15144 1593 15147
rect 1544 15116 1593 15144
rect 1544 15104 1550 15116
rect 1581 15113 1593 15116
rect 1627 15113 1639 15147
rect 1581 15107 1639 15113
rect 2501 15147 2559 15153
rect 2501 15113 2513 15147
rect 2547 15144 2559 15147
rect 2958 15144 2964 15156
rect 2547 15116 2964 15144
rect 2547 15113 2559 15116
rect 2501 15107 2559 15113
rect 2958 15104 2964 15116
rect 3016 15144 3022 15156
rect 3973 15147 4031 15153
rect 3973 15144 3985 15147
rect 3016 15116 3985 15144
rect 3016 15104 3022 15116
rect 3973 15113 3985 15116
rect 4019 15113 4031 15147
rect 3973 15107 4031 15113
rect 6270 15104 6276 15156
rect 6328 15144 6334 15156
rect 6641 15147 6699 15153
rect 6641 15144 6653 15147
rect 6328 15116 6653 15144
rect 6328 15104 6334 15116
rect 6641 15113 6653 15116
rect 6687 15144 6699 15147
rect 7282 15144 7288 15156
rect 6687 15116 7288 15144
rect 6687 15113 6699 15116
rect 6641 15107 6699 15113
rect 7282 15104 7288 15116
rect 7340 15104 7346 15156
rect 8110 15104 8116 15156
rect 8168 15144 8174 15156
rect 8481 15147 8539 15153
rect 8481 15144 8493 15147
rect 8168 15116 8493 15144
rect 8168 15104 8174 15116
rect 8481 15113 8493 15116
rect 8527 15113 8539 15147
rect 9950 15144 9956 15156
rect 9911 15116 9956 15144
rect 8481 15107 8539 15113
rect 1946 15036 1952 15088
rect 2004 15076 2010 15088
rect 2004 15048 4154 15076
rect 2004 15036 2010 15048
rect 4126 15008 4154 15048
rect 5905 15011 5963 15017
rect 5905 15008 5917 15011
rect 4126 14980 5917 15008
rect 5905 14977 5917 14980
rect 5951 15008 5963 15011
rect 6178 15008 6184 15020
rect 5951 14980 6184 15008
rect 5951 14977 5963 14980
rect 5905 14971 5963 14977
rect 6178 14968 6184 14980
rect 6236 14968 6242 15020
rect 7834 15008 7840 15020
rect 7795 14980 7840 15008
rect 7834 14968 7840 14980
rect 7892 14968 7898 15020
rect 8496 15008 8524 15107
rect 9950 15104 9956 15116
rect 10008 15104 10014 15156
rect 10318 15104 10324 15156
rect 10376 15144 10382 15156
rect 11701 15147 11759 15153
rect 11701 15144 11713 15147
rect 10376 15116 11713 15144
rect 10376 15104 10382 15116
rect 11701 15113 11713 15116
rect 11747 15144 11759 15147
rect 13354 15144 13360 15156
rect 11747 15116 13360 15144
rect 11747 15113 11759 15116
rect 11701 15107 11759 15113
rect 13354 15104 13360 15116
rect 13412 15104 13418 15156
rect 25130 15144 25136 15156
rect 25091 15116 25136 15144
rect 25130 15104 25136 15116
rect 25188 15104 25194 15156
rect 9585 15079 9643 15085
rect 9585 15045 9597 15079
rect 9631 15076 9643 15079
rect 10134 15076 10140 15088
rect 9631 15048 10140 15076
rect 9631 15045 9643 15048
rect 9585 15039 9643 15045
rect 10134 15036 10140 15048
rect 10192 15036 10198 15088
rect 10042 15008 10048 15020
rect 8496 14980 10048 15008
rect 1394 14940 1400 14952
rect 1355 14912 1400 14940
rect 1394 14900 1400 14912
rect 1452 14940 1458 14952
rect 1949 14943 2007 14949
rect 1949 14940 1961 14943
rect 1452 14912 1961 14940
rect 1452 14900 1458 14912
rect 1949 14909 1961 14912
rect 1995 14909 2007 14943
rect 3050 14940 3056 14952
rect 3011 14912 3056 14940
rect 1949 14903 2007 14909
rect 3050 14900 3056 14912
rect 3108 14900 3114 14952
rect 7098 14940 7104 14952
rect 7059 14912 7104 14940
rect 7098 14900 7104 14912
rect 7156 14900 7162 14952
rect 7190 14900 7196 14952
rect 7248 14940 7254 14952
rect 7561 14943 7619 14949
rect 7561 14940 7573 14943
rect 7248 14912 7573 14940
rect 7248 14900 7254 14912
rect 7561 14909 7573 14912
rect 7607 14940 7619 14943
rect 8110 14940 8116 14952
rect 7607 14912 8116 14940
rect 7607 14909 7619 14912
rect 7561 14903 7619 14909
rect 8110 14900 8116 14912
rect 8168 14900 8174 14952
rect 8386 14900 8392 14952
rect 8444 14940 8450 14952
rect 8665 14943 8723 14949
rect 8665 14940 8677 14943
rect 8444 14912 8677 14940
rect 8444 14900 8450 14912
rect 8665 14909 8677 14912
rect 8711 14909 8723 14943
rect 8665 14903 8723 14909
rect 3374 14875 3432 14881
rect 3374 14841 3386 14875
rect 3420 14841 3432 14875
rect 3374 14835 3432 14841
rect 4709 14875 4767 14881
rect 4709 14841 4721 14875
rect 4755 14872 4767 14875
rect 5258 14872 5264 14884
rect 4755 14844 5264 14872
rect 4755 14841 4767 14844
rect 4709 14835 4767 14841
rect 2958 14804 2964 14816
rect 2919 14776 2964 14804
rect 2958 14764 2964 14776
rect 3016 14804 3022 14816
rect 3389 14804 3417 14835
rect 5258 14832 5264 14844
rect 5316 14832 5322 14884
rect 5353 14875 5411 14881
rect 5353 14841 5365 14875
rect 5399 14872 5411 14875
rect 6822 14872 6828 14884
rect 5399 14844 6828 14872
rect 5399 14841 5411 14844
rect 5353 14835 5411 14841
rect 4246 14804 4252 14816
rect 3016 14776 4252 14804
rect 3016 14764 3022 14776
rect 4246 14764 4252 14776
rect 4304 14764 4310 14816
rect 5077 14807 5135 14813
rect 5077 14773 5089 14807
rect 5123 14804 5135 14807
rect 5368 14804 5396 14835
rect 6822 14832 6828 14844
rect 6880 14832 6886 14884
rect 7116 14872 7144 14900
rect 8205 14875 8263 14881
rect 8205 14872 8217 14875
rect 7116 14844 8217 14872
rect 8205 14841 8217 14844
rect 8251 14841 8263 14875
rect 8772 14872 8800 14980
rect 10042 14968 10048 14980
rect 10100 15008 10106 15020
rect 10229 15011 10287 15017
rect 10229 15008 10241 15011
rect 10100 14980 10241 15008
rect 10100 14968 10106 14980
rect 10229 14977 10241 14980
rect 10275 14977 10287 15011
rect 10229 14971 10287 14977
rect 8986 14875 9044 14881
rect 8986 14872 8998 14875
rect 8772 14844 8998 14872
rect 8205 14835 8263 14841
rect 8986 14841 8998 14844
rect 9032 14841 9044 14875
rect 10244 14872 10272 14971
rect 10962 14968 10968 15020
rect 11020 15008 11026 15020
rect 11020 14980 13814 15008
rect 11020 14968 11026 14980
rect 10413 14943 10471 14949
rect 10413 14909 10425 14943
rect 10459 14940 10471 14943
rect 11238 14940 11244 14952
rect 10459 14912 11244 14940
rect 10459 14909 10471 14912
rect 10413 14903 10471 14909
rect 11238 14900 11244 14912
rect 11296 14900 11302 14952
rect 11333 14943 11391 14949
rect 11333 14909 11345 14943
rect 11379 14940 11391 14943
rect 12069 14943 12127 14949
rect 12069 14940 12081 14943
rect 11379 14912 12081 14940
rect 11379 14909 11391 14912
rect 11333 14903 11391 14909
rect 12069 14909 12081 14912
rect 12115 14940 12127 14943
rect 12802 14940 12808 14952
rect 12115 14912 12808 14940
rect 12115 14909 12127 14912
rect 12069 14903 12127 14909
rect 12802 14900 12808 14912
rect 12860 14900 12866 14952
rect 13786 14940 13814 14980
rect 19004 14943 19062 14949
rect 19004 14940 19016 14943
rect 13786 14912 19016 14940
rect 19004 14909 19016 14912
rect 19050 14940 19062 14943
rect 19429 14943 19487 14949
rect 19429 14940 19441 14943
rect 19050 14912 19441 14940
rect 19050 14909 19062 14912
rect 19004 14903 19062 14909
rect 19429 14909 19441 14912
rect 19475 14909 19487 14943
rect 19429 14903 19487 14909
rect 24648 14943 24706 14949
rect 24648 14909 24660 14943
rect 24694 14940 24706 14943
rect 25130 14940 25136 14952
rect 24694 14912 25136 14940
rect 24694 14909 24706 14912
rect 24648 14903 24706 14909
rect 25130 14900 25136 14912
rect 25188 14900 25194 14952
rect 10734 14875 10792 14881
rect 10734 14872 10746 14875
rect 10244 14844 10746 14872
rect 8986 14835 9044 14841
rect 10734 14841 10746 14844
rect 10780 14841 10792 14875
rect 12434 14872 12440 14884
rect 12395 14844 12440 14872
rect 10734 14835 10792 14841
rect 12434 14832 12440 14844
rect 12492 14832 12498 14884
rect 5123 14776 5396 14804
rect 6273 14807 6331 14813
rect 5123 14773 5135 14776
rect 5077 14767 5135 14773
rect 6273 14773 6285 14807
rect 6319 14804 6331 14807
rect 6362 14804 6368 14816
rect 6319 14776 6368 14804
rect 6319 14773 6331 14776
rect 6273 14767 6331 14773
rect 6362 14764 6368 14776
rect 6420 14764 6426 14816
rect 12158 14764 12164 14816
rect 12216 14804 12222 14816
rect 14001 14807 14059 14813
rect 14001 14804 14013 14807
rect 12216 14776 14013 14804
rect 12216 14764 12222 14776
rect 14001 14773 14013 14776
rect 14047 14773 14059 14807
rect 14001 14767 14059 14773
rect 19107 14807 19165 14813
rect 19107 14773 19119 14807
rect 19153 14804 19165 14807
rect 19242 14804 19248 14816
rect 19153 14776 19248 14804
rect 19153 14773 19165 14776
rect 19107 14767 19165 14773
rect 19242 14764 19248 14776
rect 19300 14764 19306 14816
rect 24210 14764 24216 14816
rect 24268 14804 24274 14816
rect 24719 14807 24777 14813
rect 24719 14804 24731 14807
rect 24268 14776 24731 14804
rect 24268 14764 24274 14776
rect 24719 14773 24731 14776
rect 24765 14773 24777 14807
rect 24719 14767 24777 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 3050 14560 3056 14612
rect 3108 14600 3114 14612
rect 3421 14603 3479 14609
rect 3421 14600 3433 14603
rect 3108 14572 3433 14600
rect 3108 14560 3114 14572
rect 3421 14569 3433 14572
rect 3467 14600 3479 14603
rect 3510 14600 3516 14612
rect 3467 14572 3516 14600
rect 3467 14569 3479 14572
rect 3421 14563 3479 14569
rect 3510 14560 3516 14572
rect 3568 14560 3574 14612
rect 3605 14603 3663 14609
rect 3605 14569 3617 14603
rect 3651 14600 3663 14603
rect 5350 14600 5356 14612
rect 3651 14572 5356 14600
rect 3651 14569 3663 14572
rect 3605 14563 3663 14569
rect 5350 14560 5356 14572
rect 5408 14560 5414 14612
rect 6638 14560 6644 14612
rect 6696 14600 6702 14612
rect 6733 14603 6791 14609
rect 6733 14600 6745 14603
rect 6696 14572 6745 14600
rect 6696 14560 6702 14572
rect 6733 14569 6745 14572
rect 6779 14569 6791 14603
rect 6733 14563 6791 14569
rect 9766 14560 9772 14612
rect 9824 14600 9830 14612
rect 10042 14600 10048 14612
rect 9824 14572 10048 14600
rect 9824 14560 9830 14572
rect 10042 14560 10048 14572
rect 10100 14560 10106 14612
rect 10597 14603 10655 14609
rect 10597 14569 10609 14603
rect 10643 14600 10655 14603
rect 10686 14600 10692 14612
rect 10643 14572 10692 14600
rect 10643 14569 10655 14572
rect 10597 14563 10655 14569
rect 10686 14560 10692 14572
rect 10744 14560 10750 14612
rect 11238 14600 11244 14612
rect 11199 14572 11244 14600
rect 11238 14560 11244 14572
rect 11296 14560 11302 14612
rect 11606 14560 11612 14612
rect 11664 14600 11670 14612
rect 11793 14603 11851 14609
rect 11793 14600 11805 14603
rect 11664 14572 11805 14600
rect 11664 14560 11670 14572
rect 11793 14569 11805 14572
rect 11839 14569 11851 14603
rect 11793 14563 11851 14569
rect 3145 14535 3203 14541
rect 3145 14501 3157 14535
rect 3191 14532 3203 14535
rect 5442 14532 5448 14544
rect 3191 14504 5448 14532
rect 3191 14501 3203 14504
rect 3145 14495 3203 14501
rect 5442 14492 5448 14504
rect 5500 14492 5506 14544
rect 5807 14535 5865 14541
rect 5807 14501 5819 14535
rect 5853 14532 5865 14535
rect 5994 14532 6000 14544
rect 5853 14504 6000 14532
rect 5853 14501 5865 14504
rect 5807 14495 5865 14501
rect 5994 14492 6000 14504
rect 6052 14492 6058 14544
rect 8386 14532 8392 14544
rect 8347 14504 8392 14532
rect 8386 14492 8392 14504
rect 8444 14492 8450 14544
rect 12158 14532 12164 14544
rect 12119 14504 12164 14532
rect 12158 14492 12164 14504
rect 12216 14492 12222 14544
rect 12253 14535 12311 14541
rect 12253 14501 12265 14535
rect 12299 14532 12311 14535
rect 12434 14532 12440 14544
rect 12299 14504 12440 14532
rect 12299 14501 12311 14504
rect 12253 14495 12311 14501
rect 12434 14492 12440 14504
rect 12492 14492 12498 14544
rect 1464 14467 1522 14473
rect 1464 14433 1476 14467
rect 1510 14464 1522 14467
rect 2314 14464 2320 14476
rect 1510 14436 2320 14464
rect 1510 14433 1522 14436
rect 1464 14427 1522 14433
rect 2314 14424 2320 14436
rect 2372 14424 2378 14476
rect 2682 14464 2688 14476
rect 2643 14436 2688 14464
rect 2682 14424 2688 14436
rect 2740 14424 2746 14476
rect 2961 14467 3019 14473
rect 2961 14433 2973 14467
rect 3007 14464 3019 14467
rect 3418 14464 3424 14476
rect 3007 14436 3424 14464
rect 3007 14433 3019 14436
rect 2961 14427 3019 14433
rect 3418 14424 3424 14436
rect 3476 14424 3482 14476
rect 4430 14464 4436 14476
rect 4391 14436 4436 14464
rect 4430 14424 4436 14436
rect 4488 14424 4494 14476
rect 4985 14467 5043 14473
rect 4985 14433 4997 14467
rect 5031 14464 5043 14467
rect 5534 14464 5540 14476
rect 5031 14436 5540 14464
rect 5031 14433 5043 14436
rect 4985 14427 5043 14433
rect 5534 14424 5540 14436
rect 5592 14424 5598 14476
rect 7650 14464 7656 14476
rect 7611 14436 7656 14464
rect 7650 14424 7656 14436
rect 7708 14424 7714 14476
rect 7834 14424 7840 14476
rect 7892 14464 7898 14476
rect 8110 14464 8116 14476
rect 7892 14436 8116 14464
rect 7892 14424 7898 14436
rect 8110 14424 8116 14436
rect 8168 14424 8174 14476
rect 13170 14424 13176 14476
rect 13228 14464 13234 14476
rect 13725 14467 13783 14473
rect 13725 14464 13737 14467
rect 13228 14436 13737 14464
rect 13228 14424 13234 14436
rect 13725 14433 13737 14436
rect 13771 14433 13783 14467
rect 13725 14427 13783 14433
rect 15324 14467 15382 14473
rect 15324 14433 15336 14467
rect 15370 14433 15382 14467
rect 15324 14427 15382 14433
rect 4338 14356 4344 14408
rect 4396 14396 4402 14408
rect 5442 14396 5448 14408
rect 4396 14368 5349 14396
rect 5403 14368 5448 14396
rect 4396 14356 4402 14368
rect 1394 14288 1400 14340
rect 1452 14328 1458 14340
rect 1535 14331 1593 14337
rect 1535 14328 1547 14331
rect 1452 14300 1547 14328
rect 1452 14288 1458 14300
rect 1535 14297 1547 14300
rect 1581 14328 1593 14331
rect 3605 14331 3663 14337
rect 3605 14328 3617 14331
rect 1581 14300 3617 14328
rect 1581 14297 1593 14300
rect 1535 14291 1593 14297
rect 3605 14297 3617 14300
rect 3651 14297 3663 14331
rect 5321 14328 5349 14368
rect 5442 14356 5448 14368
rect 5500 14356 5506 14408
rect 9677 14399 9735 14405
rect 9677 14396 9689 14399
rect 9508 14368 9689 14396
rect 7098 14328 7104 14340
rect 5321 14300 7104 14328
rect 3605 14291 3663 14297
rect 7098 14288 7104 14300
rect 7156 14288 7162 14340
rect 9508 14272 9536 14368
rect 9677 14365 9689 14368
rect 9723 14365 9735 14399
rect 12526 14396 12532 14408
rect 12487 14368 12532 14396
rect 9677 14359 9735 14365
rect 12526 14356 12532 14368
rect 12584 14356 12590 14408
rect 13630 14396 13636 14408
rect 13591 14368 13636 14396
rect 13630 14356 13636 14368
rect 13688 14356 13694 14408
rect 15339 14396 15367 14427
rect 15654 14396 15660 14408
rect 13786 14368 15660 14396
rect 12544 14328 12572 14356
rect 13786 14328 13814 14368
rect 15654 14356 15660 14368
rect 15712 14356 15718 14408
rect 12544 14300 13814 14328
rect 1854 14260 1860 14272
rect 1815 14232 1860 14260
rect 1854 14220 1860 14232
rect 1912 14220 1918 14272
rect 2314 14260 2320 14272
rect 2275 14232 2320 14260
rect 2314 14220 2320 14232
rect 2372 14220 2378 14272
rect 3786 14260 3792 14272
rect 3747 14232 3792 14260
rect 3786 14220 3792 14232
rect 3844 14220 3850 14272
rect 4341 14263 4399 14269
rect 4341 14229 4353 14263
rect 4387 14260 4399 14263
rect 4522 14260 4528 14272
rect 4387 14232 4528 14260
rect 4387 14229 4399 14232
rect 4341 14223 4399 14229
rect 4522 14220 4528 14232
rect 4580 14220 4586 14272
rect 4617 14263 4675 14269
rect 4617 14229 4629 14263
rect 4663 14260 4675 14263
rect 5166 14260 5172 14272
rect 4663 14232 5172 14260
rect 4663 14229 4675 14232
rect 4617 14223 4675 14229
rect 5166 14220 5172 14232
rect 5224 14220 5230 14272
rect 5350 14260 5356 14272
rect 5311 14232 5356 14260
rect 5350 14220 5356 14232
rect 5408 14220 5414 14272
rect 6362 14260 6368 14272
rect 6323 14232 6368 14260
rect 6362 14220 6368 14232
rect 6420 14220 6426 14272
rect 7561 14263 7619 14269
rect 7561 14229 7573 14263
rect 7607 14260 7619 14263
rect 7926 14260 7932 14272
rect 7607 14232 7932 14260
rect 7607 14229 7619 14232
rect 7561 14223 7619 14229
rect 7926 14220 7932 14232
rect 7984 14220 7990 14272
rect 8754 14260 8760 14272
rect 8715 14232 8760 14260
rect 8754 14220 8760 14232
rect 8812 14220 8818 14272
rect 8846 14220 8852 14272
rect 8904 14260 8910 14272
rect 9033 14263 9091 14269
rect 9033 14260 9045 14263
rect 8904 14232 9045 14260
rect 8904 14220 8910 14232
rect 9033 14229 9045 14232
rect 9079 14229 9091 14263
rect 9490 14260 9496 14272
rect 9451 14232 9496 14260
rect 9033 14223 9091 14229
rect 9490 14220 9496 14232
rect 9548 14220 9554 14272
rect 10870 14260 10876 14272
rect 10831 14232 10876 14260
rect 10870 14220 10876 14232
rect 10928 14220 10934 14272
rect 15286 14220 15292 14272
rect 15344 14260 15350 14272
rect 15427 14263 15485 14269
rect 15427 14260 15439 14263
rect 15344 14232 15439 14260
rect 15344 14220 15350 14232
rect 15427 14229 15439 14232
rect 15473 14229 15485 14263
rect 15427 14223 15485 14229
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1578 14056 1584 14068
rect 1539 14028 1584 14056
rect 1578 14016 1584 14028
rect 1636 14016 1642 14068
rect 4157 14059 4215 14065
rect 4157 14025 4169 14059
rect 4203 14056 4215 14059
rect 4430 14056 4436 14068
rect 4203 14028 4436 14056
rect 4203 14025 4215 14028
rect 4157 14019 4215 14025
rect 4430 14016 4436 14028
rect 4488 14016 4494 14068
rect 9490 14016 9496 14068
rect 9548 14056 9554 14068
rect 12161 14059 12219 14065
rect 9548 14028 9593 14056
rect 9548 14016 9554 14028
rect 12161 14025 12173 14059
rect 12207 14056 12219 14059
rect 12434 14056 12440 14068
rect 12207 14028 12440 14056
rect 12207 14025 12219 14028
rect 12161 14019 12219 14025
rect 12434 14016 12440 14028
rect 12492 14016 12498 14068
rect 13170 14056 13176 14068
rect 13131 14028 13176 14056
rect 13170 14016 13176 14028
rect 13228 14016 13234 14068
rect 13541 14059 13599 14065
rect 13541 14025 13553 14059
rect 13587 14056 13599 14059
rect 13630 14056 13636 14068
rect 13587 14028 13636 14056
rect 13587 14025 13599 14028
rect 13541 14019 13599 14025
rect 13630 14016 13636 14028
rect 13688 14016 13694 14068
rect 15654 14056 15660 14068
rect 15615 14028 15660 14056
rect 15654 14016 15660 14028
rect 15712 14016 15718 14068
rect 5350 13948 5356 14000
rect 5408 13988 5414 14000
rect 11238 13988 11244 14000
rect 5408 13960 5580 13988
rect 5408 13948 5414 13960
rect 2501 13923 2559 13929
rect 2501 13889 2513 13923
rect 2547 13920 2559 13923
rect 2682 13920 2688 13932
rect 2547 13892 2688 13920
rect 2547 13889 2559 13892
rect 2501 13883 2559 13889
rect 2682 13880 2688 13892
rect 2740 13920 2746 13932
rect 5552 13920 5580 13960
rect 6288 13960 8800 13988
rect 11199 13960 11244 13988
rect 2740 13892 5488 13920
rect 5552 13892 5672 13920
rect 2740 13880 2746 13892
rect 1397 13855 1455 13861
rect 1397 13821 1409 13855
rect 1443 13852 1455 13855
rect 1670 13852 1676 13864
rect 1443 13824 1676 13852
rect 1443 13821 1455 13824
rect 1397 13815 1455 13821
rect 1670 13812 1676 13824
rect 1728 13852 1734 13864
rect 2038 13852 2044 13864
rect 1728 13824 2044 13852
rect 1728 13812 1734 13824
rect 2038 13812 2044 13824
rect 2096 13812 2102 13864
rect 2961 13855 3019 13861
rect 2961 13821 2973 13855
rect 3007 13852 3019 13855
rect 3326 13852 3332 13864
rect 3007 13824 3332 13852
rect 3007 13821 3019 13824
rect 2961 13815 3019 13821
rect 3326 13812 3332 13824
rect 3384 13812 3390 13864
rect 3418 13812 3424 13864
rect 3476 13852 3482 13864
rect 3513 13855 3571 13861
rect 3513 13852 3525 13855
rect 3476 13824 3525 13852
rect 3476 13812 3482 13824
rect 3513 13821 3525 13824
rect 3559 13852 3571 13855
rect 3602 13852 3608 13864
rect 3559 13824 3608 13852
rect 3559 13821 3571 13824
rect 3513 13815 3571 13821
rect 3602 13812 3608 13824
rect 3660 13812 3666 13864
rect 4525 13855 4583 13861
rect 4525 13821 4537 13855
rect 4571 13852 4583 13855
rect 4614 13852 4620 13864
rect 4571 13824 4620 13852
rect 4571 13821 4583 13824
rect 4525 13815 4583 13821
rect 4614 13812 4620 13824
rect 4672 13812 4678 13864
rect 5460 13861 5488 13892
rect 5445 13855 5503 13861
rect 5445 13821 5457 13855
rect 5491 13852 5503 13855
rect 5534 13852 5540 13864
rect 5491 13824 5540 13852
rect 5491 13821 5503 13824
rect 5445 13815 5503 13821
rect 5534 13812 5540 13824
rect 5592 13812 5598 13864
rect 5644 13861 5672 13892
rect 5629 13855 5687 13861
rect 5629 13821 5641 13855
rect 5675 13852 5687 13855
rect 6288 13852 6316 13960
rect 8772 13932 8800 13960
rect 11238 13948 11244 13960
rect 11296 13948 11302 14000
rect 12342 13948 12348 14000
rect 12400 13988 12406 14000
rect 12621 13991 12679 13997
rect 12621 13988 12633 13991
rect 12400 13960 12633 13988
rect 12400 13948 12406 13960
rect 12621 13957 12633 13960
rect 12667 13957 12679 13991
rect 12621 13951 12679 13957
rect 6362 13880 6368 13932
rect 6420 13920 6426 13932
rect 6641 13923 6699 13929
rect 6641 13920 6653 13923
rect 6420 13892 6653 13920
rect 6420 13880 6426 13892
rect 6641 13889 6653 13892
rect 6687 13920 6699 13923
rect 6687 13892 6960 13920
rect 6687 13889 6699 13892
rect 6641 13883 6699 13889
rect 6822 13852 6828 13864
rect 5675 13824 6316 13852
rect 6783 13824 6828 13852
rect 5675 13821 5687 13824
rect 5629 13815 5687 13821
rect 6822 13812 6828 13824
rect 6880 13812 6886 13864
rect 6932 13861 6960 13892
rect 8754 13880 8760 13932
rect 8812 13920 8818 13932
rect 9309 13923 9367 13929
rect 9309 13920 9321 13923
rect 8812 13892 9321 13920
rect 8812 13880 8818 13892
rect 9309 13889 9321 13892
rect 9355 13920 9367 13923
rect 11793 13923 11851 13929
rect 9355 13892 10916 13920
rect 9355 13889 9367 13892
rect 9309 13883 9367 13889
rect 10888 13864 10916 13892
rect 11793 13889 11805 13923
rect 11839 13920 11851 13923
rect 12158 13920 12164 13932
rect 11839 13892 12164 13920
rect 11839 13889 11851 13892
rect 11793 13883 11851 13889
rect 12158 13880 12164 13892
rect 12216 13880 12222 13932
rect 13722 13920 13728 13932
rect 13635 13892 13728 13920
rect 13722 13880 13728 13892
rect 13780 13920 13786 13932
rect 14645 13923 14703 13929
rect 14645 13920 14657 13923
rect 13780 13892 14657 13920
rect 13780 13880 13786 13892
rect 14645 13889 14657 13892
rect 14691 13889 14703 13923
rect 14645 13883 14703 13889
rect 6917 13855 6975 13861
rect 6917 13821 6929 13855
rect 6963 13821 6975 13855
rect 6917 13815 6975 13821
rect 8205 13855 8263 13861
rect 8205 13821 8217 13855
rect 8251 13821 8263 13855
rect 8205 13815 8263 13821
rect 8573 13855 8631 13861
rect 8573 13821 8585 13855
rect 8619 13821 8631 13855
rect 8573 13815 8631 13821
rect 2133 13787 2191 13793
rect 2133 13753 2145 13787
rect 2179 13784 2191 13787
rect 3620 13784 3648 13812
rect 2179 13756 3648 13784
rect 3789 13787 3847 13793
rect 2179 13753 2191 13756
rect 2133 13747 2191 13753
rect 3789 13753 3801 13787
rect 3835 13784 3847 13787
rect 5350 13784 5356 13796
rect 3835 13756 5356 13784
rect 3835 13753 3847 13756
rect 3789 13747 3847 13753
rect 5350 13744 5356 13756
rect 5408 13744 5414 13796
rect 7190 13784 7196 13796
rect 5822 13756 7196 13784
rect 4522 13676 4528 13728
rect 4580 13716 4586 13728
rect 4709 13719 4767 13725
rect 4709 13716 4721 13719
rect 4580 13688 4721 13716
rect 4580 13676 4586 13688
rect 4709 13685 4721 13688
rect 4755 13685 4767 13719
rect 4709 13679 4767 13685
rect 5166 13676 5172 13728
rect 5224 13716 5230 13728
rect 5822 13716 5850 13756
rect 7190 13744 7196 13756
rect 7248 13784 7254 13796
rect 8220 13784 8248 13815
rect 7248 13756 8340 13784
rect 7248 13744 7254 13756
rect 5994 13716 6000 13728
rect 5224 13688 5850 13716
rect 5955 13688 6000 13716
rect 5224 13676 5230 13688
rect 5994 13676 6000 13688
rect 6052 13676 6058 13728
rect 7650 13676 7656 13728
rect 7708 13716 7714 13728
rect 7929 13719 7987 13725
rect 7929 13716 7941 13719
rect 7708 13688 7941 13716
rect 7708 13676 7714 13688
rect 7929 13685 7941 13688
rect 7975 13716 7987 13719
rect 8202 13716 8208 13728
rect 7975 13688 8208 13716
rect 7975 13685 7987 13688
rect 7929 13679 7987 13685
rect 8202 13676 8208 13688
rect 8260 13676 8266 13728
rect 8312 13716 8340 13756
rect 8588 13716 8616 13815
rect 9122 13812 9128 13864
rect 9180 13852 9186 13864
rect 9217 13855 9275 13861
rect 9217 13852 9229 13855
rect 9180 13824 9229 13852
rect 9180 13812 9186 13824
rect 9217 13821 9229 13824
rect 9263 13821 9275 13855
rect 10321 13855 10379 13861
rect 10321 13852 10333 13855
rect 9217 13815 9275 13821
rect 10152 13824 10333 13852
rect 10152 13793 10180 13824
rect 10321 13821 10333 13824
rect 10367 13821 10379 13855
rect 10870 13852 10876 13864
rect 10831 13824 10876 13852
rect 10321 13815 10379 13821
rect 10870 13812 10876 13824
rect 10928 13812 10934 13864
rect 10962 13812 10968 13864
rect 11020 13852 11026 13864
rect 11149 13855 11207 13861
rect 11149 13852 11161 13855
rect 11020 13824 11161 13852
rect 11020 13812 11026 13824
rect 11149 13821 11161 13824
rect 11195 13821 11207 13855
rect 11149 13815 11207 13821
rect 12437 13855 12495 13861
rect 12437 13821 12449 13855
rect 12483 13852 12495 13855
rect 12526 13852 12532 13864
rect 12483 13824 12532 13852
rect 12483 13821 12495 13824
rect 12437 13815 12495 13821
rect 12526 13812 12532 13824
rect 12584 13812 12590 13864
rect 10137 13787 10195 13793
rect 10137 13784 10149 13787
rect 9646 13756 10149 13784
rect 9646 13716 9674 13756
rect 10137 13753 10149 13756
rect 10183 13753 10195 13787
rect 10137 13747 10195 13753
rect 13817 13787 13875 13793
rect 13817 13753 13829 13787
rect 13863 13753 13875 13787
rect 14366 13784 14372 13796
rect 14327 13756 14372 13784
rect 13817 13747 13875 13753
rect 8312 13688 9674 13716
rect 9766 13676 9772 13728
rect 9824 13716 9830 13728
rect 9861 13719 9919 13725
rect 9861 13716 9873 13719
rect 9824 13688 9873 13716
rect 9824 13676 9830 13688
rect 9861 13685 9873 13688
rect 9907 13716 9919 13719
rect 9950 13716 9956 13728
rect 9907 13688 9956 13716
rect 9907 13685 9919 13688
rect 9861 13679 9919 13685
rect 9950 13676 9956 13688
rect 10008 13676 10014 13728
rect 13630 13676 13636 13728
rect 13688 13716 13694 13728
rect 13832 13716 13860 13747
rect 14366 13744 14372 13756
rect 14424 13744 14430 13796
rect 13688 13688 13860 13716
rect 13688 13676 13694 13688
rect 14458 13676 14464 13728
rect 14516 13716 14522 13728
rect 15197 13719 15255 13725
rect 15197 13716 15209 13719
rect 14516 13688 15209 13716
rect 14516 13676 14522 13688
rect 15197 13685 15209 13688
rect 15243 13685 15255 13719
rect 15197 13679 15255 13685
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1949 13515 2007 13521
rect 1949 13481 1961 13515
rect 1995 13512 2007 13515
rect 2038 13512 2044 13524
rect 1995 13484 2044 13512
rect 1995 13481 2007 13484
rect 1949 13475 2007 13481
rect 2038 13472 2044 13484
rect 2096 13472 2102 13524
rect 2130 13472 2136 13524
rect 2188 13512 2194 13524
rect 3050 13512 3056 13524
rect 2188 13484 3056 13512
rect 2188 13472 2194 13484
rect 3050 13472 3056 13484
rect 3108 13472 3114 13524
rect 3510 13472 3516 13524
rect 3568 13512 3574 13524
rect 4709 13515 4767 13521
rect 4709 13512 4721 13515
rect 3568 13484 4721 13512
rect 3568 13472 3574 13484
rect 4709 13481 4721 13484
rect 4755 13481 4767 13515
rect 4709 13475 4767 13481
rect 5442 13472 5448 13524
rect 5500 13512 5506 13524
rect 5997 13515 6055 13521
rect 5997 13512 6009 13515
rect 5500 13484 6009 13512
rect 5500 13472 5506 13484
rect 5997 13481 6009 13484
rect 6043 13481 6055 13515
rect 6730 13512 6736 13524
rect 5997 13475 6055 13481
rect 6564 13484 6736 13512
rect 6564 13453 6592 13484
rect 6730 13472 6736 13484
rect 6788 13512 6794 13524
rect 8570 13512 8576 13524
rect 6788 13484 7328 13512
rect 8531 13484 8576 13512
rect 6788 13472 6794 13484
rect 6549 13447 6607 13453
rect 6549 13444 6561 13447
rect 3068 13416 6561 13444
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 1946 13376 1952 13388
rect 1443 13348 1952 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 1946 13336 1952 13348
rect 2004 13336 2010 13388
rect 2498 13336 2504 13388
rect 2556 13376 2562 13388
rect 3068 13385 3096 13416
rect 6549 13413 6561 13416
rect 6595 13413 6607 13447
rect 6549 13407 6607 13413
rect 6638 13404 6644 13456
rect 6696 13444 6702 13456
rect 7300 13453 7328 13484
rect 8570 13472 8576 13484
rect 8628 13472 8634 13524
rect 9122 13472 9128 13524
rect 9180 13512 9186 13524
rect 9401 13515 9459 13521
rect 9401 13512 9413 13515
rect 9180 13484 9413 13512
rect 9180 13472 9186 13484
rect 9401 13481 9413 13484
rect 9447 13481 9459 13515
rect 12621 13515 12679 13521
rect 12621 13512 12633 13515
rect 9401 13475 9459 13481
rect 11624 13484 12633 13512
rect 7193 13447 7251 13453
rect 7193 13444 7205 13447
rect 6696 13416 7205 13444
rect 6696 13404 6702 13416
rect 7193 13413 7205 13416
rect 7239 13413 7251 13447
rect 7193 13407 7251 13413
rect 7285 13447 7343 13453
rect 7285 13413 7297 13447
rect 7331 13413 7343 13447
rect 7285 13407 7343 13413
rect 3053 13379 3111 13385
rect 3053 13376 3065 13379
rect 2556 13348 3065 13376
rect 2556 13336 2562 13348
rect 3053 13345 3065 13348
rect 3099 13345 3111 13379
rect 4614 13376 4620 13388
rect 4575 13348 4620 13376
rect 3053 13339 3111 13345
rect 4614 13336 4620 13348
rect 4672 13336 4678 13388
rect 5258 13376 5264 13388
rect 5219 13348 5264 13376
rect 5258 13336 5264 13348
rect 5316 13336 5322 13388
rect 5442 13376 5448 13388
rect 5403 13348 5448 13376
rect 5442 13336 5448 13348
rect 5500 13336 5506 13388
rect 9416 13376 9444 13475
rect 11624 13453 11652 13484
rect 12621 13481 12633 13484
rect 12667 13512 12679 13515
rect 12667 13484 14412 13512
rect 12667 13481 12679 13484
rect 12621 13475 12679 13481
rect 14384 13456 14412 13484
rect 24578 13472 24584 13524
rect 24636 13512 24642 13524
rect 24719 13515 24777 13521
rect 24719 13512 24731 13515
rect 24636 13484 24731 13512
rect 24636 13472 24642 13484
rect 24719 13481 24731 13484
rect 24765 13481 24777 13515
rect 24719 13475 24777 13481
rect 11609 13447 11667 13453
rect 11609 13413 11621 13447
rect 11655 13413 11667 13447
rect 11609 13407 11667 13413
rect 11701 13447 11759 13453
rect 11701 13413 11713 13447
rect 11747 13444 11759 13447
rect 11974 13444 11980 13456
rect 11747 13416 11980 13444
rect 11747 13413 11759 13416
rect 11701 13407 11759 13413
rect 11974 13404 11980 13416
rect 12032 13404 12038 13456
rect 12526 13404 12532 13456
rect 12584 13444 12590 13456
rect 12897 13447 12955 13453
rect 12897 13444 12909 13447
rect 12584 13416 12909 13444
rect 12584 13404 12590 13416
rect 12897 13413 12909 13416
rect 12943 13413 12955 13447
rect 12897 13407 12955 13413
rect 9769 13379 9827 13385
rect 9769 13376 9781 13379
rect 9416 13348 9781 13376
rect 9769 13345 9781 13348
rect 9815 13345 9827 13379
rect 9769 13339 9827 13345
rect 10134 13336 10140 13388
rect 10192 13376 10198 13388
rect 10229 13379 10287 13385
rect 10229 13376 10241 13379
rect 10192 13348 10241 13376
rect 10192 13336 10198 13348
rect 10229 13345 10241 13348
rect 10275 13345 10287 13379
rect 10229 13339 10287 13345
rect 12250 13336 12256 13388
rect 12308 13376 12314 13388
rect 12308 13348 12353 13376
rect 12308 13336 12314 13348
rect 3142 13308 3148 13320
rect 3103 13280 3148 13308
rect 3142 13268 3148 13280
rect 3200 13268 3206 13320
rect 3326 13268 3332 13320
rect 3384 13308 3390 13320
rect 4522 13308 4528 13320
rect 3384 13280 4528 13308
rect 3384 13268 3390 13280
rect 4522 13268 4528 13280
rect 4580 13268 4586 13320
rect 5276 13308 5304 13336
rect 7558 13308 7564 13320
rect 4908 13280 5304 13308
rect 7519 13280 7564 13308
rect 3418 13200 3424 13252
rect 3476 13240 3482 13252
rect 3789 13243 3847 13249
rect 3789 13240 3801 13243
rect 3476 13212 3801 13240
rect 3476 13200 3482 13212
rect 3789 13209 3801 13212
rect 3835 13240 3847 13243
rect 4908 13240 4936 13280
rect 7558 13268 7564 13280
rect 7616 13268 7622 13320
rect 10505 13311 10563 13317
rect 10505 13277 10517 13311
rect 10551 13308 10563 13311
rect 12434 13308 12440 13320
rect 10551 13280 12440 13308
rect 10551 13277 10563 13280
rect 10505 13271 10563 13277
rect 12434 13268 12440 13280
rect 12492 13268 12498 13320
rect 3835 13212 4936 13240
rect 12912 13240 12940 13407
rect 13170 13404 13176 13456
rect 13228 13444 13234 13456
rect 13817 13447 13875 13453
rect 13817 13444 13829 13447
rect 13228 13416 13829 13444
rect 13228 13404 13234 13416
rect 13817 13413 13829 13416
rect 13863 13413 13875 13447
rect 14366 13444 14372 13456
rect 14327 13416 14372 13444
rect 13817 13407 13875 13413
rect 14366 13404 14372 13416
rect 14424 13404 14430 13456
rect 15286 13376 15292 13388
rect 15247 13348 15292 13376
rect 15286 13336 15292 13348
rect 15344 13336 15350 13388
rect 24648 13379 24706 13385
rect 24648 13345 24660 13379
rect 24694 13376 24706 13379
rect 24854 13376 24860 13388
rect 24694 13348 24860 13376
rect 24694 13345 24706 13348
rect 24648 13339 24706 13345
rect 24854 13336 24860 13348
rect 24912 13336 24918 13388
rect 13722 13308 13728 13320
rect 13683 13280 13728 13308
rect 13722 13268 13728 13280
rect 13780 13268 13786 13320
rect 15746 13240 15752 13252
rect 12912 13212 15752 13240
rect 3835 13209 3847 13212
rect 3789 13203 3847 13209
rect 15746 13200 15752 13212
rect 15804 13200 15810 13252
rect 1581 13175 1639 13181
rect 1581 13141 1593 13175
rect 1627 13172 1639 13175
rect 2130 13172 2136 13184
rect 1627 13144 2136 13172
rect 1627 13141 1639 13144
rect 1581 13135 1639 13141
rect 2130 13132 2136 13144
rect 2188 13132 2194 13184
rect 2314 13172 2320 13184
rect 2275 13144 2320 13172
rect 2314 13132 2320 13144
rect 2372 13132 2378 13184
rect 3510 13172 3516 13184
rect 3471 13144 3516 13172
rect 3510 13132 3516 13144
rect 3568 13132 3574 13184
rect 4522 13172 4528 13184
rect 4435 13144 4528 13172
rect 4522 13132 4528 13144
rect 4580 13172 4586 13184
rect 4982 13172 4988 13184
rect 4580 13144 4988 13172
rect 4580 13132 4586 13144
rect 4982 13132 4988 13144
rect 5040 13132 5046 13184
rect 6546 13132 6552 13184
rect 6604 13172 6610 13184
rect 6917 13175 6975 13181
rect 6917 13172 6929 13175
rect 6604 13144 6929 13172
rect 6604 13132 6610 13144
rect 6917 13141 6929 13144
rect 6963 13141 6975 13175
rect 6917 13135 6975 13141
rect 7834 13132 7840 13184
rect 7892 13172 7898 13184
rect 8113 13175 8171 13181
rect 8113 13172 8125 13175
rect 7892 13144 8125 13172
rect 7892 13132 7898 13144
rect 8113 13141 8125 13144
rect 8159 13141 8171 13175
rect 8113 13135 8171 13141
rect 8570 13132 8576 13184
rect 8628 13172 8634 13184
rect 8849 13175 8907 13181
rect 8849 13172 8861 13175
rect 8628 13144 8861 13172
rect 8628 13132 8634 13144
rect 8849 13141 8861 13144
rect 8895 13141 8907 13175
rect 8849 13135 8907 13141
rect 9674 13132 9680 13184
rect 9732 13172 9738 13184
rect 10781 13175 10839 13181
rect 10781 13172 10793 13175
rect 9732 13144 10793 13172
rect 9732 13132 9738 13144
rect 10781 13141 10793 13144
rect 10827 13172 10839 13175
rect 10962 13172 10968 13184
rect 10827 13144 10968 13172
rect 10827 13141 10839 13144
rect 10781 13135 10839 13141
rect 10962 13132 10968 13144
rect 11020 13132 11026 13184
rect 11146 13172 11152 13184
rect 11107 13144 11152 13172
rect 11146 13132 11152 13144
rect 11204 13132 11210 13184
rect 15473 13175 15531 13181
rect 15473 13141 15485 13175
rect 15519 13172 15531 13175
rect 15838 13172 15844 13184
rect 15519 13144 15844 13172
rect 15519 13141 15531 13144
rect 15473 13135 15531 13141
rect 15838 13132 15844 13144
rect 15896 13132 15902 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 106 12928 112 12980
rect 164 12968 170 12980
rect 1581 12971 1639 12977
rect 1581 12968 1593 12971
rect 164 12940 1593 12968
rect 164 12928 170 12940
rect 1581 12937 1593 12940
rect 1627 12937 1639 12971
rect 1946 12968 1952 12980
rect 1907 12940 1952 12968
rect 1581 12931 1639 12937
rect 1946 12928 1952 12940
rect 2004 12928 2010 12980
rect 2498 12968 2504 12980
rect 2459 12940 2504 12968
rect 2498 12928 2504 12940
rect 2556 12928 2562 12980
rect 3142 12928 3148 12980
rect 3200 12968 3206 12980
rect 7101 12971 7159 12977
rect 7101 12968 7113 12971
rect 3200 12940 7113 12968
rect 3200 12928 3206 12940
rect 7101 12937 7113 12940
rect 7147 12968 7159 12971
rect 7466 12968 7472 12980
rect 7147 12940 7472 12968
rect 7147 12937 7159 12940
rect 7101 12931 7159 12937
rect 7466 12928 7472 12940
rect 7524 12928 7530 12980
rect 9306 12968 9312 12980
rect 9267 12940 9312 12968
rect 9306 12928 9312 12940
rect 9364 12928 9370 12980
rect 13170 12928 13176 12980
rect 13228 12968 13234 12980
rect 13357 12971 13415 12977
rect 13357 12968 13369 12971
rect 13228 12940 13369 12968
rect 13228 12928 13234 12940
rect 13357 12937 13369 12940
rect 13403 12968 13415 12971
rect 13633 12971 13691 12977
rect 13633 12968 13645 12971
rect 13403 12940 13645 12968
rect 13403 12937 13415 12940
rect 13357 12931 13415 12937
rect 13633 12937 13645 12940
rect 13679 12937 13691 12971
rect 15286 12968 15292 12980
rect 15247 12940 15292 12968
rect 13633 12931 13691 12937
rect 15286 12928 15292 12940
rect 15344 12928 15350 12980
rect 24673 12971 24731 12977
rect 24673 12937 24685 12971
rect 24719 12968 24731 12971
rect 24854 12968 24860 12980
rect 24719 12940 24860 12968
rect 24719 12937 24731 12940
rect 24673 12931 24731 12937
rect 24854 12928 24860 12940
rect 24912 12928 24918 12980
rect 4338 12900 4344 12912
rect 4299 12872 4344 12900
rect 4338 12860 4344 12872
rect 4396 12860 4402 12912
rect 5074 12860 5080 12912
rect 5132 12900 5138 12912
rect 5442 12900 5448 12912
rect 5132 12872 5448 12900
rect 5132 12860 5138 12872
rect 5442 12860 5448 12872
rect 5500 12860 5506 12912
rect 8662 12860 8668 12912
rect 8720 12900 8726 12912
rect 9125 12903 9183 12909
rect 9125 12900 9137 12903
rect 8720 12872 9137 12900
rect 8720 12860 8726 12872
rect 9125 12869 9137 12872
rect 9171 12869 9183 12903
rect 9125 12863 9183 12869
rect 3053 12835 3111 12841
rect 3053 12801 3065 12835
rect 3099 12832 3111 12835
rect 3786 12832 3792 12844
rect 3099 12804 3792 12832
rect 3099 12801 3111 12804
rect 3053 12795 3111 12801
rect 3786 12792 3792 12804
rect 3844 12832 3850 12844
rect 7558 12832 7564 12844
rect 3844 12804 7564 12832
rect 3844 12792 3850 12804
rect 7558 12792 7564 12804
rect 7616 12832 7622 12844
rect 7653 12835 7711 12841
rect 7653 12832 7665 12835
rect 7616 12804 7665 12832
rect 7616 12792 7622 12804
rect 7653 12801 7665 12804
rect 7699 12801 7711 12835
rect 7653 12795 7711 12801
rect 8481 12835 8539 12841
rect 8481 12801 8493 12835
rect 8527 12832 8539 12835
rect 9217 12835 9275 12841
rect 9217 12832 9229 12835
rect 8527 12804 9229 12832
rect 8527 12801 8539 12804
rect 8481 12795 8539 12801
rect 9217 12801 9229 12804
rect 9263 12801 9275 12835
rect 9217 12795 9275 12801
rect 10413 12835 10471 12841
rect 10413 12801 10425 12835
rect 10459 12832 10471 12835
rect 10686 12832 10692 12844
rect 10459 12804 10692 12832
rect 10459 12801 10471 12804
rect 10413 12795 10471 12801
rect 10686 12792 10692 12804
rect 10744 12832 10750 12844
rect 11146 12832 11152 12844
rect 10744 12804 11152 12832
rect 10744 12792 10750 12804
rect 11146 12792 11152 12804
rect 11204 12792 11210 12844
rect 12434 12832 12440 12844
rect 12395 12804 12440 12832
rect 12434 12792 12440 12804
rect 12492 12792 12498 12844
rect 1394 12764 1400 12776
rect 1355 12736 1400 12764
rect 1394 12724 1400 12736
rect 1452 12724 1458 12776
rect 4338 12724 4344 12776
rect 4396 12764 4402 12776
rect 4798 12764 4804 12776
rect 4396 12736 4804 12764
rect 4396 12724 4402 12736
rect 4798 12724 4804 12736
rect 4856 12764 4862 12776
rect 4893 12767 4951 12773
rect 4893 12764 4905 12767
rect 4856 12736 4905 12764
rect 4856 12724 4862 12736
rect 4893 12733 4905 12736
rect 4939 12733 4951 12767
rect 4893 12727 4951 12733
rect 4982 12724 4988 12776
rect 5040 12764 5046 12776
rect 5445 12767 5503 12773
rect 5445 12764 5457 12767
rect 5040 12736 5457 12764
rect 5040 12724 5046 12736
rect 5445 12733 5457 12736
rect 5491 12764 5503 12767
rect 5905 12767 5963 12773
rect 5905 12764 5917 12767
rect 5491 12736 5917 12764
rect 5491 12733 5503 12736
rect 5445 12727 5503 12733
rect 5905 12733 5917 12736
rect 5951 12733 5963 12767
rect 5905 12727 5963 12733
rect 8570 12724 8576 12776
rect 8628 12764 8634 12776
rect 8849 12767 8907 12773
rect 8849 12764 8861 12767
rect 8628 12736 8861 12764
rect 8628 12724 8634 12736
rect 8849 12733 8861 12736
rect 8895 12733 8907 12767
rect 8849 12727 8907 12733
rect 8938 12724 8944 12776
rect 8996 12773 9002 12776
rect 8996 12767 9054 12773
rect 8996 12733 9008 12767
rect 9042 12733 9054 12767
rect 8996 12727 9054 12733
rect 14093 12767 14151 12773
rect 14093 12733 14105 12767
rect 14139 12764 14151 12767
rect 14274 12764 14280 12776
rect 14139 12736 14280 12764
rect 14139 12733 14151 12736
rect 14093 12727 14151 12733
rect 8996 12724 9002 12727
rect 14274 12724 14280 12736
rect 14332 12724 14338 12776
rect 2869 12699 2927 12705
rect 2869 12665 2881 12699
rect 2915 12696 2927 12699
rect 3145 12699 3203 12705
rect 3145 12696 3157 12699
rect 2915 12668 3157 12696
rect 2915 12665 2927 12668
rect 2869 12659 2927 12665
rect 3145 12665 3157 12668
rect 3191 12696 3203 12699
rect 3326 12696 3332 12708
rect 3191 12668 3332 12696
rect 3191 12665 3203 12668
rect 3145 12659 3203 12665
rect 3326 12656 3332 12668
rect 3384 12656 3390 12708
rect 3694 12696 3700 12708
rect 3655 12668 3700 12696
rect 3694 12656 3700 12668
rect 3752 12656 3758 12708
rect 4062 12656 4068 12708
rect 4120 12696 4126 12708
rect 7377 12699 7435 12705
rect 4120 12668 5028 12696
rect 4120 12656 4126 12668
rect 4614 12628 4620 12640
rect 4575 12600 4620 12628
rect 4614 12588 4620 12600
rect 4672 12588 4678 12640
rect 5000 12637 5028 12668
rect 7377 12665 7389 12699
rect 7423 12665 7435 12699
rect 7377 12659 7435 12665
rect 4985 12631 5043 12637
rect 4985 12597 4997 12631
rect 5031 12628 5043 12631
rect 5810 12628 5816 12640
rect 5031 12600 5816 12628
rect 5031 12597 5043 12600
rect 4985 12591 5043 12597
rect 5810 12588 5816 12600
rect 5868 12588 5874 12640
rect 6546 12628 6552 12640
rect 6507 12600 6552 12628
rect 6546 12588 6552 12600
rect 6604 12588 6610 12640
rect 7392 12628 7420 12659
rect 7466 12656 7472 12708
rect 7524 12696 7530 12708
rect 8754 12696 8760 12708
rect 7524 12668 7569 12696
rect 7668 12668 8760 12696
rect 7524 12656 7530 12668
rect 7668 12628 7696 12668
rect 8754 12656 8760 12668
rect 8812 12656 8818 12708
rect 9950 12656 9956 12708
rect 10008 12696 10014 12708
rect 10321 12699 10379 12705
rect 10321 12696 10333 12699
rect 10008 12668 10333 12696
rect 10008 12656 10014 12668
rect 10321 12665 10333 12668
rect 10367 12696 10379 12699
rect 10775 12699 10833 12705
rect 10775 12696 10787 12699
rect 10367 12668 10787 12696
rect 10367 12665 10379 12668
rect 10321 12659 10379 12665
rect 10775 12665 10787 12668
rect 10821 12696 10833 12699
rect 12758 12699 12816 12705
rect 12758 12696 12770 12699
rect 10821 12668 12770 12696
rect 10821 12665 10833 12668
rect 10775 12659 10833 12665
rect 12268 12640 12296 12668
rect 12758 12665 12770 12668
rect 12804 12665 12816 12699
rect 14182 12696 14188 12708
rect 14143 12668 14188 12696
rect 12758 12659 12816 12665
rect 14182 12656 14188 12668
rect 14240 12656 14246 12708
rect 7392 12600 7696 12628
rect 8018 12588 8024 12640
rect 8076 12628 8082 12640
rect 8297 12631 8355 12637
rect 8297 12628 8309 12631
rect 8076 12600 8309 12628
rect 8076 12588 8082 12600
rect 8297 12597 8309 12600
rect 8343 12628 8355 12631
rect 8481 12631 8539 12637
rect 8481 12628 8493 12631
rect 8343 12600 8493 12628
rect 8343 12597 8355 12600
rect 8297 12591 8355 12597
rect 8481 12597 8493 12600
rect 8527 12597 8539 12631
rect 8662 12628 8668 12640
rect 8623 12600 8668 12628
rect 8481 12591 8539 12597
rect 8662 12588 8668 12600
rect 8720 12588 8726 12640
rect 9674 12588 9680 12640
rect 9732 12628 9738 12640
rect 9861 12631 9919 12637
rect 9861 12628 9873 12631
rect 9732 12600 9873 12628
rect 9732 12588 9738 12600
rect 9861 12597 9873 12600
rect 9907 12597 9919 12631
rect 9861 12591 9919 12597
rect 11333 12631 11391 12637
rect 11333 12597 11345 12631
rect 11379 12628 11391 12631
rect 11701 12631 11759 12637
rect 11701 12628 11713 12631
rect 11379 12600 11713 12628
rect 11379 12597 11391 12600
rect 11333 12591 11391 12597
rect 11701 12597 11713 12600
rect 11747 12628 11759 12631
rect 11974 12628 11980 12640
rect 11747 12600 11980 12628
rect 11747 12597 11759 12600
rect 11701 12591 11759 12597
rect 11974 12588 11980 12600
rect 12032 12588 12038 12640
rect 12250 12628 12256 12640
rect 12211 12600 12256 12628
rect 12250 12588 12256 12600
rect 12308 12588 12314 12640
rect 15378 12588 15384 12640
rect 15436 12628 15442 12640
rect 15749 12631 15807 12637
rect 15749 12628 15761 12631
rect 15436 12600 15761 12628
rect 15436 12588 15442 12600
rect 15749 12597 15761 12600
rect 15795 12597 15807 12631
rect 15749 12591 15807 12597
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1581 12427 1639 12433
rect 1581 12393 1593 12427
rect 1627 12424 1639 12427
rect 3418 12424 3424 12436
rect 1627 12396 3424 12424
rect 1627 12393 1639 12396
rect 1581 12387 1639 12393
rect 3418 12384 3424 12396
rect 3476 12384 3482 12436
rect 3513 12427 3571 12433
rect 3513 12393 3525 12427
rect 3559 12424 3571 12427
rect 4062 12424 4068 12436
rect 3559 12396 4068 12424
rect 3559 12393 3571 12396
rect 3513 12387 3571 12393
rect 4062 12384 4068 12396
rect 4120 12384 4126 12436
rect 4338 12424 4344 12436
rect 4299 12396 4344 12424
rect 4338 12384 4344 12396
rect 4396 12384 4402 12436
rect 6730 12424 6736 12436
rect 6691 12396 6736 12424
rect 6730 12384 6736 12396
rect 6788 12384 6794 12436
rect 8846 12424 8852 12436
rect 8807 12396 8852 12424
rect 8846 12384 8852 12396
rect 8904 12384 8910 12436
rect 10134 12424 10140 12436
rect 9646 12396 10140 12424
rect 2498 12316 2504 12368
rect 2556 12356 2562 12368
rect 2593 12359 2651 12365
rect 2593 12356 2605 12359
rect 2556 12328 2605 12356
rect 2556 12316 2562 12328
rect 2593 12325 2605 12328
rect 2639 12325 2651 12359
rect 2593 12319 2651 12325
rect 2682 12316 2688 12368
rect 2740 12356 2746 12368
rect 3145 12359 3203 12365
rect 3145 12356 3157 12359
rect 2740 12328 3157 12356
rect 2740 12316 2746 12328
rect 3145 12325 3157 12328
rect 3191 12356 3203 12359
rect 3694 12356 3700 12368
rect 3191 12328 3700 12356
rect 3191 12325 3203 12328
rect 3145 12319 3203 12325
rect 3694 12316 3700 12328
rect 3752 12316 3758 12368
rect 5994 12316 6000 12368
rect 6052 12356 6058 12368
rect 6134 12359 6192 12365
rect 6134 12356 6146 12359
rect 6052 12328 6146 12356
rect 6052 12316 6058 12328
rect 6134 12325 6146 12328
rect 6180 12325 6192 12359
rect 6134 12319 6192 12325
rect 8297 12359 8355 12365
rect 8297 12325 8309 12359
rect 8343 12356 8355 12359
rect 9646 12356 9674 12396
rect 10134 12384 10140 12396
rect 10192 12424 10198 12436
rect 10781 12427 10839 12433
rect 10192 12396 10272 12424
rect 10192 12384 10198 12396
rect 8343 12328 9674 12356
rect 8343 12325 8355 12328
rect 8297 12319 8355 12325
rect 1397 12291 1455 12297
rect 1397 12257 1409 12291
rect 1443 12288 1455 12291
rect 1946 12288 1952 12300
rect 1443 12260 1952 12288
rect 1443 12257 1455 12260
rect 1397 12251 1455 12257
rect 1946 12248 1952 12260
rect 2004 12248 2010 12300
rect 4246 12288 4252 12300
rect 4207 12260 4252 12288
rect 4246 12248 4252 12260
rect 4304 12248 4310 12300
rect 4617 12291 4675 12297
rect 4617 12257 4629 12291
rect 4663 12288 4675 12291
rect 4982 12288 4988 12300
rect 4663 12260 4988 12288
rect 4663 12257 4675 12260
rect 4617 12251 4675 12257
rect 2501 12223 2559 12229
rect 2501 12220 2513 12223
rect 2240 12192 2513 12220
rect 2240 12096 2268 12192
rect 2501 12189 2513 12192
rect 2547 12189 2559 12223
rect 2501 12183 2559 12189
rect 3881 12223 3939 12229
rect 3881 12189 3893 12223
rect 3927 12220 3939 12223
rect 4632 12220 4660 12251
rect 4982 12248 4988 12260
rect 5040 12248 5046 12300
rect 5810 12288 5816 12300
rect 5771 12260 5816 12288
rect 5810 12248 5816 12260
rect 5868 12248 5874 12300
rect 7098 12248 7104 12300
rect 7156 12288 7162 12300
rect 7561 12291 7619 12297
rect 7561 12288 7573 12291
rect 7156 12260 7573 12288
rect 7156 12248 7162 12260
rect 7561 12257 7573 12260
rect 7607 12257 7619 12291
rect 9674 12288 9680 12300
rect 9635 12260 9680 12288
rect 7561 12251 7619 12257
rect 9674 12248 9680 12260
rect 9732 12248 9738 12300
rect 10244 12297 10272 12396
rect 10781 12393 10793 12427
rect 10827 12424 10839 12427
rect 11057 12427 11115 12433
rect 11057 12424 11069 12427
rect 10827 12396 11069 12424
rect 10827 12393 10839 12396
rect 10781 12387 10839 12393
rect 11057 12393 11069 12396
rect 11103 12393 11115 12427
rect 12434 12424 12440 12436
rect 12395 12396 12440 12424
rect 11057 12387 11115 12393
rect 10413 12359 10471 12365
rect 10413 12325 10425 12359
rect 10459 12356 10471 12359
rect 10686 12356 10692 12368
rect 10459 12328 10692 12356
rect 10459 12325 10471 12328
rect 10413 12319 10471 12325
rect 10686 12316 10692 12328
rect 10744 12316 10750 12368
rect 10229 12291 10287 12297
rect 10229 12257 10241 12291
rect 10275 12288 10287 12291
rect 10796 12288 10824 12387
rect 12434 12384 12440 12396
rect 12492 12384 12498 12436
rect 13722 12384 13728 12436
rect 13780 12424 13786 12436
rect 13780 12396 13952 12424
rect 13780 12384 13786 12396
rect 11422 12356 11428 12368
rect 11383 12328 11428 12356
rect 11422 12316 11428 12328
rect 11480 12316 11486 12368
rect 10275 12260 10824 12288
rect 10275 12257 10287 12260
rect 10229 12251 10287 12257
rect 11974 12248 11980 12300
rect 12032 12288 12038 12300
rect 13449 12291 13507 12297
rect 13449 12288 13461 12291
rect 12032 12260 13461 12288
rect 12032 12248 12038 12260
rect 13449 12257 13461 12260
rect 13495 12288 13507 12291
rect 13814 12288 13820 12300
rect 13495 12260 13820 12288
rect 13495 12257 13507 12260
rect 13449 12251 13507 12257
rect 13814 12248 13820 12260
rect 13872 12248 13878 12300
rect 3927 12192 4660 12220
rect 3927 12189 3939 12192
rect 3881 12183 3939 12189
rect 7650 12180 7656 12232
rect 7708 12220 7714 12232
rect 7929 12223 7987 12229
rect 7708 12192 7880 12220
rect 7708 12180 7714 12192
rect 3510 12112 3516 12164
rect 3568 12152 3574 12164
rect 5258 12152 5264 12164
rect 3568 12124 5264 12152
rect 3568 12112 3574 12124
rect 5258 12112 5264 12124
rect 5316 12112 5322 12164
rect 7852 12161 7880 12192
rect 7929 12189 7941 12223
rect 7975 12220 7987 12223
rect 8018 12220 8024 12232
rect 7975 12192 8024 12220
rect 7975 12189 7987 12192
rect 7929 12183 7987 12189
rect 8018 12180 8024 12192
rect 8076 12180 8082 12232
rect 11330 12220 11336 12232
rect 11243 12192 11336 12220
rect 11330 12180 11336 12192
rect 11388 12220 11394 12232
rect 12802 12220 12808 12232
rect 11388 12192 12112 12220
rect 12763 12192 12808 12220
rect 11388 12180 11394 12192
rect 7837 12155 7895 12161
rect 7837 12121 7849 12155
rect 7883 12121 7895 12155
rect 7837 12115 7895 12121
rect 8570 12112 8576 12164
rect 8628 12152 8634 12164
rect 9217 12155 9275 12161
rect 9217 12152 9229 12155
rect 8628 12124 9229 12152
rect 8628 12112 8634 12124
rect 9217 12121 9229 12124
rect 9263 12121 9275 12155
rect 11882 12152 11888 12164
rect 11843 12124 11888 12152
rect 9217 12115 9275 12121
rect 11882 12112 11888 12124
rect 11940 12112 11946 12164
rect 12084 12152 12112 12192
rect 12802 12180 12808 12192
rect 12860 12180 12866 12232
rect 13924 12161 13952 12396
rect 15286 12384 15292 12436
rect 15344 12424 15350 12436
rect 15344 12396 15516 12424
rect 15344 12384 15350 12396
rect 15488 12365 15516 12396
rect 15473 12359 15531 12365
rect 15473 12325 15485 12359
rect 15519 12325 15531 12359
rect 15473 12319 15531 12325
rect 15381 12223 15439 12229
rect 15381 12189 15393 12223
rect 15427 12220 15439 12223
rect 15470 12220 15476 12232
rect 15427 12192 15476 12220
rect 15427 12189 15439 12192
rect 15381 12183 15439 12189
rect 15470 12180 15476 12192
rect 15528 12180 15534 12232
rect 16022 12220 16028 12232
rect 15983 12192 16028 12220
rect 16022 12180 16028 12192
rect 16080 12180 16086 12232
rect 13909 12155 13967 12161
rect 12084 12124 13814 12152
rect 1946 12084 1952 12096
rect 1907 12056 1952 12084
rect 1946 12044 1952 12056
rect 2004 12044 2010 12096
rect 2222 12084 2228 12096
rect 2183 12056 2228 12084
rect 2222 12044 2228 12056
rect 2280 12044 2286 12096
rect 4890 12044 4896 12096
rect 4948 12084 4954 12096
rect 5077 12087 5135 12093
rect 5077 12084 5089 12087
rect 4948 12056 5089 12084
rect 4948 12044 4954 12056
rect 5077 12053 5089 12056
rect 5123 12084 5135 12087
rect 5445 12087 5503 12093
rect 5445 12084 5457 12087
rect 5123 12056 5457 12084
rect 5123 12053 5135 12056
rect 5077 12047 5135 12053
rect 5445 12053 5457 12056
rect 5491 12084 5503 12087
rect 6546 12084 6552 12096
rect 5491 12056 6552 12084
rect 5491 12053 5503 12056
rect 5445 12047 5503 12053
rect 6546 12044 6552 12056
rect 6604 12044 6610 12096
rect 7285 12087 7343 12093
rect 7285 12053 7297 12087
rect 7331 12084 7343 12087
rect 7466 12084 7472 12096
rect 7331 12056 7472 12084
rect 7331 12053 7343 12056
rect 7285 12047 7343 12053
rect 7466 12044 7472 12056
rect 7524 12044 7530 12096
rect 7558 12044 7564 12096
rect 7616 12084 7622 12096
rect 7699 12087 7757 12093
rect 7699 12084 7711 12087
rect 7616 12056 7711 12084
rect 7616 12044 7622 12056
rect 7699 12053 7711 12056
rect 7745 12084 7757 12087
rect 10134 12084 10140 12096
rect 7745 12056 10140 12084
rect 7745 12053 7757 12056
rect 7699 12047 7757 12053
rect 10134 12044 10140 12056
rect 10192 12044 10198 12096
rect 13786 12084 13814 12124
rect 13909 12121 13921 12155
rect 13955 12152 13967 12155
rect 17451 12155 17509 12161
rect 17451 12152 17463 12155
rect 13955 12124 17463 12152
rect 13955 12121 13967 12124
rect 13909 12115 13967 12121
rect 17451 12121 17463 12124
rect 17497 12121 17509 12155
rect 17451 12115 17509 12121
rect 14458 12084 14464 12096
rect 13786 12056 14464 12084
rect 14458 12044 14464 12056
rect 14516 12044 14522 12096
rect 17218 12084 17224 12096
rect 17179 12056 17224 12084
rect 17218 12044 17224 12056
rect 17276 12044 17282 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 4249 11883 4307 11889
rect 4249 11849 4261 11883
rect 4295 11880 4307 11883
rect 4706 11880 4712 11892
rect 4295 11852 4712 11880
rect 4295 11849 4307 11852
rect 4249 11843 4307 11849
rect 4706 11840 4712 11852
rect 4764 11880 4770 11892
rect 4985 11883 5043 11889
rect 4985 11880 4997 11883
rect 4764 11852 4997 11880
rect 4764 11840 4770 11852
rect 4985 11849 4997 11852
rect 5031 11849 5043 11883
rect 7558 11880 7564 11892
rect 4985 11843 5043 11849
rect 7346 11852 7564 11880
rect 4890 11821 4896 11824
rect 4874 11815 4896 11821
rect 4874 11781 4886 11815
rect 4874 11775 4896 11781
rect 4890 11772 4896 11775
rect 4948 11772 4954 11824
rect 5166 11812 5172 11824
rect 5127 11784 5172 11812
rect 5166 11772 5172 11784
rect 5224 11772 5230 11824
rect 6546 11772 6552 11824
rect 6604 11812 6610 11824
rect 6914 11812 6920 11824
rect 6604 11784 6920 11812
rect 6604 11772 6610 11784
rect 6914 11772 6920 11784
rect 6972 11812 6978 11824
rect 7346 11821 7374 11852
rect 7558 11840 7564 11852
rect 7616 11840 7622 11892
rect 7834 11880 7840 11892
rect 7795 11852 7840 11880
rect 7834 11840 7840 11852
rect 7892 11840 7898 11892
rect 8110 11840 8116 11892
rect 8168 11880 8174 11892
rect 9217 11883 9275 11889
rect 9217 11880 9229 11883
rect 8168 11852 9229 11880
rect 8168 11840 8174 11852
rect 9217 11849 9229 11852
rect 9263 11849 9275 11883
rect 10134 11880 10140 11892
rect 10095 11852 10140 11880
rect 9217 11843 9275 11849
rect 10134 11840 10140 11852
rect 10192 11840 10198 11892
rect 10689 11883 10747 11889
rect 10689 11849 10701 11883
rect 10735 11880 10747 11883
rect 10778 11880 10784 11892
rect 10735 11852 10784 11880
rect 10735 11849 10747 11852
rect 10689 11843 10747 11849
rect 10778 11840 10784 11852
rect 10836 11840 10842 11892
rect 11422 11840 11428 11892
rect 11480 11880 11486 11892
rect 11885 11883 11943 11889
rect 11885 11880 11897 11883
rect 11480 11852 11897 11880
rect 11480 11840 11486 11852
rect 11885 11849 11897 11852
rect 11931 11880 11943 11883
rect 12802 11880 12808 11892
rect 11931 11852 12808 11880
rect 11931 11849 11943 11852
rect 11885 11843 11943 11849
rect 12802 11840 12808 11852
rect 12860 11840 12866 11892
rect 13541 11883 13599 11889
rect 13541 11849 13553 11883
rect 13587 11880 13599 11883
rect 14274 11880 14280 11892
rect 13587 11852 14280 11880
rect 13587 11849 13599 11852
rect 13541 11843 13599 11849
rect 14274 11840 14280 11852
rect 14332 11840 14338 11892
rect 7331 11815 7389 11821
rect 7331 11812 7343 11815
rect 6972 11784 7343 11812
rect 6972 11772 6978 11784
rect 7331 11781 7343 11784
rect 7377 11781 7389 11815
rect 7466 11812 7472 11824
rect 7427 11784 7472 11812
rect 7331 11775 7389 11781
rect 7466 11772 7472 11784
rect 7524 11772 7530 11824
rect 8846 11772 8852 11824
rect 8904 11821 8910 11824
rect 8904 11815 8953 11821
rect 8904 11781 8907 11815
rect 8941 11781 8953 11815
rect 8904 11775 8953 11781
rect 9033 11815 9091 11821
rect 9033 11781 9045 11815
rect 9079 11781 9091 11815
rect 9033 11775 9091 11781
rect 8904 11772 8910 11775
rect 2314 11704 2320 11756
rect 2372 11744 2378 11756
rect 2961 11747 3019 11753
rect 2961 11744 2973 11747
rect 2372 11716 2973 11744
rect 2372 11704 2378 11716
rect 2961 11713 2973 11716
rect 3007 11744 3019 11747
rect 4338 11744 4344 11756
rect 3007 11716 4344 11744
rect 3007 11713 3019 11716
rect 2961 11707 3019 11713
rect 4338 11704 4344 11716
rect 4396 11704 4402 11756
rect 5077 11747 5135 11753
rect 5077 11713 5089 11747
rect 5123 11713 5135 11747
rect 5077 11707 5135 11713
rect 1394 11676 1400 11688
rect 1355 11648 1400 11676
rect 1394 11636 1400 11648
rect 1452 11676 1458 11688
rect 1854 11676 1860 11688
rect 1452 11648 1860 11676
rect 1452 11636 1458 11648
rect 1854 11636 1860 11648
rect 1912 11636 1918 11688
rect 2498 11636 2504 11688
rect 2556 11676 2562 11688
rect 4617 11679 4675 11685
rect 4617 11676 4629 11679
rect 2556 11648 4629 11676
rect 2556 11636 2562 11648
rect 4617 11645 4629 11648
rect 4663 11676 4675 11679
rect 5092 11676 5120 11707
rect 7006 11704 7012 11756
rect 7064 11744 7070 11756
rect 7561 11747 7619 11753
rect 7561 11744 7573 11747
rect 7064 11716 7573 11744
rect 7064 11704 7070 11716
rect 7561 11713 7573 11716
rect 7607 11744 7619 11747
rect 8573 11747 8631 11753
rect 8573 11744 8585 11747
rect 7607 11716 8585 11744
rect 7607 11713 7619 11716
rect 7561 11707 7619 11713
rect 8573 11713 8585 11716
rect 8619 11713 8631 11747
rect 8573 11707 8631 11713
rect 5166 11676 5172 11688
rect 4663 11648 5172 11676
rect 4663 11645 4675 11648
rect 4617 11639 4675 11645
rect 5166 11636 5172 11648
rect 5224 11636 5230 11688
rect 8588 11676 8616 11707
rect 8754 11704 8760 11756
rect 8812 11744 8818 11756
rect 9048 11744 9076 11775
rect 13814 11772 13820 11824
rect 13872 11812 13878 11824
rect 19978 11812 19984 11824
rect 13872 11784 13917 11812
rect 14476 11784 19984 11812
rect 13872 11772 13878 11784
rect 14476 11756 14504 11784
rect 19978 11772 19984 11784
rect 20036 11772 20042 11824
rect 8812 11716 9076 11744
rect 9125 11747 9183 11753
rect 8812 11704 8818 11716
rect 9125 11713 9137 11747
rect 9171 11713 9183 11747
rect 14458 11744 14464 11756
rect 14371 11716 14464 11744
rect 9125 11707 9183 11713
rect 9140 11676 9168 11707
rect 14458 11704 14464 11716
rect 14516 11704 14522 11756
rect 14826 11704 14832 11756
rect 14884 11744 14890 11756
rect 15105 11747 15163 11753
rect 15105 11744 15117 11747
rect 14884 11716 15117 11744
rect 14884 11704 14890 11716
rect 15105 11713 15117 11716
rect 15151 11744 15163 11747
rect 15470 11744 15476 11756
rect 15151 11716 15476 11744
rect 15151 11713 15163 11716
rect 15105 11707 15163 11713
rect 15470 11704 15476 11716
rect 15528 11744 15534 11756
rect 16945 11747 17003 11753
rect 16945 11744 16957 11747
rect 15528 11716 16957 11744
rect 15528 11704 15534 11716
rect 16945 11713 16957 11716
rect 16991 11713 17003 11747
rect 16945 11707 17003 11713
rect 10778 11676 10784 11688
rect 8588 11648 9168 11676
rect 10739 11648 10784 11676
rect 10778 11636 10784 11648
rect 10836 11636 10842 11688
rect 11333 11679 11391 11685
rect 11333 11645 11345 11679
rect 11379 11676 11391 11679
rect 12158 11676 12164 11688
rect 11379 11648 12164 11676
rect 11379 11645 11391 11648
rect 11333 11639 11391 11645
rect 12158 11636 12164 11648
rect 12216 11636 12222 11688
rect 12618 11676 12624 11688
rect 12579 11648 12624 11676
rect 12618 11636 12624 11648
rect 12676 11636 12682 11688
rect 16025 11679 16083 11685
rect 16025 11645 16037 11679
rect 16071 11645 16083 11679
rect 16025 11639 16083 11645
rect 2869 11611 2927 11617
rect 2869 11577 2881 11611
rect 2915 11608 2927 11611
rect 2958 11608 2964 11620
rect 2915 11580 2964 11608
rect 2915 11577 2927 11580
rect 2869 11571 2927 11577
rect 2958 11568 2964 11580
rect 3016 11608 3022 11620
rect 3282 11611 3340 11617
rect 3282 11608 3294 11611
rect 3016 11580 3294 11608
rect 3016 11568 3022 11580
rect 3282 11577 3294 11580
rect 3328 11608 3340 11611
rect 3328 11580 4476 11608
rect 3328 11577 3340 11580
rect 3282 11571 3340 11577
rect 106 11500 112 11552
rect 164 11540 170 11552
rect 1581 11543 1639 11549
rect 1581 11540 1593 11543
rect 164 11512 1593 11540
rect 164 11500 170 11512
rect 1581 11509 1593 11512
rect 1627 11509 1639 11543
rect 2038 11540 2044 11552
rect 1999 11512 2044 11540
rect 1581 11503 1639 11509
rect 2038 11500 2044 11512
rect 2096 11500 2102 11552
rect 2406 11540 2412 11552
rect 2367 11512 2412 11540
rect 2406 11500 2412 11512
rect 2464 11500 2470 11552
rect 3418 11500 3424 11552
rect 3476 11540 3482 11552
rect 3881 11543 3939 11549
rect 3881 11540 3893 11543
rect 3476 11512 3893 11540
rect 3476 11500 3482 11512
rect 3881 11509 3893 11512
rect 3927 11509 3939 11543
rect 4448 11540 4476 11580
rect 4522 11568 4528 11620
rect 4580 11608 4586 11620
rect 4709 11611 4767 11617
rect 4709 11608 4721 11611
rect 4580 11580 4721 11608
rect 4580 11568 4586 11580
rect 4709 11577 4721 11580
rect 4755 11577 4767 11611
rect 4709 11571 4767 11577
rect 5350 11568 5356 11620
rect 5408 11608 5414 11620
rect 6549 11611 6607 11617
rect 6549 11608 6561 11611
rect 5408 11580 6561 11608
rect 5408 11568 5414 11580
rect 6549 11577 6561 11580
rect 6595 11608 6607 11611
rect 7193 11611 7251 11617
rect 7193 11608 7205 11611
rect 6595 11580 7205 11608
rect 6595 11577 6607 11580
rect 6549 11571 6607 11577
rect 7193 11577 7205 11580
rect 7239 11608 7251 11611
rect 7282 11608 7288 11620
rect 7239 11580 7288 11608
rect 7239 11577 7251 11580
rect 7193 11571 7251 11577
rect 7282 11568 7288 11580
rect 7340 11568 7346 11620
rect 8570 11568 8576 11620
rect 8628 11608 8634 11620
rect 8757 11611 8815 11617
rect 8757 11608 8769 11611
rect 8628 11580 8769 11608
rect 8628 11568 8634 11580
rect 8757 11577 8769 11580
rect 8803 11577 8815 11611
rect 8757 11571 8815 11577
rect 11517 11611 11575 11617
rect 11517 11577 11529 11611
rect 11563 11608 11575 11611
rect 12802 11608 12808 11620
rect 11563 11580 12808 11608
rect 11563 11577 11575 11580
rect 11517 11571 11575 11577
rect 12802 11568 12808 11580
rect 12860 11568 12866 11620
rect 12983 11611 13041 11617
rect 12983 11577 12995 11611
rect 13029 11577 13041 11611
rect 12983 11571 13041 11577
rect 14553 11611 14611 11617
rect 14553 11577 14565 11611
rect 14599 11577 14611 11611
rect 14553 11571 14611 11577
rect 5813 11543 5871 11549
rect 5813 11540 5825 11543
rect 4448 11512 5825 11540
rect 3881 11503 3939 11509
rect 5813 11509 5825 11512
rect 5859 11540 5871 11543
rect 5994 11540 6000 11552
rect 5859 11512 6000 11540
rect 5859 11509 5871 11512
rect 5813 11503 5871 11509
rect 5994 11500 6000 11512
rect 6052 11500 6058 11552
rect 6178 11540 6184 11552
rect 6139 11512 6184 11540
rect 6178 11500 6184 11512
rect 6236 11500 6242 11552
rect 7006 11540 7012 11552
rect 6967 11512 7012 11540
rect 7006 11500 7012 11512
rect 7064 11500 7070 11552
rect 7650 11500 7656 11552
rect 7708 11540 7714 11552
rect 8205 11543 8263 11549
rect 8205 11540 8217 11543
rect 7708 11512 8217 11540
rect 7708 11500 7714 11512
rect 8205 11509 8217 11512
rect 8251 11509 8263 11543
rect 8205 11503 8263 11509
rect 9861 11543 9919 11549
rect 9861 11509 9873 11543
rect 9907 11540 9919 11543
rect 9950 11540 9956 11552
rect 9907 11512 9956 11540
rect 9907 11509 9919 11512
rect 9861 11503 9919 11509
rect 9950 11500 9956 11512
rect 10008 11500 10014 11552
rect 12250 11540 12256 11552
rect 12163 11512 12256 11540
rect 12250 11500 12256 11512
rect 12308 11540 12314 11552
rect 13004 11540 13032 11571
rect 13446 11540 13452 11552
rect 12308 11512 13452 11540
rect 12308 11500 12314 11512
rect 13446 11500 13452 11512
rect 13504 11500 13510 11552
rect 14274 11500 14280 11552
rect 14332 11540 14338 11552
rect 14568 11540 14596 11571
rect 15470 11568 15476 11620
rect 15528 11608 15534 11620
rect 15933 11611 15991 11617
rect 15933 11608 15945 11611
rect 15528 11580 15945 11608
rect 15528 11568 15534 11580
rect 15933 11577 15945 11580
rect 15979 11577 15991 11611
rect 15933 11571 15991 11577
rect 14332 11512 14596 11540
rect 14332 11500 14338 11512
rect 15286 11500 15292 11552
rect 15344 11540 15350 11552
rect 15381 11543 15439 11549
rect 15381 11540 15393 11543
rect 15344 11512 15393 11540
rect 15344 11500 15350 11512
rect 15381 11509 15393 11512
rect 15427 11540 15439 11543
rect 15749 11543 15807 11549
rect 15749 11540 15761 11543
rect 15427 11512 15761 11540
rect 15427 11509 15439 11512
rect 15381 11503 15439 11509
rect 15749 11509 15761 11512
rect 15795 11540 15807 11543
rect 16040 11540 16068 11639
rect 15795 11512 16068 11540
rect 15795 11509 15807 11512
rect 15749 11503 15807 11509
rect 17218 11500 17224 11552
rect 17276 11540 17282 11552
rect 17405 11543 17463 11549
rect 17405 11540 17417 11543
rect 17276 11512 17417 11540
rect 17276 11500 17282 11512
rect 17405 11509 17417 11512
rect 17451 11540 17463 11543
rect 19426 11540 19432 11552
rect 17451 11512 19432 11540
rect 17451 11509 17463 11512
rect 17405 11503 17463 11509
rect 19426 11500 19432 11512
rect 19484 11500 19490 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1397 11339 1455 11345
rect 1397 11305 1409 11339
rect 1443 11336 1455 11339
rect 2222 11336 2228 11348
rect 1443 11308 2228 11336
rect 1443 11305 1455 11308
rect 1397 11299 1455 11305
rect 2222 11296 2228 11308
rect 2280 11296 2286 11348
rect 4522 11296 4528 11348
rect 4580 11336 4586 11348
rect 4709 11339 4767 11345
rect 4709 11336 4721 11339
rect 4580 11308 4721 11336
rect 4580 11296 4586 11308
rect 4709 11305 4721 11308
rect 4755 11305 4767 11339
rect 4709 11299 4767 11305
rect 2406 11268 2412 11280
rect 2367 11240 2412 11268
rect 2406 11228 2412 11240
rect 2464 11228 2470 11280
rect 4724 11268 4752 11299
rect 4982 11296 4988 11348
rect 5040 11336 5046 11348
rect 5537 11339 5595 11345
rect 5537 11336 5549 11339
rect 5040 11308 5549 11336
rect 5040 11296 5046 11308
rect 5537 11305 5549 11308
rect 5583 11305 5595 11339
rect 7926 11336 7932 11348
rect 7887 11308 7932 11336
rect 5537 11299 5595 11305
rect 7926 11296 7932 11308
rect 7984 11296 7990 11348
rect 8846 11296 8852 11348
rect 8904 11336 8910 11348
rect 9125 11339 9183 11345
rect 9125 11336 9137 11339
rect 8904 11308 9137 11336
rect 8904 11296 8910 11308
rect 9125 11305 9137 11308
rect 9171 11305 9183 11339
rect 9125 11299 9183 11305
rect 11241 11339 11299 11345
rect 11241 11305 11253 11339
rect 11287 11336 11299 11339
rect 11330 11336 11336 11348
rect 11287 11308 11336 11336
rect 11287 11305 11299 11308
rect 11241 11299 11299 11305
rect 7098 11268 7104 11280
rect 4724 11240 7104 11268
rect 7098 11228 7104 11240
rect 7156 11268 7162 11280
rect 8297 11271 8355 11277
rect 8297 11268 8309 11271
rect 7156 11240 8309 11268
rect 7156 11228 7162 11240
rect 8297 11237 8309 11240
rect 8343 11237 8355 11271
rect 9140 11268 9168 11299
rect 11330 11296 11336 11308
rect 11388 11296 11394 11348
rect 13817 11339 13875 11345
rect 13817 11305 13829 11339
rect 13863 11336 13875 11339
rect 15286 11336 15292 11348
rect 13863 11308 15292 11336
rect 13863 11305 13875 11308
rect 13817 11299 13875 11305
rect 15286 11296 15292 11308
rect 15344 11296 15350 11348
rect 12069 11271 12127 11277
rect 9140 11240 9867 11268
rect 8297 11231 8355 11237
rect 3053 11203 3111 11209
rect 3053 11169 3065 11203
rect 3099 11200 3111 11203
rect 3418 11200 3424 11212
rect 3099 11172 3424 11200
rect 3099 11169 3111 11172
rect 3053 11163 3111 11169
rect 3418 11160 3424 11172
rect 3476 11160 3482 11212
rect 4893 11203 4951 11209
rect 4893 11169 4905 11203
rect 4939 11200 4951 11203
rect 5350 11200 5356 11212
rect 4939 11172 5356 11200
rect 4939 11169 4951 11172
rect 4893 11163 4951 11169
rect 5350 11160 5356 11172
rect 5408 11160 5414 11212
rect 6822 11160 6828 11212
rect 6880 11200 6886 11212
rect 7190 11200 7196 11212
rect 6880 11172 7196 11200
rect 6880 11160 6886 11172
rect 7190 11160 7196 11172
rect 7248 11200 7254 11212
rect 7285 11203 7343 11209
rect 7285 11200 7297 11203
rect 7248 11172 7297 11200
rect 7248 11160 7254 11172
rect 7285 11169 7297 11172
rect 7331 11200 7343 11203
rect 8662 11200 8668 11212
rect 7331 11172 8668 11200
rect 7331 11169 7343 11172
rect 7285 11163 7343 11169
rect 8662 11160 8668 11172
rect 8720 11200 8726 11212
rect 9677 11203 9735 11209
rect 9677 11200 9689 11203
rect 8720 11172 9689 11200
rect 8720 11160 8726 11172
rect 9677 11169 9689 11172
rect 9723 11169 9735 11203
rect 9677 11163 9735 11169
rect 5166 11092 5172 11144
rect 5224 11132 5230 11144
rect 5261 11135 5319 11141
rect 5261 11132 5273 11135
rect 5224 11104 5273 11132
rect 5224 11092 5230 11104
rect 5261 11101 5273 11104
rect 5307 11101 5319 11135
rect 5261 11095 5319 11101
rect 5442 11092 5448 11144
rect 5500 11132 5506 11144
rect 6178 11132 6184 11144
rect 5500 11104 6184 11132
rect 5500 11092 5506 11104
rect 6178 11092 6184 11104
rect 6236 11132 6242 11144
rect 6365 11135 6423 11141
rect 6365 11132 6377 11135
rect 6236 11104 6377 11132
rect 6236 11092 6242 11104
rect 6365 11101 6377 11104
rect 6411 11132 6423 11135
rect 7653 11135 7711 11141
rect 7653 11132 7665 11135
rect 6411 11104 7665 11132
rect 6411 11101 6423 11104
rect 6365 11095 6423 11101
rect 7653 11101 7665 11104
rect 7699 11132 7711 11135
rect 7926 11132 7932 11144
rect 7699 11104 7932 11132
rect 7699 11101 7711 11104
rect 7653 11095 7711 11101
rect 7926 11092 7932 11104
rect 7984 11092 7990 11144
rect 9839 11141 9867 11240
rect 12069 11237 12081 11271
rect 12115 11268 12127 11271
rect 12345 11271 12403 11277
rect 12345 11268 12357 11271
rect 12115 11240 12357 11268
rect 12115 11237 12127 11240
rect 12069 11231 12127 11237
rect 12345 11237 12357 11240
rect 12391 11268 12403 11271
rect 12618 11268 12624 11280
rect 12391 11240 12624 11268
rect 12391 11237 12403 11240
rect 12345 11231 12403 11237
rect 12618 11228 12624 11240
rect 12676 11228 12682 11280
rect 13259 11271 13317 11277
rect 13259 11237 13271 11271
rect 13305 11268 13317 11271
rect 13446 11268 13452 11280
rect 13305 11240 13452 11268
rect 13305 11237 13317 11240
rect 13259 11231 13317 11237
rect 13446 11228 13452 11240
rect 13504 11228 13510 11280
rect 14458 11268 14464 11280
rect 14419 11240 14464 11268
rect 14458 11228 14464 11240
rect 14516 11228 14522 11280
rect 15378 11268 15384 11280
rect 15339 11240 15384 11268
rect 15378 11228 15384 11240
rect 15436 11228 15442 11280
rect 15470 11228 15476 11280
rect 15528 11268 15534 11280
rect 16022 11268 16028 11280
rect 15528 11240 15573 11268
rect 15983 11240 16028 11268
rect 15528 11228 15534 11240
rect 16022 11228 16028 11240
rect 16080 11268 16086 11280
rect 16080 11240 16931 11268
rect 16080 11228 16086 11240
rect 16903 11212 16931 11240
rect 11422 11200 11428 11212
rect 11383 11172 11428 11200
rect 11422 11160 11428 11172
rect 11480 11160 11486 11212
rect 11885 11203 11943 11209
rect 11885 11169 11897 11203
rect 11931 11200 11943 11203
rect 12158 11200 12164 11212
rect 11931 11172 12164 11200
rect 11931 11169 11943 11172
rect 11885 11163 11943 11169
rect 9824 11135 9882 11141
rect 9824 11101 9836 11135
rect 9870 11101 9882 11135
rect 10042 11132 10048 11144
rect 10003 11104 10048 11132
rect 9824 11095 9882 11101
rect 10042 11092 10048 11104
rect 10100 11092 10106 11144
rect 10413 11135 10471 11141
rect 10413 11101 10425 11135
rect 10459 11132 10471 11135
rect 10873 11135 10931 11141
rect 10873 11132 10885 11135
rect 10459 11104 10885 11132
rect 10459 11101 10471 11104
rect 10413 11095 10471 11101
rect 10873 11101 10885 11104
rect 10919 11132 10931 11135
rect 11900 11132 11928 11163
rect 12158 11160 12164 11172
rect 12216 11160 12222 11212
rect 12802 11160 12808 11212
rect 12860 11200 12866 11212
rect 12897 11203 12955 11209
rect 12897 11200 12909 11203
rect 12860 11172 12909 11200
rect 12860 11160 12866 11172
rect 12897 11169 12909 11172
rect 12943 11169 12955 11203
rect 16850 11200 16856 11212
rect 16908 11209 16931 11212
rect 16908 11203 16946 11209
rect 16798 11172 16856 11200
rect 12897 11163 12955 11169
rect 16850 11160 16856 11172
rect 16934 11169 16946 11203
rect 16908 11163 16946 11169
rect 16908 11160 16914 11163
rect 10919 11104 11928 11132
rect 10919 11101 10931 11104
rect 10873 11095 10931 11101
rect 14 11024 20 11076
rect 72 11064 78 11076
rect 2406 11064 2412 11076
rect 72 11036 2412 11064
rect 72 11024 78 11036
rect 2406 11024 2412 11036
rect 2464 11024 2470 11076
rect 3697 11067 3755 11073
rect 3697 11033 3709 11067
rect 3743 11064 3755 11067
rect 3878 11064 3884 11076
rect 3743 11036 3884 11064
rect 3743 11033 3755 11036
rect 3697 11027 3755 11033
rect 3878 11024 3884 11036
rect 3936 11064 3942 11076
rect 4154 11064 4160 11076
rect 3936 11036 4160 11064
rect 3936 11024 3942 11036
rect 4154 11024 4160 11036
rect 4212 11064 4218 11076
rect 4706 11064 4712 11076
rect 4212 11036 4712 11064
rect 4212 11024 4218 11036
rect 4706 11024 4712 11036
rect 4764 11064 4770 11076
rect 6270 11064 6276 11076
rect 4764 11036 6276 11064
rect 4764 11024 4770 11036
rect 2133 10999 2191 11005
rect 2133 10965 2145 10999
rect 2179 10996 2191 10999
rect 2222 10996 2228 11008
rect 2179 10968 2228 10996
rect 2179 10965 2191 10968
rect 2133 10959 2191 10965
rect 2222 10956 2228 10968
rect 2280 10996 2286 11008
rect 2774 10996 2780 11008
rect 2280 10968 2780 10996
rect 2280 10956 2286 10968
rect 2774 10956 2780 10968
rect 2832 10956 2838 11008
rect 4338 10996 4344 11008
rect 4251 10968 4344 10996
rect 4338 10956 4344 10968
rect 4396 10956 4402 11008
rect 4890 10956 4896 11008
rect 4948 10996 4954 11008
rect 5184 11005 5212 11036
rect 6270 11024 6276 11036
rect 6328 11064 6334 11076
rect 6825 11067 6883 11073
rect 6825 11064 6837 11067
rect 6328 11036 6837 11064
rect 6328 11024 6334 11036
rect 6825 11033 6837 11036
rect 6871 11064 6883 11067
rect 7558 11064 7564 11076
rect 6871 11036 7564 11064
rect 6871 11033 6883 11036
rect 6825 11027 6883 11033
rect 7558 11024 7564 11036
rect 7616 11064 7622 11076
rect 9950 11064 9956 11076
rect 7616 11036 9956 11064
rect 7616 11024 7622 11036
rect 9950 11024 9956 11036
rect 10008 11024 10014 11076
rect 5031 10999 5089 11005
rect 5031 10996 5043 10999
rect 4948 10968 5043 10996
rect 4948 10956 4954 10968
rect 5031 10965 5043 10968
rect 5077 10965 5089 10999
rect 5031 10959 5089 10965
rect 5169 10999 5227 11005
rect 5169 10965 5181 10999
rect 5215 10965 5227 10999
rect 5994 10996 6000 11008
rect 5955 10968 6000 10996
rect 5169 10959 5227 10965
rect 5994 10956 6000 10968
rect 6052 10956 6058 11008
rect 7190 10956 7196 11008
rect 7248 10996 7254 11008
rect 7423 10999 7481 11005
rect 7423 10996 7435 10999
rect 7248 10968 7435 10996
rect 7248 10956 7254 10968
rect 7423 10965 7435 10968
rect 7469 10965 7481 10999
rect 8754 10996 8760 11008
rect 8715 10968 8760 10996
rect 7423 10959 7481 10965
rect 8754 10956 8760 10968
rect 8812 10956 8818 11008
rect 12805 10999 12863 11005
rect 12805 10965 12817 10999
rect 12851 10996 12863 10999
rect 13078 10996 13084 11008
rect 12851 10968 13084 10996
rect 12851 10965 12863 10968
rect 12805 10959 12863 10965
rect 13078 10956 13084 10968
rect 13136 10956 13142 11008
rect 16991 10999 17049 11005
rect 16991 10965 17003 10999
rect 17037 10996 17049 10999
rect 20254 10996 20260 11008
rect 17037 10968 20260 10996
rect 17037 10965 17049 10968
rect 16991 10959 17049 10965
rect 20254 10956 20260 10968
rect 20312 10956 20318 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1946 10752 1952 10804
rect 2004 10792 2010 10804
rect 2501 10795 2559 10801
rect 2501 10792 2513 10795
rect 2004 10764 2513 10792
rect 2004 10752 2010 10764
rect 2501 10761 2513 10764
rect 2547 10761 2559 10795
rect 3878 10792 3884 10804
rect 3839 10764 3884 10792
rect 2501 10755 2559 10761
rect 3878 10752 3884 10764
rect 3936 10752 3942 10804
rect 6549 10795 6607 10801
rect 6549 10792 6561 10795
rect 3988 10764 6561 10792
rect 2222 10733 2228 10736
rect 2206 10727 2228 10733
rect 2206 10693 2218 10727
rect 2206 10687 2228 10693
rect 2222 10684 2228 10687
rect 2280 10684 2286 10736
rect 2317 10727 2375 10733
rect 2317 10693 2329 10727
rect 2363 10724 2375 10727
rect 2363 10696 2728 10724
rect 2363 10693 2375 10696
rect 2317 10687 2375 10693
rect 2406 10656 2412 10668
rect 2367 10628 2412 10656
rect 2406 10616 2412 10628
rect 2464 10616 2470 10668
rect 1949 10591 2007 10597
rect 1949 10557 1961 10591
rect 1995 10588 2007 10591
rect 2700 10588 2728 10696
rect 3326 10684 3332 10736
rect 3384 10724 3390 10736
rect 3743 10727 3801 10733
rect 3743 10724 3755 10727
rect 3384 10696 3755 10724
rect 3384 10684 3390 10696
rect 3743 10693 3755 10696
rect 3789 10724 3801 10727
rect 3988 10724 4016 10764
rect 6549 10761 6561 10764
rect 6595 10792 6607 10795
rect 7190 10792 7196 10804
rect 6595 10764 7196 10792
rect 6595 10761 6607 10764
rect 6549 10755 6607 10761
rect 7190 10752 7196 10764
rect 7248 10752 7254 10804
rect 8754 10752 8760 10804
rect 8812 10792 8818 10804
rect 9033 10795 9091 10801
rect 9033 10792 9045 10795
rect 8812 10764 9045 10792
rect 8812 10752 8818 10764
rect 9033 10761 9045 10764
rect 9079 10761 9091 10795
rect 9033 10755 9091 10761
rect 9401 10795 9459 10801
rect 9401 10761 9413 10795
rect 9447 10792 9459 10795
rect 9582 10792 9588 10804
rect 9447 10764 9588 10792
rect 9447 10761 9459 10764
rect 9401 10755 9459 10761
rect 9582 10752 9588 10764
rect 9640 10752 9646 10804
rect 12158 10792 12164 10804
rect 12119 10764 12164 10792
rect 12158 10752 12164 10764
rect 12216 10752 12222 10804
rect 14182 10792 14188 10804
rect 14143 10764 14188 10792
rect 14182 10752 14188 10764
rect 14240 10752 14246 10804
rect 15378 10752 15384 10804
rect 15436 10792 15442 10804
rect 15657 10795 15715 10801
rect 15657 10792 15669 10795
rect 15436 10764 15669 10792
rect 15436 10752 15442 10764
rect 15657 10761 15669 10764
rect 15703 10761 15715 10795
rect 15657 10755 15715 10761
rect 15746 10752 15752 10804
rect 15804 10792 15810 10804
rect 15979 10795 16037 10801
rect 15979 10792 15991 10795
rect 15804 10764 15991 10792
rect 15804 10752 15810 10764
rect 15979 10761 15991 10764
rect 16025 10761 16037 10795
rect 16850 10792 16856 10804
rect 16811 10764 16856 10792
rect 15979 10755 16037 10761
rect 16850 10752 16856 10764
rect 16908 10752 16914 10804
rect 24765 10795 24823 10801
rect 24765 10761 24777 10795
rect 24811 10792 24823 10795
rect 25130 10792 25136 10804
rect 24811 10764 25136 10792
rect 24811 10761 24823 10764
rect 24765 10755 24823 10761
rect 25130 10752 25136 10764
rect 25188 10752 25194 10804
rect 3789 10696 4016 10724
rect 4985 10727 5043 10733
rect 3789 10693 3801 10696
rect 3743 10687 3801 10693
rect 4985 10693 4997 10727
rect 5031 10724 5043 10727
rect 5166 10724 5172 10736
rect 5031 10696 5172 10724
rect 5031 10693 5043 10696
rect 4985 10687 5043 10693
rect 5166 10684 5172 10696
rect 5224 10684 5230 10736
rect 6270 10724 6276 10736
rect 6231 10696 6276 10724
rect 6270 10684 6276 10696
rect 6328 10684 6334 10736
rect 6638 10684 6644 10736
rect 6696 10724 6702 10736
rect 6914 10724 6920 10736
rect 6696 10696 6920 10724
rect 6696 10684 6702 10696
rect 6914 10684 6920 10696
rect 6972 10724 6978 10736
rect 7331 10727 7389 10733
rect 7331 10724 7343 10727
rect 6972 10696 7343 10724
rect 6972 10684 6978 10696
rect 7331 10693 7343 10696
rect 7377 10693 7389 10727
rect 7466 10724 7472 10736
rect 7427 10696 7472 10724
rect 7331 10687 7389 10693
rect 7466 10684 7472 10696
rect 7524 10684 7530 10736
rect 7742 10684 7748 10736
rect 7800 10724 7806 10736
rect 8297 10727 8355 10733
rect 8297 10724 8309 10727
rect 7800 10696 8309 10724
rect 7800 10684 7806 10696
rect 8297 10693 8309 10696
rect 8343 10724 8355 10727
rect 8846 10724 8852 10736
rect 8343 10696 8852 10724
rect 8343 10693 8355 10696
rect 8297 10687 8355 10693
rect 8846 10684 8852 10696
rect 8904 10733 8910 10736
rect 8904 10727 8953 10733
rect 8904 10693 8907 10727
rect 8941 10724 8953 10727
rect 10137 10727 10195 10733
rect 10137 10724 10149 10727
rect 8941 10696 10149 10724
rect 8941 10693 8953 10696
rect 8904 10687 8953 10693
rect 10137 10693 10149 10696
rect 10183 10693 10195 10727
rect 10137 10687 10195 10693
rect 8904 10684 8910 10687
rect 14826 10684 14832 10736
rect 14884 10724 14890 10736
rect 14921 10727 14979 10733
rect 14921 10724 14933 10727
rect 14884 10696 14933 10724
rect 14884 10684 14890 10696
rect 14921 10693 14933 10696
rect 14967 10693 14979 10727
rect 14921 10687 14979 10693
rect 15289 10727 15347 10733
rect 15289 10693 15301 10727
rect 15335 10724 15347 10727
rect 15470 10724 15476 10736
rect 15335 10696 15476 10724
rect 15335 10693 15347 10696
rect 15289 10687 15347 10693
rect 15470 10684 15476 10696
rect 15528 10684 15534 10736
rect 3145 10659 3203 10665
rect 3145 10625 3157 10659
rect 3191 10656 3203 10659
rect 3973 10659 4031 10665
rect 3973 10656 3985 10659
rect 3191 10628 3985 10656
rect 3191 10625 3203 10628
rect 3145 10619 3203 10625
rect 3973 10625 3985 10628
rect 4019 10656 4031 10659
rect 4801 10659 4859 10665
rect 4801 10656 4813 10659
rect 4019 10628 4813 10656
rect 4019 10625 4031 10628
rect 3973 10619 4031 10625
rect 4801 10625 4813 10628
rect 4847 10625 4859 10659
rect 4801 10619 4859 10625
rect 4062 10588 4068 10600
rect 1995 10560 4068 10588
rect 1995 10557 2007 10560
rect 1949 10551 2007 10557
rect 4062 10548 4068 10560
rect 4120 10548 4126 10600
rect 5184 10588 5212 10684
rect 7006 10616 7012 10668
rect 7064 10656 7070 10668
rect 7561 10659 7619 10665
rect 7561 10656 7573 10659
rect 7064 10628 7573 10656
rect 7064 10616 7070 10628
rect 7561 10625 7573 10628
rect 7607 10656 7619 10659
rect 8573 10659 8631 10665
rect 8573 10656 8585 10659
rect 7607 10628 8585 10656
rect 7607 10625 7619 10628
rect 7561 10619 7619 10625
rect 8573 10625 8585 10628
rect 8619 10656 8631 10659
rect 9125 10659 9183 10665
rect 9125 10656 9137 10659
rect 8619 10628 9137 10656
rect 8619 10625 8631 10628
rect 8573 10619 8631 10625
rect 9125 10625 9137 10628
rect 9171 10656 9183 10659
rect 9769 10659 9827 10665
rect 9769 10656 9781 10659
rect 9171 10628 9781 10656
rect 9171 10625 9183 10628
rect 9125 10619 9183 10625
rect 9769 10625 9781 10628
rect 9815 10656 9827 10659
rect 10042 10656 10048 10668
rect 9815 10628 10048 10656
rect 9815 10625 9827 10628
rect 9769 10619 9827 10625
rect 10042 10616 10048 10628
rect 10100 10616 10106 10668
rect 13262 10656 13268 10668
rect 13223 10628 13268 10656
rect 13262 10616 13268 10628
rect 13320 10656 13326 10668
rect 13320 10628 15919 10656
rect 13320 10616 13326 10628
rect 5261 10591 5319 10597
rect 5261 10588 5273 10591
rect 5184 10560 5273 10588
rect 5261 10557 5273 10560
rect 5307 10557 5319 10591
rect 5261 10551 5319 10557
rect 7098 10548 7104 10600
rect 7156 10588 7162 10600
rect 7193 10591 7251 10597
rect 7193 10588 7205 10591
rect 7156 10560 7205 10588
rect 7156 10548 7162 10560
rect 7193 10557 7205 10560
rect 7239 10557 7251 10591
rect 7193 10551 7251 10557
rect 8662 10548 8668 10600
rect 8720 10588 8726 10600
rect 8757 10591 8815 10597
rect 8757 10588 8769 10591
rect 8720 10560 8769 10588
rect 8720 10548 8726 10560
rect 8757 10557 8769 10560
rect 8803 10557 8815 10591
rect 8757 10551 8815 10557
rect 10781 10591 10839 10597
rect 10781 10557 10793 10591
rect 10827 10557 10839 10591
rect 11330 10588 11336 10600
rect 11291 10560 11336 10588
rect 10781 10551 10839 10557
rect 2038 10520 2044 10532
rect 1999 10492 2044 10520
rect 2038 10480 2044 10492
rect 2096 10480 2102 10532
rect 3605 10523 3663 10529
rect 3605 10489 3617 10523
rect 3651 10520 3663 10523
rect 4341 10523 4399 10529
rect 3651 10492 3832 10520
rect 3651 10489 3663 10492
rect 3605 10483 3663 10489
rect 3804 10464 3832 10492
rect 4341 10489 4353 10523
rect 4387 10520 4399 10523
rect 6914 10520 6920 10532
rect 4387 10492 6920 10520
rect 4387 10489 4399 10492
rect 4341 10483 4399 10489
rect 6914 10480 6920 10492
rect 6972 10480 6978 10532
rect 3326 10412 3332 10464
rect 3384 10452 3390 10464
rect 3421 10455 3479 10461
rect 3421 10452 3433 10455
rect 3384 10424 3433 10452
rect 3384 10412 3390 10424
rect 3421 10421 3433 10424
rect 3467 10421 3479 10455
rect 3421 10415 3479 10421
rect 3786 10412 3792 10464
rect 3844 10452 3850 10464
rect 4614 10452 4620 10464
rect 3844 10424 4620 10452
rect 3844 10412 3850 10424
rect 4614 10412 4620 10424
rect 4672 10412 4678 10464
rect 4801 10455 4859 10461
rect 4801 10421 4813 10455
rect 4847 10452 4859 10455
rect 5442 10452 5448 10464
rect 4847 10424 5448 10452
rect 4847 10421 4859 10424
rect 4801 10415 4859 10421
rect 5442 10412 5448 10424
rect 5500 10412 5506 10464
rect 5534 10412 5540 10464
rect 5592 10452 5598 10464
rect 5629 10455 5687 10461
rect 5629 10452 5641 10455
rect 5592 10424 5641 10452
rect 5592 10412 5598 10424
rect 5629 10421 5641 10424
rect 5675 10421 5687 10455
rect 7006 10452 7012 10464
rect 6967 10424 7012 10452
rect 5629 10415 5687 10421
rect 7006 10412 7012 10424
rect 7064 10412 7070 10464
rect 7834 10452 7840 10464
rect 7795 10424 7840 10452
rect 7834 10412 7840 10424
rect 7892 10412 7898 10464
rect 10689 10455 10747 10461
rect 10689 10421 10701 10455
rect 10735 10452 10747 10455
rect 10796 10452 10824 10551
rect 11330 10548 11336 10560
rect 11388 10548 11394 10600
rect 15891 10597 15919 10628
rect 15876 10591 15934 10597
rect 15876 10557 15888 10591
rect 15922 10588 15934 10591
rect 16301 10591 16359 10597
rect 16301 10588 16313 10591
rect 15922 10560 16313 10588
rect 15922 10557 15934 10560
rect 15876 10551 15934 10557
rect 16301 10557 16313 10560
rect 16347 10557 16359 10591
rect 16301 10551 16359 10557
rect 24118 10548 24124 10600
rect 24176 10588 24182 10600
rect 24581 10591 24639 10597
rect 24581 10588 24593 10591
rect 24176 10560 24593 10588
rect 24176 10548 24182 10560
rect 24581 10557 24593 10560
rect 24627 10588 24639 10591
rect 25133 10591 25191 10597
rect 25133 10588 25145 10591
rect 24627 10560 25145 10588
rect 24627 10557 24639 10560
rect 24581 10551 24639 10557
rect 25133 10557 25145 10560
rect 25179 10557 25191 10591
rect 25133 10551 25191 10557
rect 11517 10523 11575 10529
rect 11517 10489 11529 10523
rect 11563 10520 11575 10523
rect 12618 10520 12624 10532
rect 11563 10492 12624 10520
rect 11563 10489 11575 10492
rect 11517 10483 11575 10489
rect 12618 10480 12624 10492
rect 12676 10480 12682 10532
rect 12805 10523 12863 10529
rect 12805 10489 12817 10523
rect 12851 10489 12863 10523
rect 12805 10483 12863 10489
rect 12897 10523 12955 10529
rect 12897 10489 12909 10523
rect 12943 10520 12955 10523
rect 13078 10520 13084 10532
rect 12943 10492 13084 10520
rect 12943 10489 12955 10492
rect 12897 10483 12955 10489
rect 10870 10452 10876 10464
rect 10735 10424 10876 10452
rect 10735 10421 10747 10424
rect 10689 10415 10747 10421
rect 10870 10412 10876 10424
rect 10928 10452 10934 10464
rect 11422 10452 11428 10464
rect 10928 10424 11428 10452
rect 10928 10412 10934 10424
rect 11422 10412 11428 10424
rect 11480 10452 11486 10464
rect 11793 10455 11851 10461
rect 11793 10452 11805 10455
rect 11480 10424 11805 10452
rect 11480 10412 11486 10424
rect 11793 10421 11805 10424
rect 11839 10421 11851 10455
rect 11793 10415 11851 10421
rect 12710 10412 12716 10464
rect 12768 10452 12774 10464
rect 12820 10452 12848 10483
rect 13078 10480 13084 10492
rect 13136 10480 13142 10532
rect 14366 10520 14372 10532
rect 14327 10492 14372 10520
rect 14366 10480 14372 10492
rect 14424 10480 14430 10532
rect 14461 10523 14519 10529
rect 14461 10489 14473 10523
rect 14507 10489 14519 10523
rect 14461 10483 14519 10489
rect 12768 10424 12848 10452
rect 12768 10412 12774 10424
rect 13446 10412 13452 10464
rect 13504 10452 13510 10464
rect 13725 10455 13783 10461
rect 13725 10452 13737 10455
rect 13504 10424 13737 10452
rect 13504 10412 13510 10424
rect 13725 10421 13737 10424
rect 13771 10421 13783 10455
rect 13725 10415 13783 10421
rect 14182 10412 14188 10464
rect 14240 10452 14246 10464
rect 14476 10452 14504 10483
rect 14240 10424 14504 10452
rect 14240 10412 14246 10424
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 1578 10248 1584 10260
rect 1539 10220 1584 10248
rect 1578 10208 1584 10220
rect 1636 10208 1642 10260
rect 2130 10208 2136 10260
rect 2188 10248 2194 10260
rect 2869 10251 2927 10257
rect 2869 10248 2881 10251
rect 2188 10220 2881 10248
rect 2188 10208 2194 10220
rect 2869 10217 2881 10220
rect 2915 10248 2927 10251
rect 3326 10248 3332 10260
rect 2915 10220 3332 10248
rect 2915 10217 2927 10220
rect 2869 10211 2927 10217
rect 3326 10208 3332 10220
rect 3384 10208 3390 10260
rect 5166 10248 5172 10260
rect 5127 10220 5172 10248
rect 5166 10208 5172 10220
rect 5224 10208 5230 10260
rect 6822 10248 6828 10260
rect 6783 10220 6828 10248
rect 6822 10208 6828 10220
rect 6880 10208 6886 10260
rect 7466 10248 7472 10260
rect 7208 10220 7472 10248
rect 2038 10140 2044 10192
rect 2096 10180 2102 10192
rect 3694 10180 3700 10192
rect 2096 10152 3700 10180
rect 2096 10140 2102 10152
rect 3694 10140 3700 10152
rect 3752 10180 3758 10192
rect 3752 10152 4200 10180
rect 3752 10140 3758 10152
rect 1397 10115 1455 10121
rect 1397 10081 1409 10115
rect 1443 10112 1455 10115
rect 1486 10112 1492 10124
rect 1443 10084 1492 10112
rect 1443 10081 1455 10084
rect 1397 10075 1455 10081
rect 1486 10072 1492 10084
rect 1544 10072 1550 10124
rect 2133 10115 2191 10121
rect 2133 10081 2145 10115
rect 2179 10112 2191 10115
rect 2406 10112 2412 10124
rect 2179 10084 2412 10112
rect 2179 10081 2191 10084
rect 2133 10075 2191 10081
rect 2406 10072 2412 10084
rect 2464 10072 2470 10124
rect 2590 10112 2596 10124
rect 2551 10084 2596 10112
rect 2590 10072 2596 10084
rect 2648 10072 2654 10124
rect 2774 10112 2780 10124
rect 2735 10084 2780 10112
rect 2774 10072 2780 10084
rect 2832 10072 2838 10124
rect 4172 10121 4200 10152
rect 4540 10152 5911 10180
rect 4540 10124 4568 10152
rect 4157 10115 4215 10121
rect 4157 10081 4169 10115
rect 4203 10081 4215 10115
rect 4522 10112 4528 10124
rect 4435 10084 4528 10112
rect 4157 10075 4215 10081
rect 4522 10072 4528 10084
rect 4580 10072 4586 10124
rect 4709 10115 4767 10121
rect 4709 10081 4721 10115
rect 4755 10081 4767 10115
rect 4709 10075 4767 10081
rect 2792 10044 2820 10072
rect 4614 10044 4620 10056
rect 2792 10016 4620 10044
rect 4614 10004 4620 10016
rect 4672 10044 4678 10056
rect 4724 10044 4752 10075
rect 5350 10072 5356 10124
rect 5408 10112 5414 10124
rect 5883 10121 5911 10152
rect 5721 10115 5779 10121
rect 5721 10112 5733 10115
rect 5408 10084 5733 10112
rect 5408 10072 5414 10084
rect 5721 10081 5733 10084
rect 5767 10081 5779 10115
rect 5721 10075 5779 10081
rect 5868 10115 5926 10121
rect 5868 10081 5880 10115
rect 5914 10112 5926 10115
rect 5994 10112 6000 10124
rect 5914 10084 6000 10112
rect 5914 10081 5926 10084
rect 5868 10075 5926 10081
rect 5994 10072 6000 10084
rect 6052 10072 6058 10124
rect 4672 10016 4752 10044
rect 4672 10004 4678 10016
rect 5534 10004 5540 10056
rect 5592 10044 5598 10056
rect 6089 10047 6147 10053
rect 6089 10044 6101 10047
rect 5592 10016 6101 10044
rect 5592 10004 5598 10016
rect 6089 10013 6101 10016
rect 6135 10013 6147 10047
rect 6089 10007 6147 10013
rect 1578 9936 1584 9988
rect 1636 9976 1642 9988
rect 2409 9979 2467 9985
rect 2409 9976 2421 9979
rect 1636 9948 2421 9976
rect 1636 9936 1642 9948
rect 2409 9945 2421 9948
rect 2455 9945 2467 9979
rect 2409 9939 2467 9945
rect 5442 9936 5448 9988
rect 5500 9976 5506 9988
rect 5997 9979 6055 9985
rect 5997 9976 6009 9979
rect 5500 9948 6009 9976
rect 5500 9936 5506 9948
rect 5997 9945 6009 9948
rect 6043 9945 6055 9979
rect 5997 9939 6055 9945
rect 6730 9936 6736 9988
rect 6788 9976 6794 9988
rect 7208 9985 7236 10220
rect 7466 10208 7472 10220
rect 7524 10248 7530 10260
rect 8754 10248 8760 10260
rect 7524 10220 8760 10248
rect 7524 10208 7530 10220
rect 8754 10208 8760 10220
rect 8812 10208 8818 10260
rect 12345 10251 12403 10257
rect 12345 10217 12357 10251
rect 12391 10248 12403 10251
rect 12802 10248 12808 10260
rect 12391 10220 12808 10248
rect 12391 10217 12403 10220
rect 12345 10211 12403 10217
rect 12802 10208 12808 10220
rect 12860 10208 12866 10260
rect 14366 10248 14372 10260
rect 14327 10220 14372 10248
rect 14366 10208 14372 10220
rect 14424 10208 14430 10260
rect 7282 10140 7288 10192
rect 7340 10180 7346 10192
rect 7377 10183 7435 10189
rect 7377 10180 7389 10183
rect 7340 10152 7389 10180
rect 7340 10140 7346 10152
rect 7377 10149 7389 10152
rect 7423 10149 7435 10183
rect 7377 10143 7435 10149
rect 8481 10183 8539 10189
rect 8481 10149 8493 10183
rect 8527 10180 8539 10183
rect 8662 10180 8668 10192
rect 8527 10152 8668 10180
rect 8527 10149 8539 10152
rect 8481 10143 8539 10149
rect 8662 10140 8668 10152
rect 8720 10180 8726 10192
rect 9401 10183 9459 10189
rect 9401 10180 9413 10183
rect 8720 10152 9413 10180
rect 8720 10140 8726 10152
rect 9401 10149 9413 10152
rect 9447 10149 9459 10183
rect 9401 10143 9459 10149
rect 9861 10183 9919 10189
rect 9861 10149 9873 10183
rect 9907 10180 9919 10183
rect 9950 10180 9956 10192
rect 9907 10152 9956 10180
rect 9907 10149 9919 10152
rect 9861 10143 9919 10149
rect 9950 10140 9956 10152
rect 10008 10140 10014 10192
rect 13167 10183 13225 10189
rect 13167 10149 13179 10183
rect 13213 10180 13225 10183
rect 13446 10180 13452 10192
rect 13213 10152 13452 10180
rect 13213 10149 13225 10152
rect 13167 10143 13225 10149
rect 13446 10140 13452 10152
rect 13504 10140 13510 10192
rect 14826 10140 14832 10192
rect 14884 10180 14890 10192
rect 15473 10183 15531 10189
rect 15473 10180 15485 10183
rect 14884 10152 15485 10180
rect 14884 10140 14890 10152
rect 15473 10149 15485 10152
rect 15519 10149 15531 10183
rect 15473 10143 15531 10149
rect 24210 10140 24216 10192
rect 24268 10180 24274 10192
rect 24305 10183 24363 10189
rect 24305 10180 24317 10183
rect 24268 10152 24317 10180
rect 24268 10140 24274 10152
rect 24305 10149 24317 10152
rect 24351 10149 24363 10183
rect 24305 10143 24363 10149
rect 10778 10072 10784 10124
rect 10836 10112 10842 10124
rect 11241 10115 11299 10121
rect 11241 10112 11253 10115
rect 10836 10084 11253 10112
rect 10836 10072 10842 10084
rect 11241 10081 11253 10084
rect 11287 10112 11299 10115
rect 11606 10112 11612 10124
rect 11287 10084 11612 10112
rect 11287 10081 11299 10084
rect 11241 10075 11299 10081
rect 11606 10072 11612 10084
rect 11664 10072 11670 10124
rect 11701 10115 11759 10121
rect 11701 10081 11713 10115
rect 11747 10081 11759 10115
rect 11701 10075 11759 10081
rect 7745 10047 7803 10053
rect 7745 10013 7757 10047
rect 7791 10044 7803 10047
rect 7926 10044 7932 10056
rect 7791 10016 7932 10044
rect 7791 10013 7803 10016
rect 7745 10007 7803 10013
rect 7926 10004 7932 10016
rect 7984 10004 7990 10056
rect 9398 10004 9404 10056
rect 9456 10044 9462 10056
rect 9769 10047 9827 10053
rect 9769 10044 9781 10047
rect 9456 10016 9781 10044
rect 9456 10004 9462 10016
rect 9769 10013 9781 10016
rect 9815 10013 9827 10047
rect 10042 10044 10048 10056
rect 10003 10016 10048 10044
rect 9769 10007 9827 10013
rect 10042 10004 10048 10016
rect 10100 10004 10106 10056
rect 11330 10044 11336 10056
rect 10796 10016 11336 10044
rect 7193 9979 7251 9985
rect 7193 9976 7205 9979
rect 6788 9948 7205 9976
rect 6788 9936 6794 9948
rect 7193 9945 7205 9948
rect 7239 9945 7251 9979
rect 7650 9976 7656 9988
rect 7611 9948 7656 9976
rect 7193 9939 7251 9945
rect 7650 9936 7656 9948
rect 7708 9936 7714 9988
rect 10796 9920 10824 10016
rect 11330 10004 11336 10016
rect 11388 10044 11394 10056
rect 11716 10044 11744 10075
rect 12618 10072 12624 10124
rect 12676 10112 12682 10124
rect 12805 10115 12863 10121
rect 12805 10112 12817 10115
rect 12676 10084 12817 10112
rect 12676 10072 12682 10084
rect 12805 10081 12817 10084
rect 12851 10081 12863 10115
rect 12805 10075 12863 10081
rect 11388 10016 11744 10044
rect 11977 10047 12035 10053
rect 11388 10004 11394 10016
rect 11977 10013 11989 10047
rect 12023 10044 12035 10047
rect 12986 10044 12992 10056
rect 12023 10016 12992 10044
rect 12023 10013 12035 10016
rect 11977 10007 12035 10013
rect 12986 10004 12992 10016
rect 13044 10004 13050 10056
rect 15381 10047 15439 10053
rect 15381 10013 15393 10047
rect 15427 10044 15439 10047
rect 15562 10044 15568 10056
rect 15427 10016 15568 10044
rect 15427 10013 15439 10016
rect 15381 10007 15439 10013
rect 15562 10004 15568 10016
rect 15620 10004 15626 10056
rect 15657 10047 15715 10053
rect 15657 10013 15669 10047
rect 15703 10013 15715 10047
rect 15657 10007 15715 10013
rect 24213 10047 24271 10053
rect 24213 10013 24225 10047
rect 24259 10044 24271 10047
rect 24302 10044 24308 10056
rect 24259 10016 24308 10044
rect 24259 10013 24271 10016
rect 24213 10007 24271 10013
rect 13722 9976 13728 9988
rect 13683 9948 13728 9976
rect 13722 9936 13728 9948
rect 13780 9936 13786 9988
rect 15286 9936 15292 9988
rect 15344 9976 15350 9988
rect 15672 9976 15700 10007
rect 24302 10004 24308 10016
rect 24360 10044 24366 10056
rect 25038 10044 25044 10056
rect 24360 10016 25044 10044
rect 24360 10004 24366 10016
rect 25038 10004 25044 10016
rect 25096 10004 25102 10056
rect 24762 9976 24768 9988
rect 15344 9948 15700 9976
rect 24723 9948 24768 9976
rect 15344 9936 15350 9948
rect 24762 9936 24768 9948
rect 24820 9936 24826 9988
rect 3697 9911 3755 9917
rect 3697 9877 3709 9911
rect 3743 9908 3755 9911
rect 3786 9908 3792 9920
rect 3743 9880 3792 9908
rect 3743 9877 3755 9880
rect 3697 9871 3755 9877
rect 3786 9868 3792 9880
rect 3844 9868 3850 9920
rect 5350 9868 5356 9920
rect 5408 9908 5414 9920
rect 5537 9911 5595 9917
rect 5537 9908 5549 9911
rect 5408 9880 5549 9908
rect 5408 9868 5414 9880
rect 5537 9877 5549 9880
rect 5583 9877 5595 9911
rect 6362 9908 6368 9920
rect 6323 9880 6368 9908
rect 5537 9871 5595 9877
rect 6362 9868 6368 9880
rect 6420 9868 6426 9920
rect 6638 9868 6644 9920
rect 6696 9908 6702 9920
rect 7466 9908 7472 9920
rect 6696 9880 7472 9908
rect 6696 9868 6702 9880
rect 7466 9868 7472 9880
rect 7524 9917 7530 9920
rect 7524 9911 7573 9917
rect 7524 9877 7527 9911
rect 7561 9877 7573 9911
rect 7524 9871 7573 9877
rect 8021 9911 8079 9917
rect 8021 9877 8033 9911
rect 8067 9908 8079 9911
rect 8294 9908 8300 9920
rect 8067 9880 8300 9908
rect 8067 9877 8079 9880
rect 8021 9871 8079 9877
rect 7524 9868 7530 9871
rect 8294 9868 8300 9880
rect 8352 9868 8358 9920
rect 10778 9908 10784 9920
rect 10739 9880 10784 9908
rect 10778 9868 10784 9880
rect 10836 9868 10842 9920
rect 12710 9908 12716 9920
rect 12671 9880 12716 9908
rect 12710 9868 12716 9880
rect 12768 9868 12774 9920
rect 13538 9868 13544 9920
rect 13596 9908 13602 9920
rect 14366 9908 14372 9920
rect 13596 9880 14372 9908
rect 13596 9868 13602 9880
rect 14366 9868 14372 9880
rect 14424 9868 14430 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 3694 9664 3700 9716
rect 3752 9704 3758 9716
rect 3881 9707 3939 9713
rect 3881 9704 3893 9707
rect 3752 9676 3893 9704
rect 3752 9664 3758 9676
rect 3881 9673 3893 9676
rect 3927 9673 3939 9707
rect 4614 9704 4620 9716
rect 4575 9676 4620 9704
rect 3881 9667 3939 9673
rect 4614 9664 4620 9676
rect 4672 9664 4678 9716
rect 7469 9707 7527 9713
rect 7469 9673 7481 9707
rect 7515 9704 7527 9707
rect 7558 9704 7564 9716
rect 7515 9676 7564 9704
rect 7515 9673 7527 9676
rect 7469 9667 7527 9673
rect 7558 9664 7564 9676
rect 7616 9664 7622 9716
rect 7837 9707 7895 9713
rect 7837 9673 7849 9707
rect 7883 9704 7895 9707
rect 10778 9704 10784 9716
rect 7883 9676 10784 9704
rect 7883 9673 7895 9676
rect 7837 9667 7895 9673
rect 10778 9664 10784 9676
rect 10836 9664 10842 9716
rect 11606 9664 11612 9716
rect 11664 9704 11670 9716
rect 11701 9707 11759 9713
rect 11701 9704 11713 9707
rect 11664 9676 11713 9704
rect 11664 9664 11670 9676
rect 11701 9673 11713 9676
rect 11747 9673 11759 9707
rect 11701 9667 11759 9673
rect 13722 9664 13728 9716
rect 13780 9704 13786 9716
rect 14826 9704 14832 9716
rect 13780 9676 14832 9704
rect 13780 9664 13786 9676
rect 14826 9664 14832 9676
rect 14884 9704 14890 9716
rect 15013 9707 15071 9713
rect 15013 9704 15025 9707
rect 14884 9676 15025 9704
rect 14884 9664 14890 9676
rect 15013 9673 15025 9676
rect 15059 9673 15071 9707
rect 15013 9667 15071 9673
rect 15562 9664 15568 9716
rect 15620 9704 15626 9716
rect 16209 9707 16267 9713
rect 16209 9704 16221 9707
rect 15620 9676 16221 9704
rect 15620 9664 15626 9676
rect 16209 9673 16221 9676
rect 16255 9673 16267 9707
rect 25038 9704 25044 9716
rect 24999 9676 25044 9704
rect 16209 9667 16267 9673
rect 25038 9664 25044 9676
rect 25096 9664 25102 9716
rect 3970 9596 3976 9648
rect 4028 9636 4034 9648
rect 6638 9636 6644 9648
rect 4028 9608 5120 9636
rect 6551 9608 6644 9636
rect 4028 9596 4034 9608
rect 1765 9571 1823 9577
rect 1765 9537 1777 9571
rect 1811 9568 1823 9571
rect 4430 9568 4436 9580
rect 1811 9540 4436 9568
rect 1811 9537 1823 9540
rect 1765 9531 1823 9537
rect 4430 9528 4436 9540
rect 4488 9528 4494 9580
rect 1578 9500 1584 9512
rect 1539 9472 1584 9500
rect 1578 9460 1584 9472
rect 1636 9460 1642 9512
rect 2133 9503 2191 9509
rect 2133 9469 2145 9503
rect 2179 9500 2191 9503
rect 3513 9503 3571 9509
rect 2179 9472 2452 9500
rect 2179 9469 2191 9472
rect 2133 9463 2191 9469
rect 2424 9376 2452 9472
rect 3513 9469 3525 9503
rect 3559 9500 3571 9503
rect 3694 9500 3700 9512
rect 3559 9472 3700 9500
rect 3559 9469 3571 9472
rect 3513 9463 3571 9469
rect 3694 9460 3700 9472
rect 3752 9460 3758 9512
rect 5092 9509 5120 9608
rect 6638 9596 6644 9608
rect 6696 9636 6702 9648
rect 7358 9639 7416 9645
rect 7358 9636 7370 9639
rect 6696 9608 7370 9636
rect 6696 9596 6702 9608
rect 7358 9605 7370 9608
rect 7404 9636 7416 9639
rect 7742 9636 7748 9648
rect 7404 9608 7748 9636
rect 7404 9605 7416 9608
rect 7358 9599 7416 9605
rect 7742 9596 7748 9608
rect 7800 9596 7806 9648
rect 12618 9596 12624 9648
rect 12676 9636 12682 9648
rect 14001 9639 14059 9645
rect 14001 9636 14013 9639
rect 12676 9608 14013 9636
rect 12676 9596 12682 9608
rect 14001 9605 14013 9608
rect 14047 9605 14059 9639
rect 14001 9599 14059 9605
rect 7006 9528 7012 9580
rect 7064 9568 7070 9580
rect 7561 9571 7619 9577
rect 7561 9568 7573 9571
rect 7064 9540 7573 9568
rect 7064 9528 7070 9540
rect 7561 9537 7573 9540
rect 7607 9537 7619 9571
rect 7561 9531 7619 9537
rect 12710 9528 12716 9580
rect 12768 9568 12774 9580
rect 14185 9571 14243 9577
rect 14185 9568 14197 9571
rect 12768 9540 14197 9568
rect 12768 9528 12774 9540
rect 14185 9537 14197 9540
rect 14231 9537 14243 9571
rect 14185 9531 14243 9537
rect 15286 9528 15292 9580
rect 15344 9568 15350 9580
rect 16577 9571 16635 9577
rect 16577 9568 16589 9571
rect 15344 9540 16589 9568
rect 15344 9528 15350 9540
rect 16577 9537 16589 9540
rect 16623 9537 16635 9571
rect 16577 9531 16635 9537
rect 24210 9528 24216 9580
rect 24268 9568 24274 9580
rect 24397 9571 24455 9577
rect 24397 9568 24409 9571
rect 24268 9540 24409 9568
rect 24268 9528 24274 9540
rect 24397 9537 24409 9540
rect 24443 9568 24455 9571
rect 24673 9571 24731 9577
rect 24673 9568 24685 9571
rect 24443 9540 24685 9568
rect 24443 9537 24455 9540
rect 24397 9531 24455 9537
rect 24673 9537 24685 9540
rect 24719 9537 24731 9571
rect 24673 9531 24731 9537
rect 5077 9503 5135 9509
rect 5077 9469 5089 9503
rect 5123 9500 5135 9503
rect 5813 9503 5871 9509
rect 5813 9500 5825 9503
rect 5123 9472 5825 9500
rect 5123 9469 5135 9472
rect 5077 9463 5135 9469
rect 5813 9469 5825 9472
rect 5859 9500 5871 9503
rect 7650 9500 7656 9512
rect 5859 9472 7656 9500
rect 5859 9469 5871 9472
rect 5813 9463 5871 9469
rect 7650 9460 7656 9472
rect 7708 9460 7714 9512
rect 8754 9500 8760 9512
rect 8715 9472 8760 9500
rect 8754 9460 8760 9472
rect 8812 9460 8818 9512
rect 10505 9503 10563 9509
rect 10505 9469 10517 9503
rect 10551 9500 10563 9503
rect 10686 9500 10692 9512
rect 10551 9472 10692 9500
rect 10551 9469 10563 9472
rect 10505 9463 10563 9469
rect 10686 9460 10692 9472
rect 10744 9460 10750 9512
rect 12434 9500 12440 9512
rect 12395 9472 12440 9500
rect 12434 9460 12440 9472
rect 12492 9460 12498 9512
rect 23753 9503 23811 9509
rect 23753 9469 23765 9503
rect 23799 9469 23811 9503
rect 23753 9463 23811 9469
rect 4338 9432 4344 9444
rect 4299 9404 4344 9432
rect 4338 9392 4344 9404
rect 4396 9392 4402 9444
rect 5350 9432 5356 9444
rect 4908 9404 5356 9432
rect 2406 9364 2412 9376
rect 2367 9336 2412 9364
rect 2406 9324 2412 9336
rect 2464 9324 2470 9376
rect 2774 9364 2780 9376
rect 2735 9336 2780 9364
rect 2774 9324 2780 9336
rect 2832 9324 2838 9376
rect 3970 9324 3976 9376
rect 4028 9364 4034 9376
rect 4908 9364 4936 9404
rect 5350 9392 5356 9404
rect 5408 9432 5414 9444
rect 6181 9435 6239 9441
rect 6181 9432 6193 9435
rect 5408 9404 6193 9432
rect 5408 9392 5414 9404
rect 6181 9401 6193 9404
rect 6227 9401 6239 9435
rect 7190 9432 7196 9444
rect 7151 9404 7196 9432
rect 6181 9395 6239 9401
rect 7190 9392 7196 9404
rect 7248 9392 7254 9444
rect 9078 9435 9136 9441
rect 9078 9401 9090 9435
rect 9124 9432 9136 9435
rect 10321 9435 10379 9441
rect 10321 9432 10333 9435
rect 9124 9404 10333 9432
rect 9124 9401 9136 9404
rect 9078 9395 9136 9401
rect 10321 9401 10333 9404
rect 10367 9432 10379 9435
rect 10826 9435 10884 9441
rect 10826 9432 10838 9435
rect 10367 9404 10838 9432
rect 10367 9401 10379 9404
rect 10321 9395 10379 9401
rect 10826 9401 10838 9404
rect 10872 9432 10884 9435
rect 11974 9432 11980 9444
rect 10872 9404 11980 9432
rect 10872 9401 10884 9404
rect 10826 9395 10884 9401
rect 5442 9364 5448 9376
rect 4028 9336 4936 9364
rect 5403 9336 5448 9364
rect 4028 9324 4034 9336
rect 5442 9324 5448 9336
rect 5500 9324 5506 9376
rect 7006 9364 7012 9376
rect 6967 9336 7012 9364
rect 7006 9324 7012 9336
rect 7064 9324 7070 9376
rect 7650 9324 7656 9376
rect 7708 9364 7714 9376
rect 8205 9367 8263 9373
rect 8205 9364 8217 9367
rect 7708 9336 8217 9364
rect 7708 9324 7714 9336
rect 8205 9333 8217 9336
rect 8251 9333 8263 9367
rect 8205 9327 8263 9333
rect 8386 9324 8392 9376
rect 8444 9364 8450 9376
rect 8573 9367 8631 9373
rect 8573 9364 8585 9367
rect 8444 9336 8585 9364
rect 8444 9324 8450 9336
rect 8573 9333 8585 9336
rect 8619 9364 8631 9367
rect 9093 9364 9121 9395
rect 11974 9392 11980 9404
rect 12032 9432 12038 9444
rect 12161 9435 12219 9441
rect 12161 9432 12173 9435
rect 12032 9404 12173 9432
rect 12032 9392 12038 9404
rect 12161 9401 12173 9404
rect 12207 9432 12219 9435
rect 12758 9435 12816 9441
rect 12758 9432 12770 9435
rect 12207 9404 12770 9432
rect 12207 9401 12219 9404
rect 12161 9395 12219 9401
rect 12758 9401 12770 9404
rect 12804 9432 12816 9435
rect 13446 9432 13452 9444
rect 12804 9404 13452 9432
rect 12804 9401 12816 9404
rect 12758 9395 12816 9401
rect 13446 9392 13452 9404
rect 13504 9432 13510 9444
rect 13633 9435 13691 9441
rect 13633 9432 13645 9435
rect 13504 9404 13645 9432
rect 13504 9392 13510 9404
rect 13633 9401 13645 9404
rect 13679 9401 13691 9435
rect 13633 9395 13691 9401
rect 13906 9392 13912 9444
rect 13964 9432 13970 9444
rect 14737 9435 14795 9441
rect 14737 9432 14749 9435
rect 13964 9404 14749 9432
rect 13964 9392 13970 9404
rect 14737 9401 14749 9404
rect 14783 9432 14795 9435
rect 15286 9432 15292 9444
rect 14783 9404 15148 9432
rect 15247 9404 15292 9432
rect 14783 9401 14795 9404
rect 14737 9395 14795 9401
rect 8619 9336 9121 9364
rect 9677 9367 9735 9373
rect 8619 9333 8631 9336
rect 8573 9327 8631 9333
rect 9677 9333 9689 9367
rect 9723 9364 9735 9367
rect 9766 9364 9772 9376
rect 9723 9336 9772 9364
rect 9723 9333 9735 9336
rect 9677 9327 9735 9333
rect 9766 9324 9772 9336
rect 9824 9324 9830 9376
rect 9950 9364 9956 9376
rect 9911 9336 9956 9364
rect 9950 9324 9956 9336
rect 10008 9324 10014 9376
rect 11422 9364 11428 9376
rect 11383 9336 11428 9364
rect 11422 9324 11428 9336
rect 11480 9324 11486 9376
rect 13354 9364 13360 9376
rect 13315 9336 13360 9364
rect 13354 9324 13360 9336
rect 13412 9324 13418 9376
rect 15120 9364 15148 9404
rect 15286 9392 15292 9404
rect 15344 9392 15350 9444
rect 15381 9435 15439 9441
rect 15381 9401 15393 9435
rect 15427 9401 15439 9435
rect 15930 9432 15936 9444
rect 15891 9404 15936 9432
rect 15381 9395 15439 9401
rect 15396 9364 15424 9395
rect 15930 9392 15936 9404
rect 15988 9392 15994 9444
rect 16298 9364 16304 9376
rect 15120 9336 16304 9364
rect 16298 9324 16304 9336
rect 16356 9324 16362 9376
rect 16758 9364 16764 9376
rect 16719 9336 16764 9364
rect 16758 9324 16764 9336
rect 16816 9324 16822 9376
rect 23477 9367 23535 9373
rect 23477 9333 23489 9367
rect 23523 9364 23535 9367
rect 23768 9364 23796 9463
rect 24026 9364 24032 9376
rect 23523 9336 24032 9364
rect 23523 9333 23535 9336
rect 23477 9327 23535 9333
rect 24026 9324 24032 9336
rect 24084 9324 24090 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 3142 9160 3148 9172
rect 3103 9132 3148 9160
rect 3142 9120 3148 9132
rect 3200 9120 3206 9172
rect 3418 9160 3424 9172
rect 3379 9132 3424 9160
rect 3418 9120 3424 9132
rect 3476 9120 3482 9172
rect 4338 9160 4344 9172
rect 4299 9132 4344 9160
rect 4338 9120 4344 9132
rect 4396 9120 4402 9172
rect 6270 9160 6276 9172
rect 6231 9132 6276 9160
rect 6270 9120 6276 9132
rect 6328 9120 6334 9172
rect 7282 9120 7288 9172
rect 7340 9160 7346 9172
rect 7469 9163 7527 9169
rect 7469 9160 7481 9163
rect 7340 9132 7481 9160
rect 7340 9120 7346 9132
rect 7469 9129 7481 9132
rect 7515 9129 7527 9163
rect 12253 9163 12311 9169
rect 12253 9160 12265 9163
rect 7469 9123 7527 9129
rect 9048 9132 12265 9160
rect 4706 9052 4712 9104
rect 4764 9092 4770 9104
rect 5074 9092 5080 9104
rect 4764 9064 5080 9092
rect 4764 9052 4770 9064
rect 5074 9052 5080 9064
rect 5132 9092 5138 9104
rect 6457 9095 6515 9101
rect 5132 9064 6177 9092
rect 5132 9052 5138 9064
rect 1578 9024 1584 9036
rect 1539 8996 1584 9024
rect 1578 8984 1584 8996
rect 1636 8984 1642 9036
rect 2958 9024 2964 9036
rect 2919 8996 2964 9024
rect 2958 8984 2964 8996
rect 3016 8984 3022 9036
rect 4982 9024 4988 9036
rect 4943 8996 4988 9024
rect 4982 8984 4988 8996
rect 5040 8984 5046 9036
rect 6149 9024 6177 9064
rect 6457 9061 6469 9095
rect 6503 9092 6515 9095
rect 6822 9092 6828 9104
rect 6503 9064 6828 9092
rect 6503 9061 6515 9064
rect 6457 9055 6515 9061
rect 6822 9052 6828 9064
rect 6880 9052 6886 9104
rect 7190 9052 7196 9104
rect 7248 9092 7254 9104
rect 7837 9095 7895 9101
rect 7837 9092 7849 9095
rect 7248 9064 7849 9092
rect 7248 9052 7254 9064
rect 7837 9061 7849 9064
rect 7883 9092 7895 9095
rect 8570 9092 8576 9104
rect 7883 9064 8576 9092
rect 7883 9061 7895 9064
rect 7837 9055 7895 9061
rect 8570 9052 8576 9064
rect 8628 9052 8634 9104
rect 8021 9027 8079 9033
rect 8021 9024 8033 9027
rect 6149 8996 8033 9024
rect 8021 8993 8033 8996
rect 8067 9024 8079 9027
rect 8110 9024 8116 9036
rect 8067 8996 8116 9024
rect 8067 8993 8079 8996
rect 8021 8987 8079 8993
rect 8110 8984 8116 8996
rect 8168 8984 8174 9036
rect 8294 8984 8300 9036
rect 8352 9024 8358 9036
rect 8481 9027 8539 9033
rect 8481 9024 8493 9027
rect 8352 8996 8493 9024
rect 8352 8984 8358 8996
rect 8481 8993 8493 8996
rect 8527 8993 8539 9027
rect 8754 9024 8760 9036
rect 8715 8996 8760 9024
rect 8481 8987 8539 8993
rect 8754 8984 8760 8996
rect 8812 9024 8818 9036
rect 9048 9024 9076 9132
rect 12253 9129 12265 9132
rect 12299 9129 12311 9163
rect 13906 9160 13912 9172
rect 13867 9132 13912 9160
rect 12253 9123 12311 9129
rect 13906 9120 13912 9132
rect 13964 9120 13970 9172
rect 16224 9132 17172 9160
rect 9766 9052 9772 9104
rect 9824 9092 9830 9104
rect 9861 9095 9919 9101
rect 9861 9092 9873 9095
rect 9824 9064 9873 9092
rect 9824 9052 9830 9064
rect 9861 9061 9873 9064
rect 9907 9061 9919 9095
rect 9861 9055 9919 9061
rect 10778 9052 10784 9104
rect 10836 9092 10842 9104
rect 11057 9095 11115 9101
rect 11057 9092 11069 9095
rect 10836 9064 11069 9092
rect 10836 9052 10842 9064
rect 11057 9061 11069 9064
rect 11103 9061 11115 9095
rect 11606 9092 11612 9104
rect 11057 9055 11115 9061
rect 11532 9064 11612 9092
rect 11532 9033 11560 9064
rect 11606 9052 11612 9064
rect 11664 9052 11670 9104
rect 11977 9095 12035 9101
rect 11977 9061 11989 9095
rect 12023 9092 12035 9095
rect 12434 9092 12440 9104
rect 12023 9064 12440 9092
rect 12023 9061 12035 9064
rect 11977 9055 12035 9061
rect 12434 9052 12440 9064
rect 12492 9092 12498 9104
rect 12621 9095 12679 9101
rect 12621 9092 12633 9095
rect 12492 9064 12633 9092
rect 12492 9052 12498 9064
rect 12621 9061 12633 9064
rect 12667 9061 12679 9095
rect 12621 9055 12679 9061
rect 13351 9095 13409 9101
rect 13351 9061 13363 9095
rect 13397 9092 13409 9095
rect 13446 9092 13452 9104
rect 13397 9064 13452 9092
rect 13397 9061 13409 9064
rect 13351 9055 13409 9061
rect 13446 9052 13452 9064
rect 13504 9052 13510 9104
rect 15654 9092 15660 9104
rect 15615 9064 15660 9092
rect 15654 9052 15660 9064
rect 15712 9052 15718 9104
rect 15930 9052 15936 9104
rect 15988 9092 15994 9104
rect 16224 9101 16252 9132
rect 16209 9095 16267 9101
rect 16209 9092 16221 9095
rect 15988 9064 16221 9092
rect 15988 9052 15994 9064
rect 16209 9061 16221 9064
rect 16255 9061 16267 9095
rect 16209 9055 16267 9061
rect 17144 9036 17172 9132
rect 24118 9052 24124 9104
rect 24176 9092 24182 9104
rect 24213 9095 24271 9101
rect 24213 9092 24225 9095
rect 24176 9064 24225 9092
rect 24176 9052 24182 9064
rect 24213 9061 24225 9064
rect 24259 9061 24271 9095
rect 24213 9055 24271 9061
rect 8812 8996 9076 9024
rect 11517 9027 11575 9033
rect 8812 8984 8818 8996
rect 11517 8993 11529 9027
rect 11563 8993 11575 9027
rect 11517 8987 11575 8993
rect 11793 9027 11851 9033
rect 11793 8993 11805 9027
rect 11839 9024 11851 9027
rect 11882 9024 11888 9036
rect 11839 8996 11888 9024
rect 11839 8993 11851 8996
rect 11793 8987 11851 8993
rect 11882 8984 11888 8996
rect 11940 8984 11946 9036
rect 12986 9024 12992 9036
rect 12947 8996 12992 9024
rect 12986 8984 12992 8996
rect 13044 8984 13050 9036
rect 17126 9033 17132 9036
rect 17104 9027 17132 9033
rect 17104 8993 17116 9027
rect 17184 9024 17190 9036
rect 17184 8996 17277 9024
rect 17104 8987 17132 8993
rect 17126 8984 17132 8987
rect 17184 8984 17190 8996
rect 24762 8984 24768 9036
rect 24820 9024 24826 9036
rect 24820 8996 24865 9024
rect 24820 8984 24826 8996
rect 1486 8916 1492 8968
rect 1544 8956 1550 8968
rect 3789 8959 3847 8965
rect 3789 8956 3801 8959
rect 1544 8928 3801 8956
rect 1544 8916 1550 8928
rect 3789 8925 3801 8928
rect 3835 8925 3847 8959
rect 3789 8919 3847 8925
rect 4062 8916 4068 8968
rect 4120 8956 4126 8968
rect 4893 8959 4951 8965
rect 4893 8956 4905 8959
rect 4120 8928 4905 8956
rect 4120 8916 4126 8928
rect 4893 8925 4905 8928
rect 4939 8925 4951 8959
rect 4893 8919 4951 8925
rect 5074 8916 5080 8968
rect 5132 8956 5138 8968
rect 5132 8928 6177 8956
rect 5132 8916 5138 8928
rect 2590 8848 2596 8900
rect 2648 8888 2654 8900
rect 2685 8891 2743 8897
rect 2685 8888 2697 8891
rect 2648 8860 2697 8888
rect 2648 8848 2654 8860
rect 2685 8857 2697 8860
rect 2731 8888 2743 8891
rect 3694 8888 3700 8900
rect 2731 8860 3700 8888
rect 2731 8857 2743 8860
rect 2685 8851 2743 8857
rect 3694 8848 3700 8860
rect 3752 8848 3758 8900
rect 5442 8848 5448 8900
rect 5500 8888 5506 8900
rect 5905 8891 5963 8897
rect 5905 8888 5917 8891
rect 5500 8860 5917 8888
rect 5500 8848 5506 8860
rect 5905 8857 5917 8860
rect 5951 8857 5963 8891
rect 6149 8888 6177 8928
rect 6270 8916 6276 8968
rect 6328 8956 6334 8968
rect 6825 8959 6883 8965
rect 6825 8956 6837 8959
rect 6328 8928 6837 8956
rect 6328 8916 6334 8928
rect 6825 8925 6837 8928
rect 6871 8956 6883 8959
rect 7098 8956 7104 8968
rect 6871 8928 7104 8956
rect 6871 8925 6883 8928
rect 6825 8919 6883 8925
rect 7098 8916 7104 8928
rect 7156 8956 7162 8968
rect 7745 8959 7803 8965
rect 7745 8956 7757 8959
rect 7156 8928 7757 8956
rect 7156 8916 7162 8928
rect 7745 8925 7757 8928
rect 7791 8925 7803 8959
rect 9769 8959 9827 8965
rect 7745 8919 7803 8925
rect 8128 8928 9536 8956
rect 8128 8888 8156 8928
rect 6149 8860 8156 8888
rect 5905 8851 5963 8857
rect 8202 8848 8208 8900
rect 8260 8888 8266 8900
rect 9398 8888 9404 8900
rect 8260 8860 9404 8888
rect 8260 8848 8266 8860
rect 9398 8848 9404 8860
rect 9456 8848 9462 8900
rect 9508 8888 9536 8928
rect 9769 8925 9781 8959
rect 9815 8956 9827 8959
rect 11606 8956 11612 8968
rect 9815 8928 11612 8956
rect 9815 8925 9827 8928
rect 9769 8919 9827 8925
rect 11606 8916 11612 8928
rect 11664 8916 11670 8968
rect 15565 8959 15623 8965
rect 15565 8925 15577 8959
rect 15611 8956 15623 8959
rect 16758 8956 16764 8968
rect 15611 8928 16764 8956
rect 15611 8925 15623 8928
rect 15565 8919 15623 8925
rect 16758 8916 16764 8928
rect 16816 8916 16822 8968
rect 24121 8959 24179 8965
rect 24121 8925 24133 8959
rect 24167 8956 24179 8959
rect 24854 8956 24860 8968
rect 24167 8928 24860 8956
rect 24167 8925 24179 8928
rect 24121 8919 24179 8925
rect 24854 8916 24860 8928
rect 24912 8916 24918 8968
rect 10042 8888 10048 8900
rect 9508 8860 10048 8888
rect 10042 8848 10048 8860
rect 10100 8888 10106 8900
rect 10321 8891 10379 8897
rect 10321 8888 10333 8891
rect 10100 8860 10333 8888
rect 10100 8848 10106 8860
rect 10321 8857 10333 8860
rect 10367 8857 10379 8891
rect 10321 8851 10379 8857
rect 1670 8820 1676 8832
rect 1631 8792 1676 8820
rect 1670 8780 1676 8792
rect 1728 8780 1734 8832
rect 4801 8823 4859 8829
rect 4801 8789 4813 8823
rect 4847 8820 4859 8823
rect 5534 8820 5540 8832
rect 4847 8792 5540 8820
rect 4847 8789 4859 8792
rect 4801 8783 4859 8789
rect 5534 8780 5540 8792
rect 5592 8780 5598 8832
rect 6546 8780 6552 8832
rect 6604 8829 6610 8832
rect 6604 8823 6653 8829
rect 6604 8789 6607 8823
rect 6641 8789 6653 8823
rect 6730 8820 6736 8832
rect 6691 8792 6736 8820
rect 6604 8783 6653 8789
rect 6604 8780 6610 8783
rect 6730 8780 6736 8792
rect 6788 8780 6794 8832
rect 7098 8820 7104 8832
rect 7059 8792 7104 8820
rect 7098 8780 7104 8792
rect 7156 8780 7162 8832
rect 7745 8823 7803 8829
rect 7745 8789 7757 8823
rect 7791 8820 7803 8823
rect 9033 8823 9091 8829
rect 9033 8820 9045 8823
rect 7791 8792 9045 8820
rect 7791 8789 7803 8792
rect 7745 8783 7803 8789
rect 9033 8789 9045 8792
rect 9079 8789 9091 8823
rect 9033 8783 9091 8789
rect 9766 8780 9772 8832
rect 9824 8820 9830 8832
rect 10686 8820 10692 8832
rect 9824 8792 10692 8820
rect 9824 8780 9830 8792
rect 10686 8780 10692 8792
rect 10744 8780 10750 8832
rect 14274 8820 14280 8832
rect 14235 8792 14280 8820
rect 14274 8780 14280 8792
rect 14332 8780 14338 8832
rect 14366 8780 14372 8832
rect 14424 8820 14430 8832
rect 14553 8823 14611 8829
rect 14553 8820 14565 8823
rect 14424 8792 14565 8820
rect 14424 8780 14430 8792
rect 14553 8789 14565 8792
rect 14599 8789 14611 8823
rect 14553 8783 14611 8789
rect 17175 8823 17233 8829
rect 17175 8789 17187 8823
rect 17221 8820 17233 8823
rect 17310 8820 17316 8832
rect 17221 8792 17316 8820
rect 17221 8789 17233 8792
rect 17175 8783 17233 8789
rect 17310 8780 17316 8792
rect 17368 8780 17374 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 4341 8619 4399 8625
rect 4341 8585 4353 8619
rect 4387 8616 4399 8619
rect 4706 8616 4712 8628
rect 4387 8588 4712 8616
rect 4387 8585 4399 8588
rect 4341 8579 4399 8585
rect 4706 8576 4712 8588
rect 4764 8576 4770 8628
rect 5442 8616 5448 8628
rect 5184 8588 5448 8616
rect 3329 8551 3387 8557
rect 3329 8517 3341 8551
rect 3375 8548 3387 8551
rect 4154 8548 4160 8560
rect 3375 8520 4160 8548
rect 3375 8517 3387 8520
rect 3329 8511 3387 8517
rect 4154 8508 4160 8520
rect 4212 8508 4218 8560
rect 3697 8483 3755 8489
rect 3697 8449 3709 8483
rect 3743 8480 3755 8483
rect 5184 8480 5212 8588
rect 5442 8576 5448 8588
rect 5500 8576 5506 8628
rect 6362 8576 6368 8628
rect 6420 8616 6426 8628
rect 10042 8616 10048 8628
rect 6420 8588 10048 8616
rect 6420 8576 6426 8588
rect 10042 8576 10048 8588
rect 10100 8576 10106 8628
rect 11701 8619 11759 8625
rect 11701 8585 11713 8619
rect 11747 8616 11759 8619
rect 11790 8616 11796 8628
rect 11747 8588 11796 8616
rect 11747 8585 11759 8588
rect 11701 8579 11759 8585
rect 11790 8576 11796 8588
rect 11848 8576 11854 8628
rect 13446 8576 13452 8628
rect 13504 8616 13510 8628
rect 13633 8619 13691 8625
rect 13633 8616 13645 8619
rect 13504 8588 13645 8616
rect 13504 8576 13510 8588
rect 13633 8585 13645 8588
rect 13679 8585 13691 8619
rect 16758 8616 16764 8628
rect 16719 8588 16764 8616
rect 13633 8579 13691 8585
rect 16758 8576 16764 8588
rect 16816 8576 16822 8628
rect 17126 8616 17132 8628
rect 17087 8588 17132 8616
rect 17126 8576 17132 8588
rect 17184 8576 17190 8628
rect 5258 8508 5264 8560
rect 5316 8548 5322 8560
rect 5629 8551 5687 8557
rect 5629 8548 5641 8551
rect 5316 8520 5641 8548
rect 5316 8508 5322 8520
rect 5629 8517 5641 8520
rect 5675 8517 5687 8551
rect 5629 8511 5687 8517
rect 6638 8508 6644 8560
rect 6696 8548 6702 8560
rect 7009 8551 7067 8557
rect 7009 8548 7021 8551
rect 6696 8520 7021 8548
rect 6696 8508 6702 8520
rect 7009 8517 7021 8520
rect 7055 8517 7067 8551
rect 7009 8511 7067 8517
rect 7098 8508 7104 8560
rect 7156 8548 7162 8560
rect 11238 8548 11244 8560
rect 7156 8520 11244 8548
rect 7156 8508 7162 8520
rect 11238 8508 11244 8520
rect 11296 8548 11302 8560
rect 11882 8548 11888 8560
rect 11296 8520 11888 8548
rect 11296 8508 11302 8520
rect 11882 8508 11888 8520
rect 11940 8548 11946 8560
rect 11977 8551 12035 8557
rect 11977 8548 11989 8551
rect 11940 8520 11989 8548
rect 11940 8508 11946 8520
rect 11977 8517 11989 8520
rect 12023 8517 12035 8551
rect 13262 8548 13268 8560
rect 13223 8520 13268 8548
rect 11977 8511 12035 8517
rect 13262 8508 13268 8520
rect 13320 8508 13326 8560
rect 24762 8548 24768 8560
rect 24723 8520 24768 8548
rect 24762 8508 24768 8520
rect 24820 8508 24826 8560
rect 5534 8480 5540 8492
rect 3743 8452 5212 8480
rect 5495 8452 5540 8480
rect 3743 8449 3755 8452
rect 3697 8443 3755 8449
rect 1581 8415 1639 8421
rect 1581 8381 1593 8415
rect 1627 8412 1639 8415
rect 1670 8412 1676 8424
rect 1627 8384 1676 8412
rect 1627 8381 1639 8384
rect 1581 8375 1639 8381
rect 1670 8372 1676 8384
rect 1728 8372 1734 8424
rect 1762 8372 1768 8424
rect 1820 8412 1826 8424
rect 2406 8412 2412 8424
rect 1820 8384 2412 8412
rect 1820 8372 1826 8384
rect 2406 8372 2412 8384
rect 2464 8372 2470 8424
rect 3145 8415 3203 8421
rect 3145 8381 3157 8415
rect 3191 8412 3203 8415
rect 3712 8412 3740 8443
rect 5534 8440 5540 8452
rect 5592 8440 5598 8492
rect 7926 8440 7932 8492
rect 7984 8480 7990 8492
rect 8297 8483 8355 8489
rect 8297 8480 8309 8483
rect 7984 8452 8309 8480
rect 7984 8440 7990 8452
rect 8297 8449 8309 8452
rect 8343 8449 8355 8483
rect 9766 8480 9772 8492
rect 9727 8452 9772 8480
rect 8297 8443 8355 8449
rect 9766 8440 9772 8452
rect 9824 8440 9830 8492
rect 14921 8483 14979 8489
rect 14921 8449 14933 8483
rect 14967 8480 14979 8483
rect 15286 8480 15292 8492
rect 14967 8452 15292 8480
rect 14967 8449 14979 8452
rect 14921 8443 14979 8449
rect 15286 8440 15292 8452
rect 15344 8440 15350 8492
rect 15565 8483 15623 8489
rect 15565 8449 15577 8483
rect 15611 8480 15623 8483
rect 15654 8480 15660 8492
rect 15611 8452 15660 8480
rect 15611 8449 15623 8452
rect 15565 8443 15623 8449
rect 15654 8440 15660 8452
rect 15712 8480 15718 8492
rect 15749 8483 15807 8489
rect 15749 8480 15761 8483
rect 15712 8452 15761 8480
rect 15712 8440 15718 8452
rect 15749 8449 15761 8452
rect 15795 8449 15807 8483
rect 15749 8443 15807 8449
rect 4062 8412 4068 8424
rect 3191 8384 3740 8412
rect 3975 8384 4068 8412
rect 3191 8381 3203 8384
rect 3145 8375 3203 8381
rect 2133 8347 2191 8353
rect 2133 8313 2145 8347
rect 2179 8344 2191 8347
rect 3878 8344 3884 8356
rect 2179 8316 3884 8344
rect 2179 8313 2191 8316
rect 2133 8307 2191 8313
rect 3878 8304 3884 8316
rect 3936 8304 3942 8356
rect 2958 8276 2964 8288
rect 2919 8248 2964 8276
rect 2958 8236 2964 8248
rect 3016 8276 3022 8288
rect 3988 8285 4016 8384
rect 4062 8372 4068 8384
rect 4120 8412 4126 8424
rect 4157 8415 4215 8421
rect 4157 8412 4169 8415
rect 4120 8384 4169 8412
rect 4120 8372 4126 8384
rect 4157 8381 4169 8384
rect 4203 8381 4215 8415
rect 4157 8375 4215 8381
rect 4522 8372 4528 8424
rect 4580 8412 4586 8424
rect 5350 8421 5356 8424
rect 5316 8415 5356 8421
rect 5316 8412 5328 8415
rect 4580 8384 5328 8412
rect 4580 8372 4586 8384
rect 5316 8381 5328 8384
rect 5316 8375 5356 8381
rect 5350 8372 5356 8375
rect 5408 8372 5414 8424
rect 7282 8412 7288 8424
rect 7243 8384 7288 8412
rect 7282 8372 7288 8384
rect 7340 8372 7346 8424
rect 7834 8412 7840 8424
rect 7795 8384 7840 8412
rect 7834 8372 7840 8384
rect 7892 8412 7898 8424
rect 8665 8415 8723 8421
rect 8665 8412 8677 8415
rect 7892 8384 8677 8412
rect 7892 8372 7898 8384
rect 8665 8381 8677 8384
rect 8711 8381 8723 8415
rect 9122 8412 9128 8424
rect 9083 8384 9128 8412
rect 8665 8375 8723 8381
rect 9122 8372 9128 8384
rect 9180 8372 9186 8424
rect 9490 8412 9496 8424
rect 9451 8384 9496 8412
rect 9490 8372 9496 8384
rect 9548 8372 9554 8424
rect 10321 8415 10379 8421
rect 10321 8381 10333 8415
rect 10367 8412 10379 8415
rect 10597 8415 10655 8421
rect 10597 8412 10609 8415
rect 10367 8384 10609 8412
rect 10367 8381 10379 8384
rect 10321 8375 10379 8381
rect 10597 8381 10609 8384
rect 10643 8381 10655 8415
rect 10597 8375 10655 8381
rect 11057 8415 11115 8421
rect 11057 8381 11069 8415
rect 11103 8381 11115 8415
rect 16298 8412 16304 8424
rect 16259 8384 16304 8412
rect 11057 8375 11115 8381
rect 4430 8304 4436 8356
rect 4488 8344 4494 8356
rect 5169 8347 5227 8353
rect 5169 8344 5181 8347
rect 4488 8316 5181 8344
rect 4488 8304 4494 8316
rect 5169 8313 5181 8316
rect 5215 8344 5227 8347
rect 5626 8344 5632 8356
rect 5215 8316 5632 8344
rect 5215 8313 5227 8316
rect 5169 8307 5227 8313
rect 5626 8304 5632 8316
rect 5684 8304 5690 8356
rect 8018 8344 8024 8356
rect 7979 8316 8024 8344
rect 8018 8304 8024 8316
rect 8076 8304 8082 8356
rect 10042 8304 10048 8356
rect 10100 8344 10106 8356
rect 11072 8344 11100 8375
rect 16298 8372 16304 8384
rect 16356 8372 16362 8424
rect 24118 8372 24124 8424
rect 24176 8412 24182 8424
rect 24581 8415 24639 8421
rect 24581 8412 24593 8415
rect 24176 8384 24593 8412
rect 24176 8372 24182 8384
rect 24581 8381 24593 8384
rect 24627 8412 24639 8415
rect 25133 8415 25191 8421
rect 25133 8412 25145 8415
rect 24627 8384 25145 8412
rect 24627 8381 24639 8384
rect 24581 8375 24639 8381
rect 25133 8381 25145 8384
rect 25179 8381 25191 8415
rect 25133 8375 25191 8381
rect 11330 8344 11336 8356
rect 10100 8316 11100 8344
rect 11291 8316 11336 8344
rect 10100 8304 10106 8316
rect 11330 8304 11336 8316
rect 11388 8304 11394 8356
rect 12710 8344 12716 8356
rect 12671 8316 12716 8344
rect 12710 8304 12716 8316
rect 12768 8304 12774 8356
rect 12805 8347 12863 8353
rect 12805 8313 12817 8347
rect 12851 8344 12863 8347
rect 13354 8344 13360 8356
rect 12851 8316 13360 8344
rect 12851 8313 12863 8316
rect 12805 8307 12863 8313
rect 13354 8304 13360 8316
rect 13412 8304 13418 8356
rect 14274 8344 14280 8356
rect 14235 8316 14280 8344
rect 14274 8304 14280 8316
rect 14332 8304 14338 8356
rect 14369 8347 14427 8353
rect 14369 8313 14381 8347
rect 14415 8344 14427 8347
rect 14458 8344 14464 8356
rect 14415 8316 14464 8344
rect 14415 8313 14427 8316
rect 14369 8307 14427 8313
rect 3973 8279 4031 8285
rect 3973 8276 3985 8279
rect 3016 8248 3985 8276
rect 3016 8236 3022 8248
rect 3973 8245 3985 8248
rect 4019 8245 4031 8279
rect 4982 8276 4988 8288
rect 4943 8248 4988 8276
rect 3973 8239 4031 8245
rect 4982 8236 4988 8248
rect 5040 8236 5046 8288
rect 6546 8276 6552 8288
rect 6507 8248 6552 8276
rect 6546 8236 6552 8248
rect 6604 8236 6610 8288
rect 8110 8236 8116 8288
rect 8168 8276 8174 8288
rect 9674 8276 9680 8288
rect 8168 8248 9680 8276
rect 8168 8236 8174 8248
rect 9674 8236 9680 8248
rect 9732 8276 9738 8288
rect 10321 8279 10379 8285
rect 10321 8276 10333 8279
rect 9732 8248 10333 8276
rect 9732 8236 9738 8248
rect 10321 8245 10333 8248
rect 10367 8276 10379 8279
rect 10413 8279 10471 8285
rect 10413 8276 10425 8279
rect 10367 8248 10425 8276
rect 10367 8245 10379 8248
rect 10321 8239 10379 8245
rect 10413 8245 10425 8248
rect 10459 8245 10471 8279
rect 10413 8239 10471 8245
rect 14093 8279 14151 8285
rect 14093 8245 14105 8279
rect 14139 8276 14151 8279
rect 14384 8276 14412 8307
rect 14458 8304 14464 8316
rect 14516 8304 14522 8356
rect 24026 8276 24032 8288
rect 14139 8248 14412 8276
rect 23987 8248 24032 8276
rect 14139 8245 14151 8248
rect 14093 8239 14151 8245
rect 24026 8236 24032 8248
rect 24084 8236 24090 8288
rect 24489 8279 24547 8285
rect 24489 8245 24501 8279
rect 24535 8276 24547 8279
rect 24854 8276 24860 8288
rect 24535 8248 24860 8276
rect 24535 8245 24547 8248
rect 24489 8239 24547 8245
rect 24854 8236 24860 8248
rect 24912 8236 24918 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1670 8032 1676 8084
rect 1728 8072 1734 8084
rect 2225 8075 2283 8081
rect 2225 8072 2237 8075
rect 1728 8044 2237 8072
rect 1728 8032 1734 8044
rect 2225 8041 2237 8044
rect 2271 8041 2283 8075
rect 2225 8035 2283 8041
rect 2866 8032 2872 8084
rect 2924 8072 2930 8084
rect 3145 8075 3203 8081
rect 3145 8072 3157 8075
rect 2924 8044 3157 8072
rect 2924 8032 2930 8044
rect 3145 8041 3157 8044
rect 3191 8041 3203 8075
rect 4522 8072 4528 8084
rect 4483 8044 4528 8072
rect 3145 8035 3203 8041
rect 4522 8032 4528 8044
rect 4580 8032 4586 8084
rect 5442 8032 5448 8084
rect 5500 8072 5506 8084
rect 5813 8075 5871 8081
rect 5813 8072 5825 8075
rect 5500 8044 5825 8072
rect 5500 8032 5506 8044
rect 5813 8041 5825 8044
rect 5859 8041 5871 8075
rect 5813 8035 5871 8041
rect 6549 8075 6607 8081
rect 6549 8041 6561 8075
rect 6595 8072 6607 8075
rect 8202 8072 8208 8084
rect 6595 8044 8208 8072
rect 6595 8041 6607 8044
rect 6549 8035 6607 8041
rect 8202 8032 8208 8044
rect 8260 8032 8266 8084
rect 8294 8032 8300 8084
rect 8352 8072 8358 8084
rect 9033 8075 9091 8081
rect 9033 8072 9045 8075
rect 8352 8044 9045 8072
rect 8352 8032 8358 8044
rect 9033 8041 9045 8044
rect 9079 8072 9091 8075
rect 9490 8072 9496 8084
rect 9079 8044 9496 8072
rect 9079 8041 9091 8044
rect 9033 8035 9091 8041
rect 9490 8032 9496 8044
rect 9548 8032 9554 8084
rect 9858 8032 9864 8084
rect 9916 8072 9922 8084
rect 10781 8075 10839 8081
rect 10781 8072 10793 8075
rect 9916 8044 10793 8072
rect 9916 8032 9922 8044
rect 10781 8041 10793 8044
rect 10827 8041 10839 8075
rect 10781 8035 10839 8041
rect 11241 8075 11299 8081
rect 11241 8041 11253 8075
rect 11287 8072 11299 8075
rect 11330 8072 11336 8084
rect 11287 8044 11336 8072
rect 11287 8041 11299 8044
rect 11241 8035 11299 8041
rect 11330 8032 11336 8044
rect 11388 8032 11394 8084
rect 12986 8032 12992 8084
rect 13044 8072 13050 8084
rect 14093 8075 14151 8081
rect 14093 8072 14105 8075
rect 13044 8044 14105 8072
rect 13044 8032 13050 8044
rect 14093 8041 14105 8044
rect 14139 8041 14151 8075
rect 14550 8072 14556 8084
rect 14511 8044 14556 8072
rect 14093 8035 14151 8041
rect 14550 8032 14556 8044
rect 14608 8032 14614 8084
rect 16298 8072 16304 8084
rect 16259 8044 16304 8072
rect 16298 8032 16304 8044
rect 16356 8032 16362 8084
rect 1535 8007 1593 8013
rect 1535 7973 1547 8007
rect 1581 8004 1593 8007
rect 8938 8004 8944 8016
rect 1581 7976 8944 8004
rect 1581 7973 1593 7976
rect 1535 7967 1593 7973
rect 8938 7964 8944 7976
rect 8996 7964 9002 8016
rect 9122 7964 9128 8016
rect 9180 8004 9186 8016
rect 9401 8007 9459 8013
rect 9401 8004 9413 8007
rect 9180 7976 9413 8004
rect 9180 7964 9186 7976
rect 9401 7973 9413 7976
rect 9447 8004 9459 8007
rect 9447 7976 9812 8004
rect 9447 7973 9459 7976
rect 9401 7967 9459 7973
rect 106 7896 112 7948
rect 164 7936 170 7948
rect 1432 7939 1490 7945
rect 1432 7936 1444 7939
rect 164 7908 1444 7936
rect 164 7896 170 7908
rect 1432 7905 1444 7908
rect 1478 7936 1490 7939
rect 2130 7936 2136 7948
rect 1478 7908 2136 7936
rect 1478 7905 1490 7908
rect 1432 7899 1490 7905
rect 2130 7896 2136 7908
rect 2188 7896 2194 7948
rect 2958 7936 2964 7948
rect 2919 7908 2964 7936
rect 2958 7896 2964 7908
rect 3016 7896 3022 7948
rect 4982 7936 4988 7948
rect 4943 7908 4988 7936
rect 4982 7896 4988 7908
rect 5040 7896 5046 7948
rect 5537 7939 5595 7945
rect 5537 7905 5549 7939
rect 5583 7936 5595 7939
rect 5626 7936 5632 7948
rect 5583 7908 5632 7936
rect 5583 7905 5595 7908
rect 5537 7899 5595 7905
rect 5626 7896 5632 7908
rect 5684 7896 5690 7948
rect 6822 7896 6828 7948
rect 6880 7936 6886 7948
rect 7009 7939 7067 7945
rect 7009 7936 7021 7939
rect 6880 7908 7021 7936
rect 6880 7896 6886 7908
rect 7009 7905 7021 7908
rect 7055 7905 7067 7939
rect 7009 7899 7067 7905
rect 7282 7896 7288 7948
rect 7340 7936 7346 7948
rect 7377 7939 7435 7945
rect 7377 7936 7389 7939
rect 7340 7908 7389 7936
rect 7340 7896 7346 7908
rect 7377 7905 7389 7908
rect 7423 7905 7435 7939
rect 7377 7899 7435 7905
rect 7466 7896 7472 7948
rect 7524 7936 7530 7948
rect 7561 7939 7619 7945
rect 7561 7936 7573 7939
rect 7524 7908 7573 7936
rect 7524 7896 7530 7908
rect 7561 7905 7573 7908
rect 7607 7905 7619 7939
rect 7561 7899 7619 7905
rect 7834 7896 7840 7948
rect 7892 7936 7898 7948
rect 8021 7939 8079 7945
rect 8021 7936 8033 7939
rect 7892 7908 8033 7936
rect 7892 7896 7898 7908
rect 8021 7905 8033 7908
rect 8067 7905 8079 7939
rect 9140 7936 9168 7964
rect 9784 7948 9812 7976
rect 9766 7936 9772 7948
rect 8021 7899 8079 7905
rect 8220 7908 9168 7936
rect 9679 7908 9772 7936
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7868 5319 7871
rect 8220 7868 8248 7908
rect 9766 7896 9772 7908
rect 9824 7896 9830 7948
rect 10042 7896 10048 7948
rect 10100 7936 10106 7948
rect 11348 7945 11376 8032
rect 11695 8007 11753 8013
rect 11695 7973 11707 8007
rect 11741 8004 11753 8007
rect 11974 8004 11980 8016
rect 11741 7976 11980 8004
rect 11741 7973 11753 7976
rect 11695 7967 11753 7973
rect 11974 7964 11980 7976
rect 12032 7964 12038 8016
rect 13078 8004 13084 8016
rect 13039 7976 13084 8004
rect 13078 7964 13084 7976
rect 13136 7964 13142 8016
rect 14458 7964 14464 8016
rect 14516 8004 14522 8016
rect 15289 8007 15347 8013
rect 15289 8004 15301 8007
rect 14516 7976 15301 8004
rect 14516 7964 14522 7976
rect 15289 7973 15301 7976
rect 15335 7973 15347 8007
rect 15289 7967 15347 7973
rect 10229 7939 10287 7945
rect 10229 7936 10241 7939
rect 10100 7908 10241 7936
rect 10100 7896 10106 7908
rect 10229 7905 10241 7908
rect 10275 7905 10287 7939
rect 10229 7899 10287 7905
rect 11333 7939 11391 7945
rect 11333 7905 11345 7939
rect 11379 7905 11391 7939
rect 11333 7899 11391 7905
rect 12713 7939 12771 7945
rect 12713 7905 12725 7939
rect 12759 7936 12771 7939
rect 13354 7936 13360 7948
rect 12759 7908 13360 7936
rect 12759 7905 12771 7908
rect 12713 7899 12771 7905
rect 13354 7896 13360 7908
rect 13412 7896 13418 7948
rect 14826 7896 14832 7948
rect 14884 7936 14890 7948
rect 15378 7936 15384 7948
rect 14884 7908 15384 7936
rect 14884 7896 14890 7908
rect 15378 7896 15384 7908
rect 15436 7896 15442 7948
rect 5307 7840 8248 7868
rect 8297 7871 8355 7877
rect 5307 7837 5319 7840
rect 5261 7831 5319 7837
rect 8297 7837 8309 7871
rect 8343 7868 8355 7871
rect 8478 7868 8484 7880
rect 8343 7840 8484 7868
rect 8343 7837 8355 7840
rect 8297 7831 8355 7837
rect 8478 7828 8484 7840
rect 8536 7828 8542 7880
rect 10502 7868 10508 7880
rect 10463 7840 10508 7868
rect 10502 7828 10508 7840
rect 10560 7828 10566 7880
rect 4893 7803 4951 7809
rect 4893 7769 4905 7803
rect 4939 7800 4951 7803
rect 5534 7800 5540 7812
rect 4939 7772 5540 7800
rect 4939 7769 4951 7772
rect 4893 7763 4951 7769
rect 5534 7760 5540 7772
rect 5592 7800 5598 7812
rect 6178 7800 6184 7812
rect 5592 7772 6184 7800
rect 5592 7760 5598 7772
rect 6178 7760 6184 7772
rect 6236 7760 6242 7812
rect 8110 7760 8116 7812
rect 8168 7800 8174 7812
rect 8573 7803 8631 7809
rect 8573 7800 8585 7803
rect 8168 7772 8585 7800
rect 8168 7760 8174 7772
rect 8573 7769 8585 7772
rect 8619 7769 8631 7803
rect 8573 7763 8631 7769
rect 1026 7692 1032 7744
rect 1084 7732 1090 7744
rect 1578 7732 1584 7744
rect 1084 7704 1584 7732
rect 1084 7692 1090 7704
rect 1578 7692 1584 7704
rect 1636 7732 1642 7744
rect 1857 7735 1915 7741
rect 1857 7732 1869 7735
rect 1636 7704 1869 7732
rect 1636 7692 1642 7704
rect 1857 7701 1869 7704
rect 1903 7701 1915 7735
rect 1857 7695 1915 7701
rect 5169 7735 5227 7741
rect 5169 7701 5181 7735
rect 5215 7732 5227 7735
rect 5261 7735 5319 7741
rect 5261 7732 5273 7735
rect 5215 7704 5273 7732
rect 5215 7701 5227 7704
rect 5169 7695 5227 7701
rect 5261 7701 5273 7704
rect 5307 7701 5319 7735
rect 5261 7695 5319 7701
rect 6270 7692 6276 7744
rect 6328 7732 6334 7744
rect 6365 7735 6423 7741
rect 6365 7732 6377 7735
rect 6328 7704 6377 7732
rect 6328 7692 6334 7704
rect 6365 7701 6377 7704
rect 6411 7701 6423 7735
rect 6365 7695 6423 7701
rect 12253 7735 12311 7741
rect 12253 7701 12265 7735
rect 12299 7732 12311 7735
rect 13170 7732 13176 7744
rect 12299 7704 13176 7732
rect 12299 7701 12311 7704
rect 12253 7695 12311 7701
rect 13170 7692 13176 7704
rect 13228 7692 13234 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1486 7488 1492 7540
rect 1544 7528 1550 7540
rect 1811 7531 1869 7537
rect 1811 7528 1823 7531
rect 1544 7500 1823 7528
rect 1544 7488 1550 7500
rect 1811 7497 1823 7500
rect 1857 7497 1869 7531
rect 2130 7528 2136 7540
rect 2091 7500 2136 7528
rect 1811 7491 1869 7497
rect 2130 7488 2136 7500
rect 2188 7488 2194 7540
rect 2958 7528 2964 7540
rect 2919 7500 2964 7528
rect 2958 7488 2964 7500
rect 3016 7488 3022 7540
rect 3786 7488 3792 7540
rect 3844 7528 3850 7540
rect 4065 7531 4123 7537
rect 4065 7528 4077 7531
rect 3844 7500 4077 7528
rect 3844 7488 3850 7500
rect 4065 7497 4077 7500
rect 4111 7497 4123 7531
rect 4065 7491 4123 7497
rect 4890 7488 4896 7540
rect 4948 7528 4954 7540
rect 5077 7531 5135 7537
rect 5077 7528 5089 7531
rect 4948 7500 5089 7528
rect 4948 7488 4954 7500
rect 5077 7497 5089 7500
rect 5123 7497 5135 7531
rect 5077 7491 5135 7497
rect 5350 7488 5356 7540
rect 5408 7528 5414 7540
rect 5721 7531 5779 7537
rect 5721 7528 5733 7531
rect 5408 7500 5733 7528
rect 5408 7488 5414 7500
rect 5721 7497 5733 7500
rect 5767 7497 5779 7531
rect 5721 7491 5779 7497
rect 8294 7488 8300 7540
rect 8352 7528 8358 7540
rect 8481 7531 8539 7537
rect 8481 7528 8493 7531
rect 8352 7500 8493 7528
rect 8352 7488 8358 7500
rect 8481 7497 8493 7500
rect 8527 7497 8539 7531
rect 9766 7528 9772 7540
rect 9727 7500 9772 7528
rect 8481 7491 8539 7497
rect 9766 7488 9772 7500
rect 9824 7488 9830 7540
rect 10042 7488 10048 7540
rect 10100 7528 10106 7540
rect 10137 7531 10195 7537
rect 10137 7528 10149 7531
rect 10100 7500 10149 7528
rect 10100 7488 10106 7500
rect 10137 7497 10149 7500
rect 10183 7497 10195 7531
rect 10137 7491 10195 7497
rect 11885 7531 11943 7537
rect 11885 7497 11897 7531
rect 11931 7528 11943 7531
rect 11974 7528 11980 7540
rect 11931 7500 11980 7528
rect 11931 7497 11943 7500
rect 11885 7491 11943 7497
rect 11974 7488 11980 7500
rect 12032 7528 12038 7540
rect 12161 7531 12219 7537
rect 12161 7528 12173 7531
rect 12032 7500 12173 7528
rect 12032 7488 12038 7500
rect 12161 7497 12173 7500
rect 12207 7497 12219 7531
rect 12161 7491 12219 7497
rect 13354 7488 13360 7540
rect 13412 7528 13418 7540
rect 13633 7531 13691 7537
rect 13633 7528 13645 7531
rect 13412 7500 13645 7528
rect 13412 7488 13418 7500
rect 13633 7497 13645 7500
rect 13679 7497 13691 7531
rect 15378 7528 15384 7540
rect 15339 7500 15384 7528
rect 13633 7491 13691 7497
rect 15378 7488 15384 7500
rect 15436 7488 15442 7540
rect 24719 7531 24777 7537
rect 24719 7497 24731 7531
rect 24765 7528 24777 7531
rect 24854 7528 24860 7540
rect 24765 7500 24860 7528
rect 24765 7497 24777 7500
rect 24719 7491 24777 7497
rect 24854 7488 24860 7500
rect 24912 7488 24918 7540
rect 2593 7395 2651 7401
rect 2593 7392 2605 7395
rect 1755 7364 2605 7392
rect 1755 7333 1783 7364
rect 2593 7361 2605 7364
rect 2639 7392 2651 7395
rect 5074 7392 5080 7404
rect 2639 7364 5080 7392
rect 2639 7361 2651 7364
rect 2593 7355 2651 7361
rect 5074 7352 5080 7364
rect 5132 7352 5138 7404
rect 1740 7327 1798 7333
rect 1740 7293 1752 7327
rect 1786 7293 1798 7327
rect 3878 7324 3884 7336
rect 3839 7296 3884 7324
rect 1740 7287 1798 7293
rect 3878 7284 3884 7296
rect 3936 7324 3942 7336
rect 4341 7327 4399 7333
rect 4341 7324 4353 7327
rect 3936 7296 4353 7324
rect 3936 7284 3942 7296
rect 4341 7293 4353 7296
rect 4387 7293 4399 7327
rect 4341 7287 4399 7293
rect 4893 7327 4951 7333
rect 4893 7293 4905 7327
rect 4939 7324 4951 7327
rect 5368 7324 5396 7488
rect 6914 7352 6920 7404
rect 6972 7392 6978 7404
rect 6972 7364 7604 7392
rect 6972 7352 6978 7364
rect 7101 7327 7159 7333
rect 7101 7324 7113 7327
rect 4939 7296 5396 7324
rect 6564 7296 7113 7324
rect 4939 7293 4951 7296
rect 4893 7287 4951 7293
rect 4614 7216 4620 7268
rect 4672 7256 4678 7268
rect 4982 7256 4988 7268
rect 4672 7228 4988 7256
rect 4672 7216 4678 7228
rect 4982 7216 4988 7228
rect 5040 7256 5046 7268
rect 5353 7259 5411 7265
rect 5353 7256 5365 7259
rect 5040 7228 5365 7256
rect 5040 7216 5046 7228
rect 5353 7225 5365 7228
rect 5399 7225 5411 7259
rect 5353 7219 5411 7225
rect 6454 7148 6460 7200
rect 6512 7188 6518 7200
rect 6564 7197 6592 7296
rect 7101 7293 7113 7296
rect 7147 7324 7159 7327
rect 7282 7324 7288 7336
rect 7147 7296 7288 7324
rect 7147 7293 7159 7296
rect 7101 7287 7159 7293
rect 7282 7284 7288 7296
rect 7340 7284 7346 7336
rect 7576 7333 7604 7364
rect 10502 7352 10508 7404
rect 10560 7392 10566 7404
rect 12434 7392 12440 7404
rect 10560 7364 12440 7392
rect 10560 7352 10566 7364
rect 12434 7352 12440 7364
rect 12492 7352 12498 7404
rect 14277 7395 14335 7401
rect 14277 7361 14289 7395
rect 14323 7392 14335 7395
rect 14366 7392 14372 7404
rect 14323 7364 14372 7392
rect 14323 7361 14335 7364
rect 14277 7355 14335 7361
rect 14366 7352 14372 7364
rect 14424 7352 14430 7404
rect 14550 7392 14556 7404
rect 14511 7364 14556 7392
rect 14550 7352 14556 7364
rect 14608 7352 14614 7404
rect 7561 7327 7619 7333
rect 7561 7293 7573 7327
rect 7607 7324 7619 7327
rect 7926 7324 7932 7336
rect 7607 7296 7932 7324
rect 7607 7293 7619 7296
rect 7561 7287 7619 7293
rect 7926 7284 7932 7296
rect 7984 7284 7990 7336
rect 10781 7327 10839 7333
rect 10781 7324 10793 7327
rect 10612 7296 10793 7324
rect 7466 7216 7472 7268
rect 7524 7256 7530 7268
rect 8113 7259 8171 7265
rect 8113 7256 8125 7259
rect 7524 7228 8125 7256
rect 7524 7216 7530 7228
rect 8113 7225 8125 7228
rect 8159 7225 8171 7259
rect 8754 7256 8760 7268
rect 8715 7228 8760 7256
rect 8113 7219 8171 7225
rect 8754 7216 8760 7228
rect 8812 7216 8818 7268
rect 8846 7216 8852 7268
rect 8904 7256 8910 7268
rect 9398 7256 9404 7268
rect 8904 7228 8949 7256
rect 9359 7228 9404 7256
rect 8904 7216 8910 7228
rect 9398 7216 9404 7228
rect 9456 7216 9462 7268
rect 6549 7191 6607 7197
rect 6549 7188 6561 7191
rect 6512 7160 6561 7188
rect 6512 7148 6518 7160
rect 6549 7157 6561 7160
rect 6595 7157 6607 7191
rect 6549 7151 6607 7157
rect 7377 7191 7435 7197
rect 7377 7157 7389 7191
rect 7423 7188 7435 7191
rect 7558 7188 7564 7200
rect 7423 7160 7564 7188
rect 7423 7157 7435 7160
rect 7377 7151 7435 7157
rect 7558 7148 7564 7160
rect 7616 7148 7622 7200
rect 9306 7148 9312 7200
rect 9364 7188 9370 7200
rect 10612 7197 10640 7296
rect 10781 7293 10793 7296
rect 10827 7324 10839 7327
rect 10870 7324 10876 7336
rect 10827 7296 10876 7324
rect 10827 7293 10839 7296
rect 10781 7287 10839 7293
rect 10870 7284 10876 7296
rect 10928 7284 10934 7336
rect 11238 7324 11244 7336
rect 11199 7296 11244 7324
rect 11238 7284 11244 7296
rect 11296 7284 11302 7336
rect 11974 7284 11980 7336
rect 12032 7324 12038 7336
rect 24648 7327 24706 7333
rect 12032 7296 12801 7324
rect 12032 7284 12038 7296
rect 11517 7259 11575 7265
rect 11517 7225 11529 7259
rect 11563 7256 11575 7259
rect 12250 7256 12256 7268
rect 11563 7228 12256 7256
rect 11563 7225 11575 7228
rect 11517 7219 11575 7225
rect 12250 7216 12256 7228
rect 12308 7216 12314 7268
rect 12773 7265 12801 7296
rect 24648 7293 24660 7327
rect 24694 7324 24706 7327
rect 24694 7296 25176 7324
rect 24694 7293 24706 7296
rect 24648 7287 24706 7293
rect 12758 7259 12816 7265
rect 12758 7225 12770 7259
rect 12804 7225 12816 7259
rect 12758 7219 12816 7225
rect 14369 7259 14427 7265
rect 14369 7225 14381 7259
rect 14415 7256 14427 7259
rect 14642 7256 14648 7268
rect 14415 7228 14648 7256
rect 14415 7225 14427 7228
rect 14369 7219 14427 7225
rect 10597 7191 10655 7197
rect 10597 7188 10609 7191
rect 9364 7160 10609 7188
rect 9364 7148 9370 7160
rect 10597 7157 10609 7160
rect 10643 7157 10655 7191
rect 13354 7188 13360 7200
rect 13315 7160 13360 7188
rect 10597 7151 10655 7157
rect 13354 7148 13360 7160
rect 13412 7148 13418 7200
rect 14093 7191 14151 7197
rect 14093 7157 14105 7191
rect 14139 7188 14151 7191
rect 14384 7188 14412 7219
rect 14642 7216 14648 7228
rect 14700 7216 14706 7268
rect 25148 7200 25176 7296
rect 25130 7188 25136 7200
rect 14139 7160 14412 7188
rect 25091 7160 25136 7188
rect 14139 7157 14151 7160
rect 14093 7151 14151 7157
rect 25130 7148 25136 7160
rect 25188 7148 25194 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 1394 6944 1400 6996
rect 1452 6984 1458 6996
rect 1903 6987 1961 6993
rect 1903 6984 1915 6987
rect 1452 6956 1915 6984
rect 1452 6944 1458 6956
rect 1903 6953 1915 6956
rect 1949 6953 1961 6987
rect 4798 6984 4804 6996
rect 4759 6956 4804 6984
rect 1903 6947 1961 6953
rect 4798 6944 4804 6956
rect 4856 6984 4862 6996
rect 6454 6984 6460 6996
rect 4856 6956 6460 6984
rect 4856 6944 4862 6956
rect 6454 6944 6460 6956
rect 6512 6944 6518 6996
rect 6914 6944 6920 6996
rect 6972 6984 6978 6996
rect 7101 6987 7159 6993
rect 7101 6984 7113 6987
rect 6972 6956 7113 6984
rect 6972 6944 6978 6956
rect 7101 6953 7113 6956
rect 7147 6953 7159 6987
rect 7101 6947 7159 6953
rect 7653 6987 7711 6993
rect 7653 6953 7665 6987
rect 7699 6984 7711 6987
rect 7834 6984 7840 6996
rect 7699 6956 7840 6984
rect 7699 6953 7711 6956
rect 7653 6947 7711 6953
rect 7834 6944 7840 6956
rect 7892 6944 7898 6996
rect 8202 6984 8208 6996
rect 8163 6956 8208 6984
rect 8202 6944 8208 6956
rect 8260 6944 8266 6996
rect 8754 6944 8760 6996
rect 8812 6984 8818 6996
rect 9401 6987 9459 6993
rect 9401 6984 9413 6987
rect 8812 6956 9413 6984
rect 8812 6944 8818 6956
rect 9401 6953 9413 6956
rect 9447 6953 9459 6987
rect 9950 6984 9956 6996
rect 9911 6956 9956 6984
rect 9401 6947 9459 6953
rect 9950 6944 9956 6956
rect 10008 6944 10014 6996
rect 10873 6987 10931 6993
rect 10873 6953 10885 6987
rect 10919 6984 10931 6987
rect 11238 6984 11244 6996
rect 10919 6956 11244 6984
rect 10919 6953 10931 6956
rect 10873 6947 10931 6953
rect 11238 6944 11244 6956
rect 11296 6944 11302 6996
rect 12434 6984 12440 6996
rect 12395 6956 12440 6984
rect 12434 6944 12440 6956
rect 12492 6944 12498 6996
rect 12710 6944 12716 6996
rect 12768 6984 12774 6996
rect 12805 6987 12863 6993
rect 12805 6984 12817 6987
rect 12768 6956 12817 6984
rect 12768 6944 12774 6956
rect 12805 6953 12817 6956
rect 12851 6953 12863 6987
rect 12805 6947 12863 6953
rect 13354 6876 13360 6928
rect 13412 6916 13418 6928
rect 13814 6916 13820 6928
rect 13412 6888 13820 6916
rect 13412 6876 13418 6888
rect 13814 6876 13820 6888
rect 13872 6916 13878 6928
rect 14369 6919 14427 6925
rect 13872 6888 13917 6916
rect 13872 6876 13878 6888
rect 14369 6885 14381 6919
rect 14415 6916 14427 6919
rect 14550 6916 14556 6928
rect 14415 6888 14556 6916
rect 14415 6885 14427 6888
rect 14369 6879 14427 6885
rect 1832 6851 1890 6857
rect 1832 6817 1844 6851
rect 1878 6848 1890 6851
rect 2682 6848 2688 6860
rect 1878 6820 2688 6848
rect 1878 6817 1890 6820
rect 1832 6811 1890 6817
rect 2682 6808 2688 6820
rect 2740 6808 2746 6860
rect 4614 6848 4620 6860
rect 4575 6820 4620 6848
rect 4614 6808 4620 6820
rect 4672 6808 4678 6860
rect 6089 6851 6147 6857
rect 6089 6817 6101 6851
rect 6135 6848 6147 6851
rect 6178 6848 6184 6860
rect 6135 6820 6184 6848
rect 6135 6817 6147 6820
rect 6089 6811 6147 6817
rect 6178 6808 6184 6820
rect 6236 6808 6242 6860
rect 9858 6848 9864 6860
rect 9819 6820 9864 6848
rect 9858 6808 9864 6820
rect 9916 6808 9922 6860
rect 11330 6848 11336 6860
rect 11291 6820 11336 6848
rect 11330 6808 11336 6820
rect 11388 6808 11394 6860
rect 7837 6783 7895 6789
rect 7837 6749 7849 6783
rect 7883 6780 7895 6783
rect 8018 6780 8024 6792
rect 7883 6752 8024 6780
rect 7883 6749 7895 6752
rect 7837 6743 7895 6749
rect 8018 6740 8024 6752
rect 8076 6740 8082 6792
rect 11238 6780 11244 6792
rect 11199 6752 11244 6780
rect 11238 6740 11244 6752
rect 11296 6740 11302 6792
rect 13722 6780 13728 6792
rect 13683 6752 13728 6780
rect 13722 6740 13728 6752
rect 13780 6740 13786 6792
rect 6270 6712 6276 6724
rect 6231 6684 6276 6712
rect 6270 6672 6276 6684
rect 6328 6672 6334 6724
rect 13446 6712 13452 6724
rect 13359 6684 13452 6712
rect 13446 6672 13452 6684
rect 13504 6712 13510 6724
rect 14384 6712 14412 6879
rect 14550 6876 14556 6888
rect 14608 6876 14614 6928
rect 14642 6876 14648 6928
rect 14700 6916 14706 6928
rect 15289 6919 15347 6925
rect 15289 6916 15301 6919
rect 14700 6888 15301 6916
rect 14700 6876 14706 6888
rect 15289 6885 15301 6888
rect 15335 6885 15347 6919
rect 15289 6879 15347 6885
rect 15930 6848 15936 6860
rect 15891 6820 15936 6848
rect 15930 6808 15936 6820
rect 15988 6808 15994 6860
rect 13504 6684 14412 6712
rect 13504 6672 13510 6684
rect 8294 6604 8300 6656
rect 8352 6644 8358 6656
rect 8757 6647 8815 6653
rect 8757 6644 8769 6647
rect 8352 6616 8769 6644
rect 8352 6604 8358 6616
rect 8757 6613 8769 6616
rect 8803 6644 8815 6647
rect 8846 6644 8852 6656
rect 8803 6616 8852 6644
rect 8803 6613 8815 6616
rect 8757 6607 8815 6613
rect 8846 6604 8852 6616
rect 8904 6644 8910 6656
rect 9033 6647 9091 6653
rect 9033 6644 9045 6647
rect 8904 6616 9045 6644
rect 8904 6604 8910 6616
rect 9033 6613 9045 6616
rect 9079 6613 9091 6647
rect 9033 6607 9091 6613
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 2317 6443 2375 6449
rect 2317 6409 2329 6443
rect 2363 6440 2375 6443
rect 2682 6440 2688 6452
rect 2363 6412 2688 6440
rect 2363 6409 2375 6412
rect 2317 6403 2375 6409
rect 2682 6400 2688 6412
rect 2740 6400 2746 6452
rect 6178 6440 6184 6452
rect 6139 6412 6184 6440
rect 6178 6400 6184 6412
rect 6236 6400 6242 6452
rect 9401 6443 9459 6449
rect 9401 6409 9413 6443
rect 9447 6440 9459 6443
rect 9858 6440 9864 6452
rect 9447 6412 9864 6440
rect 9447 6409 9459 6412
rect 9401 6403 9459 6409
rect 9858 6400 9864 6412
rect 9916 6440 9922 6452
rect 11330 6440 11336 6452
rect 9916 6412 11336 6440
rect 9916 6400 9922 6412
rect 11330 6400 11336 6412
rect 11388 6400 11394 6452
rect 13170 6440 13176 6452
rect 13131 6412 13176 6440
rect 13170 6400 13176 6412
rect 13228 6400 13234 6452
rect 13814 6400 13820 6452
rect 13872 6440 13878 6452
rect 14461 6443 14519 6449
rect 14461 6440 14473 6443
rect 13872 6412 14473 6440
rect 13872 6400 13878 6412
rect 14461 6409 14473 6412
rect 14507 6440 14519 6443
rect 15930 6440 15936 6452
rect 14507 6412 15936 6440
rect 14507 6409 14519 6412
rect 14461 6403 14519 6409
rect 15930 6400 15936 6412
rect 15988 6400 15994 6452
rect 1535 6375 1593 6381
rect 1535 6341 1547 6375
rect 1581 6372 1593 6375
rect 3234 6372 3240 6384
rect 1581 6344 3240 6372
rect 1581 6341 1593 6344
rect 1535 6335 1593 6341
rect 3234 6332 3240 6344
rect 3292 6332 3298 6384
rect 5353 6375 5411 6381
rect 5353 6341 5365 6375
rect 5399 6372 5411 6375
rect 9306 6372 9312 6384
rect 5399 6344 9312 6372
rect 5399 6341 5411 6344
rect 5353 6335 5411 6341
rect 9306 6332 9312 6344
rect 9364 6332 9370 6384
rect 9490 6332 9496 6384
rect 9548 6372 9554 6384
rect 10873 6375 10931 6381
rect 10873 6372 10885 6375
rect 9548 6344 10885 6372
rect 9548 6332 9554 6344
rect 10873 6341 10885 6344
rect 10919 6372 10931 6375
rect 11146 6372 11152 6384
rect 10919 6344 11152 6372
rect 10919 6341 10931 6344
rect 10873 6335 10931 6341
rect 11146 6332 11152 6344
rect 11204 6332 11210 6384
rect 7653 6307 7711 6313
rect 7653 6273 7665 6307
rect 7699 6304 7711 6307
rect 10045 6307 10103 6313
rect 10045 6304 10057 6307
rect 7699 6276 10057 6304
rect 7699 6273 7711 6276
rect 7653 6267 7711 6273
rect 10045 6273 10057 6276
rect 10091 6273 10103 6307
rect 10045 6267 10103 6273
rect 10321 6307 10379 6313
rect 10321 6273 10333 6307
rect 10367 6304 10379 6307
rect 10778 6304 10784 6316
rect 10367 6276 10784 6304
rect 10367 6273 10379 6276
rect 10321 6267 10379 6273
rect 1432 6239 1490 6245
rect 1432 6205 1444 6239
rect 1478 6205 1490 6239
rect 5169 6239 5227 6245
rect 5169 6236 5181 6239
rect 1432 6199 1490 6205
rect 4632 6208 5181 6236
rect 106 6128 112 6180
rect 164 6168 170 6180
rect 1447 6168 1475 6199
rect 1857 6171 1915 6177
rect 1857 6168 1869 6171
rect 164 6140 1869 6168
rect 164 6128 170 6140
rect 1857 6137 1869 6140
rect 1903 6137 1915 6171
rect 1857 6131 1915 6137
rect 4632 6112 4660 6208
rect 5169 6205 5181 6208
rect 5215 6236 5227 6239
rect 5629 6239 5687 6245
rect 5629 6236 5641 6239
rect 5215 6208 5641 6236
rect 5215 6205 5227 6208
rect 5169 6199 5227 6205
rect 5629 6205 5641 6208
rect 5675 6205 5687 6239
rect 5629 6199 5687 6205
rect 6641 6239 6699 6245
rect 6641 6205 6653 6239
rect 6687 6236 6699 6239
rect 7009 6239 7067 6245
rect 7009 6236 7021 6239
rect 6687 6208 7021 6236
rect 6687 6205 6699 6208
rect 6641 6199 6699 6205
rect 7009 6205 7021 6208
rect 7055 6236 7067 6239
rect 8294 6236 8300 6248
rect 7055 6208 8300 6236
rect 7055 6205 7067 6208
rect 7009 6199 7067 6205
rect 8294 6196 8300 6208
rect 8352 6196 8358 6248
rect 8478 6236 8484 6248
rect 8439 6208 8484 6236
rect 8478 6196 8484 6208
rect 8536 6196 8542 6248
rect 9766 6236 9772 6248
rect 9727 6208 9772 6236
rect 9766 6196 9772 6208
rect 9824 6196 9830 6248
rect 8802 6171 8860 6177
rect 8802 6168 8814 6171
rect 8312 6140 8814 6168
rect 8312 6112 8340 6140
rect 8802 6137 8814 6140
rect 8848 6137 8860 6171
rect 8802 6131 8860 6137
rect 4614 6100 4620 6112
rect 4575 6072 4620 6100
rect 4614 6060 4620 6072
rect 4672 6060 4678 6112
rect 8021 6103 8079 6109
rect 8021 6069 8033 6103
rect 8067 6100 8079 6103
rect 8294 6100 8300 6112
rect 8067 6072 8300 6100
rect 8067 6069 8079 6072
rect 8021 6063 8079 6069
rect 8294 6060 8300 6072
rect 8352 6060 8358 6112
rect 10060 6100 10088 6267
rect 10778 6264 10784 6276
rect 10836 6264 10842 6316
rect 13446 6304 13452 6316
rect 13407 6276 13452 6304
rect 13446 6264 13452 6276
rect 13504 6264 13510 6316
rect 14093 6307 14151 6313
rect 14093 6273 14105 6307
rect 14139 6304 14151 6307
rect 14642 6304 14648 6316
rect 14139 6276 14648 6304
rect 14139 6273 14151 6276
rect 14093 6267 14151 6273
rect 14642 6264 14648 6276
rect 14700 6304 14706 6316
rect 15289 6307 15347 6313
rect 15289 6304 15301 6307
rect 14700 6276 15301 6304
rect 14700 6264 14706 6276
rect 15289 6273 15301 6276
rect 15335 6273 15347 6307
rect 15289 6267 15347 6273
rect 10413 6171 10471 6177
rect 10413 6137 10425 6171
rect 10459 6137 10471 6171
rect 10413 6131 10471 6137
rect 10428 6100 10456 6131
rect 13170 6128 13176 6180
rect 13228 6168 13234 6180
rect 13541 6171 13599 6177
rect 13541 6168 13553 6171
rect 13228 6140 13553 6168
rect 13228 6128 13234 6140
rect 13541 6137 13553 6140
rect 13587 6168 13599 6171
rect 14734 6168 14740 6180
rect 13587 6140 14740 6168
rect 13587 6137 13599 6140
rect 13541 6131 13599 6137
rect 14734 6128 14740 6140
rect 14792 6128 14798 6180
rect 15010 6168 15016 6180
rect 14971 6140 15016 6168
rect 15010 6128 15016 6140
rect 15068 6128 15074 6180
rect 15102 6128 15108 6180
rect 15160 6168 15166 6180
rect 15160 6140 15205 6168
rect 15160 6128 15166 6140
rect 10060 6072 10456 6100
rect 14829 6103 14887 6109
rect 14829 6069 14841 6103
rect 14875 6100 14887 6103
rect 15120 6100 15148 6128
rect 14875 6072 15148 6100
rect 14875 6069 14887 6072
rect 14829 6063 14887 6069
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 6181 5899 6239 5905
rect 6181 5865 6193 5899
rect 6227 5896 6239 5899
rect 7006 5896 7012 5908
rect 6227 5868 7012 5896
rect 6227 5865 6239 5868
rect 6181 5859 6239 5865
rect 7006 5856 7012 5868
rect 7064 5856 7070 5908
rect 8478 5856 8484 5908
rect 8536 5896 8542 5908
rect 8849 5899 8907 5905
rect 8849 5896 8861 5899
rect 8536 5868 8861 5896
rect 8536 5856 8542 5868
rect 8849 5865 8861 5868
rect 8895 5865 8907 5899
rect 13722 5896 13728 5908
rect 13683 5868 13728 5896
rect 8849 5859 8907 5865
rect 13722 5856 13728 5868
rect 13780 5856 13786 5908
rect 9858 5828 9864 5840
rect 9819 5800 9864 5828
rect 9858 5788 9864 5800
rect 9916 5788 9922 5840
rect 10226 5788 10232 5840
rect 10284 5828 10290 5840
rect 11241 5831 11299 5837
rect 11241 5828 11253 5831
rect 10284 5800 11253 5828
rect 10284 5788 10290 5800
rect 11241 5797 11253 5800
rect 11287 5797 11299 5831
rect 11241 5791 11299 5797
rect 11974 5788 11980 5840
rect 12032 5828 12038 5840
rect 12574 5831 12632 5837
rect 12574 5828 12586 5831
rect 12032 5800 12586 5828
rect 12032 5788 12038 5800
rect 12574 5797 12586 5800
rect 12620 5828 12632 5831
rect 12986 5828 12992 5840
rect 12620 5800 12992 5828
rect 12620 5797 12632 5800
rect 12574 5791 12632 5797
rect 12986 5788 12992 5800
rect 13044 5788 13050 5840
rect 15102 5788 15108 5840
rect 15160 5828 15166 5840
rect 15289 5831 15347 5837
rect 15289 5828 15301 5831
rect 15160 5800 15301 5828
rect 15160 5788 15166 5800
rect 15289 5797 15301 5800
rect 15335 5797 15347 5831
rect 15289 5791 15347 5797
rect 5166 5720 5172 5772
rect 5224 5760 5230 5772
rect 5994 5760 6000 5772
rect 5224 5732 6000 5760
rect 5224 5720 5230 5732
rect 5994 5720 6000 5732
rect 6052 5720 6058 5772
rect 7466 5760 7472 5772
rect 7427 5732 7472 5760
rect 7466 5720 7472 5732
rect 7524 5720 7530 5772
rect 7926 5760 7932 5772
rect 7887 5732 7932 5760
rect 7926 5720 7932 5732
rect 7984 5720 7990 5772
rect 8018 5720 8024 5772
rect 8076 5760 8082 5772
rect 8481 5763 8539 5769
rect 8481 5760 8493 5763
rect 8076 5732 8493 5760
rect 8076 5720 8082 5732
rect 8481 5729 8493 5732
rect 8527 5729 8539 5763
rect 12250 5760 12256 5772
rect 12211 5732 12256 5760
rect 8481 5723 8539 5729
rect 12250 5720 12256 5732
rect 12308 5720 12314 5772
rect 14068 5763 14126 5769
rect 14068 5729 14080 5763
rect 14114 5760 14126 5763
rect 14642 5760 14648 5772
rect 14114 5732 14648 5760
rect 14114 5729 14126 5732
rect 14068 5723 14126 5729
rect 14642 5720 14648 5732
rect 14700 5720 14706 5772
rect 14734 5720 14740 5772
rect 14792 5760 14798 5772
rect 15381 5763 15439 5769
rect 15381 5760 15393 5763
rect 14792 5732 15393 5760
rect 14792 5720 14798 5732
rect 15381 5729 15393 5732
rect 15427 5760 15439 5763
rect 16022 5760 16028 5772
rect 15427 5732 16028 5760
rect 15427 5729 15439 5732
rect 15381 5723 15439 5729
rect 16022 5720 16028 5732
rect 16080 5720 16086 5772
rect 8202 5692 8208 5704
rect 8163 5664 8208 5692
rect 8202 5652 8208 5664
rect 8260 5652 8266 5704
rect 9398 5652 9404 5704
rect 9456 5692 9462 5704
rect 9769 5695 9827 5701
rect 9769 5692 9781 5695
rect 9456 5664 9781 5692
rect 9456 5652 9462 5664
rect 9769 5661 9781 5664
rect 9815 5661 9827 5695
rect 9769 5655 9827 5661
rect 10413 5695 10471 5701
rect 10413 5661 10425 5695
rect 10459 5692 10471 5695
rect 10502 5692 10508 5704
rect 10459 5664 10508 5692
rect 10459 5661 10471 5664
rect 10413 5655 10471 5661
rect 10502 5652 10508 5664
rect 10560 5652 10566 5704
rect 12526 5652 12532 5704
rect 12584 5692 12590 5704
rect 14921 5695 14979 5701
rect 14921 5692 14933 5695
rect 12584 5664 14933 5692
rect 12584 5652 12590 5664
rect 14921 5661 14933 5664
rect 14967 5692 14979 5695
rect 15010 5692 15016 5704
rect 14967 5664 15016 5692
rect 14967 5661 14979 5664
rect 14921 5655 14979 5661
rect 15010 5652 15016 5664
rect 15068 5652 15074 5704
rect 13722 5584 13728 5636
rect 13780 5624 13786 5636
rect 15470 5624 15476 5636
rect 13780 5596 15476 5624
rect 13780 5584 13786 5596
rect 15470 5584 15476 5596
rect 15528 5584 15534 5636
rect 10778 5556 10784 5568
rect 10739 5528 10784 5556
rect 10778 5516 10784 5528
rect 10836 5516 10842 5568
rect 13170 5556 13176 5568
rect 13131 5528 13176 5556
rect 13170 5516 13176 5528
rect 13228 5516 13234 5568
rect 14139 5559 14197 5565
rect 14139 5525 14151 5559
rect 14185 5556 14197 5559
rect 14366 5556 14372 5568
rect 14185 5528 14372 5556
rect 14185 5525 14197 5528
rect 14139 5519 14197 5525
rect 14366 5516 14372 5528
rect 14424 5516 14430 5568
rect 14550 5556 14556 5568
rect 14511 5528 14556 5556
rect 14550 5516 14556 5528
rect 14608 5516 14614 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 5994 5352 6000 5364
rect 5955 5324 6000 5352
rect 5994 5312 6000 5324
rect 6052 5312 6058 5364
rect 6546 5312 6552 5364
rect 6604 5352 6610 5364
rect 7285 5355 7343 5361
rect 7285 5352 7297 5355
rect 6604 5324 7297 5352
rect 6604 5312 6610 5324
rect 7285 5321 7297 5324
rect 7331 5321 7343 5355
rect 7285 5315 7343 5321
rect 9677 5355 9735 5361
rect 9677 5321 9689 5355
rect 9723 5352 9735 5355
rect 9858 5352 9864 5364
rect 9723 5324 9864 5352
rect 9723 5321 9735 5324
rect 9677 5315 9735 5321
rect 9858 5312 9864 5324
rect 9916 5312 9922 5364
rect 11146 5352 11152 5364
rect 11107 5324 11152 5352
rect 11146 5312 11152 5324
rect 11204 5312 11210 5364
rect 12250 5352 12256 5364
rect 12211 5324 12256 5352
rect 12250 5312 12256 5324
rect 12308 5312 12314 5364
rect 12986 5352 12992 5364
rect 12947 5324 12992 5352
rect 12986 5312 12992 5324
rect 13044 5312 13050 5364
rect 13170 5312 13176 5364
rect 13228 5352 13234 5364
rect 13449 5355 13507 5361
rect 13449 5352 13461 5355
rect 13228 5324 13461 5352
rect 13228 5312 13234 5324
rect 13449 5321 13461 5324
rect 13495 5352 13507 5355
rect 13814 5352 13820 5364
rect 13495 5324 13820 5352
rect 13495 5321 13507 5324
rect 13449 5315 13507 5321
rect 13814 5312 13820 5324
rect 13872 5312 13878 5364
rect 13906 5312 13912 5364
rect 13964 5352 13970 5364
rect 22235 5355 22293 5361
rect 22235 5352 22247 5355
rect 13964 5324 22247 5352
rect 13964 5312 13970 5324
rect 22235 5321 22247 5324
rect 22281 5321 22293 5355
rect 22235 5315 22293 5321
rect 12710 5244 12716 5296
rect 12768 5284 12774 5296
rect 13998 5284 14004 5296
rect 12768 5256 14004 5284
rect 12768 5244 12774 5256
rect 13998 5244 14004 5256
rect 14056 5284 14062 5296
rect 14277 5287 14335 5293
rect 14277 5284 14289 5287
rect 14056 5256 14289 5284
rect 14056 5244 14062 5256
rect 14277 5253 14289 5256
rect 14323 5253 14335 5287
rect 14642 5284 14648 5296
rect 14603 5256 14648 5284
rect 14277 5247 14335 5253
rect 14642 5244 14648 5256
rect 14700 5244 14706 5296
rect 15470 5284 15476 5296
rect 15431 5256 15476 5284
rect 15470 5244 15476 5256
rect 15528 5244 15534 5296
rect 16022 5284 16028 5296
rect 15983 5256 16028 5284
rect 16022 5244 16028 5256
rect 16080 5244 16086 5296
rect 8202 5176 8208 5228
rect 8260 5216 8266 5228
rect 8389 5219 8447 5225
rect 8389 5216 8401 5219
rect 8260 5188 8401 5216
rect 8260 5176 8266 5188
rect 8389 5185 8401 5188
rect 8435 5185 8447 5219
rect 10226 5216 10232 5228
rect 10187 5188 10232 5216
rect 8389 5179 8447 5185
rect 10226 5176 10232 5188
rect 10284 5176 10290 5228
rect 10502 5216 10508 5228
rect 10463 5188 10508 5216
rect 10502 5176 10508 5188
rect 10560 5176 10566 5228
rect 12526 5216 12532 5228
rect 12487 5188 12532 5216
rect 12526 5176 12532 5188
rect 12584 5176 12590 5228
rect 7101 5151 7159 5157
rect 7101 5117 7113 5151
rect 7147 5148 7159 5151
rect 15264 5151 15322 5157
rect 7147 5120 7696 5148
rect 7147 5117 7159 5120
rect 7101 5111 7159 5117
rect 7668 5024 7696 5120
rect 15264 5117 15276 5151
rect 15310 5117 15322 5151
rect 15264 5111 15322 5117
rect 22164 5151 22222 5157
rect 22164 5117 22176 5151
rect 22210 5148 22222 5151
rect 22210 5120 22692 5148
rect 22210 5117 22222 5120
rect 22164 5111 22222 5117
rect 8710 5083 8768 5089
rect 8710 5049 8722 5083
rect 8756 5049 8768 5083
rect 8710 5043 8768 5049
rect 10045 5083 10103 5089
rect 10045 5049 10057 5083
rect 10091 5080 10103 5083
rect 10321 5083 10379 5089
rect 10321 5080 10333 5083
rect 10091 5052 10333 5080
rect 10091 5049 10103 5052
rect 10045 5043 10103 5049
rect 10321 5049 10333 5052
rect 10367 5080 10379 5083
rect 11238 5080 11244 5092
rect 10367 5052 11244 5080
rect 10367 5049 10379 5052
rect 10321 5043 10379 5049
rect 7650 5012 7656 5024
rect 7611 4984 7656 5012
rect 7650 4972 7656 4984
rect 7708 4972 7714 5024
rect 8294 5012 8300 5024
rect 8255 4984 8300 5012
rect 8294 4972 8300 4984
rect 8352 5012 8358 5024
rect 8725 5012 8753 5043
rect 11238 5040 11244 5052
rect 11296 5040 11302 5092
rect 13725 5083 13783 5089
rect 13725 5049 13737 5083
rect 13771 5049 13783 5083
rect 13725 5043 13783 5049
rect 9306 5012 9312 5024
rect 8352 4984 8753 5012
rect 9267 4984 9312 5012
rect 8352 4972 8358 4984
rect 9306 4972 9312 4984
rect 9364 4972 9370 5024
rect 13740 5012 13768 5043
rect 13814 5040 13820 5092
rect 13872 5080 13878 5092
rect 15279 5080 15307 5111
rect 15749 5083 15807 5089
rect 15749 5080 15761 5083
rect 13872 5052 13917 5080
rect 15279 5052 15761 5080
rect 13872 5040 13878 5052
rect 15749 5049 15761 5052
rect 15795 5080 15807 5083
rect 17494 5080 17500 5092
rect 15795 5052 17500 5080
rect 15795 5049 15807 5052
rect 15749 5043 15807 5049
rect 17494 5040 17500 5052
rect 17552 5040 17558 5092
rect 14550 5012 14556 5024
rect 13740 4984 14556 5012
rect 14550 4972 14556 4984
rect 14608 4972 14614 5024
rect 22664 5021 22692 5120
rect 22649 5015 22707 5021
rect 22649 4981 22661 5015
rect 22695 5012 22707 5015
rect 23750 5012 23756 5024
rect 22695 4984 23756 5012
rect 22695 4981 22707 4984
rect 22649 4975 22707 4981
rect 23750 4972 23756 4984
rect 23808 4972 23814 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 7466 4808 7472 4820
rect 7427 4780 7472 4808
rect 7466 4768 7472 4780
rect 7524 4768 7530 4820
rect 7926 4808 7932 4820
rect 7887 4780 7932 4808
rect 7926 4768 7932 4780
rect 7984 4768 7990 4820
rect 8202 4768 8208 4820
rect 8260 4808 8266 4820
rect 8389 4811 8447 4817
rect 8389 4808 8401 4811
rect 8260 4780 8401 4808
rect 8260 4768 8266 4780
rect 8389 4777 8401 4780
rect 8435 4777 8447 4811
rect 10134 4808 10140 4820
rect 10095 4780 10140 4808
rect 8389 4771 8447 4777
rect 10134 4768 10140 4780
rect 10192 4768 10198 4820
rect 23658 4768 23664 4820
rect 23716 4808 23722 4820
rect 23799 4811 23857 4817
rect 23799 4808 23811 4811
rect 23716 4780 23811 4808
rect 23716 4768 23722 4780
rect 23799 4777 23811 4780
rect 23845 4777 23857 4811
rect 23799 4771 23857 4777
rect 10686 4740 10692 4752
rect 10463 4712 10692 4740
rect 10463 4681 10491 4712
rect 10686 4700 10692 4712
rect 10744 4700 10750 4752
rect 13814 4700 13820 4752
rect 13872 4740 13878 4752
rect 13872 4712 13917 4740
rect 13872 4700 13878 4712
rect 10448 4675 10506 4681
rect 10448 4641 10460 4675
rect 10494 4641 10506 4675
rect 10448 4635 10506 4641
rect 10551 4675 10609 4681
rect 10551 4641 10563 4675
rect 10597 4672 10609 4675
rect 11422 4672 11428 4684
rect 10597 4644 11428 4672
rect 10597 4641 10609 4644
rect 10551 4635 10609 4641
rect 11422 4632 11428 4644
rect 11480 4632 11486 4684
rect 14366 4632 14372 4684
rect 14424 4672 14430 4684
rect 15286 4672 15292 4684
rect 14424 4644 15292 4672
rect 14424 4632 14430 4644
rect 15286 4632 15292 4644
rect 15344 4632 15350 4684
rect 23728 4675 23786 4681
rect 23728 4641 23740 4675
rect 23774 4672 23786 4675
rect 23934 4672 23940 4684
rect 23774 4644 23940 4672
rect 23774 4641 23786 4644
rect 23728 4635 23786 4641
rect 23934 4632 23940 4644
rect 23992 4632 23998 4684
rect 13722 4604 13728 4616
rect 13683 4576 13728 4604
rect 13722 4564 13728 4576
rect 13780 4564 13786 4616
rect 13998 4604 14004 4616
rect 13959 4576 14004 4604
rect 13998 4564 14004 4576
rect 14056 4564 14062 4616
rect 11609 4471 11667 4477
rect 11609 4437 11621 4471
rect 11655 4468 11667 4471
rect 12894 4468 12900 4480
rect 11655 4440 12900 4468
rect 11655 4437 11667 4440
rect 11609 4431 11667 4437
rect 12894 4428 12900 4440
rect 12952 4428 12958 4480
rect 14826 4428 14832 4480
rect 14884 4468 14890 4480
rect 15473 4471 15531 4477
rect 15473 4468 15485 4471
rect 14884 4440 15485 4468
rect 14884 4428 14890 4440
rect 15473 4437 15485 4440
rect 15519 4437 15531 4471
rect 15473 4431 15531 4437
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 7558 4264 7564 4276
rect 7519 4236 7564 4264
rect 7558 4224 7564 4236
rect 7616 4264 7622 4276
rect 7616 4236 8156 4264
rect 7616 4224 7622 4236
rect 8128 4137 8156 4236
rect 10686 4224 10692 4276
rect 10744 4264 10750 4276
rect 10873 4267 10931 4273
rect 10873 4264 10885 4267
rect 10744 4236 10885 4264
rect 10744 4224 10750 4236
rect 10873 4233 10885 4236
rect 10919 4233 10931 4267
rect 11422 4264 11428 4276
rect 11383 4236 11428 4264
rect 10873 4227 10931 4233
rect 11422 4224 11428 4236
rect 11480 4224 11486 4276
rect 13170 4264 13176 4276
rect 13131 4236 13176 4264
rect 13170 4224 13176 4236
rect 13228 4224 13234 4276
rect 15286 4264 15292 4276
rect 15247 4236 15292 4264
rect 15286 4224 15292 4236
rect 15344 4224 15350 4276
rect 8113 4131 8171 4137
rect 8113 4097 8125 4131
rect 8159 4097 8171 4131
rect 8113 4091 8171 4097
rect 9953 4063 10011 4069
rect 9953 4029 9965 4063
rect 9999 4029 10011 4063
rect 9953 4023 10011 4029
rect 8294 3992 8300 4004
rect 7944 3964 8300 3992
rect 2498 3884 2504 3936
rect 2556 3924 2562 3936
rect 7944 3933 7972 3964
rect 8294 3952 8300 3964
rect 8352 3992 8358 4004
rect 8434 3995 8492 4001
rect 8434 3992 8446 3995
rect 8352 3964 8446 3992
rect 8352 3952 8358 3964
rect 8434 3961 8446 3964
rect 8480 3961 8492 3995
rect 9858 3992 9864 4004
rect 9819 3964 9864 3992
rect 8434 3955 8492 3961
rect 9858 3952 9864 3964
rect 9916 3952 9922 4004
rect 9968 3936 9996 4023
rect 13170 4020 13176 4072
rect 13228 4060 13234 4072
rect 13449 4063 13507 4069
rect 13449 4060 13461 4063
rect 13228 4032 13461 4060
rect 13228 4020 13234 4032
rect 13449 4029 13461 4032
rect 13495 4029 13507 4063
rect 13449 4023 13507 4029
rect 24648 4063 24706 4069
rect 24648 4029 24660 4063
rect 24694 4060 24706 4063
rect 24694 4032 25176 4060
rect 24694 4029 24706 4032
rect 24648 4023 24706 4029
rect 13814 3952 13820 4004
rect 13872 3992 13878 4004
rect 14093 3995 14151 4001
rect 14093 3992 14105 3995
rect 13872 3964 14105 3992
rect 13872 3952 13878 3964
rect 14093 3961 14105 3964
rect 14139 3992 14151 3995
rect 14369 3995 14427 4001
rect 14369 3992 14381 3995
rect 14139 3964 14381 3992
rect 14139 3961 14151 3964
rect 14093 3955 14151 3961
rect 14369 3961 14381 3964
rect 14415 3961 14427 3995
rect 14369 3955 14427 3961
rect 7929 3927 7987 3933
rect 7929 3924 7941 3927
rect 2556 3896 7941 3924
rect 2556 3884 2562 3896
rect 7929 3893 7941 3896
rect 7975 3893 7987 3927
rect 9030 3924 9036 3936
rect 8991 3896 9036 3924
rect 7929 3887 7987 3893
rect 9030 3884 9036 3896
rect 9088 3884 9094 3936
rect 9306 3884 9312 3936
rect 9364 3924 9370 3936
rect 9769 3927 9827 3933
rect 9769 3924 9781 3927
rect 9364 3896 9781 3924
rect 9364 3884 9370 3896
rect 9769 3893 9781 3896
rect 9815 3924 9827 3927
rect 9950 3924 9956 3936
rect 9815 3896 9956 3924
rect 9815 3893 9827 3896
rect 9769 3887 9827 3893
rect 9950 3884 9956 3896
rect 10008 3884 10014 3936
rect 23934 3924 23940 3936
rect 23895 3896 23940 3924
rect 23934 3884 23940 3896
rect 23992 3884 23998 3936
rect 24026 3884 24032 3936
rect 24084 3924 24090 3936
rect 25148 3933 25176 4032
rect 24719 3927 24777 3933
rect 24719 3924 24731 3927
rect 24084 3896 24731 3924
rect 24084 3884 24090 3896
rect 24719 3893 24731 3896
rect 24765 3893 24777 3927
rect 24719 3887 24777 3893
rect 25133 3927 25191 3933
rect 25133 3893 25145 3927
rect 25179 3924 25191 3927
rect 27614 3924 27620 3936
rect 25179 3896 27620 3924
rect 25179 3893 25191 3896
rect 25133 3887 25191 3893
rect 27614 3884 27620 3896
rect 27672 3884 27678 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 13722 3720 13728 3732
rect 13683 3692 13728 3720
rect 13722 3680 13728 3692
rect 13780 3680 13786 3732
rect 9858 3612 9864 3664
rect 9916 3652 9922 3664
rect 9953 3655 10011 3661
rect 9953 3652 9965 3655
rect 9916 3624 9965 3652
rect 9916 3612 9922 3624
rect 9953 3621 9965 3624
rect 9999 3621 10011 3655
rect 9953 3615 10011 3621
rect 8665 3587 8723 3593
rect 8665 3553 8677 3587
rect 8711 3584 8723 3587
rect 9030 3584 9036 3596
rect 8711 3556 9036 3584
rect 8711 3553 8723 3556
rect 8665 3547 8723 3553
rect 9030 3544 9036 3556
rect 9088 3544 9094 3596
rect 8018 3516 8024 3528
rect 7979 3488 8024 3516
rect 8018 3476 8024 3488
rect 8076 3476 8082 3528
rect 9214 3476 9220 3528
rect 9272 3516 9278 3528
rect 9861 3519 9919 3525
rect 9861 3516 9873 3519
rect 9272 3488 9873 3516
rect 9272 3476 9278 3488
rect 9861 3485 9873 3488
rect 9907 3516 9919 3519
rect 11333 3519 11391 3525
rect 11333 3516 11345 3519
rect 9907 3488 11345 3516
rect 9907 3485 9919 3488
rect 9861 3479 9919 3485
rect 11333 3485 11345 3488
rect 11379 3485 11391 3519
rect 11333 3479 11391 3485
rect 10410 3448 10416 3460
rect 10371 3420 10416 3448
rect 10410 3408 10416 3420
rect 10468 3408 10474 3460
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 8018 3176 8024 3188
rect 7979 3148 8024 3176
rect 8018 3136 8024 3148
rect 8076 3136 8082 3188
rect 9214 3176 9220 3188
rect 9175 3148 9220 3176
rect 9214 3136 9220 3148
rect 9272 3136 9278 3188
rect 9585 3179 9643 3185
rect 9585 3145 9597 3179
rect 9631 3176 9643 3179
rect 9858 3176 9864 3188
rect 9631 3148 9864 3176
rect 9631 3145 9643 3148
rect 9585 3139 9643 3145
rect 9858 3136 9864 3148
rect 9916 3136 9922 3188
rect 9950 3068 9956 3120
rect 10008 3108 10014 3120
rect 10689 3111 10747 3117
rect 10689 3108 10701 3111
rect 10008 3080 10701 3108
rect 10008 3068 10014 3080
rect 10689 3077 10701 3080
rect 10735 3077 10747 3111
rect 10689 3071 10747 3077
rect 7653 3043 7711 3049
rect 7653 3009 7665 3043
rect 7699 3040 7711 3043
rect 9030 3040 9036 3052
rect 7699 3012 9036 3040
rect 7699 3009 7711 3012
rect 7653 3003 7711 3009
rect 9030 3000 9036 3012
rect 9088 3000 9094 3052
rect 10410 3040 10416 3052
rect 10371 3012 10416 3040
rect 10410 3000 10416 3012
rect 10468 3000 10474 3052
rect 10428 2972 10456 3000
rect 11276 2975 11334 2981
rect 11276 2972 11288 2975
rect 10428 2944 11288 2972
rect 11276 2941 11288 2944
rect 11322 2972 11334 2975
rect 11701 2975 11759 2981
rect 11701 2972 11713 2975
rect 11322 2944 11713 2972
rect 11322 2941 11334 2944
rect 11276 2935 11334 2941
rect 11701 2941 11713 2944
rect 11747 2941 11759 2975
rect 11701 2935 11759 2941
rect 7285 2907 7343 2913
rect 7285 2873 7297 2907
rect 7331 2904 7343 2907
rect 8202 2904 8208 2916
rect 7331 2876 8208 2904
rect 7331 2873 7343 2876
rect 7285 2867 7343 2873
rect 8202 2864 8208 2876
rect 8260 2864 8266 2916
rect 8297 2907 8355 2913
rect 8297 2873 8309 2907
rect 8343 2873 8355 2907
rect 8297 2867 8355 2873
rect 8849 2907 8907 2913
rect 8849 2873 8861 2907
rect 8895 2904 8907 2907
rect 9769 2907 9827 2913
rect 9769 2904 9781 2907
rect 8895 2876 9781 2904
rect 8895 2873 8907 2876
rect 8849 2867 8907 2873
rect 9769 2873 9781 2876
rect 9815 2873 9827 2907
rect 9769 2867 9827 2873
rect 9861 2907 9919 2913
rect 9861 2873 9873 2907
rect 9907 2904 9919 2907
rect 9950 2904 9956 2916
rect 9907 2876 9956 2904
rect 9907 2873 9919 2876
rect 9861 2867 9919 2873
rect 8018 2796 8024 2848
rect 8076 2836 8082 2848
rect 8312 2836 8340 2867
rect 8076 2808 8340 2836
rect 9784 2836 9812 2867
rect 9950 2864 9956 2876
rect 10008 2864 10014 2916
rect 11057 2907 11115 2913
rect 11057 2904 11069 2907
rect 10152 2876 11069 2904
rect 10152 2848 10180 2876
rect 11057 2873 11069 2876
rect 11103 2873 11115 2907
rect 11057 2867 11115 2873
rect 11379 2907 11437 2913
rect 11379 2873 11391 2907
rect 11425 2904 11437 2907
rect 18782 2904 18788 2916
rect 11425 2876 18788 2904
rect 11425 2873 11437 2876
rect 11379 2867 11437 2873
rect 18782 2864 18788 2876
rect 18840 2864 18846 2916
rect 10134 2836 10140 2848
rect 9784 2808 10140 2836
rect 8076 2796 8082 2808
rect 10134 2796 10140 2808
rect 10192 2796 10198 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 5675 2635 5733 2641
rect 5675 2601 5687 2635
rect 5721 2632 5733 2635
rect 6086 2632 6092 2644
rect 5721 2604 6092 2632
rect 5721 2601 5733 2604
rect 5675 2595 5733 2601
rect 6086 2592 6092 2604
rect 6144 2592 6150 2644
rect 7055 2635 7113 2641
rect 7055 2601 7067 2635
rect 7101 2632 7113 2635
rect 7282 2632 7288 2644
rect 7101 2604 7288 2632
rect 7101 2601 7113 2604
rect 7055 2595 7113 2601
rect 7282 2592 7288 2604
rect 7340 2592 7346 2644
rect 8067 2635 8125 2641
rect 8067 2601 8079 2635
rect 8113 2632 8125 2635
rect 8202 2632 8208 2644
rect 8113 2604 8208 2632
rect 8113 2601 8125 2604
rect 8067 2595 8125 2601
rect 8202 2592 8208 2604
rect 8260 2592 8266 2644
rect 11514 2592 11520 2644
rect 11572 2632 11578 2644
rect 11609 2635 11667 2641
rect 11609 2632 11621 2635
rect 11572 2604 11621 2632
rect 11572 2592 11578 2604
rect 11609 2601 11621 2604
rect 11655 2601 11667 2635
rect 11609 2595 11667 2601
rect 13035 2635 13093 2641
rect 13035 2601 13047 2635
rect 13081 2632 13093 2635
rect 13538 2632 13544 2644
rect 13081 2604 13544 2632
rect 13081 2601 13093 2604
rect 13035 2595 13093 2601
rect 13538 2592 13544 2604
rect 13596 2592 13602 2644
rect 23934 2592 23940 2644
rect 23992 2632 23998 2644
rect 25222 2632 25228 2644
rect 23992 2604 25228 2632
rect 23992 2592 23998 2604
rect 25222 2592 25228 2604
rect 25280 2592 25286 2644
rect 9030 2524 9036 2576
rect 9088 2564 9094 2576
rect 9585 2567 9643 2573
rect 9585 2564 9597 2567
rect 9088 2536 9597 2564
rect 9088 2524 9094 2536
rect 9585 2533 9597 2536
rect 9631 2564 9643 2567
rect 9953 2567 10011 2573
rect 9953 2564 9965 2567
rect 9631 2536 9965 2564
rect 9631 2533 9643 2536
rect 9585 2527 9643 2533
rect 9953 2533 9965 2536
rect 9999 2533 10011 2567
rect 9953 2527 10011 2533
rect 19242 2524 19248 2576
rect 19300 2564 19306 2576
rect 20533 2567 20591 2573
rect 20533 2564 20545 2567
rect 19300 2536 20545 2564
rect 19300 2524 19306 2536
rect 5572 2499 5630 2505
rect 5572 2496 5584 2499
rect 5552 2465 5584 2496
rect 5618 2465 5630 2499
rect 5552 2459 5630 2465
rect 6984 2499 7042 2505
rect 6984 2465 6996 2499
rect 7030 2496 7042 2499
rect 7190 2496 7196 2508
rect 7030 2468 7196 2496
rect 7030 2465 7042 2468
rect 6984 2459 7042 2465
rect 5552 2304 5580 2459
rect 7190 2456 7196 2468
rect 7248 2496 7254 2508
rect 7377 2499 7435 2505
rect 7377 2496 7389 2499
rect 7248 2468 7389 2496
rect 7248 2456 7254 2468
rect 7377 2465 7389 2468
rect 7423 2465 7435 2499
rect 7377 2459 7435 2465
rect 7996 2499 8054 2505
rect 7996 2465 8008 2499
rect 8042 2496 8054 2499
rect 11400 2499 11458 2505
rect 8042 2468 8524 2496
rect 8042 2465 8054 2468
rect 7996 2459 8054 2465
rect 5534 2252 5540 2304
rect 5592 2292 5598 2304
rect 8496 2301 8524 2468
rect 11400 2465 11412 2499
rect 11446 2496 11458 2499
rect 11790 2496 11796 2508
rect 11446 2468 11796 2496
rect 11446 2465 11458 2468
rect 11400 2459 11458 2465
rect 11790 2456 11796 2468
rect 11848 2456 11854 2508
rect 12932 2499 12990 2505
rect 12932 2465 12944 2499
rect 12978 2465 12990 2499
rect 18782 2496 18788 2508
rect 18743 2468 18788 2496
rect 12932 2459 12990 2465
rect 9217 2431 9275 2437
rect 9217 2397 9229 2431
rect 9263 2428 9275 2431
rect 9858 2428 9864 2440
rect 9263 2400 9864 2428
rect 9263 2397 9275 2400
rect 9217 2391 9275 2397
rect 9858 2388 9864 2400
rect 9916 2388 9922 2440
rect 10134 2428 10140 2440
rect 10095 2400 10140 2428
rect 10134 2388 10140 2400
rect 10192 2388 10198 2440
rect 10318 2388 10324 2440
rect 10376 2428 10382 2440
rect 12947 2428 12975 2459
rect 18782 2456 18788 2468
rect 18840 2496 18846 2508
rect 19996 2505 20024 2536
rect 20533 2533 20545 2536
rect 20579 2533 20591 2567
rect 20533 2527 20591 2533
rect 19337 2499 19395 2505
rect 19337 2496 19349 2499
rect 18840 2468 19349 2496
rect 18840 2456 18846 2468
rect 19337 2465 19349 2468
rect 19383 2465 19395 2499
rect 19337 2459 19395 2465
rect 19981 2499 20039 2505
rect 19981 2465 19993 2499
rect 20027 2465 20039 2499
rect 19981 2459 20039 2465
rect 24648 2499 24706 2505
rect 24648 2465 24660 2499
rect 24694 2496 24706 2499
rect 24694 2468 25176 2496
rect 24694 2465 24706 2468
rect 24648 2459 24706 2465
rect 13357 2431 13415 2437
rect 13357 2428 13369 2431
rect 10376 2400 13369 2428
rect 10376 2388 10382 2400
rect 13357 2397 13369 2400
rect 13403 2397 13415 2431
rect 13357 2391 13415 2397
rect 20165 2363 20223 2369
rect 20165 2329 20177 2363
rect 20211 2360 20223 2363
rect 22554 2360 22560 2372
rect 20211 2332 22560 2360
rect 20211 2329 20223 2332
rect 20165 2323 20223 2329
rect 22554 2320 22560 2332
rect 22612 2320 22618 2372
rect 5997 2295 6055 2301
rect 5997 2292 6009 2295
rect 5592 2264 6009 2292
rect 5592 2252 5598 2264
rect 5997 2261 6009 2264
rect 6043 2261 6055 2295
rect 5997 2255 6055 2261
rect 8481 2295 8539 2301
rect 8481 2261 8493 2295
rect 8527 2292 8539 2295
rect 8570 2292 8576 2304
rect 8527 2264 8576 2292
rect 8527 2261 8539 2264
rect 8481 2255 8539 2261
rect 8570 2252 8576 2264
rect 8628 2252 8634 2304
rect 11790 2292 11796 2304
rect 11751 2264 11796 2292
rect 11790 2252 11796 2264
rect 11848 2252 11854 2304
rect 18969 2295 19027 2301
rect 18969 2261 18981 2295
rect 19015 2292 19027 2295
rect 20622 2292 20628 2304
rect 19015 2264 20628 2292
rect 19015 2261 19027 2264
rect 18969 2255 19027 2261
rect 20622 2252 20628 2264
rect 20680 2252 20686 2304
rect 20714 2252 20720 2304
rect 20772 2292 20778 2304
rect 25148 2301 25176 2468
rect 24719 2295 24777 2301
rect 24719 2292 24731 2295
rect 20772 2264 24731 2292
rect 20772 2252 20778 2264
rect 24719 2261 24731 2264
rect 24765 2261 24777 2295
rect 24719 2255 24777 2261
rect 25133 2295 25191 2301
rect 25133 2261 25145 2295
rect 25179 2292 25191 2295
rect 26878 2292 26884 2304
rect 25179 2264 26884 2292
rect 25179 2261 25191 2264
rect 25133 2255 25191 2261
rect 26878 2252 26884 2264
rect 26936 2252 26942 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
<< via1 >>
rect 20 27072 72 27124
rect 756 27072 808 27124
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 6276 24259 6328 24268
rect 6276 24225 6294 24259
rect 6294 24225 6328 24259
rect 6276 24216 6328 24225
rect 7012 24216 7064 24268
rect 8208 24216 8260 24268
rect 11612 24216 11664 24268
rect 23940 24284 23992 24336
rect 25412 24284 25464 24336
rect 25136 24216 25188 24268
rect 22192 24080 22244 24132
rect 6736 24012 6788 24064
rect 6828 24012 6880 24064
rect 10232 24055 10284 24064
rect 10232 24021 10241 24055
rect 10241 24021 10275 24055
rect 10275 24021 10284 24055
rect 10232 24012 10284 24021
rect 11336 24012 11388 24064
rect 20628 24012 20680 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 2504 23851 2556 23860
rect 2504 23817 2513 23851
rect 2513 23817 2547 23851
rect 2547 23817 2556 23851
rect 2504 23808 2556 23817
rect 6276 23851 6328 23860
rect 6276 23817 6285 23851
rect 6285 23817 6319 23851
rect 6319 23817 6328 23851
rect 6276 23808 6328 23817
rect 7748 23740 7800 23792
rect 2504 23604 2556 23656
rect 8944 23808 8996 23860
rect 11612 23851 11664 23860
rect 11612 23817 11621 23851
rect 11621 23817 11655 23851
rect 11655 23817 11664 23851
rect 11612 23808 11664 23817
rect 8208 23715 8260 23724
rect 8208 23681 8217 23715
rect 8217 23681 8251 23715
rect 8251 23681 8260 23715
rect 8208 23672 8260 23681
rect 10232 23715 10284 23724
rect 10232 23681 10241 23715
rect 10241 23681 10275 23715
rect 10275 23681 10284 23715
rect 10232 23672 10284 23681
rect 15476 23808 15528 23860
rect 18788 23808 18840 23860
rect 23756 23808 23808 23860
rect 23940 23851 23992 23860
rect 23940 23817 23949 23851
rect 23949 23817 23983 23851
rect 23983 23817 23992 23851
rect 23940 23808 23992 23817
rect 25136 23851 25188 23860
rect 25136 23817 25145 23851
rect 25145 23817 25179 23851
rect 25179 23817 25188 23851
rect 25136 23808 25188 23817
rect 27068 23808 27120 23860
rect 6000 23536 6052 23588
rect 6644 23468 6696 23520
rect 9956 23468 10008 23520
rect 11612 23536 11664 23588
rect 13728 23468 13780 23520
rect 15752 23468 15804 23520
rect 19984 23468 20036 23520
rect 23940 23468 23992 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 1584 23307 1636 23316
rect 1584 23273 1593 23307
rect 1593 23273 1627 23307
rect 1627 23273 1636 23307
rect 1584 23264 1636 23273
rect 3976 23264 4028 23316
rect 6920 23239 6972 23248
rect 6920 23205 6929 23239
rect 6929 23205 6963 23239
rect 6963 23205 6972 23239
rect 6920 23196 6972 23205
rect 9772 23196 9824 23248
rect 11428 23239 11480 23248
rect 11428 23205 11437 23239
rect 11437 23205 11471 23239
rect 11471 23205 11480 23239
rect 11428 23196 11480 23205
rect 1400 23171 1452 23180
rect 1400 23137 1409 23171
rect 1409 23137 1443 23171
rect 1443 23137 1452 23171
rect 1400 23128 1452 23137
rect 2504 23128 2556 23180
rect 6552 23060 6604 23112
rect 6828 23103 6880 23112
rect 6828 23069 6837 23103
rect 6837 23069 6871 23103
rect 6871 23069 6880 23103
rect 6828 23060 6880 23069
rect 10140 23060 10192 23112
rect 10232 23103 10284 23112
rect 10232 23069 10241 23103
rect 10241 23069 10275 23103
rect 10275 23069 10284 23103
rect 11336 23103 11388 23112
rect 10232 23060 10284 23069
rect 11336 23069 11345 23103
rect 11345 23069 11379 23103
rect 11379 23069 11388 23103
rect 11336 23060 11388 23069
rect 11612 23103 11664 23112
rect 11612 23069 11621 23103
rect 11621 23069 11655 23103
rect 11655 23069 11664 23103
rect 11612 23060 11664 23069
rect 7380 23035 7432 23044
rect 7380 23001 7389 23035
rect 7389 23001 7423 23035
rect 7423 23001 7432 23035
rect 7380 22992 7432 23001
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 6552 22720 6604 22772
rect 6920 22720 6972 22772
rect 11336 22720 11388 22772
rect 6736 22584 6788 22636
rect 7380 22627 7432 22636
rect 7380 22593 7389 22627
rect 7389 22593 7423 22627
rect 7423 22593 7432 22627
rect 7380 22584 7432 22593
rect 7748 22584 7800 22636
rect 8852 22627 8904 22636
rect 8852 22593 8861 22627
rect 8861 22593 8895 22627
rect 8895 22593 8904 22627
rect 8852 22584 8904 22593
rect 9496 22627 9548 22636
rect 9496 22593 9505 22627
rect 9505 22593 9539 22627
rect 9539 22593 9548 22627
rect 9496 22584 9548 22593
rect 10232 22584 10284 22636
rect 11428 22584 11480 22636
rect 2780 22516 2832 22568
rect 9956 22516 10008 22568
rect 10784 22559 10836 22568
rect 10784 22525 10793 22559
rect 10793 22525 10827 22559
rect 10827 22525 10836 22559
rect 10784 22516 10836 22525
rect 15844 22516 15896 22568
rect 1400 22448 1452 22500
rect 3332 22448 3384 22500
rect 2504 22423 2556 22432
rect 2504 22389 2513 22423
rect 2513 22389 2547 22423
rect 2547 22389 2556 22423
rect 2504 22380 2556 22389
rect 2780 22423 2832 22432
rect 2780 22389 2789 22423
rect 2789 22389 2823 22423
rect 2823 22389 2832 22423
rect 2780 22380 2832 22389
rect 3240 22423 3292 22432
rect 3240 22389 3249 22423
rect 3249 22389 3283 22423
rect 3283 22389 3292 22423
rect 3240 22380 3292 22389
rect 6736 22380 6788 22432
rect 8668 22423 8720 22432
rect 8668 22389 8677 22423
rect 8677 22389 8711 22423
rect 8711 22389 8720 22423
rect 8668 22380 8720 22389
rect 9128 22380 9180 22432
rect 9772 22423 9824 22432
rect 9772 22389 9781 22423
rect 9781 22389 9815 22423
rect 9815 22389 9824 22423
rect 9772 22380 9824 22389
rect 15568 22380 15620 22432
rect 15844 22423 15896 22432
rect 15844 22389 15853 22423
rect 15853 22389 15887 22423
rect 15887 22389 15896 22423
rect 15844 22380 15896 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 2504 22176 2556 22228
rect 3332 22176 3384 22228
rect 6920 22176 6972 22228
rect 8852 22219 8904 22228
rect 8852 22185 8861 22219
rect 8861 22185 8895 22219
rect 8895 22185 8904 22219
rect 8852 22176 8904 22185
rect 10692 22176 10744 22228
rect 1492 22040 1544 22092
rect 3056 22040 3108 22092
rect 4436 22040 4488 22092
rect 6736 22083 6788 22092
rect 6736 22049 6745 22083
rect 6745 22049 6779 22083
rect 6779 22049 6788 22083
rect 6736 22040 6788 22049
rect 9680 22083 9732 22092
rect 9680 22049 9689 22083
rect 9689 22049 9723 22083
rect 9723 22049 9732 22083
rect 9680 22040 9732 22049
rect 5080 22015 5132 22024
rect 5080 21981 5089 22015
rect 5089 21981 5123 22015
rect 5123 21981 5132 22015
rect 5080 21972 5132 21981
rect 10324 22015 10376 22024
rect 10324 21981 10333 22015
rect 10333 21981 10367 22015
rect 10367 21981 10376 22015
rect 10324 21972 10376 21981
rect 1860 21879 1912 21888
rect 1860 21845 1869 21879
rect 1869 21845 1903 21879
rect 1903 21845 1912 21879
rect 1860 21836 1912 21845
rect 1952 21836 2004 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 1492 21632 1544 21684
rect 3240 21675 3292 21684
rect 3240 21641 3249 21675
rect 3249 21641 3283 21675
rect 3283 21641 3292 21675
rect 3240 21632 3292 21641
rect 4436 21675 4488 21684
rect 4436 21641 4445 21675
rect 4445 21641 4479 21675
rect 4479 21641 4488 21675
rect 4436 21632 4488 21641
rect 9680 21675 9732 21684
rect 9680 21641 9689 21675
rect 9689 21641 9723 21675
rect 9723 21641 9732 21675
rect 9680 21632 9732 21641
rect 9864 21632 9916 21684
rect 1952 21539 2004 21548
rect 1952 21505 1961 21539
rect 1961 21505 1995 21539
rect 1995 21505 2004 21539
rect 1952 21496 2004 21505
rect 3056 21496 3108 21548
rect 8668 21539 8720 21548
rect 8668 21505 8677 21539
rect 8677 21505 8711 21539
rect 8711 21505 8720 21539
rect 8668 21496 8720 21505
rect 9128 21471 9180 21480
rect 1952 21360 2004 21412
rect 2688 21360 2740 21412
rect 3516 21403 3568 21412
rect 3516 21369 3525 21403
rect 3525 21369 3559 21403
rect 3559 21369 3568 21403
rect 3516 21360 3568 21369
rect 4988 21403 5040 21412
rect 3056 21292 3108 21344
rect 3240 21292 3292 21344
rect 4988 21369 4997 21403
rect 4997 21369 5031 21403
rect 5031 21369 5040 21403
rect 4988 21360 5040 21369
rect 4896 21335 4948 21344
rect 4896 21301 4905 21335
rect 4905 21301 4939 21335
rect 4939 21301 4948 21335
rect 9128 21437 9137 21471
rect 9137 21437 9171 21471
rect 9171 21437 9180 21471
rect 9128 21428 9180 21437
rect 4896 21292 4948 21301
rect 6736 21292 6788 21344
rect 11060 21335 11112 21344
rect 11060 21301 11069 21335
rect 11069 21301 11103 21335
rect 11103 21301 11112 21335
rect 11060 21292 11112 21301
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 3516 21131 3568 21140
rect 3516 21097 3525 21131
rect 3525 21097 3559 21131
rect 3559 21097 3568 21131
rect 3516 21088 3568 21097
rect 9680 21088 9732 21140
rect 2320 21020 2372 21072
rect 2688 21063 2740 21072
rect 2688 21029 2697 21063
rect 2697 21029 2731 21063
rect 2731 21029 2740 21063
rect 2688 21020 2740 21029
rect 5356 21063 5408 21072
rect 5356 21029 5365 21063
rect 5365 21029 5399 21063
rect 5399 21029 5408 21063
rect 5356 21020 5408 21029
rect 7564 20995 7616 21004
rect 7564 20961 7573 20995
rect 7573 20961 7607 20995
rect 7607 20961 7616 20995
rect 7564 20952 7616 20961
rect 9220 20952 9272 21004
rect 2044 20927 2096 20936
rect 2044 20893 2053 20927
rect 2053 20893 2087 20927
rect 2087 20893 2096 20927
rect 2044 20884 2096 20893
rect 5540 20927 5592 20936
rect 5540 20893 5549 20927
rect 5549 20893 5583 20927
rect 5583 20893 5592 20927
rect 5540 20884 5592 20893
rect 7288 20927 7340 20936
rect 7288 20893 7297 20927
rect 7297 20893 7331 20927
rect 7331 20893 7340 20927
rect 7288 20884 7340 20893
rect 11428 20927 11480 20936
rect 11428 20893 11437 20927
rect 11437 20893 11471 20927
rect 11471 20893 11480 20927
rect 11428 20884 11480 20893
rect 6000 20816 6052 20868
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 2044 20544 2096 20596
rect 6000 20587 6052 20596
rect 6000 20553 6009 20587
rect 6009 20553 6043 20587
rect 6043 20553 6052 20587
rect 6000 20544 6052 20553
rect 9220 20587 9272 20596
rect 9220 20553 9229 20587
rect 9229 20553 9263 20587
rect 9263 20553 9272 20587
rect 9220 20544 9272 20553
rect 11060 20544 11112 20596
rect 13912 20544 13964 20596
rect 4436 20476 4488 20528
rect 5172 20519 5224 20528
rect 5172 20485 5181 20519
rect 5181 20485 5215 20519
rect 5215 20485 5224 20519
rect 5172 20476 5224 20485
rect 8760 20519 8812 20528
rect 8760 20485 8769 20519
rect 8769 20485 8803 20519
rect 8803 20485 8812 20519
rect 8760 20476 8812 20485
rect 2688 20408 2740 20460
rect 3056 20408 3108 20460
rect 4620 20451 4672 20460
rect 4620 20417 4629 20451
rect 4629 20417 4663 20451
rect 4663 20417 4672 20451
rect 4620 20408 4672 20417
rect 5080 20408 5132 20460
rect 1124 20340 1176 20392
rect 9588 20383 9640 20392
rect 9588 20349 9597 20383
rect 9597 20349 9631 20383
rect 9631 20349 9640 20383
rect 9588 20340 9640 20349
rect 2780 20315 2832 20324
rect 2780 20281 2789 20315
rect 2789 20281 2823 20315
rect 2823 20281 2832 20315
rect 3056 20315 3108 20324
rect 2780 20272 2832 20281
rect 3056 20281 3065 20315
rect 3065 20281 3099 20315
rect 3099 20281 3108 20315
rect 3056 20272 3108 20281
rect 2320 20247 2372 20256
rect 2320 20213 2329 20247
rect 2329 20213 2363 20247
rect 2363 20213 2372 20247
rect 2320 20204 2372 20213
rect 4988 20272 5040 20324
rect 5356 20272 5408 20324
rect 6000 20272 6052 20324
rect 12348 20340 12400 20392
rect 22100 20544 22152 20596
rect 25136 20587 25188 20596
rect 25136 20553 25145 20587
rect 25145 20553 25179 20587
rect 25179 20553 25188 20587
rect 25136 20544 25188 20553
rect 25136 20340 25188 20392
rect 11796 20247 11848 20256
rect 11796 20213 11805 20247
rect 11805 20213 11839 20247
rect 11839 20213 11848 20247
rect 11796 20204 11848 20213
rect 12900 20204 12952 20256
rect 17132 20204 17184 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 2044 20000 2096 20052
rect 2688 20000 2740 20052
rect 4620 20043 4672 20052
rect 4620 20009 4629 20043
rect 4629 20009 4663 20043
rect 4663 20009 4672 20043
rect 4620 20000 4672 20009
rect 7564 20043 7616 20052
rect 7564 20009 7573 20043
rect 7573 20009 7607 20043
rect 7607 20009 7616 20043
rect 7564 20000 7616 20009
rect 1952 19975 2004 19984
rect 1952 19941 1961 19975
rect 1961 19941 1995 19975
rect 1995 19941 2004 19975
rect 1952 19932 2004 19941
rect 4988 19975 5040 19984
rect 4988 19941 4997 19975
rect 4997 19941 5031 19975
rect 5031 19941 5040 19975
rect 4988 19932 5040 19941
rect 5172 19932 5224 19984
rect 6552 19932 6604 19984
rect 7288 19932 7340 19984
rect 8208 19975 8260 19984
rect 8208 19941 8217 19975
rect 8217 19941 8251 19975
rect 8251 19941 8260 19975
rect 8208 19932 8260 19941
rect 8760 19975 8812 19984
rect 8760 19941 8769 19975
rect 8769 19941 8803 19975
rect 8803 19941 8812 19975
rect 8760 19932 8812 19941
rect 9772 19932 9824 19984
rect 11428 19932 11480 19984
rect 11888 19932 11940 19984
rect 2320 19907 2372 19916
rect 2320 19873 2329 19907
rect 2329 19873 2363 19907
rect 2363 19873 2372 19907
rect 2320 19864 2372 19873
rect 13452 19907 13504 19916
rect 13452 19873 13461 19907
rect 13461 19873 13495 19907
rect 13495 19873 13504 19907
rect 13452 19864 13504 19873
rect 5540 19796 5592 19848
rect 6092 19796 6144 19848
rect 10876 19796 10928 19848
rect 11796 19796 11848 19848
rect 12808 19796 12860 19848
rect 8484 19728 8536 19780
rect 7840 19703 7892 19712
rect 7840 19669 7849 19703
rect 7849 19669 7883 19703
rect 7883 19669 7892 19703
rect 7840 19660 7892 19669
rect 12624 19703 12676 19712
rect 12624 19669 12633 19703
rect 12633 19669 12667 19703
rect 12667 19669 12676 19703
rect 12624 19660 12676 19669
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 5540 19456 5592 19508
rect 6552 19499 6604 19508
rect 6552 19465 6561 19499
rect 6561 19465 6595 19499
rect 6595 19465 6604 19499
rect 6552 19456 6604 19465
rect 8208 19456 8260 19508
rect 9588 19456 9640 19508
rect 11428 19456 11480 19508
rect 13452 19499 13504 19508
rect 13452 19465 13461 19499
rect 13461 19465 13495 19499
rect 13495 19465 13504 19499
rect 13452 19456 13504 19465
rect 11888 19431 11940 19440
rect 11888 19397 11897 19431
rect 11897 19397 11931 19431
rect 11931 19397 11940 19431
rect 11888 19388 11940 19397
rect 7840 19320 7892 19372
rect 10876 19363 10928 19372
rect 10876 19329 10885 19363
rect 10885 19329 10919 19363
rect 10919 19329 10928 19363
rect 10876 19320 10928 19329
rect 12348 19320 12400 19372
rect 12624 19320 12676 19372
rect 12808 19363 12860 19372
rect 12808 19329 12817 19363
rect 12817 19329 12851 19363
rect 12851 19329 12860 19363
rect 12808 19320 12860 19329
rect 3332 19295 3384 19304
rect 3332 19261 3341 19295
rect 3341 19261 3375 19295
rect 3375 19261 3384 19295
rect 3332 19252 3384 19261
rect 2320 19116 2372 19168
rect 3240 19116 3292 19168
rect 9864 19295 9916 19304
rect 9864 19261 9873 19295
rect 9873 19261 9907 19295
rect 9907 19261 9916 19295
rect 9864 19252 9916 19261
rect 10784 19252 10836 19304
rect 4344 19227 4396 19236
rect 4344 19193 4353 19227
rect 4353 19193 4387 19227
rect 4387 19193 4396 19227
rect 4344 19184 4396 19193
rect 5264 19184 5316 19236
rect 7472 19184 7524 19236
rect 4988 19116 5040 19168
rect 5908 19116 5960 19168
rect 6092 19159 6144 19168
rect 6092 19125 6101 19159
rect 6101 19125 6135 19159
rect 6135 19125 6144 19159
rect 6092 19116 6144 19125
rect 7564 19116 7616 19168
rect 9772 19116 9824 19168
rect 10048 19159 10100 19168
rect 10048 19125 10057 19159
rect 10057 19125 10091 19159
rect 10091 19125 10100 19159
rect 10048 19116 10100 19125
rect 12532 19116 12584 19168
rect 13452 19116 13504 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 4344 18955 4396 18964
rect 4344 18921 4353 18955
rect 4353 18921 4387 18955
rect 4387 18921 4396 18955
rect 4344 18912 4396 18921
rect 5264 18912 5316 18964
rect 5908 18955 5960 18964
rect 5908 18921 5917 18955
rect 5917 18921 5951 18955
rect 5951 18921 5960 18955
rect 5908 18912 5960 18921
rect 7472 18912 7524 18964
rect 7656 18912 7708 18964
rect 8484 18955 8536 18964
rect 8484 18921 8493 18955
rect 8493 18921 8527 18955
rect 8527 18921 8536 18955
rect 8484 18912 8536 18921
rect 11152 18912 11204 18964
rect 12532 18955 12584 18964
rect 12532 18921 12541 18955
rect 12541 18921 12575 18955
rect 12575 18921 12584 18955
rect 12532 18912 12584 18921
rect 12900 18887 12952 18896
rect 12900 18853 12909 18887
rect 12909 18853 12943 18887
rect 12943 18853 12952 18887
rect 12900 18844 12952 18853
rect 12992 18887 13044 18896
rect 12992 18853 13001 18887
rect 13001 18853 13035 18887
rect 13035 18853 13044 18887
rect 12992 18844 13044 18853
rect 1400 18819 1452 18828
rect 1400 18785 1409 18819
rect 1409 18785 1443 18819
rect 1443 18785 1452 18819
rect 1400 18776 1452 18785
rect 2688 18819 2740 18828
rect 2688 18785 2697 18819
rect 2697 18785 2731 18819
rect 2731 18785 2740 18819
rect 2688 18776 2740 18785
rect 2872 18819 2924 18828
rect 2872 18785 2881 18819
rect 2881 18785 2915 18819
rect 2915 18785 2924 18819
rect 2872 18776 2924 18785
rect 3332 18776 3384 18828
rect 6000 18776 6052 18828
rect 3148 18751 3200 18760
rect 3148 18717 3157 18751
rect 3157 18717 3191 18751
rect 3191 18717 3200 18751
rect 3148 18708 3200 18717
rect 5356 18708 5408 18760
rect 7196 18751 7248 18760
rect 7196 18717 7205 18751
rect 7205 18717 7239 18751
rect 7239 18717 7248 18751
rect 7196 18708 7248 18717
rect 9956 18751 10008 18760
rect 9956 18717 9965 18751
rect 9965 18717 9999 18751
rect 9999 18717 10008 18751
rect 9956 18708 10008 18717
rect 11428 18708 11480 18760
rect 12624 18640 12676 18692
rect 2136 18572 2188 18624
rect 3332 18572 3384 18624
rect 4344 18572 4396 18624
rect 7012 18615 7064 18624
rect 7012 18581 7021 18615
rect 7021 18581 7055 18615
rect 7055 18581 7064 18615
rect 7012 18572 7064 18581
rect 8852 18615 8904 18624
rect 8852 18581 8861 18615
rect 8861 18581 8895 18615
rect 8895 18581 8904 18615
rect 8852 18572 8904 18581
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 112 18368 164 18420
rect 1400 18368 1452 18420
rect 2688 18368 2740 18420
rect 3976 18368 4028 18420
rect 6000 18368 6052 18420
rect 7472 18368 7524 18420
rect 3240 18343 3292 18352
rect 3240 18309 3249 18343
rect 3249 18309 3283 18343
rect 3283 18309 3292 18343
rect 3240 18300 3292 18309
rect 3148 18232 3200 18284
rect 2320 18207 2372 18216
rect 2320 18173 2329 18207
rect 2329 18173 2363 18207
rect 2363 18173 2372 18207
rect 2320 18164 2372 18173
rect 2872 18164 2924 18216
rect 4068 18164 4120 18216
rect 7840 18232 7892 18284
rect 4252 18096 4304 18148
rect 5080 18164 5132 18216
rect 6920 18207 6972 18216
rect 6920 18173 6929 18207
rect 6929 18173 6963 18207
rect 6963 18173 6972 18207
rect 6920 18164 6972 18173
rect 7012 18164 7064 18216
rect 3976 18028 4028 18080
rect 4344 18028 4396 18080
rect 5264 18028 5316 18080
rect 8852 18368 8904 18420
rect 10048 18368 10100 18420
rect 11152 18411 11204 18420
rect 11152 18377 11161 18411
rect 11161 18377 11195 18411
rect 11195 18377 11204 18411
rect 11152 18368 11204 18377
rect 12992 18368 13044 18420
rect 8852 18275 8904 18284
rect 8852 18241 8861 18275
rect 8861 18241 8895 18275
rect 8895 18241 8904 18275
rect 8852 18232 8904 18241
rect 9956 18232 10008 18284
rect 12624 18232 12676 18284
rect 8668 18139 8720 18148
rect 8668 18105 8677 18139
rect 8677 18105 8711 18139
rect 8711 18105 8720 18139
rect 8668 18096 8720 18105
rect 10140 18096 10192 18148
rect 10784 18139 10836 18148
rect 10784 18105 10793 18139
rect 10793 18105 10827 18139
rect 10827 18105 10836 18139
rect 10784 18096 10836 18105
rect 9312 18028 9364 18080
rect 11428 18071 11480 18080
rect 11428 18037 11437 18071
rect 11437 18037 11471 18071
rect 11471 18037 11480 18071
rect 11428 18028 11480 18037
rect 11520 18028 11572 18080
rect 12624 18139 12676 18148
rect 12624 18105 12633 18139
rect 12633 18105 12667 18139
rect 12667 18105 12676 18139
rect 12624 18096 12676 18105
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 3056 17824 3108 17876
rect 5080 17824 5132 17876
rect 5356 17824 5408 17876
rect 11796 17824 11848 17876
rect 4068 17756 4120 17808
rect 4252 17756 4304 17808
rect 1308 17688 1360 17740
rect 2688 17731 2740 17740
rect 2688 17697 2697 17731
rect 2697 17697 2731 17731
rect 2731 17697 2740 17731
rect 2688 17688 2740 17697
rect 2872 17731 2924 17740
rect 2872 17697 2881 17731
rect 2881 17697 2915 17731
rect 2915 17697 2924 17731
rect 2872 17688 2924 17697
rect 7196 17799 7248 17808
rect 7196 17765 7205 17799
rect 7205 17765 7239 17799
rect 7239 17765 7248 17799
rect 7196 17756 7248 17765
rect 7748 17756 7800 17808
rect 8852 17756 8904 17808
rect 9404 17756 9456 17808
rect 9956 17799 10008 17808
rect 9956 17765 9965 17799
rect 9965 17765 9999 17799
rect 9999 17765 10008 17799
rect 9956 17756 10008 17765
rect 10784 17756 10836 17808
rect 11152 17756 11204 17808
rect 11336 17756 11388 17808
rect 12900 17799 12952 17808
rect 12900 17765 12909 17799
rect 12909 17765 12943 17799
rect 12943 17765 12952 17799
rect 12900 17756 12952 17765
rect 7012 17731 7064 17740
rect 4068 17663 4120 17672
rect 4068 17629 4077 17663
rect 4077 17629 4111 17663
rect 4111 17629 4120 17663
rect 4068 17620 4120 17629
rect 4344 17620 4396 17672
rect 7012 17697 7021 17731
rect 7021 17697 7055 17731
rect 7055 17697 7064 17731
rect 7012 17688 7064 17697
rect 12256 17731 12308 17740
rect 12256 17697 12265 17731
rect 12265 17697 12299 17731
rect 12299 17697 12308 17731
rect 12256 17688 12308 17697
rect 12992 17688 13044 17740
rect 13544 17731 13596 17740
rect 6828 17620 6880 17672
rect 1768 17484 1820 17536
rect 1952 17527 2004 17536
rect 1952 17493 1961 17527
rect 1961 17493 1995 17527
rect 1995 17493 2004 17527
rect 1952 17484 2004 17493
rect 2320 17527 2372 17536
rect 2320 17493 2329 17527
rect 2329 17493 2363 17527
rect 2363 17493 2372 17527
rect 2320 17484 2372 17493
rect 4620 17484 4672 17536
rect 7380 17484 7432 17536
rect 11796 17620 11848 17672
rect 13544 17697 13553 17731
rect 13553 17697 13587 17731
rect 13587 17697 13596 17731
rect 13544 17688 13596 17697
rect 15384 17688 15436 17740
rect 9220 17552 9272 17604
rect 11152 17552 11204 17604
rect 13452 17620 13504 17672
rect 14556 17484 14608 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 1308 17280 1360 17332
rect 2872 17323 2924 17332
rect 2872 17289 2881 17323
rect 2881 17289 2915 17323
rect 2915 17289 2924 17323
rect 2872 17280 2924 17289
rect 6828 17280 6880 17332
rect 9220 17280 9272 17332
rect 9864 17280 9916 17332
rect 11336 17323 11388 17332
rect 11336 17289 11345 17323
rect 11345 17289 11379 17323
rect 11379 17289 11388 17323
rect 11336 17280 11388 17289
rect 11796 17323 11848 17332
rect 11796 17289 11805 17323
rect 11805 17289 11839 17323
rect 11839 17289 11848 17323
rect 11796 17280 11848 17289
rect 12256 17323 12308 17332
rect 12256 17289 12265 17323
rect 12265 17289 12299 17323
rect 12299 17289 12308 17323
rect 12256 17280 12308 17289
rect 12624 17280 12676 17332
rect 13452 17323 13504 17332
rect 13452 17289 13461 17323
rect 13461 17289 13495 17323
rect 13495 17289 13504 17323
rect 13452 17280 13504 17289
rect 8668 17212 8720 17264
rect 11980 17212 12032 17264
rect 10876 17144 10928 17196
rect 13544 17144 13596 17196
rect 15384 17187 15436 17196
rect 15384 17153 15393 17187
rect 15393 17153 15427 17187
rect 15427 17153 15436 17187
rect 15384 17144 15436 17153
rect 1952 17076 2004 17128
rect 3516 17119 3568 17128
rect 3516 17085 3525 17119
rect 3525 17085 3559 17119
rect 3559 17085 3568 17119
rect 3516 17076 3568 17085
rect 4988 17076 5040 17128
rect 5080 17119 5132 17128
rect 5080 17085 5089 17119
rect 5089 17085 5123 17119
rect 5123 17085 5132 17119
rect 5080 17076 5132 17085
rect 7012 17076 7064 17128
rect 8024 17076 8076 17128
rect 8300 17076 8352 17128
rect 9956 17119 10008 17128
rect 9956 17085 9965 17119
rect 9965 17085 9999 17119
rect 9999 17085 10008 17119
rect 9956 17076 10008 17085
rect 12256 17076 12308 17128
rect 3792 17051 3844 17060
rect 3792 17017 3801 17051
rect 3801 17017 3835 17051
rect 3835 17017 3844 17051
rect 3792 17008 3844 17017
rect 11336 17008 11388 17060
rect 1676 16940 1728 16992
rect 2688 16940 2740 16992
rect 2872 16940 2924 16992
rect 4252 16940 4304 16992
rect 4712 16983 4764 16992
rect 4712 16949 4721 16983
rect 4721 16949 4755 16983
rect 4755 16949 4764 16983
rect 4712 16940 4764 16949
rect 7748 16983 7800 16992
rect 7748 16949 7757 16983
rect 7757 16949 7791 16983
rect 7791 16949 7800 16983
rect 7748 16940 7800 16949
rect 8116 16983 8168 16992
rect 8116 16949 8125 16983
rect 8125 16949 8159 16983
rect 8159 16949 8168 16983
rect 8116 16940 8168 16949
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 4068 16736 4120 16788
rect 4712 16736 4764 16788
rect 6736 16779 6788 16788
rect 6736 16745 6745 16779
rect 6745 16745 6779 16779
rect 6779 16745 6788 16779
rect 6736 16736 6788 16745
rect 9404 16779 9456 16788
rect 9404 16745 9413 16779
rect 9413 16745 9447 16779
rect 9447 16745 9456 16779
rect 9404 16736 9456 16745
rect 1768 16668 1820 16720
rect 2228 16668 2280 16720
rect 2596 16711 2648 16720
rect 2596 16677 2605 16711
rect 2605 16677 2639 16711
rect 2639 16677 2648 16711
rect 2596 16668 2648 16677
rect 3516 16668 3568 16720
rect 3792 16668 3844 16720
rect 6000 16668 6052 16720
rect 6920 16668 6972 16720
rect 2320 16600 2372 16652
rect 4988 16600 5040 16652
rect 7656 16643 7708 16652
rect 7656 16609 7665 16643
rect 7665 16609 7699 16643
rect 7699 16609 7708 16643
rect 7656 16600 7708 16609
rect 7932 16600 7984 16652
rect 9956 16711 10008 16720
rect 9956 16677 9965 16711
rect 9965 16677 9999 16711
rect 9999 16677 10008 16711
rect 9956 16668 10008 16677
rect 10968 16668 11020 16720
rect 11428 16668 11480 16720
rect 10876 16643 10928 16652
rect 10876 16609 10885 16643
rect 10885 16609 10919 16643
rect 10919 16609 10928 16643
rect 10876 16600 10928 16609
rect 11980 16643 12032 16652
rect 11980 16609 11989 16643
rect 11989 16609 12023 16643
rect 12023 16609 12032 16643
rect 11980 16600 12032 16609
rect 4160 16575 4212 16584
rect 4160 16541 4169 16575
rect 4169 16541 4203 16575
rect 4203 16541 4212 16575
rect 4160 16532 4212 16541
rect 3056 16507 3108 16516
rect 3056 16473 3065 16507
rect 3065 16473 3099 16507
rect 3099 16473 3108 16507
rect 5448 16532 5500 16584
rect 7748 16532 7800 16584
rect 3056 16464 3108 16473
rect 1400 16396 1452 16448
rect 1860 16439 1912 16448
rect 1860 16405 1869 16439
rect 1869 16405 1903 16439
rect 1903 16405 1912 16439
rect 1860 16396 1912 16405
rect 2320 16439 2372 16448
rect 2320 16405 2329 16439
rect 2329 16405 2363 16439
rect 2363 16405 2372 16439
rect 2320 16396 2372 16405
rect 3516 16439 3568 16448
rect 3516 16405 3525 16439
rect 3525 16405 3559 16439
rect 3559 16405 3568 16439
rect 3516 16396 3568 16405
rect 4344 16396 4396 16448
rect 8300 16396 8352 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 2596 16192 2648 16244
rect 3792 16192 3844 16244
rect 7656 16235 7708 16244
rect 7656 16201 7665 16235
rect 7665 16201 7699 16235
rect 7699 16201 7708 16235
rect 7656 16192 7708 16201
rect 9128 16235 9180 16244
rect 9128 16201 9137 16235
rect 9137 16201 9171 16235
rect 9171 16201 9180 16235
rect 9128 16192 9180 16201
rect 9496 16235 9548 16244
rect 9496 16201 9505 16235
rect 9505 16201 9539 16235
rect 9539 16201 9548 16235
rect 11980 16235 12032 16244
rect 9496 16192 9548 16201
rect 1860 16056 1912 16108
rect 2320 16056 2372 16108
rect 11980 16201 11989 16235
rect 11989 16201 12023 16235
rect 12023 16201 12032 16235
rect 11980 16192 12032 16201
rect 10140 16056 10192 16108
rect 4344 15988 4396 16040
rect 5080 16031 5132 16040
rect 5080 15997 5089 16031
rect 5089 15997 5123 16031
rect 5123 15997 5132 16031
rect 5080 15988 5132 15997
rect 5448 15988 5500 16040
rect 8208 16031 8260 16040
rect 8208 15997 8217 16031
rect 8217 15997 8251 16031
rect 8251 15997 8260 16031
rect 8208 15988 8260 15997
rect 10968 15988 11020 16040
rect 1584 15963 1636 15972
rect 1584 15929 1593 15963
rect 1593 15929 1627 15963
rect 1627 15929 1636 15963
rect 1584 15920 1636 15929
rect 3056 15963 3108 15972
rect 3056 15929 3065 15963
rect 3065 15929 3099 15963
rect 3099 15929 3108 15963
rect 3056 15920 3108 15929
rect 2964 15852 3016 15904
rect 5264 15920 5316 15972
rect 7932 15920 7984 15972
rect 10140 15963 10192 15972
rect 10140 15929 10149 15963
rect 10149 15929 10183 15963
rect 10183 15929 10192 15963
rect 10140 15920 10192 15929
rect 10784 15920 10836 15972
rect 4620 15895 4672 15904
rect 4620 15861 4629 15895
rect 4629 15861 4663 15895
rect 4663 15861 4672 15895
rect 4620 15852 4672 15861
rect 6000 15852 6052 15904
rect 8116 15852 8168 15904
rect 9588 15852 9640 15904
rect 10876 15852 10928 15904
rect 11060 15895 11112 15904
rect 11060 15861 11069 15895
rect 11069 15861 11103 15895
rect 11103 15861 11112 15895
rect 11060 15852 11112 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 1860 15648 1912 15700
rect 2228 15691 2280 15700
rect 2228 15657 2237 15691
rect 2237 15657 2271 15691
rect 2271 15657 2280 15691
rect 2228 15648 2280 15657
rect 3056 15648 3108 15700
rect 3516 15648 3568 15700
rect 10140 15648 10192 15700
rect 4160 15580 4212 15632
rect 4252 15580 4304 15632
rect 6368 15580 6420 15632
rect 8300 15623 8352 15632
rect 8300 15589 8309 15623
rect 8309 15589 8343 15623
rect 8343 15589 8352 15623
rect 8300 15580 8352 15589
rect 9956 15580 10008 15632
rect 10784 15580 10836 15632
rect 11612 15580 11664 15632
rect 12808 15580 12860 15632
rect 1584 15512 1636 15564
rect 2964 15555 3016 15564
rect 2964 15521 2973 15555
rect 2973 15521 3007 15555
rect 3007 15521 3016 15555
rect 2964 15512 3016 15521
rect 7104 15512 7156 15564
rect 7932 15512 7984 15564
rect 4528 15444 4580 15496
rect 6184 15444 6236 15496
rect 10324 15487 10376 15496
rect 10324 15453 10333 15487
rect 10333 15453 10367 15487
rect 10367 15453 10376 15487
rect 10324 15444 10376 15453
rect 10968 15487 11020 15496
rect 10968 15453 10977 15487
rect 10977 15453 11011 15487
rect 11011 15453 11020 15487
rect 10968 15444 11020 15453
rect 12532 15487 12584 15496
rect 12532 15453 12541 15487
rect 12541 15453 12575 15487
rect 12575 15453 12584 15487
rect 12532 15444 12584 15453
rect 13360 15487 13412 15496
rect 13360 15453 13369 15487
rect 13369 15453 13403 15487
rect 13403 15453 13412 15487
rect 13360 15444 13412 15453
rect 6276 15376 6328 15428
rect 8392 15376 8444 15428
rect 5080 15308 5132 15360
rect 5356 15308 5408 15360
rect 7196 15351 7248 15360
rect 7196 15317 7205 15351
rect 7205 15317 7239 15351
rect 7239 15317 7248 15351
rect 7196 15308 7248 15317
rect 7840 15308 7892 15360
rect 8208 15308 8260 15360
rect 12808 15351 12860 15360
rect 12808 15317 12817 15351
rect 12817 15317 12851 15351
rect 12851 15317 12860 15351
rect 12808 15308 12860 15317
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 1492 15104 1544 15156
rect 2964 15104 3016 15156
rect 6276 15104 6328 15156
rect 7288 15104 7340 15156
rect 8116 15104 8168 15156
rect 9956 15147 10008 15156
rect 1952 15036 2004 15088
rect 6184 14968 6236 15020
rect 7840 15011 7892 15020
rect 7840 14977 7849 15011
rect 7849 14977 7883 15011
rect 7883 14977 7892 15011
rect 7840 14968 7892 14977
rect 9956 15113 9965 15147
rect 9965 15113 9999 15147
rect 9999 15113 10008 15147
rect 9956 15104 10008 15113
rect 10324 15104 10376 15156
rect 13360 15104 13412 15156
rect 25136 15147 25188 15156
rect 25136 15113 25145 15147
rect 25145 15113 25179 15147
rect 25179 15113 25188 15147
rect 25136 15104 25188 15113
rect 10140 15036 10192 15088
rect 1400 14943 1452 14952
rect 1400 14909 1409 14943
rect 1409 14909 1443 14943
rect 1443 14909 1452 14943
rect 1400 14900 1452 14909
rect 3056 14943 3108 14952
rect 3056 14909 3065 14943
rect 3065 14909 3099 14943
rect 3099 14909 3108 14943
rect 3056 14900 3108 14909
rect 7104 14943 7156 14952
rect 7104 14909 7113 14943
rect 7113 14909 7147 14943
rect 7147 14909 7156 14943
rect 7104 14900 7156 14909
rect 7196 14900 7248 14952
rect 8116 14900 8168 14952
rect 8392 14900 8444 14952
rect 5264 14875 5316 14884
rect 2964 14807 3016 14816
rect 2964 14773 2973 14807
rect 2973 14773 3007 14807
rect 3007 14773 3016 14807
rect 5264 14841 5273 14875
rect 5273 14841 5307 14875
rect 5307 14841 5316 14875
rect 5264 14832 5316 14841
rect 4252 14807 4304 14816
rect 2964 14764 3016 14773
rect 4252 14773 4261 14807
rect 4261 14773 4295 14807
rect 4295 14773 4304 14807
rect 4252 14764 4304 14773
rect 6828 14832 6880 14884
rect 10048 14968 10100 15020
rect 10968 14968 11020 15020
rect 11244 14900 11296 14952
rect 12808 14943 12860 14952
rect 12808 14909 12817 14943
rect 12817 14909 12851 14943
rect 12851 14909 12860 14943
rect 12808 14900 12860 14909
rect 25136 14900 25188 14952
rect 12440 14875 12492 14884
rect 12440 14841 12449 14875
rect 12449 14841 12483 14875
rect 12483 14841 12492 14875
rect 12440 14832 12492 14841
rect 6368 14764 6420 14816
rect 12164 14764 12216 14816
rect 19248 14764 19300 14816
rect 24216 14764 24268 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 3056 14560 3108 14612
rect 3516 14560 3568 14612
rect 5356 14560 5408 14612
rect 6644 14560 6696 14612
rect 9772 14560 9824 14612
rect 10048 14603 10100 14612
rect 10048 14569 10057 14603
rect 10057 14569 10091 14603
rect 10091 14569 10100 14603
rect 10048 14560 10100 14569
rect 10692 14560 10744 14612
rect 11244 14603 11296 14612
rect 11244 14569 11253 14603
rect 11253 14569 11287 14603
rect 11287 14569 11296 14603
rect 11244 14560 11296 14569
rect 11612 14560 11664 14612
rect 5448 14492 5500 14544
rect 6000 14492 6052 14544
rect 8392 14535 8444 14544
rect 8392 14501 8401 14535
rect 8401 14501 8435 14535
rect 8435 14501 8444 14535
rect 8392 14492 8444 14501
rect 12164 14535 12216 14544
rect 12164 14501 12173 14535
rect 12173 14501 12207 14535
rect 12207 14501 12216 14535
rect 12164 14492 12216 14501
rect 12440 14492 12492 14544
rect 2320 14424 2372 14476
rect 2688 14467 2740 14476
rect 2688 14433 2697 14467
rect 2697 14433 2731 14467
rect 2731 14433 2740 14467
rect 2688 14424 2740 14433
rect 3424 14424 3476 14476
rect 4436 14467 4488 14476
rect 4436 14433 4445 14467
rect 4445 14433 4479 14467
rect 4479 14433 4488 14467
rect 4436 14424 4488 14433
rect 5540 14424 5592 14476
rect 7656 14467 7708 14476
rect 7656 14433 7665 14467
rect 7665 14433 7699 14467
rect 7699 14433 7708 14467
rect 7656 14424 7708 14433
rect 7840 14424 7892 14476
rect 8116 14467 8168 14476
rect 8116 14433 8125 14467
rect 8125 14433 8159 14467
rect 8159 14433 8168 14467
rect 8116 14424 8168 14433
rect 13176 14424 13228 14476
rect 4344 14356 4396 14408
rect 5448 14399 5500 14408
rect 1400 14288 1452 14340
rect 5448 14365 5457 14399
rect 5457 14365 5491 14399
rect 5491 14365 5500 14399
rect 5448 14356 5500 14365
rect 7104 14331 7156 14340
rect 7104 14297 7113 14331
rect 7113 14297 7147 14331
rect 7147 14297 7156 14331
rect 7104 14288 7156 14297
rect 12532 14399 12584 14408
rect 12532 14365 12541 14399
rect 12541 14365 12575 14399
rect 12575 14365 12584 14399
rect 12532 14356 12584 14365
rect 13636 14399 13688 14408
rect 13636 14365 13645 14399
rect 13645 14365 13679 14399
rect 13679 14365 13688 14399
rect 13636 14356 13688 14365
rect 15660 14356 15712 14408
rect 1860 14263 1912 14272
rect 1860 14229 1869 14263
rect 1869 14229 1903 14263
rect 1903 14229 1912 14263
rect 1860 14220 1912 14229
rect 2320 14263 2372 14272
rect 2320 14229 2329 14263
rect 2329 14229 2363 14263
rect 2363 14229 2372 14263
rect 2320 14220 2372 14229
rect 3792 14263 3844 14272
rect 3792 14229 3801 14263
rect 3801 14229 3835 14263
rect 3835 14229 3844 14263
rect 3792 14220 3844 14229
rect 4528 14220 4580 14272
rect 5172 14220 5224 14272
rect 5356 14263 5408 14272
rect 5356 14229 5365 14263
rect 5365 14229 5399 14263
rect 5399 14229 5408 14263
rect 5356 14220 5408 14229
rect 6368 14263 6420 14272
rect 6368 14229 6377 14263
rect 6377 14229 6411 14263
rect 6411 14229 6420 14263
rect 6368 14220 6420 14229
rect 7932 14220 7984 14272
rect 8760 14263 8812 14272
rect 8760 14229 8769 14263
rect 8769 14229 8803 14263
rect 8803 14229 8812 14263
rect 8760 14220 8812 14229
rect 8852 14220 8904 14272
rect 9496 14263 9548 14272
rect 9496 14229 9505 14263
rect 9505 14229 9539 14263
rect 9539 14229 9548 14263
rect 9496 14220 9548 14229
rect 10876 14263 10928 14272
rect 10876 14229 10885 14263
rect 10885 14229 10919 14263
rect 10919 14229 10928 14263
rect 10876 14220 10928 14229
rect 15292 14220 15344 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 1584 14059 1636 14068
rect 1584 14025 1593 14059
rect 1593 14025 1627 14059
rect 1627 14025 1636 14059
rect 1584 14016 1636 14025
rect 4436 14016 4488 14068
rect 9496 14059 9548 14068
rect 9496 14025 9505 14059
rect 9505 14025 9539 14059
rect 9539 14025 9548 14059
rect 9496 14016 9548 14025
rect 12440 14016 12492 14068
rect 13176 14059 13228 14068
rect 13176 14025 13185 14059
rect 13185 14025 13219 14059
rect 13219 14025 13228 14059
rect 13176 14016 13228 14025
rect 13636 14016 13688 14068
rect 15660 14059 15712 14068
rect 15660 14025 15669 14059
rect 15669 14025 15703 14059
rect 15703 14025 15712 14059
rect 15660 14016 15712 14025
rect 5356 13948 5408 14000
rect 11244 13991 11296 14000
rect 2688 13880 2740 13932
rect 1676 13812 1728 13864
rect 2044 13812 2096 13864
rect 3332 13855 3384 13864
rect 3332 13821 3341 13855
rect 3341 13821 3375 13855
rect 3375 13821 3384 13855
rect 3332 13812 3384 13821
rect 3424 13812 3476 13864
rect 3608 13812 3660 13864
rect 4620 13855 4672 13864
rect 4620 13821 4629 13855
rect 4629 13821 4663 13855
rect 4663 13821 4672 13855
rect 4620 13812 4672 13821
rect 5540 13812 5592 13864
rect 11244 13957 11253 13991
rect 11253 13957 11287 13991
rect 11287 13957 11296 13991
rect 11244 13948 11296 13957
rect 12348 13948 12400 14000
rect 6368 13880 6420 13932
rect 6828 13855 6880 13864
rect 6828 13821 6837 13855
rect 6837 13821 6871 13855
rect 6871 13821 6880 13855
rect 6828 13812 6880 13821
rect 8760 13880 8812 13932
rect 12164 13880 12216 13932
rect 13728 13923 13780 13932
rect 13728 13889 13737 13923
rect 13737 13889 13771 13923
rect 13771 13889 13780 13923
rect 13728 13880 13780 13889
rect 5356 13744 5408 13796
rect 4528 13676 4580 13728
rect 5172 13676 5224 13728
rect 7196 13744 7248 13796
rect 6000 13719 6052 13728
rect 6000 13685 6009 13719
rect 6009 13685 6043 13719
rect 6043 13685 6052 13719
rect 6000 13676 6052 13685
rect 7656 13676 7708 13728
rect 8208 13676 8260 13728
rect 9128 13812 9180 13864
rect 10876 13855 10928 13864
rect 10876 13821 10885 13855
rect 10885 13821 10919 13855
rect 10919 13821 10928 13855
rect 10876 13812 10928 13821
rect 10968 13812 11020 13864
rect 12532 13812 12584 13864
rect 14372 13787 14424 13796
rect 9772 13676 9824 13728
rect 9956 13676 10008 13728
rect 13636 13676 13688 13728
rect 14372 13753 14381 13787
rect 14381 13753 14415 13787
rect 14415 13753 14424 13787
rect 14372 13744 14424 13753
rect 14464 13676 14516 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 2044 13472 2096 13524
rect 2136 13472 2188 13524
rect 3056 13472 3108 13524
rect 3516 13472 3568 13524
rect 5448 13472 5500 13524
rect 6736 13472 6788 13524
rect 8576 13515 8628 13524
rect 1952 13336 2004 13388
rect 2504 13336 2556 13388
rect 6644 13404 6696 13456
rect 8576 13481 8585 13515
rect 8585 13481 8619 13515
rect 8619 13481 8628 13515
rect 8576 13472 8628 13481
rect 9128 13472 9180 13524
rect 4620 13379 4672 13388
rect 4620 13345 4629 13379
rect 4629 13345 4663 13379
rect 4663 13345 4672 13379
rect 4620 13336 4672 13345
rect 5264 13379 5316 13388
rect 5264 13345 5273 13379
rect 5273 13345 5307 13379
rect 5307 13345 5316 13379
rect 5264 13336 5316 13345
rect 5448 13379 5500 13388
rect 5448 13345 5457 13379
rect 5457 13345 5491 13379
rect 5491 13345 5500 13379
rect 5448 13336 5500 13345
rect 24584 13472 24636 13524
rect 11980 13404 12032 13456
rect 12532 13404 12584 13456
rect 10140 13336 10192 13388
rect 12256 13379 12308 13388
rect 12256 13345 12265 13379
rect 12265 13345 12299 13379
rect 12299 13345 12308 13379
rect 12256 13336 12308 13345
rect 3148 13311 3200 13320
rect 3148 13277 3157 13311
rect 3157 13277 3191 13311
rect 3191 13277 3200 13311
rect 3148 13268 3200 13277
rect 3332 13268 3384 13320
rect 4528 13268 4580 13320
rect 7564 13311 7616 13320
rect 3424 13200 3476 13252
rect 7564 13277 7573 13311
rect 7573 13277 7607 13311
rect 7607 13277 7616 13311
rect 7564 13268 7616 13277
rect 12440 13268 12492 13320
rect 13176 13404 13228 13456
rect 14372 13447 14424 13456
rect 14372 13413 14381 13447
rect 14381 13413 14415 13447
rect 14415 13413 14424 13447
rect 14372 13404 14424 13413
rect 15292 13379 15344 13388
rect 15292 13345 15301 13379
rect 15301 13345 15335 13379
rect 15335 13345 15344 13379
rect 15292 13336 15344 13345
rect 24860 13336 24912 13388
rect 13728 13311 13780 13320
rect 13728 13277 13737 13311
rect 13737 13277 13771 13311
rect 13771 13277 13780 13311
rect 13728 13268 13780 13277
rect 15752 13200 15804 13252
rect 2136 13132 2188 13184
rect 2320 13175 2372 13184
rect 2320 13141 2329 13175
rect 2329 13141 2363 13175
rect 2363 13141 2372 13175
rect 2320 13132 2372 13141
rect 3516 13175 3568 13184
rect 3516 13141 3525 13175
rect 3525 13141 3559 13175
rect 3559 13141 3568 13175
rect 3516 13132 3568 13141
rect 4528 13175 4580 13184
rect 4528 13141 4537 13175
rect 4537 13141 4571 13175
rect 4571 13141 4580 13175
rect 4528 13132 4580 13141
rect 4988 13132 5040 13184
rect 6552 13132 6604 13184
rect 7840 13132 7892 13184
rect 8576 13132 8628 13184
rect 9680 13132 9732 13184
rect 10968 13132 11020 13184
rect 11152 13175 11204 13184
rect 11152 13141 11161 13175
rect 11161 13141 11195 13175
rect 11195 13141 11204 13175
rect 11152 13132 11204 13141
rect 15844 13132 15896 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 112 12928 164 12980
rect 1952 12971 2004 12980
rect 1952 12937 1961 12971
rect 1961 12937 1995 12971
rect 1995 12937 2004 12971
rect 1952 12928 2004 12937
rect 2504 12971 2556 12980
rect 2504 12937 2513 12971
rect 2513 12937 2547 12971
rect 2547 12937 2556 12971
rect 2504 12928 2556 12937
rect 3148 12928 3200 12980
rect 7472 12928 7524 12980
rect 9312 12971 9364 12980
rect 9312 12937 9321 12971
rect 9321 12937 9355 12971
rect 9355 12937 9364 12971
rect 9312 12928 9364 12937
rect 13176 12928 13228 12980
rect 15292 12971 15344 12980
rect 15292 12937 15301 12971
rect 15301 12937 15335 12971
rect 15335 12937 15344 12971
rect 15292 12928 15344 12937
rect 24860 12928 24912 12980
rect 4344 12903 4396 12912
rect 4344 12869 4353 12903
rect 4353 12869 4387 12903
rect 4387 12869 4396 12903
rect 4344 12860 4396 12869
rect 5080 12860 5132 12912
rect 5448 12860 5500 12912
rect 8668 12860 8720 12912
rect 3792 12792 3844 12844
rect 7564 12792 7616 12844
rect 10692 12792 10744 12844
rect 11152 12792 11204 12844
rect 12440 12835 12492 12844
rect 12440 12801 12449 12835
rect 12449 12801 12483 12835
rect 12483 12801 12492 12835
rect 12440 12792 12492 12801
rect 1400 12767 1452 12776
rect 1400 12733 1409 12767
rect 1409 12733 1443 12767
rect 1443 12733 1452 12767
rect 1400 12724 1452 12733
rect 4344 12724 4396 12776
rect 4804 12724 4856 12776
rect 4988 12724 5040 12776
rect 8576 12724 8628 12776
rect 8944 12724 8996 12776
rect 14280 12767 14332 12776
rect 14280 12733 14289 12767
rect 14289 12733 14323 12767
rect 14323 12733 14332 12767
rect 14280 12724 14332 12733
rect 3332 12656 3384 12708
rect 3700 12699 3752 12708
rect 3700 12665 3709 12699
rect 3709 12665 3743 12699
rect 3743 12665 3752 12699
rect 3700 12656 3752 12665
rect 4068 12656 4120 12708
rect 4620 12631 4672 12640
rect 4620 12597 4629 12631
rect 4629 12597 4663 12631
rect 4663 12597 4672 12631
rect 4620 12588 4672 12597
rect 5816 12588 5868 12640
rect 6552 12631 6604 12640
rect 6552 12597 6561 12631
rect 6561 12597 6595 12631
rect 6595 12597 6604 12631
rect 6552 12588 6604 12597
rect 7472 12699 7524 12708
rect 7472 12665 7481 12699
rect 7481 12665 7515 12699
rect 7515 12665 7524 12699
rect 7472 12656 7524 12665
rect 8760 12656 8812 12708
rect 9956 12656 10008 12708
rect 14188 12699 14240 12708
rect 14188 12665 14197 12699
rect 14197 12665 14231 12699
rect 14231 12665 14240 12699
rect 14188 12656 14240 12665
rect 8024 12588 8076 12640
rect 8668 12631 8720 12640
rect 8668 12597 8677 12631
rect 8677 12597 8711 12631
rect 8711 12597 8720 12631
rect 8668 12588 8720 12597
rect 9680 12588 9732 12640
rect 11980 12588 12032 12640
rect 12256 12631 12308 12640
rect 12256 12597 12265 12631
rect 12265 12597 12299 12631
rect 12299 12597 12308 12631
rect 12256 12588 12308 12597
rect 15384 12588 15436 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 3424 12384 3476 12436
rect 4068 12384 4120 12436
rect 4344 12427 4396 12436
rect 4344 12393 4353 12427
rect 4353 12393 4387 12427
rect 4387 12393 4396 12427
rect 4344 12384 4396 12393
rect 6736 12427 6788 12436
rect 6736 12393 6745 12427
rect 6745 12393 6779 12427
rect 6779 12393 6788 12427
rect 6736 12384 6788 12393
rect 8852 12427 8904 12436
rect 8852 12393 8861 12427
rect 8861 12393 8895 12427
rect 8895 12393 8904 12427
rect 8852 12384 8904 12393
rect 2504 12316 2556 12368
rect 2688 12316 2740 12368
rect 3700 12316 3752 12368
rect 6000 12316 6052 12368
rect 10140 12384 10192 12436
rect 1952 12248 2004 12300
rect 4252 12291 4304 12300
rect 4252 12257 4261 12291
rect 4261 12257 4295 12291
rect 4295 12257 4304 12291
rect 4252 12248 4304 12257
rect 4988 12248 5040 12300
rect 5816 12291 5868 12300
rect 5816 12257 5825 12291
rect 5825 12257 5859 12291
rect 5859 12257 5868 12291
rect 5816 12248 5868 12257
rect 7104 12248 7156 12300
rect 9680 12291 9732 12300
rect 9680 12257 9689 12291
rect 9689 12257 9723 12291
rect 9723 12257 9732 12291
rect 9680 12248 9732 12257
rect 12440 12427 12492 12436
rect 10692 12316 10744 12368
rect 12440 12393 12449 12427
rect 12449 12393 12483 12427
rect 12483 12393 12492 12427
rect 12440 12384 12492 12393
rect 13728 12384 13780 12436
rect 11428 12359 11480 12368
rect 11428 12325 11437 12359
rect 11437 12325 11471 12359
rect 11471 12325 11480 12359
rect 11428 12316 11480 12325
rect 11980 12248 12032 12300
rect 13820 12248 13872 12300
rect 7656 12180 7708 12232
rect 3516 12112 3568 12164
rect 5264 12112 5316 12164
rect 8024 12180 8076 12232
rect 11336 12223 11388 12232
rect 11336 12189 11345 12223
rect 11345 12189 11379 12223
rect 11379 12189 11388 12223
rect 12808 12223 12860 12232
rect 11336 12180 11388 12189
rect 8576 12112 8628 12164
rect 11888 12155 11940 12164
rect 11888 12121 11897 12155
rect 11897 12121 11931 12155
rect 11931 12121 11940 12155
rect 11888 12112 11940 12121
rect 12808 12189 12817 12223
rect 12817 12189 12851 12223
rect 12851 12189 12860 12223
rect 12808 12180 12860 12189
rect 15292 12384 15344 12436
rect 15476 12180 15528 12232
rect 16028 12223 16080 12232
rect 16028 12189 16037 12223
rect 16037 12189 16071 12223
rect 16071 12189 16080 12223
rect 16028 12180 16080 12189
rect 1952 12087 2004 12096
rect 1952 12053 1961 12087
rect 1961 12053 1995 12087
rect 1995 12053 2004 12087
rect 1952 12044 2004 12053
rect 2228 12087 2280 12096
rect 2228 12053 2237 12087
rect 2237 12053 2271 12087
rect 2271 12053 2280 12087
rect 2228 12044 2280 12053
rect 4896 12044 4948 12096
rect 6552 12044 6604 12096
rect 7472 12044 7524 12096
rect 7564 12044 7616 12096
rect 10140 12044 10192 12096
rect 14464 12044 14516 12096
rect 17224 12087 17276 12096
rect 17224 12053 17233 12087
rect 17233 12053 17267 12087
rect 17267 12053 17276 12087
rect 17224 12044 17276 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 4712 11840 4764 11892
rect 4896 11815 4948 11824
rect 4896 11781 4920 11815
rect 4920 11781 4948 11815
rect 4896 11772 4948 11781
rect 5172 11815 5224 11824
rect 5172 11781 5181 11815
rect 5181 11781 5215 11815
rect 5215 11781 5224 11815
rect 5172 11772 5224 11781
rect 6552 11772 6604 11824
rect 6920 11772 6972 11824
rect 7564 11840 7616 11892
rect 7840 11883 7892 11892
rect 7840 11849 7849 11883
rect 7849 11849 7883 11883
rect 7883 11849 7892 11883
rect 7840 11840 7892 11849
rect 8116 11840 8168 11892
rect 10140 11883 10192 11892
rect 10140 11849 10149 11883
rect 10149 11849 10183 11883
rect 10183 11849 10192 11883
rect 10140 11840 10192 11849
rect 10784 11840 10836 11892
rect 11428 11840 11480 11892
rect 12808 11840 12860 11892
rect 14280 11883 14332 11892
rect 14280 11849 14289 11883
rect 14289 11849 14323 11883
rect 14323 11849 14332 11883
rect 14280 11840 14332 11849
rect 7472 11815 7524 11824
rect 7472 11781 7481 11815
rect 7481 11781 7515 11815
rect 7515 11781 7524 11815
rect 7472 11772 7524 11781
rect 8852 11772 8904 11824
rect 2320 11704 2372 11756
rect 4344 11704 4396 11756
rect 1400 11679 1452 11688
rect 1400 11645 1409 11679
rect 1409 11645 1443 11679
rect 1443 11645 1452 11679
rect 1400 11636 1452 11645
rect 1860 11636 1912 11688
rect 2504 11636 2556 11688
rect 7012 11704 7064 11756
rect 5172 11636 5224 11688
rect 8760 11704 8812 11756
rect 13820 11815 13872 11824
rect 13820 11781 13829 11815
rect 13829 11781 13863 11815
rect 13863 11781 13872 11815
rect 13820 11772 13872 11781
rect 19984 11772 20036 11824
rect 14464 11747 14516 11756
rect 14464 11713 14473 11747
rect 14473 11713 14507 11747
rect 14507 11713 14516 11747
rect 14464 11704 14516 11713
rect 14832 11704 14884 11756
rect 15476 11704 15528 11756
rect 10784 11679 10836 11688
rect 10784 11645 10793 11679
rect 10793 11645 10827 11679
rect 10827 11645 10836 11679
rect 10784 11636 10836 11645
rect 12164 11636 12216 11688
rect 12624 11679 12676 11688
rect 12624 11645 12633 11679
rect 12633 11645 12667 11679
rect 12667 11645 12676 11679
rect 12624 11636 12676 11645
rect 2964 11568 3016 11620
rect 112 11500 164 11552
rect 2044 11543 2096 11552
rect 2044 11509 2053 11543
rect 2053 11509 2087 11543
rect 2087 11509 2096 11543
rect 2044 11500 2096 11509
rect 2412 11543 2464 11552
rect 2412 11509 2421 11543
rect 2421 11509 2455 11543
rect 2455 11509 2464 11543
rect 2412 11500 2464 11509
rect 3424 11500 3476 11552
rect 4528 11568 4580 11620
rect 5356 11568 5408 11620
rect 7288 11568 7340 11620
rect 8576 11568 8628 11620
rect 12808 11568 12860 11620
rect 6000 11500 6052 11552
rect 6184 11543 6236 11552
rect 6184 11509 6193 11543
rect 6193 11509 6227 11543
rect 6227 11509 6236 11543
rect 6184 11500 6236 11509
rect 7012 11543 7064 11552
rect 7012 11509 7021 11543
rect 7021 11509 7055 11543
rect 7055 11509 7064 11543
rect 7012 11500 7064 11509
rect 7656 11500 7708 11552
rect 9956 11500 10008 11552
rect 12256 11543 12308 11552
rect 12256 11509 12265 11543
rect 12265 11509 12299 11543
rect 12299 11509 12308 11543
rect 12256 11500 12308 11509
rect 13452 11500 13504 11552
rect 14280 11500 14332 11552
rect 15476 11568 15528 11620
rect 15292 11500 15344 11552
rect 17224 11500 17276 11552
rect 19432 11500 19484 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 2228 11296 2280 11348
rect 4528 11296 4580 11348
rect 2412 11271 2464 11280
rect 2412 11237 2421 11271
rect 2421 11237 2455 11271
rect 2455 11237 2464 11271
rect 2412 11228 2464 11237
rect 4988 11296 5040 11348
rect 7932 11339 7984 11348
rect 7932 11305 7941 11339
rect 7941 11305 7975 11339
rect 7975 11305 7984 11339
rect 7932 11296 7984 11305
rect 8852 11296 8904 11348
rect 7104 11271 7156 11280
rect 7104 11237 7113 11271
rect 7113 11237 7147 11271
rect 7147 11237 7156 11271
rect 7104 11228 7156 11237
rect 11336 11296 11388 11348
rect 15292 11296 15344 11348
rect 3424 11160 3476 11212
rect 5356 11160 5408 11212
rect 6828 11160 6880 11212
rect 7196 11160 7248 11212
rect 8668 11160 8720 11212
rect 5172 11092 5224 11144
rect 5448 11092 5500 11144
rect 6184 11092 6236 11144
rect 7932 11092 7984 11144
rect 12624 11228 12676 11280
rect 13452 11228 13504 11280
rect 14464 11271 14516 11280
rect 14464 11237 14473 11271
rect 14473 11237 14507 11271
rect 14507 11237 14516 11271
rect 14464 11228 14516 11237
rect 15384 11271 15436 11280
rect 15384 11237 15393 11271
rect 15393 11237 15427 11271
rect 15427 11237 15436 11271
rect 15384 11228 15436 11237
rect 15476 11271 15528 11280
rect 15476 11237 15485 11271
rect 15485 11237 15519 11271
rect 15519 11237 15528 11271
rect 16028 11271 16080 11280
rect 15476 11228 15528 11237
rect 16028 11237 16037 11271
rect 16037 11237 16071 11271
rect 16071 11237 16080 11271
rect 16028 11228 16080 11237
rect 11428 11203 11480 11212
rect 11428 11169 11437 11203
rect 11437 11169 11471 11203
rect 11471 11169 11480 11203
rect 11428 11160 11480 11169
rect 10048 11135 10100 11144
rect 10048 11101 10057 11135
rect 10057 11101 10091 11135
rect 10091 11101 10100 11135
rect 10048 11092 10100 11101
rect 12164 11160 12216 11212
rect 12808 11160 12860 11212
rect 16856 11203 16908 11212
rect 16856 11169 16900 11203
rect 16900 11169 16908 11203
rect 16856 11160 16908 11169
rect 20 11024 72 11076
rect 2412 11024 2464 11076
rect 3884 11024 3936 11076
rect 4160 11024 4212 11076
rect 4712 11024 4764 11076
rect 2228 10956 2280 11008
rect 2780 10956 2832 11008
rect 4344 10999 4396 11008
rect 4344 10965 4353 10999
rect 4353 10965 4387 10999
rect 4387 10965 4396 10999
rect 4344 10956 4396 10965
rect 4896 10956 4948 11008
rect 6276 11024 6328 11076
rect 7564 11067 7616 11076
rect 7564 11033 7573 11067
rect 7573 11033 7607 11067
rect 7607 11033 7616 11067
rect 9956 11067 10008 11076
rect 7564 11024 7616 11033
rect 9956 11033 9965 11067
rect 9965 11033 9999 11067
rect 9999 11033 10008 11067
rect 9956 11024 10008 11033
rect 6000 10999 6052 11008
rect 6000 10965 6009 10999
rect 6009 10965 6043 10999
rect 6043 10965 6052 10999
rect 6000 10956 6052 10965
rect 7196 10956 7248 11008
rect 8760 10999 8812 11008
rect 8760 10965 8769 10999
rect 8769 10965 8803 10999
rect 8803 10965 8812 10999
rect 8760 10956 8812 10965
rect 13084 10956 13136 11008
rect 20260 10956 20312 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 1952 10752 2004 10804
rect 3884 10795 3936 10804
rect 3884 10761 3893 10795
rect 3893 10761 3927 10795
rect 3927 10761 3936 10795
rect 3884 10752 3936 10761
rect 2228 10727 2280 10736
rect 2228 10693 2252 10727
rect 2252 10693 2280 10727
rect 2228 10684 2280 10693
rect 2412 10659 2464 10668
rect 2412 10625 2421 10659
rect 2421 10625 2455 10659
rect 2455 10625 2464 10659
rect 2412 10616 2464 10625
rect 3332 10684 3384 10736
rect 7196 10752 7248 10804
rect 8760 10752 8812 10804
rect 9588 10752 9640 10804
rect 12164 10795 12216 10804
rect 12164 10761 12173 10795
rect 12173 10761 12207 10795
rect 12207 10761 12216 10795
rect 12164 10752 12216 10761
rect 14188 10795 14240 10804
rect 14188 10761 14197 10795
rect 14197 10761 14231 10795
rect 14231 10761 14240 10795
rect 14188 10752 14240 10761
rect 15384 10752 15436 10804
rect 15752 10752 15804 10804
rect 16856 10795 16908 10804
rect 16856 10761 16865 10795
rect 16865 10761 16899 10795
rect 16899 10761 16908 10795
rect 16856 10752 16908 10761
rect 25136 10752 25188 10804
rect 5172 10684 5224 10736
rect 6276 10727 6328 10736
rect 6276 10693 6285 10727
rect 6285 10693 6319 10727
rect 6319 10693 6328 10727
rect 6276 10684 6328 10693
rect 6644 10684 6696 10736
rect 6920 10684 6972 10736
rect 7472 10727 7524 10736
rect 7472 10693 7481 10727
rect 7481 10693 7515 10727
rect 7515 10693 7524 10727
rect 7472 10684 7524 10693
rect 7748 10684 7800 10736
rect 8852 10684 8904 10736
rect 14832 10684 14884 10736
rect 15476 10684 15528 10736
rect 4068 10548 4120 10600
rect 7012 10616 7064 10668
rect 10048 10616 10100 10668
rect 13268 10659 13320 10668
rect 13268 10625 13277 10659
rect 13277 10625 13311 10659
rect 13311 10625 13320 10659
rect 13268 10616 13320 10625
rect 7104 10548 7156 10600
rect 8668 10548 8720 10600
rect 11336 10591 11388 10600
rect 2044 10523 2096 10532
rect 2044 10489 2053 10523
rect 2053 10489 2087 10523
rect 2087 10489 2096 10523
rect 2044 10480 2096 10489
rect 6920 10480 6972 10532
rect 3332 10412 3384 10464
rect 3792 10412 3844 10464
rect 4620 10412 4672 10464
rect 5448 10412 5500 10464
rect 5540 10412 5592 10464
rect 7012 10455 7064 10464
rect 7012 10421 7021 10455
rect 7021 10421 7055 10455
rect 7055 10421 7064 10455
rect 7012 10412 7064 10421
rect 7840 10455 7892 10464
rect 7840 10421 7849 10455
rect 7849 10421 7883 10455
rect 7883 10421 7892 10455
rect 7840 10412 7892 10421
rect 11336 10557 11345 10591
rect 11345 10557 11379 10591
rect 11379 10557 11388 10591
rect 11336 10548 11388 10557
rect 24124 10548 24176 10600
rect 12624 10480 12676 10532
rect 10876 10412 10928 10464
rect 11428 10412 11480 10464
rect 12716 10412 12768 10464
rect 13084 10480 13136 10532
rect 14372 10523 14424 10532
rect 14372 10489 14381 10523
rect 14381 10489 14415 10523
rect 14415 10489 14424 10523
rect 14372 10480 14424 10489
rect 13452 10412 13504 10464
rect 14188 10412 14240 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 1584 10251 1636 10260
rect 1584 10217 1593 10251
rect 1593 10217 1627 10251
rect 1627 10217 1636 10251
rect 1584 10208 1636 10217
rect 2136 10208 2188 10260
rect 3332 10208 3384 10260
rect 5172 10251 5224 10260
rect 5172 10217 5181 10251
rect 5181 10217 5215 10251
rect 5215 10217 5224 10251
rect 5172 10208 5224 10217
rect 6828 10251 6880 10260
rect 6828 10217 6837 10251
rect 6837 10217 6871 10251
rect 6871 10217 6880 10251
rect 6828 10208 6880 10217
rect 2044 10140 2096 10192
rect 3700 10140 3752 10192
rect 1492 10072 1544 10124
rect 2412 10072 2464 10124
rect 2596 10115 2648 10124
rect 2596 10081 2605 10115
rect 2605 10081 2639 10115
rect 2639 10081 2648 10115
rect 2596 10072 2648 10081
rect 2780 10115 2832 10124
rect 2780 10081 2789 10115
rect 2789 10081 2823 10115
rect 2823 10081 2832 10115
rect 2780 10072 2832 10081
rect 4528 10115 4580 10124
rect 4528 10081 4537 10115
rect 4537 10081 4571 10115
rect 4571 10081 4580 10115
rect 4528 10072 4580 10081
rect 4620 10004 4672 10056
rect 5356 10072 5408 10124
rect 6000 10072 6052 10124
rect 5540 10004 5592 10056
rect 1584 9936 1636 9988
rect 5448 9936 5500 9988
rect 6736 9936 6788 9988
rect 7472 10208 7524 10260
rect 8760 10251 8812 10260
rect 8760 10217 8769 10251
rect 8769 10217 8803 10251
rect 8803 10217 8812 10251
rect 8760 10208 8812 10217
rect 12808 10208 12860 10260
rect 14372 10251 14424 10260
rect 14372 10217 14381 10251
rect 14381 10217 14415 10251
rect 14415 10217 14424 10251
rect 14372 10208 14424 10217
rect 7288 10140 7340 10192
rect 8668 10140 8720 10192
rect 9956 10140 10008 10192
rect 13452 10140 13504 10192
rect 14832 10140 14884 10192
rect 24216 10140 24268 10192
rect 10784 10072 10836 10124
rect 11612 10072 11664 10124
rect 7932 10004 7984 10056
rect 9404 10004 9456 10056
rect 10048 10047 10100 10056
rect 10048 10013 10057 10047
rect 10057 10013 10091 10047
rect 10091 10013 10100 10047
rect 10048 10004 10100 10013
rect 7656 9979 7708 9988
rect 7656 9945 7665 9979
rect 7665 9945 7699 9979
rect 7699 9945 7708 9979
rect 7656 9936 7708 9945
rect 11336 10004 11388 10056
rect 12624 10072 12676 10124
rect 12992 10004 13044 10056
rect 15568 10004 15620 10056
rect 13728 9979 13780 9988
rect 13728 9945 13737 9979
rect 13737 9945 13771 9979
rect 13771 9945 13780 9979
rect 13728 9936 13780 9945
rect 15292 9936 15344 9988
rect 24308 10004 24360 10056
rect 25044 10004 25096 10056
rect 24768 9979 24820 9988
rect 24768 9945 24777 9979
rect 24777 9945 24811 9979
rect 24811 9945 24820 9979
rect 24768 9936 24820 9945
rect 3792 9868 3844 9920
rect 5356 9868 5408 9920
rect 6368 9911 6420 9920
rect 6368 9877 6377 9911
rect 6377 9877 6411 9911
rect 6411 9877 6420 9911
rect 6368 9868 6420 9877
rect 6644 9868 6696 9920
rect 7472 9868 7524 9920
rect 8300 9868 8352 9920
rect 10784 9911 10836 9920
rect 10784 9877 10793 9911
rect 10793 9877 10827 9911
rect 10827 9877 10836 9911
rect 10784 9868 10836 9877
rect 12716 9911 12768 9920
rect 12716 9877 12725 9911
rect 12725 9877 12759 9911
rect 12759 9877 12768 9911
rect 12716 9868 12768 9877
rect 13544 9868 13596 9920
rect 14372 9868 14424 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 3700 9664 3752 9716
rect 4620 9707 4672 9716
rect 4620 9673 4629 9707
rect 4629 9673 4663 9707
rect 4663 9673 4672 9707
rect 4620 9664 4672 9673
rect 7564 9664 7616 9716
rect 10784 9664 10836 9716
rect 11612 9664 11664 9716
rect 13728 9664 13780 9716
rect 14832 9664 14884 9716
rect 15568 9664 15620 9716
rect 25044 9707 25096 9716
rect 25044 9673 25053 9707
rect 25053 9673 25087 9707
rect 25087 9673 25096 9707
rect 25044 9664 25096 9673
rect 3976 9596 4028 9648
rect 6644 9639 6696 9648
rect 4436 9528 4488 9580
rect 1584 9503 1636 9512
rect 1584 9469 1593 9503
rect 1593 9469 1627 9503
rect 1627 9469 1636 9503
rect 1584 9460 1636 9469
rect 3700 9503 3752 9512
rect 3700 9469 3709 9503
rect 3709 9469 3743 9503
rect 3743 9469 3752 9503
rect 3700 9460 3752 9469
rect 6644 9605 6653 9639
rect 6653 9605 6687 9639
rect 6687 9605 6696 9639
rect 6644 9596 6696 9605
rect 7748 9596 7800 9648
rect 12624 9596 12676 9648
rect 7012 9528 7064 9580
rect 12716 9528 12768 9580
rect 15292 9528 15344 9580
rect 24216 9528 24268 9580
rect 7656 9460 7708 9512
rect 8760 9503 8812 9512
rect 8760 9469 8769 9503
rect 8769 9469 8803 9503
rect 8803 9469 8812 9503
rect 8760 9460 8812 9469
rect 10692 9460 10744 9512
rect 12440 9503 12492 9512
rect 12440 9469 12449 9503
rect 12449 9469 12483 9503
rect 12483 9469 12492 9503
rect 12440 9460 12492 9469
rect 4344 9435 4396 9444
rect 4344 9401 4353 9435
rect 4353 9401 4387 9435
rect 4387 9401 4396 9435
rect 4344 9392 4396 9401
rect 2412 9367 2464 9376
rect 2412 9333 2421 9367
rect 2421 9333 2455 9367
rect 2455 9333 2464 9367
rect 2412 9324 2464 9333
rect 2780 9367 2832 9376
rect 2780 9333 2789 9367
rect 2789 9333 2823 9367
rect 2823 9333 2832 9367
rect 2780 9324 2832 9333
rect 3976 9324 4028 9376
rect 5356 9392 5408 9444
rect 7196 9435 7248 9444
rect 7196 9401 7205 9435
rect 7205 9401 7239 9435
rect 7239 9401 7248 9435
rect 7196 9392 7248 9401
rect 5448 9367 5500 9376
rect 5448 9333 5457 9367
rect 5457 9333 5491 9367
rect 5491 9333 5500 9367
rect 5448 9324 5500 9333
rect 7012 9367 7064 9376
rect 7012 9333 7021 9367
rect 7021 9333 7055 9367
rect 7055 9333 7064 9367
rect 7012 9324 7064 9333
rect 7656 9324 7708 9376
rect 8392 9324 8444 9376
rect 11980 9392 12032 9444
rect 13452 9392 13504 9444
rect 13912 9392 13964 9444
rect 15292 9435 15344 9444
rect 9772 9324 9824 9376
rect 9956 9367 10008 9376
rect 9956 9333 9965 9367
rect 9965 9333 9999 9367
rect 9999 9333 10008 9367
rect 9956 9324 10008 9333
rect 11428 9367 11480 9376
rect 11428 9333 11437 9367
rect 11437 9333 11471 9367
rect 11471 9333 11480 9367
rect 11428 9324 11480 9333
rect 13360 9367 13412 9376
rect 13360 9333 13369 9367
rect 13369 9333 13403 9367
rect 13403 9333 13412 9367
rect 13360 9324 13412 9333
rect 15292 9401 15301 9435
rect 15301 9401 15335 9435
rect 15335 9401 15344 9435
rect 15292 9392 15344 9401
rect 15936 9435 15988 9444
rect 15936 9401 15945 9435
rect 15945 9401 15979 9435
rect 15979 9401 15988 9435
rect 15936 9392 15988 9401
rect 16304 9324 16356 9376
rect 16764 9367 16816 9376
rect 16764 9333 16773 9367
rect 16773 9333 16807 9367
rect 16807 9333 16816 9367
rect 16764 9324 16816 9333
rect 24032 9324 24084 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 3148 9163 3200 9172
rect 3148 9129 3157 9163
rect 3157 9129 3191 9163
rect 3191 9129 3200 9163
rect 3148 9120 3200 9129
rect 3424 9163 3476 9172
rect 3424 9129 3433 9163
rect 3433 9129 3467 9163
rect 3467 9129 3476 9163
rect 3424 9120 3476 9129
rect 4344 9163 4396 9172
rect 4344 9129 4353 9163
rect 4353 9129 4387 9163
rect 4387 9129 4396 9163
rect 4344 9120 4396 9129
rect 6276 9163 6328 9172
rect 6276 9129 6285 9163
rect 6285 9129 6319 9163
rect 6319 9129 6328 9163
rect 6276 9120 6328 9129
rect 7288 9120 7340 9172
rect 4712 9052 4764 9104
rect 5080 9052 5132 9104
rect 1584 9027 1636 9036
rect 1584 8993 1593 9027
rect 1593 8993 1627 9027
rect 1627 8993 1636 9027
rect 1584 8984 1636 8993
rect 2964 9027 3016 9036
rect 2964 8993 2973 9027
rect 2973 8993 3007 9027
rect 3007 8993 3016 9027
rect 2964 8984 3016 8993
rect 4988 9027 5040 9036
rect 4988 8993 4997 9027
rect 4997 8993 5031 9027
rect 5031 8993 5040 9027
rect 4988 8984 5040 8993
rect 6828 9052 6880 9104
rect 7196 9052 7248 9104
rect 8576 9052 8628 9104
rect 8116 8984 8168 9036
rect 8300 8984 8352 9036
rect 8760 9027 8812 9036
rect 8760 8993 8769 9027
rect 8769 8993 8803 9027
rect 8803 8993 8812 9027
rect 13912 9163 13964 9172
rect 13912 9129 13921 9163
rect 13921 9129 13955 9163
rect 13955 9129 13964 9163
rect 13912 9120 13964 9129
rect 9772 9052 9824 9104
rect 10784 9052 10836 9104
rect 11612 9052 11664 9104
rect 12440 9052 12492 9104
rect 13452 9052 13504 9104
rect 15660 9095 15712 9104
rect 15660 9061 15669 9095
rect 15669 9061 15703 9095
rect 15703 9061 15712 9095
rect 15660 9052 15712 9061
rect 15936 9052 15988 9104
rect 24124 9052 24176 9104
rect 8760 8984 8812 8993
rect 11888 8984 11940 9036
rect 12992 9027 13044 9036
rect 12992 8993 13001 9027
rect 13001 8993 13035 9027
rect 13035 8993 13044 9027
rect 12992 8984 13044 8993
rect 17132 9027 17184 9036
rect 17132 8993 17150 9027
rect 17150 8993 17184 9027
rect 17132 8984 17184 8993
rect 24768 9027 24820 9036
rect 24768 8993 24777 9027
rect 24777 8993 24811 9027
rect 24811 8993 24820 9027
rect 24768 8984 24820 8993
rect 1492 8916 1544 8968
rect 4068 8916 4120 8968
rect 5080 8916 5132 8968
rect 2596 8848 2648 8900
rect 3700 8848 3752 8900
rect 5448 8848 5500 8900
rect 6276 8916 6328 8968
rect 7104 8916 7156 8968
rect 8208 8848 8260 8900
rect 9404 8891 9456 8900
rect 9404 8857 9413 8891
rect 9413 8857 9447 8891
rect 9447 8857 9456 8891
rect 9404 8848 9456 8857
rect 11612 8916 11664 8968
rect 16764 8916 16816 8968
rect 24860 8916 24912 8968
rect 10048 8848 10100 8900
rect 1676 8823 1728 8832
rect 1676 8789 1685 8823
rect 1685 8789 1719 8823
rect 1719 8789 1728 8823
rect 1676 8780 1728 8789
rect 5540 8780 5592 8832
rect 6552 8780 6604 8832
rect 6736 8823 6788 8832
rect 6736 8789 6745 8823
rect 6745 8789 6779 8823
rect 6779 8789 6788 8823
rect 6736 8780 6788 8789
rect 7104 8823 7156 8832
rect 7104 8789 7113 8823
rect 7113 8789 7147 8823
rect 7147 8789 7156 8823
rect 7104 8780 7156 8789
rect 9772 8780 9824 8832
rect 10692 8823 10744 8832
rect 10692 8789 10701 8823
rect 10701 8789 10735 8823
rect 10735 8789 10744 8823
rect 10692 8780 10744 8789
rect 14280 8823 14332 8832
rect 14280 8789 14289 8823
rect 14289 8789 14323 8823
rect 14323 8789 14332 8823
rect 14280 8780 14332 8789
rect 14372 8780 14424 8832
rect 17316 8780 17368 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 4712 8576 4764 8628
rect 5448 8619 5500 8628
rect 4160 8508 4212 8560
rect 5448 8585 5457 8619
rect 5457 8585 5491 8619
rect 5491 8585 5500 8619
rect 5448 8576 5500 8585
rect 6368 8576 6420 8628
rect 10048 8619 10100 8628
rect 10048 8585 10057 8619
rect 10057 8585 10091 8619
rect 10091 8585 10100 8619
rect 10048 8576 10100 8585
rect 11796 8576 11848 8628
rect 13452 8576 13504 8628
rect 16764 8619 16816 8628
rect 16764 8585 16773 8619
rect 16773 8585 16807 8619
rect 16807 8585 16816 8619
rect 16764 8576 16816 8585
rect 17132 8619 17184 8628
rect 17132 8585 17141 8619
rect 17141 8585 17175 8619
rect 17175 8585 17184 8619
rect 17132 8576 17184 8585
rect 5264 8508 5316 8560
rect 6644 8508 6696 8560
rect 7104 8508 7156 8560
rect 11244 8508 11296 8560
rect 11888 8508 11940 8560
rect 13268 8551 13320 8560
rect 13268 8517 13277 8551
rect 13277 8517 13311 8551
rect 13311 8517 13320 8551
rect 13268 8508 13320 8517
rect 24768 8551 24820 8560
rect 24768 8517 24777 8551
rect 24777 8517 24811 8551
rect 24811 8517 24820 8551
rect 24768 8508 24820 8517
rect 5540 8483 5592 8492
rect 1676 8372 1728 8424
rect 1768 8415 1820 8424
rect 1768 8381 1777 8415
rect 1777 8381 1811 8415
rect 1811 8381 1820 8415
rect 2412 8415 2464 8424
rect 1768 8372 1820 8381
rect 2412 8381 2421 8415
rect 2421 8381 2455 8415
rect 2455 8381 2464 8415
rect 2412 8372 2464 8381
rect 5540 8449 5549 8483
rect 5549 8449 5583 8483
rect 5583 8449 5592 8483
rect 5540 8440 5592 8449
rect 7932 8440 7984 8492
rect 9772 8483 9824 8492
rect 9772 8449 9781 8483
rect 9781 8449 9815 8483
rect 9815 8449 9824 8483
rect 9772 8440 9824 8449
rect 15292 8440 15344 8492
rect 15660 8440 15712 8492
rect 3884 8304 3936 8356
rect 2964 8279 3016 8288
rect 2964 8245 2973 8279
rect 2973 8245 3007 8279
rect 3007 8245 3016 8279
rect 4068 8372 4120 8424
rect 4528 8372 4580 8424
rect 5356 8415 5408 8424
rect 5356 8381 5362 8415
rect 5362 8381 5408 8415
rect 5356 8372 5408 8381
rect 7288 8415 7340 8424
rect 7288 8381 7297 8415
rect 7297 8381 7331 8415
rect 7331 8381 7340 8415
rect 7288 8372 7340 8381
rect 7840 8415 7892 8424
rect 7840 8381 7849 8415
rect 7849 8381 7883 8415
rect 7883 8381 7892 8415
rect 7840 8372 7892 8381
rect 9128 8415 9180 8424
rect 9128 8381 9137 8415
rect 9137 8381 9171 8415
rect 9171 8381 9180 8415
rect 9128 8372 9180 8381
rect 9496 8415 9548 8424
rect 9496 8381 9505 8415
rect 9505 8381 9539 8415
rect 9539 8381 9548 8415
rect 9496 8372 9548 8381
rect 16304 8415 16356 8424
rect 4436 8304 4488 8356
rect 5632 8304 5684 8356
rect 8024 8347 8076 8356
rect 8024 8313 8033 8347
rect 8033 8313 8067 8347
rect 8067 8313 8076 8347
rect 8024 8304 8076 8313
rect 10048 8304 10100 8356
rect 16304 8381 16313 8415
rect 16313 8381 16347 8415
rect 16347 8381 16356 8415
rect 16304 8372 16356 8381
rect 24124 8372 24176 8424
rect 11336 8347 11388 8356
rect 11336 8313 11345 8347
rect 11345 8313 11379 8347
rect 11379 8313 11388 8347
rect 11336 8304 11388 8313
rect 12716 8347 12768 8356
rect 12716 8313 12725 8347
rect 12725 8313 12759 8347
rect 12759 8313 12768 8347
rect 12716 8304 12768 8313
rect 13360 8304 13412 8356
rect 14280 8347 14332 8356
rect 14280 8313 14289 8347
rect 14289 8313 14323 8347
rect 14323 8313 14332 8347
rect 14280 8304 14332 8313
rect 2964 8236 3016 8245
rect 4988 8279 5040 8288
rect 4988 8245 4997 8279
rect 4997 8245 5031 8279
rect 5031 8245 5040 8279
rect 4988 8236 5040 8245
rect 6552 8279 6604 8288
rect 6552 8245 6561 8279
rect 6561 8245 6595 8279
rect 6595 8245 6604 8279
rect 6552 8236 6604 8245
rect 8116 8236 8168 8288
rect 9680 8236 9732 8288
rect 14464 8304 14516 8356
rect 24032 8279 24084 8288
rect 24032 8245 24041 8279
rect 24041 8245 24075 8279
rect 24075 8245 24084 8279
rect 24032 8236 24084 8245
rect 24860 8236 24912 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 1676 8032 1728 8084
rect 2872 8032 2924 8084
rect 4528 8075 4580 8084
rect 4528 8041 4537 8075
rect 4537 8041 4571 8075
rect 4571 8041 4580 8075
rect 4528 8032 4580 8041
rect 5448 8032 5500 8084
rect 8208 8032 8260 8084
rect 8300 8032 8352 8084
rect 9496 8032 9548 8084
rect 9864 8032 9916 8084
rect 11336 8032 11388 8084
rect 12992 8032 13044 8084
rect 14556 8075 14608 8084
rect 14556 8041 14565 8075
rect 14565 8041 14599 8075
rect 14599 8041 14608 8075
rect 14556 8032 14608 8041
rect 16304 8075 16356 8084
rect 16304 8041 16313 8075
rect 16313 8041 16347 8075
rect 16347 8041 16356 8075
rect 16304 8032 16356 8041
rect 8944 7964 8996 8016
rect 9128 7964 9180 8016
rect 112 7896 164 7948
rect 2136 7896 2188 7948
rect 2964 7939 3016 7948
rect 2964 7905 2973 7939
rect 2973 7905 3007 7939
rect 3007 7905 3016 7939
rect 2964 7896 3016 7905
rect 4988 7939 5040 7948
rect 4988 7905 4997 7939
rect 4997 7905 5031 7939
rect 5031 7905 5040 7939
rect 4988 7896 5040 7905
rect 5632 7896 5684 7948
rect 6828 7896 6880 7948
rect 7288 7896 7340 7948
rect 7472 7896 7524 7948
rect 7840 7896 7892 7948
rect 9772 7939 9824 7948
rect 9772 7905 9781 7939
rect 9781 7905 9815 7939
rect 9815 7905 9824 7939
rect 9772 7896 9824 7905
rect 10048 7896 10100 7948
rect 11980 7964 12032 8016
rect 13084 8007 13136 8016
rect 13084 7973 13093 8007
rect 13093 7973 13127 8007
rect 13127 7973 13136 8007
rect 13084 7964 13136 7973
rect 14464 7964 14516 8016
rect 13360 7939 13412 7948
rect 13360 7905 13369 7939
rect 13369 7905 13403 7939
rect 13403 7905 13412 7939
rect 13360 7896 13412 7905
rect 14832 7896 14884 7948
rect 15384 7939 15436 7948
rect 15384 7905 15393 7939
rect 15393 7905 15427 7939
rect 15427 7905 15436 7939
rect 15384 7896 15436 7905
rect 8484 7828 8536 7880
rect 10508 7871 10560 7880
rect 10508 7837 10517 7871
rect 10517 7837 10551 7871
rect 10551 7837 10560 7871
rect 10508 7828 10560 7837
rect 5540 7760 5592 7812
rect 6184 7760 6236 7812
rect 8116 7760 8168 7812
rect 1032 7692 1084 7744
rect 1584 7692 1636 7744
rect 6276 7692 6328 7744
rect 13176 7692 13228 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 1492 7488 1544 7540
rect 2136 7531 2188 7540
rect 2136 7497 2145 7531
rect 2145 7497 2179 7531
rect 2179 7497 2188 7531
rect 2136 7488 2188 7497
rect 2964 7531 3016 7540
rect 2964 7497 2973 7531
rect 2973 7497 3007 7531
rect 3007 7497 3016 7531
rect 2964 7488 3016 7497
rect 3792 7488 3844 7540
rect 4896 7488 4948 7540
rect 5356 7488 5408 7540
rect 8300 7488 8352 7540
rect 9772 7531 9824 7540
rect 9772 7497 9781 7531
rect 9781 7497 9815 7531
rect 9815 7497 9824 7531
rect 9772 7488 9824 7497
rect 10048 7488 10100 7540
rect 11980 7488 12032 7540
rect 13360 7488 13412 7540
rect 15384 7531 15436 7540
rect 15384 7497 15393 7531
rect 15393 7497 15427 7531
rect 15427 7497 15436 7531
rect 15384 7488 15436 7497
rect 24860 7488 24912 7540
rect 5080 7352 5132 7404
rect 3884 7327 3936 7336
rect 3884 7293 3893 7327
rect 3893 7293 3927 7327
rect 3927 7293 3936 7327
rect 3884 7284 3936 7293
rect 6920 7352 6972 7404
rect 4620 7216 4672 7268
rect 4988 7216 5040 7268
rect 6460 7148 6512 7200
rect 7288 7284 7340 7336
rect 10508 7352 10560 7404
rect 12440 7395 12492 7404
rect 12440 7361 12449 7395
rect 12449 7361 12483 7395
rect 12483 7361 12492 7395
rect 12440 7352 12492 7361
rect 14372 7352 14424 7404
rect 14556 7395 14608 7404
rect 14556 7361 14565 7395
rect 14565 7361 14599 7395
rect 14599 7361 14608 7395
rect 14556 7352 14608 7361
rect 7932 7284 7984 7336
rect 7472 7216 7524 7268
rect 8760 7259 8812 7268
rect 8760 7225 8769 7259
rect 8769 7225 8803 7259
rect 8803 7225 8812 7259
rect 8760 7216 8812 7225
rect 8852 7259 8904 7268
rect 8852 7225 8861 7259
rect 8861 7225 8895 7259
rect 8895 7225 8904 7259
rect 9404 7259 9456 7268
rect 8852 7216 8904 7225
rect 9404 7225 9413 7259
rect 9413 7225 9447 7259
rect 9447 7225 9456 7259
rect 9404 7216 9456 7225
rect 7564 7148 7616 7200
rect 9312 7148 9364 7200
rect 10876 7284 10928 7336
rect 11244 7327 11296 7336
rect 11244 7293 11253 7327
rect 11253 7293 11287 7327
rect 11287 7293 11296 7327
rect 11244 7284 11296 7293
rect 11980 7284 12032 7336
rect 12256 7216 12308 7268
rect 13360 7191 13412 7200
rect 13360 7157 13369 7191
rect 13369 7157 13403 7191
rect 13403 7157 13412 7191
rect 13360 7148 13412 7157
rect 14648 7216 14700 7268
rect 25136 7191 25188 7200
rect 25136 7157 25145 7191
rect 25145 7157 25179 7191
rect 25179 7157 25188 7191
rect 25136 7148 25188 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 1400 6944 1452 6996
rect 4804 6987 4856 6996
rect 4804 6953 4813 6987
rect 4813 6953 4847 6987
rect 4847 6953 4856 6987
rect 4804 6944 4856 6953
rect 6460 6944 6512 6996
rect 6920 6944 6972 6996
rect 7840 6944 7892 6996
rect 8208 6987 8260 6996
rect 8208 6953 8217 6987
rect 8217 6953 8251 6987
rect 8251 6953 8260 6987
rect 8208 6944 8260 6953
rect 8760 6944 8812 6996
rect 9956 6987 10008 6996
rect 9956 6953 9965 6987
rect 9965 6953 9999 6987
rect 9999 6953 10008 6987
rect 9956 6944 10008 6953
rect 11244 6944 11296 6996
rect 12440 6987 12492 6996
rect 12440 6953 12449 6987
rect 12449 6953 12483 6987
rect 12483 6953 12492 6987
rect 12440 6944 12492 6953
rect 12716 6944 12768 6996
rect 13360 6876 13412 6928
rect 13820 6919 13872 6928
rect 13820 6885 13829 6919
rect 13829 6885 13863 6919
rect 13863 6885 13872 6919
rect 13820 6876 13872 6885
rect 2688 6808 2740 6860
rect 4620 6851 4672 6860
rect 4620 6817 4629 6851
rect 4629 6817 4663 6851
rect 4663 6817 4672 6851
rect 4620 6808 4672 6817
rect 6184 6808 6236 6860
rect 9864 6851 9916 6860
rect 9864 6817 9873 6851
rect 9873 6817 9907 6851
rect 9907 6817 9916 6851
rect 9864 6808 9916 6817
rect 11336 6851 11388 6860
rect 11336 6817 11345 6851
rect 11345 6817 11379 6851
rect 11379 6817 11388 6851
rect 11336 6808 11388 6817
rect 8024 6740 8076 6792
rect 11244 6783 11296 6792
rect 11244 6749 11253 6783
rect 11253 6749 11287 6783
rect 11287 6749 11296 6783
rect 11244 6740 11296 6749
rect 13728 6783 13780 6792
rect 13728 6749 13737 6783
rect 13737 6749 13771 6783
rect 13771 6749 13780 6783
rect 13728 6740 13780 6749
rect 6276 6715 6328 6724
rect 6276 6681 6285 6715
rect 6285 6681 6319 6715
rect 6319 6681 6328 6715
rect 6276 6672 6328 6681
rect 13452 6715 13504 6724
rect 13452 6681 13461 6715
rect 13461 6681 13495 6715
rect 13495 6681 13504 6715
rect 14556 6876 14608 6928
rect 14648 6876 14700 6928
rect 15936 6851 15988 6860
rect 15936 6817 15945 6851
rect 15945 6817 15979 6851
rect 15979 6817 15988 6851
rect 15936 6808 15988 6817
rect 13452 6672 13504 6681
rect 8300 6604 8352 6656
rect 8852 6604 8904 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 2688 6400 2740 6452
rect 6184 6443 6236 6452
rect 6184 6409 6193 6443
rect 6193 6409 6227 6443
rect 6227 6409 6236 6443
rect 6184 6400 6236 6409
rect 9864 6400 9916 6452
rect 11336 6443 11388 6452
rect 11336 6409 11345 6443
rect 11345 6409 11379 6443
rect 11379 6409 11388 6443
rect 11336 6400 11388 6409
rect 13176 6443 13228 6452
rect 13176 6409 13185 6443
rect 13185 6409 13219 6443
rect 13219 6409 13228 6443
rect 13176 6400 13228 6409
rect 13820 6400 13872 6452
rect 15936 6443 15988 6452
rect 15936 6409 15945 6443
rect 15945 6409 15979 6443
rect 15979 6409 15988 6443
rect 15936 6400 15988 6409
rect 3240 6332 3292 6384
rect 9312 6332 9364 6384
rect 9496 6332 9548 6384
rect 11152 6332 11204 6384
rect 112 6128 164 6180
rect 8300 6196 8352 6248
rect 8484 6239 8536 6248
rect 8484 6205 8493 6239
rect 8493 6205 8527 6239
rect 8527 6205 8536 6239
rect 8484 6196 8536 6205
rect 9772 6239 9824 6248
rect 9772 6205 9781 6239
rect 9781 6205 9815 6239
rect 9815 6205 9824 6239
rect 9772 6196 9824 6205
rect 4620 6103 4672 6112
rect 4620 6069 4629 6103
rect 4629 6069 4663 6103
rect 4663 6069 4672 6103
rect 4620 6060 4672 6069
rect 8300 6103 8352 6112
rect 8300 6069 8309 6103
rect 8309 6069 8343 6103
rect 8343 6069 8352 6103
rect 8300 6060 8352 6069
rect 10784 6264 10836 6316
rect 13452 6307 13504 6316
rect 13452 6273 13461 6307
rect 13461 6273 13495 6307
rect 13495 6273 13504 6307
rect 13452 6264 13504 6273
rect 14648 6264 14700 6316
rect 13176 6128 13228 6180
rect 14740 6128 14792 6180
rect 15016 6171 15068 6180
rect 15016 6137 15025 6171
rect 15025 6137 15059 6171
rect 15059 6137 15068 6171
rect 15016 6128 15068 6137
rect 15108 6171 15160 6180
rect 15108 6137 15117 6171
rect 15117 6137 15151 6171
rect 15151 6137 15160 6171
rect 15108 6128 15160 6137
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 7012 5856 7064 5908
rect 8484 5856 8536 5908
rect 13728 5899 13780 5908
rect 13728 5865 13737 5899
rect 13737 5865 13771 5899
rect 13771 5865 13780 5899
rect 13728 5856 13780 5865
rect 9864 5831 9916 5840
rect 9864 5797 9873 5831
rect 9873 5797 9907 5831
rect 9907 5797 9916 5831
rect 9864 5788 9916 5797
rect 10232 5788 10284 5840
rect 11980 5788 12032 5840
rect 12992 5788 13044 5840
rect 15108 5788 15160 5840
rect 5172 5720 5224 5772
rect 6000 5763 6052 5772
rect 6000 5729 6009 5763
rect 6009 5729 6043 5763
rect 6043 5729 6052 5763
rect 6000 5720 6052 5729
rect 7472 5763 7524 5772
rect 7472 5729 7481 5763
rect 7481 5729 7515 5763
rect 7515 5729 7524 5763
rect 7472 5720 7524 5729
rect 7932 5763 7984 5772
rect 7932 5729 7941 5763
rect 7941 5729 7975 5763
rect 7975 5729 7984 5763
rect 7932 5720 7984 5729
rect 8024 5720 8076 5772
rect 12256 5763 12308 5772
rect 12256 5729 12265 5763
rect 12265 5729 12299 5763
rect 12299 5729 12308 5763
rect 12256 5720 12308 5729
rect 14648 5720 14700 5772
rect 14740 5720 14792 5772
rect 16028 5720 16080 5772
rect 8208 5695 8260 5704
rect 8208 5661 8217 5695
rect 8217 5661 8251 5695
rect 8251 5661 8260 5695
rect 8208 5652 8260 5661
rect 9404 5652 9456 5704
rect 10508 5652 10560 5704
rect 12532 5652 12584 5704
rect 15016 5652 15068 5704
rect 13728 5584 13780 5636
rect 15476 5584 15528 5636
rect 10784 5559 10836 5568
rect 10784 5525 10793 5559
rect 10793 5525 10827 5559
rect 10827 5525 10836 5559
rect 10784 5516 10836 5525
rect 13176 5559 13228 5568
rect 13176 5525 13185 5559
rect 13185 5525 13219 5559
rect 13219 5525 13228 5559
rect 13176 5516 13228 5525
rect 14372 5516 14424 5568
rect 14556 5559 14608 5568
rect 14556 5525 14565 5559
rect 14565 5525 14599 5559
rect 14599 5525 14608 5559
rect 14556 5516 14608 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 6000 5355 6052 5364
rect 6000 5321 6009 5355
rect 6009 5321 6043 5355
rect 6043 5321 6052 5355
rect 6000 5312 6052 5321
rect 6552 5312 6604 5364
rect 9864 5312 9916 5364
rect 11152 5355 11204 5364
rect 11152 5321 11161 5355
rect 11161 5321 11195 5355
rect 11195 5321 11204 5355
rect 11152 5312 11204 5321
rect 12256 5355 12308 5364
rect 12256 5321 12265 5355
rect 12265 5321 12299 5355
rect 12299 5321 12308 5355
rect 12256 5312 12308 5321
rect 12992 5355 13044 5364
rect 12992 5321 13001 5355
rect 13001 5321 13035 5355
rect 13035 5321 13044 5355
rect 12992 5312 13044 5321
rect 13176 5312 13228 5364
rect 13820 5312 13872 5364
rect 13912 5312 13964 5364
rect 12716 5244 12768 5296
rect 14004 5244 14056 5296
rect 14648 5287 14700 5296
rect 14648 5253 14657 5287
rect 14657 5253 14691 5287
rect 14691 5253 14700 5287
rect 14648 5244 14700 5253
rect 15476 5287 15528 5296
rect 15476 5253 15485 5287
rect 15485 5253 15519 5287
rect 15519 5253 15528 5287
rect 15476 5244 15528 5253
rect 16028 5287 16080 5296
rect 16028 5253 16037 5287
rect 16037 5253 16071 5287
rect 16071 5253 16080 5287
rect 16028 5244 16080 5253
rect 8208 5176 8260 5228
rect 10232 5219 10284 5228
rect 10232 5185 10241 5219
rect 10241 5185 10275 5219
rect 10275 5185 10284 5219
rect 10232 5176 10284 5185
rect 10508 5219 10560 5228
rect 10508 5185 10517 5219
rect 10517 5185 10551 5219
rect 10551 5185 10560 5219
rect 10508 5176 10560 5185
rect 12532 5219 12584 5228
rect 12532 5185 12541 5219
rect 12541 5185 12575 5219
rect 12575 5185 12584 5219
rect 12532 5176 12584 5185
rect 7656 5015 7708 5024
rect 7656 4981 7665 5015
rect 7665 4981 7699 5015
rect 7699 4981 7708 5015
rect 7656 4972 7708 4981
rect 8300 5015 8352 5024
rect 8300 4981 8309 5015
rect 8309 4981 8343 5015
rect 8343 4981 8352 5015
rect 11244 5040 11296 5092
rect 9312 5015 9364 5024
rect 8300 4972 8352 4981
rect 9312 4981 9321 5015
rect 9321 4981 9355 5015
rect 9355 4981 9364 5015
rect 9312 4972 9364 4981
rect 13820 5083 13872 5092
rect 13820 5049 13829 5083
rect 13829 5049 13863 5083
rect 13863 5049 13872 5083
rect 13820 5040 13872 5049
rect 17500 5040 17552 5092
rect 14556 4972 14608 5024
rect 23756 4972 23808 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 7472 4811 7524 4820
rect 7472 4777 7481 4811
rect 7481 4777 7515 4811
rect 7515 4777 7524 4811
rect 7472 4768 7524 4777
rect 7932 4811 7984 4820
rect 7932 4777 7941 4811
rect 7941 4777 7975 4811
rect 7975 4777 7984 4811
rect 7932 4768 7984 4777
rect 8208 4768 8260 4820
rect 10140 4811 10192 4820
rect 10140 4777 10149 4811
rect 10149 4777 10183 4811
rect 10183 4777 10192 4811
rect 10140 4768 10192 4777
rect 23664 4768 23716 4820
rect 10692 4700 10744 4752
rect 13820 4743 13872 4752
rect 13820 4709 13829 4743
rect 13829 4709 13863 4743
rect 13863 4709 13872 4743
rect 13820 4700 13872 4709
rect 11428 4675 11480 4684
rect 11428 4641 11437 4675
rect 11437 4641 11471 4675
rect 11471 4641 11480 4675
rect 11428 4632 11480 4641
rect 14372 4632 14424 4684
rect 15292 4675 15344 4684
rect 15292 4641 15301 4675
rect 15301 4641 15335 4675
rect 15335 4641 15344 4675
rect 15292 4632 15344 4641
rect 23940 4632 23992 4684
rect 13728 4607 13780 4616
rect 13728 4573 13737 4607
rect 13737 4573 13771 4607
rect 13771 4573 13780 4607
rect 13728 4564 13780 4573
rect 14004 4607 14056 4616
rect 14004 4573 14013 4607
rect 14013 4573 14047 4607
rect 14047 4573 14056 4607
rect 14004 4564 14056 4573
rect 12900 4428 12952 4480
rect 14832 4428 14884 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 7564 4267 7616 4276
rect 7564 4233 7573 4267
rect 7573 4233 7607 4267
rect 7607 4233 7616 4267
rect 7564 4224 7616 4233
rect 10692 4224 10744 4276
rect 11428 4267 11480 4276
rect 11428 4233 11437 4267
rect 11437 4233 11471 4267
rect 11471 4233 11480 4267
rect 11428 4224 11480 4233
rect 13176 4267 13228 4276
rect 13176 4233 13185 4267
rect 13185 4233 13219 4267
rect 13219 4233 13228 4267
rect 13176 4224 13228 4233
rect 15292 4267 15344 4276
rect 15292 4233 15301 4267
rect 15301 4233 15335 4267
rect 15335 4233 15344 4267
rect 15292 4224 15344 4233
rect 2504 3884 2556 3936
rect 8300 3952 8352 4004
rect 9864 3995 9916 4004
rect 9864 3961 9873 3995
rect 9873 3961 9907 3995
rect 9907 3961 9916 3995
rect 9864 3952 9916 3961
rect 13176 4020 13228 4072
rect 13820 3952 13872 4004
rect 9036 3927 9088 3936
rect 9036 3893 9045 3927
rect 9045 3893 9079 3927
rect 9079 3893 9088 3927
rect 9036 3884 9088 3893
rect 9312 3884 9364 3936
rect 9956 3884 10008 3936
rect 23940 3927 23992 3936
rect 23940 3893 23949 3927
rect 23949 3893 23983 3927
rect 23983 3893 23992 3927
rect 23940 3884 23992 3893
rect 24032 3884 24084 3936
rect 27620 3884 27672 3936
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 13728 3723 13780 3732
rect 13728 3689 13737 3723
rect 13737 3689 13771 3723
rect 13771 3689 13780 3723
rect 13728 3680 13780 3689
rect 9864 3612 9916 3664
rect 9036 3544 9088 3596
rect 8024 3519 8076 3528
rect 8024 3485 8033 3519
rect 8033 3485 8067 3519
rect 8067 3485 8076 3519
rect 8024 3476 8076 3485
rect 9220 3476 9272 3528
rect 10416 3451 10468 3460
rect 10416 3417 10425 3451
rect 10425 3417 10459 3451
rect 10459 3417 10468 3451
rect 10416 3408 10468 3417
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 8024 3179 8076 3188
rect 8024 3145 8033 3179
rect 8033 3145 8067 3179
rect 8067 3145 8076 3179
rect 8024 3136 8076 3145
rect 9220 3179 9272 3188
rect 9220 3145 9229 3179
rect 9229 3145 9263 3179
rect 9263 3145 9272 3179
rect 9220 3136 9272 3145
rect 9864 3136 9916 3188
rect 9956 3068 10008 3120
rect 9036 3000 9088 3052
rect 10416 3043 10468 3052
rect 10416 3009 10425 3043
rect 10425 3009 10459 3043
rect 10459 3009 10468 3043
rect 10416 3000 10468 3009
rect 8208 2907 8260 2916
rect 8208 2873 8217 2907
rect 8217 2873 8251 2907
rect 8251 2873 8260 2907
rect 8208 2864 8260 2873
rect 8024 2796 8076 2848
rect 9956 2864 10008 2916
rect 18788 2864 18840 2916
rect 10140 2796 10192 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 6092 2592 6144 2644
rect 7288 2592 7340 2644
rect 8208 2592 8260 2644
rect 11520 2592 11572 2644
rect 13544 2592 13596 2644
rect 23940 2592 23992 2644
rect 25228 2592 25280 2644
rect 9036 2524 9088 2576
rect 19248 2524 19300 2576
rect 7196 2456 7248 2508
rect 5540 2252 5592 2304
rect 11796 2456 11848 2508
rect 18788 2499 18840 2508
rect 9864 2431 9916 2440
rect 9864 2397 9873 2431
rect 9873 2397 9907 2431
rect 9907 2397 9916 2431
rect 9864 2388 9916 2397
rect 10140 2431 10192 2440
rect 10140 2397 10149 2431
rect 10149 2397 10183 2431
rect 10183 2397 10192 2431
rect 10140 2388 10192 2397
rect 10324 2388 10376 2440
rect 18788 2465 18797 2499
rect 18797 2465 18831 2499
rect 18831 2465 18840 2499
rect 18788 2456 18840 2465
rect 22560 2320 22612 2372
rect 8576 2252 8628 2304
rect 11796 2295 11848 2304
rect 11796 2261 11805 2295
rect 11805 2261 11839 2295
rect 11839 2261 11848 2295
rect 11796 2252 11848 2261
rect 20628 2252 20680 2304
rect 20720 2252 20772 2304
rect 26884 2252 26936 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
<< metal2 >>
rect 754 27520 810 28000
rect 2318 27554 2374 28000
rect 2318 27526 2544 27554
rect 2318 27520 2374 27526
rect 768 27130 796 27520
rect 20 27124 72 27130
rect 20 27066 72 27072
rect 756 27124 808 27130
rect 756 27066 808 27072
rect 32 11082 60 27066
rect 1490 26616 1546 26625
rect 1490 26551 1546 26560
rect 1400 23180 1452 23186
rect 1400 23122 1452 23128
rect 1412 22506 1440 23122
rect 1400 22500 1452 22506
rect 1400 22442 1452 22448
rect 1504 22098 1532 26551
rect 1582 24848 1638 24857
rect 1582 24783 1638 24792
rect 1596 23322 1624 24783
rect 2516 23866 2544 27526
rect 3974 27520 4030 28000
rect 5630 27554 5686 28000
rect 7286 27554 7342 28000
rect 5630 27526 6040 27554
rect 5630 27520 5686 27526
rect 2504 23860 2556 23866
rect 2504 23802 2556 23808
rect 2516 23662 2544 23802
rect 2504 23656 2556 23662
rect 2504 23598 2556 23604
rect 3988 23322 4016 27520
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 6012 23594 6040 27526
rect 7024 27526 7342 27554
rect 7024 24274 7052 27526
rect 7286 27520 7342 27526
rect 8942 27520 8998 28000
rect 10598 27520 10654 28000
rect 12254 27520 12310 28000
rect 13910 27520 13966 28000
rect 15474 27520 15530 28000
rect 17130 27520 17186 28000
rect 18786 27520 18842 28000
rect 20442 27520 20498 28000
rect 22098 27520 22154 28000
rect 23754 27520 23810 28000
rect 25410 27520 25466 28000
rect 27066 27520 27122 28000
rect 6276 24268 6328 24274
rect 6276 24210 6328 24216
rect 7012 24268 7064 24274
rect 7012 24210 7064 24216
rect 8208 24268 8260 24274
rect 8208 24210 8260 24216
rect 6288 23866 6316 24210
rect 6736 24064 6788 24070
rect 6736 24006 6788 24012
rect 6828 24064 6880 24070
rect 6828 24006 6880 24012
rect 6276 23860 6328 23866
rect 6276 23802 6328 23808
rect 6000 23588 6052 23594
rect 6000 23530 6052 23536
rect 6644 23520 6696 23526
rect 6644 23462 6696 23468
rect 1584 23316 1636 23322
rect 1584 23258 1636 23264
rect 3976 23316 4028 23322
rect 3976 23258 4028 23264
rect 2504 23180 2556 23186
rect 2504 23122 2556 23128
rect 2516 22438 2544 23122
rect 6552 23112 6604 23118
rect 6552 23054 6604 23060
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 6564 22778 6592 23054
rect 6552 22772 6604 22778
rect 6552 22714 6604 22720
rect 2780 22568 2832 22574
rect 2780 22510 2832 22516
rect 2792 22438 2820 22510
rect 3332 22500 3384 22506
rect 3332 22442 3384 22448
rect 2504 22432 2556 22438
rect 2504 22374 2556 22380
rect 2780 22432 2832 22438
rect 2780 22374 2832 22380
rect 3240 22432 3292 22438
rect 3240 22374 3292 22380
rect 2516 22234 2544 22374
rect 2504 22228 2556 22234
rect 2504 22170 2556 22176
rect 1492 22092 1544 22098
rect 1492 22034 1544 22040
rect 1504 21690 1532 22034
rect 1860 21888 1912 21894
rect 1860 21830 1912 21836
rect 1952 21888 2004 21894
rect 1952 21830 2004 21836
rect 1492 21684 1544 21690
rect 1492 21626 1544 21632
rect 1872 21400 1900 21830
rect 1964 21554 1992 21830
rect 1952 21548 2004 21554
rect 1952 21490 2004 21496
rect 1952 21412 2004 21418
rect 1872 21372 1952 21400
rect 1952 21354 2004 21360
rect 2688 21412 2740 21418
rect 2688 21354 2740 21360
rect 1122 21312 1178 21321
rect 1122 21247 1178 21256
rect 1136 20398 1164 21247
rect 1124 20392 1176 20398
rect 1124 20334 1176 20340
rect 1964 19990 1992 21354
rect 2700 21078 2728 21354
rect 2320 21072 2372 21078
rect 2320 21014 2372 21020
rect 2688 21072 2740 21078
rect 2688 21014 2740 21020
rect 2044 20936 2096 20942
rect 2044 20878 2096 20884
rect 2056 20602 2084 20878
rect 2044 20596 2096 20602
rect 2044 20538 2096 20544
rect 2056 20058 2084 20538
rect 2332 20262 2360 21014
rect 2700 20466 2728 21014
rect 2688 20460 2740 20466
rect 2688 20402 2740 20408
rect 2320 20256 2372 20262
rect 2320 20198 2372 20204
rect 2044 20052 2096 20058
rect 2044 19994 2096 20000
rect 1952 19984 2004 19990
rect 1952 19926 2004 19932
rect 2332 19922 2360 20198
rect 2700 20058 2728 20402
rect 2792 20330 2820 22374
rect 3056 22092 3108 22098
rect 3056 22034 3108 22040
rect 3068 21554 3096 22034
rect 3252 21690 3280 22374
rect 3344 22234 3372 22442
rect 3332 22228 3384 22234
rect 3332 22170 3384 22176
rect 4436 22092 4488 22098
rect 4436 22034 4488 22040
rect 4448 21690 4476 22034
rect 5080 22024 5132 22030
rect 5080 21966 5132 21972
rect 3240 21684 3292 21690
rect 3240 21626 3292 21632
rect 4436 21684 4488 21690
rect 4436 21626 4488 21632
rect 3056 21548 3108 21554
rect 3056 21490 3108 21496
rect 3068 21350 3096 21490
rect 3252 21350 3280 21626
rect 3516 21412 3568 21418
rect 3516 21354 3568 21360
rect 3056 21344 3108 21350
rect 3056 21286 3108 21292
rect 3240 21344 3292 21350
rect 3240 21286 3292 21292
rect 3068 20466 3096 21286
rect 3528 21146 3556 21354
rect 3516 21140 3568 21146
rect 3516 21082 3568 21088
rect 4448 20534 4476 21626
rect 4988 21412 5040 21418
rect 4988 21354 5040 21360
rect 4896 21344 4948 21350
rect 4896 21286 4948 21292
rect 4436 20528 4488 20534
rect 4436 20470 4488 20476
rect 3056 20460 3108 20466
rect 3056 20402 3108 20408
rect 4620 20460 4672 20466
rect 4620 20402 4672 20408
rect 2780 20324 2832 20330
rect 2780 20266 2832 20272
rect 3056 20324 3108 20330
rect 3056 20266 3108 20272
rect 2688 20052 2740 20058
rect 2688 19994 2740 20000
rect 2320 19916 2372 19922
rect 2320 19858 2372 19864
rect 1306 19544 1362 19553
rect 1306 19479 1362 19488
rect 112 18420 164 18426
rect 112 18362 164 18368
rect 124 18329 152 18362
rect 110 18320 166 18329
rect 110 18255 166 18264
rect 1320 17746 1348 19479
rect 2332 19174 2360 19858
rect 2320 19168 2372 19174
rect 2320 19110 2372 19116
rect 1400 18828 1452 18834
rect 1400 18770 1452 18776
rect 2688 18828 2740 18834
rect 2688 18770 2740 18776
rect 2872 18828 2924 18834
rect 2872 18770 2924 18776
rect 1412 18426 1440 18770
rect 2136 18624 2188 18630
rect 2136 18566 2188 18572
rect 1400 18420 1452 18426
rect 1400 18362 1452 18368
rect 1308 17740 1360 17746
rect 1308 17682 1360 17688
rect 1320 17338 1348 17682
rect 1768 17536 1820 17542
rect 1768 17478 1820 17484
rect 1952 17536 2004 17542
rect 1952 17478 2004 17484
rect 1308 17332 1360 17338
rect 1308 17274 1360 17280
rect 1676 16992 1728 16998
rect 1676 16934 1728 16940
rect 1400 16448 1452 16454
rect 1400 16390 1452 16396
rect 1412 14958 1440 16390
rect 1490 16008 1546 16017
rect 1490 15943 1546 15952
rect 1584 15972 1636 15978
rect 1504 15162 1532 15943
rect 1584 15914 1636 15920
rect 1596 15570 1624 15914
rect 1584 15564 1636 15570
rect 1584 15506 1636 15512
rect 1492 15156 1544 15162
rect 1492 15098 1544 15104
rect 1400 14952 1452 14958
rect 1400 14894 1452 14900
rect 1582 14512 1638 14521
rect 1582 14447 1638 14456
rect 1400 14340 1452 14346
rect 1400 14282 1452 14288
rect 110 13152 166 13161
rect 110 13087 166 13096
rect 124 12986 152 13087
rect 112 12980 164 12986
rect 112 12922 164 12928
rect 1412 12782 1440 14282
rect 1596 14074 1624 14447
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 1688 13870 1716 16934
rect 1780 16726 1808 17478
rect 1964 17134 1992 17478
rect 1952 17128 2004 17134
rect 1952 17070 2004 17076
rect 1768 16720 1820 16726
rect 1768 16662 1820 16668
rect 1860 16448 1912 16454
rect 1860 16390 1912 16396
rect 1872 16114 1900 16390
rect 1860 16108 1912 16114
rect 1860 16050 1912 16056
rect 1872 15706 1900 16050
rect 1860 15700 1912 15706
rect 1860 15642 1912 15648
rect 1964 15094 1992 17070
rect 1952 15088 2004 15094
rect 1952 15030 2004 15036
rect 1860 14272 1912 14278
rect 1860 14214 1912 14220
rect 1676 13864 1728 13870
rect 1676 13806 1728 13812
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 1872 11694 1900 14214
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 2056 13530 2084 13806
rect 2148 13530 2176 18566
rect 2700 18426 2728 18770
rect 2688 18420 2740 18426
rect 2688 18362 2740 18368
rect 2884 18222 2912 18770
rect 2320 18216 2372 18222
rect 2320 18158 2372 18164
rect 2872 18216 2924 18222
rect 2872 18158 2924 18164
rect 2332 17542 2360 18158
rect 2884 17746 2912 18158
rect 3068 17882 3096 20266
rect 4632 20058 4660 20402
rect 4620 20052 4672 20058
rect 4620 19994 4672 20000
rect 4908 19972 4936 21286
rect 5000 20330 5028 21354
rect 5092 20466 5120 21966
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5998 21448 6054 21457
rect 5998 21383 6054 21392
rect 5356 21072 5408 21078
rect 5356 21014 5408 21020
rect 5172 20528 5224 20534
rect 5172 20470 5224 20476
rect 5080 20460 5132 20466
rect 5080 20402 5132 20408
rect 4988 20324 5040 20330
rect 4988 20266 5040 20272
rect 5184 19990 5212 20470
rect 5368 20330 5396 21014
rect 5540 20936 5592 20942
rect 5540 20878 5592 20884
rect 5356 20324 5408 20330
rect 5356 20266 5408 20272
rect 4988 19984 5040 19990
rect 4908 19944 4988 19972
rect 4988 19926 5040 19932
rect 5172 19984 5224 19990
rect 5172 19926 5224 19932
rect 3332 19304 3384 19310
rect 3332 19246 3384 19252
rect 3240 19168 3292 19174
rect 3240 19110 3292 19116
rect 3148 18760 3200 18766
rect 3148 18702 3200 18708
rect 3160 18290 3188 18702
rect 3252 18358 3280 19110
rect 3344 18834 3372 19246
rect 4344 19236 4396 19242
rect 4344 19178 4396 19184
rect 4356 18970 4384 19178
rect 5000 19174 5028 19926
rect 5552 19854 5580 20878
rect 6012 20874 6040 21383
rect 6000 20868 6052 20874
rect 6000 20810 6052 20816
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 6012 20602 6040 20810
rect 6000 20596 6052 20602
rect 6000 20538 6052 20544
rect 6000 20324 6052 20330
rect 6000 20266 6052 20272
rect 5540 19848 5592 19854
rect 5540 19790 5592 19796
rect 5552 19514 5580 19790
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5540 19508 5592 19514
rect 5540 19450 5592 19456
rect 5264 19236 5316 19242
rect 5264 19178 5316 19184
rect 4988 19168 5040 19174
rect 4988 19110 5040 19116
rect 5276 18970 5304 19178
rect 5908 19168 5960 19174
rect 5908 19110 5960 19116
rect 5920 18970 5948 19110
rect 4344 18964 4396 18970
rect 4344 18906 4396 18912
rect 5264 18964 5316 18970
rect 5264 18906 5316 18912
rect 5908 18964 5960 18970
rect 5908 18906 5960 18912
rect 3332 18828 3384 18834
rect 3332 18770 3384 18776
rect 4356 18630 4384 18906
rect 3332 18624 3384 18630
rect 3332 18566 3384 18572
rect 4344 18624 4396 18630
rect 4344 18566 4396 18572
rect 3240 18352 3292 18358
rect 3240 18294 3292 18300
rect 3148 18284 3200 18290
rect 3148 18226 3200 18232
rect 3056 17876 3108 17882
rect 3056 17818 3108 17824
rect 2688 17740 2740 17746
rect 2688 17682 2740 17688
rect 2872 17740 2924 17746
rect 2872 17682 2924 17688
rect 2320 17536 2372 17542
rect 2320 17478 2372 17484
rect 2700 16998 2728 17682
rect 2884 17338 2912 17682
rect 2872 17332 2924 17338
rect 2872 17274 2924 17280
rect 2688 16992 2740 16998
rect 2688 16934 2740 16940
rect 2872 16992 2924 16998
rect 2872 16934 2924 16940
rect 2228 16720 2280 16726
rect 2228 16662 2280 16668
rect 2596 16720 2648 16726
rect 2596 16662 2648 16668
rect 2240 15706 2268 16662
rect 2320 16652 2372 16658
rect 2320 16594 2372 16600
rect 2332 16454 2360 16594
rect 2320 16448 2372 16454
rect 2320 16390 2372 16396
rect 2332 16114 2360 16390
rect 2608 16250 2636 16662
rect 2596 16244 2648 16250
rect 2596 16186 2648 16192
rect 2320 16108 2372 16114
rect 2320 16050 2372 16056
rect 2228 15700 2280 15706
rect 2228 15642 2280 15648
rect 2320 14476 2372 14482
rect 2320 14418 2372 14424
rect 2688 14476 2740 14482
rect 2688 14418 2740 14424
rect 2332 14278 2360 14418
rect 2320 14272 2372 14278
rect 2320 14214 2372 14220
rect 2044 13524 2096 13530
rect 2044 13466 2096 13472
rect 2136 13524 2188 13530
rect 2136 13466 2188 13472
rect 1952 13388 2004 13394
rect 1952 13330 2004 13336
rect 1964 12986 1992 13330
rect 2332 13297 2360 14214
rect 2700 13938 2728 14418
rect 2688 13932 2740 13938
rect 2688 13874 2740 13880
rect 2504 13388 2556 13394
rect 2504 13330 2556 13336
rect 2318 13288 2374 13297
rect 2318 13223 2374 13232
rect 2136 13184 2188 13190
rect 2136 13126 2188 13132
rect 2320 13184 2372 13190
rect 2320 13126 2372 13132
rect 1952 12980 2004 12986
rect 2004 12940 2084 12968
rect 1952 12922 2004 12928
rect 1952 12300 2004 12306
rect 1952 12242 2004 12248
rect 1964 12102 1992 12242
rect 1952 12096 2004 12102
rect 1952 12038 2004 12044
rect 1400 11688 1452 11694
rect 1400 11630 1452 11636
rect 1860 11688 1912 11694
rect 1860 11630 1912 11636
rect 112 11552 164 11558
rect 112 11494 164 11500
rect 20 11076 72 11082
rect 20 11018 72 11024
rect 124 9625 152 11494
rect 110 9616 166 9625
rect 110 9551 166 9560
rect 112 7948 164 7954
rect 112 7890 164 7896
rect 124 7857 152 7890
rect 110 7848 166 7857
rect 110 7783 166 7792
rect 1032 7744 1084 7750
rect 1032 7686 1084 7692
rect 112 6180 164 6186
rect 112 6122 164 6128
rect 124 6089 152 6122
rect 110 6080 166 6089
rect 110 6015 166 6024
rect 754 82 810 480
rect 1044 82 1072 7686
rect 1412 7002 1440 11630
rect 1582 10840 1638 10849
rect 1964 10810 1992 12038
rect 2056 11642 2084 12940
rect 2148 12617 2176 13126
rect 2134 12608 2190 12617
rect 2134 12543 2190 12552
rect 2228 12096 2280 12102
rect 2228 12038 2280 12044
rect 2056 11614 2176 11642
rect 2044 11552 2096 11558
rect 2044 11494 2096 11500
rect 1582 10775 1638 10784
rect 1952 10804 2004 10810
rect 1596 10266 1624 10775
rect 1952 10746 2004 10752
rect 2056 10538 2084 11494
rect 2044 10532 2096 10538
rect 2044 10474 2096 10480
rect 1584 10260 1636 10266
rect 1584 10202 1636 10208
rect 2056 10198 2084 10474
rect 2148 10266 2176 11614
rect 2240 11354 2268 12038
rect 2332 11762 2360 13126
rect 2516 12986 2544 13330
rect 2504 12980 2556 12986
rect 2504 12922 2556 12928
rect 2504 12368 2556 12374
rect 2424 12328 2504 12356
rect 2320 11756 2372 11762
rect 2320 11698 2372 11704
rect 2424 11558 2452 12328
rect 2504 12310 2556 12316
rect 2688 12368 2740 12374
rect 2688 12310 2740 12316
rect 2504 11688 2556 11694
rect 2504 11630 2556 11636
rect 2412 11552 2464 11558
rect 2412 11494 2464 11500
rect 2228 11348 2280 11354
rect 2228 11290 2280 11296
rect 2424 11286 2452 11494
rect 2412 11280 2464 11286
rect 2412 11222 2464 11228
rect 2412 11076 2464 11082
rect 2516 11064 2544 11630
rect 2464 11036 2544 11064
rect 2412 11018 2464 11024
rect 2228 11008 2280 11014
rect 2228 10950 2280 10956
rect 2240 10742 2268 10950
rect 2228 10736 2280 10742
rect 2228 10678 2280 10684
rect 2424 10674 2452 11018
rect 2412 10668 2464 10674
rect 2412 10610 2464 10616
rect 2136 10260 2188 10266
rect 2136 10202 2188 10208
rect 2044 10192 2096 10198
rect 2044 10134 2096 10140
rect 2424 10130 2452 10610
rect 1492 10124 1544 10130
rect 1492 10066 1544 10072
rect 2412 10124 2464 10130
rect 2412 10066 2464 10072
rect 2596 10124 2648 10130
rect 2596 10066 2648 10072
rect 1504 8974 1532 10066
rect 1584 9988 1636 9994
rect 1584 9930 1636 9936
rect 1596 9518 1624 9930
rect 1584 9512 1636 9518
rect 1584 9454 1636 9460
rect 1596 9042 1624 9454
rect 2412 9376 2464 9382
rect 2412 9318 2464 9324
rect 1584 9036 1636 9042
rect 1584 8978 1636 8984
rect 1492 8968 1544 8974
rect 1492 8910 1544 8916
rect 1504 7546 1532 8910
rect 1596 7750 1624 8978
rect 1676 8832 1728 8838
rect 1676 8774 1728 8780
rect 1688 8430 1716 8774
rect 2424 8430 2452 9318
rect 2608 8906 2636 10066
rect 2596 8900 2648 8906
rect 2596 8842 2648 8848
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1768 8424 1820 8430
rect 1768 8366 1820 8372
rect 2412 8424 2464 8430
rect 2412 8366 2464 8372
rect 1688 8090 1716 8366
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 1584 7744 1636 7750
rect 1584 7686 1636 7692
rect 1492 7540 1544 7546
rect 1492 7482 1544 7488
rect 1400 6996 1452 7002
rect 1400 6938 1452 6944
rect 1780 2961 1808 8366
rect 2136 7948 2188 7954
rect 2136 7890 2188 7896
rect 2148 7546 2176 7890
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 2700 6866 2728 12310
rect 2780 11008 2832 11014
rect 2780 10950 2832 10956
rect 2792 10130 2820 10950
rect 2780 10124 2832 10130
rect 2780 10066 2832 10072
rect 2792 9382 2820 10066
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2688 6860 2740 6866
rect 2688 6802 2740 6808
rect 2700 6458 2728 6802
rect 2688 6452 2740 6458
rect 2688 6394 2740 6400
rect 2792 4865 2820 9318
rect 2884 8090 2912 16934
rect 3056 16516 3108 16522
rect 3056 16458 3108 16464
rect 3068 15978 3096 16458
rect 3344 16232 3372 18566
rect 3976 18420 4028 18426
rect 3976 18362 4028 18368
rect 3988 18086 4016 18362
rect 4068 18216 4120 18222
rect 4068 18158 4120 18164
rect 5080 18216 5132 18222
rect 5080 18158 5132 18164
rect 3976 18080 4028 18086
rect 3976 18022 4028 18028
rect 4080 17814 4108 18158
rect 4252 18148 4304 18154
rect 4252 18090 4304 18096
rect 4264 17814 4292 18090
rect 4344 18080 4396 18086
rect 4344 18022 4396 18028
rect 4068 17808 4120 17814
rect 4068 17750 4120 17756
rect 4252 17808 4304 17814
rect 4252 17750 4304 17756
rect 4068 17672 4120 17678
rect 4068 17614 4120 17620
rect 3516 17128 3568 17134
rect 3516 17070 3568 17076
rect 3528 16726 3556 17070
rect 3792 17060 3844 17066
rect 3792 17002 3844 17008
rect 3804 16726 3832 17002
rect 4080 16794 4108 17614
rect 4264 16998 4292 17750
rect 4356 17678 4384 18022
rect 5092 17882 5120 18158
rect 5276 18086 5304 18906
rect 6012 18834 6040 20266
rect 6552 19984 6604 19990
rect 6552 19926 6604 19932
rect 6092 19848 6144 19854
rect 6092 19790 6144 19796
rect 6104 19174 6132 19790
rect 6564 19514 6592 19926
rect 6552 19508 6604 19514
rect 6552 19450 6604 19456
rect 6092 19168 6144 19174
rect 6092 19110 6144 19116
rect 6000 18828 6052 18834
rect 6000 18770 6052 18776
rect 5356 18760 5408 18766
rect 5356 18702 5408 18708
rect 5264 18080 5316 18086
rect 5264 18022 5316 18028
rect 5368 17882 5396 18702
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 6012 18426 6040 18770
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 5080 17876 5132 17882
rect 5080 17818 5132 17824
rect 5356 17876 5408 17882
rect 5356 17818 5408 17824
rect 4344 17672 4396 17678
rect 4344 17614 4396 17620
rect 4620 17536 4672 17542
rect 4620 17478 4672 17484
rect 4252 16992 4304 16998
rect 4252 16934 4304 16940
rect 4068 16788 4120 16794
rect 4068 16730 4120 16736
rect 3516 16720 3568 16726
rect 3516 16662 3568 16668
rect 3792 16720 3844 16726
rect 3792 16662 3844 16668
rect 4158 16688 4214 16697
rect 3528 16454 3556 16662
rect 3516 16448 3568 16454
rect 3516 16390 3568 16396
rect 3252 16204 3372 16232
rect 3056 15972 3108 15978
rect 3056 15914 3108 15920
rect 2964 15904 3016 15910
rect 2964 15846 3016 15852
rect 2976 15570 3004 15846
rect 3068 15706 3096 15914
rect 3056 15700 3108 15706
rect 3056 15642 3108 15648
rect 2964 15564 3016 15570
rect 2964 15506 3016 15512
rect 2976 15162 3004 15506
rect 2964 15156 3016 15162
rect 2964 15098 3016 15104
rect 3056 14952 3108 14958
rect 3056 14894 3108 14900
rect 2964 14816 3016 14822
rect 2964 14758 3016 14764
rect 2976 11626 3004 14758
rect 3068 14618 3096 14894
rect 3056 14612 3108 14618
rect 3056 14554 3108 14560
rect 3056 13524 3108 13530
rect 3056 13466 3108 13472
rect 2964 11620 3016 11626
rect 2964 11562 3016 11568
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 2976 8294 3004 8978
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2872 8084 2924 8090
rect 2872 8026 2924 8032
rect 2976 7954 3004 8230
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 2976 7546 3004 7890
rect 2964 7540 3016 7546
rect 2964 7482 3016 7488
rect 3068 7449 3096 13466
rect 3148 13320 3200 13326
rect 3148 13262 3200 13268
rect 3160 12986 3188 13262
rect 3148 12980 3200 12986
rect 3148 12922 3200 12928
rect 3146 9480 3202 9489
rect 3146 9415 3202 9424
rect 3160 9178 3188 9415
rect 3148 9172 3200 9178
rect 3148 9114 3200 9120
rect 3054 7440 3110 7449
rect 3054 7375 3110 7384
rect 3252 6390 3280 16204
rect 3528 15706 3556 16390
rect 3804 16250 3832 16662
rect 4158 16623 4214 16632
rect 4172 16590 4200 16623
rect 4160 16584 4212 16590
rect 4160 16526 4212 16532
rect 3792 16244 3844 16250
rect 3792 16186 3844 16192
rect 3516 15700 3568 15706
rect 3516 15642 3568 15648
rect 4172 15638 4200 16526
rect 4264 15638 4292 16934
rect 4344 16448 4396 16454
rect 4344 16390 4396 16396
rect 4356 16046 4384 16390
rect 4344 16040 4396 16046
rect 4344 15982 4396 15988
rect 4160 15632 4212 15638
rect 4160 15574 4212 15580
rect 4252 15632 4304 15638
rect 4252 15574 4304 15580
rect 4264 14822 4292 15574
rect 4252 14816 4304 14822
rect 4252 14758 4304 14764
rect 3516 14612 3568 14618
rect 3516 14554 3568 14560
rect 3424 14476 3476 14482
rect 3424 14418 3476 14424
rect 3436 13870 3464 14418
rect 3332 13864 3384 13870
rect 3332 13806 3384 13812
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 3344 13326 3372 13806
rect 3528 13530 3556 14554
rect 4356 14414 4384 15982
rect 4632 15910 4660 17478
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 4988 17128 5040 17134
rect 4988 17070 5040 17076
rect 5080 17128 5132 17134
rect 5080 17070 5132 17076
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4724 16794 4752 16934
rect 4712 16788 4764 16794
rect 4712 16730 4764 16736
rect 5000 16658 5028 17070
rect 4988 16652 5040 16658
rect 4988 16594 5040 16600
rect 5092 16046 5120 17070
rect 6000 16720 6052 16726
rect 6000 16662 6052 16668
rect 5448 16584 5500 16590
rect 5448 16526 5500 16532
rect 5460 16046 5488 16526
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5080 16040 5132 16046
rect 5080 15982 5132 15988
rect 5448 16040 5500 16046
rect 5448 15982 5500 15988
rect 4620 15904 4672 15910
rect 4620 15846 4672 15852
rect 4528 15496 4580 15502
rect 4528 15438 4580 15444
rect 4436 14476 4488 14482
rect 4436 14418 4488 14424
rect 4344 14408 4396 14414
rect 4344 14350 4396 14356
rect 3792 14272 3844 14278
rect 3792 14214 3844 14220
rect 3608 13864 3660 13870
rect 3608 13806 3660 13812
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 3332 13320 3384 13326
rect 3332 13262 3384 13268
rect 3424 13252 3476 13258
rect 3424 13194 3476 13200
rect 3332 12708 3384 12714
rect 3332 12650 3384 12656
rect 3344 11540 3372 12650
rect 3436 12442 3464 13194
rect 3516 13184 3568 13190
rect 3620 13172 3648 13806
rect 3568 13144 3648 13172
rect 3516 13126 3568 13132
rect 3424 12436 3476 12442
rect 3424 12378 3476 12384
rect 3528 12170 3556 13126
rect 3804 12850 3832 14214
rect 4356 12918 4384 14350
rect 4448 14074 4476 14418
rect 4540 14278 4568 15438
rect 5092 15366 5120 15982
rect 5264 15972 5316 15978
rect 5264 15914 5316 15920
rect 5080 15360 5132 15366
rect 5080 15302 5132 15308
rect 4528 14272 4580 14278
rect 4528 14214 4580 14220
rect 4436 14068 4488 14074
rect 4436 14010 4488 14016
rect 4344 12912 4396 12918
rect 4344 12854 4396 12860
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 4356 12782 4384 12854
rect 4344 12776 4396 12782
rect 4344 12718 4396 12724
rect 3700 12708 3752 12714
rect 3700 12650 3752 12656
rect 4068 12708 4120 12714
rect 4068 12650 4120 12656
rect 3712 12374 3740 12650
rect 4080 12442 4108 12650
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 4344 12436 4396 12442
rect 4344 12378 4396 12384
rect 3700 12368 3752 12374
rect 3700 12310 3752 12316
rect 4252 12300 4304 12306
rect 4252 12242 4304 12248
rect 3516 12164 3568 12170
rect 3516 12106 3568 12112
rect 3424 11552 3476 11558
rect 3344 11512 3424 11540
rect 3424 11494 3476 11500
rect 3436 11218 3464 11494
rect 3424 11212 3476 11218
rect 3424 11154 3476 11160
rect 3332 10736 3384 10742
rect 3332 10678 3384 10684
rect 3344 10470 3372 10678
rect 3332 10464 3384 10470
rect 3332 10406 3384 10412
rect 3344 10266 3372 10406
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 3436 9178 3464 11154
rect 3884 11076 3936 11082
rect 3884 11018 3936 11024
rect 4160 11076 4212 11082
rect 4160 11018 4212 11024
rect 3896 10810 3924 11018
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 3792 10464 3844 10470
rect 3792 10406 3844 10412
rect 3700 10192 3752 10198
rect 3700 10134 3752 10140
rect 3712 9722 3740 10134
rect 3804 9926 3832 10406
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 3700 9716 3752 9722
rect 3700 9658 3752 9664
rect 3700 9512 3752 9518
rect 3700 9454 3752 9460
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3712 8906 3740 9454
rect 3804 9353 3832 9862
rect 4080 9674 4108 10542
rect 3988 9654 4108 9674
rect 3976 9648 4108 9654
rect 4028 9646 4108 9648
rect 3976 9590 4028 9596
rect 3976 9376 4028 9382
rect 3790 9344 3846 9353
rect 3790 9279 3846 9288
rect 3896 9336 3976 9364
rect 3700 8900 3752 8906
rect 3700 8842 3752 8848
rect 3240 6384 3292 6390
rect 3240 6326 3292 6332
rect 2778 4856 2834 4865
rect 2778 4791 2834 4800
rect 2504 3936 2556 3942
rect 2504 3878 2556 3884
rect 1766 2952 1822 2961
rect 1766 2887 1822 2896
rect 754 54 1072 82
rect 2226 82 2282 480
rect 2516 82 2544 3878
rect 2226 54 2544 82
rect 3712 82 3740 8842
rect 3804 7546 3832 9279
rect 3896 8362 3924 9336
rect 3976 9318 4028 9324
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 4080 8430 4108 8910
rect 4172 8566 4200 11018
rect 4264 10996 4292 12242
rect 4356 11762 4384 12378
rect 4344 11756 4396 11762
rect 4344 11698 4396 11704
rect 4448 11608 4476 14010
rect 4540 13734 4568 14214
rect 4620 13864 4672 13870
rect 4620 13806 4672 13812
rect 4528 13728 4580 13734
rect 4528 13670 4580 13676
rect 4632 13394 4660 13806
rect 5092 13546 5120 15302
rect 5276 14890 5304 15914
rect 5356 15360 5408 15366
rect 5356 15302 5408 15308
rect 5264 14884 5316 14890
rect 5264 14826 5316 14832
rect 5368 14618 5396 15302
rect 5356 14612 5408 14618
rect 5356 14554 5408 14560
rect 5460 14550 5488 15982
rect 6012 15910 6040 16662
rect 6000 15904 6052 15910
rect 6000 15846 6052 15852
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 6012 14550 6040 15846
rect 5448 14544 5500 14550
rect 5448 14486 5500 14492
rect 6000 14544 6052 14550
rect 6000 14486 6052 14492
rect 5540 14476 5592 14482
rect 5540 14418 5592 14424
rect 5448 14408 5500 14414
rect 5448 14350 5500 14356
rect 5172 14272 5224 14278
rect 5172 14214 5224 14220
rect 5356 14272 5408 14278
rect 5356 14214 5408 14220
rect 5184 13734 5212 14214
rect 5368 14006 5396 14214
rect 5356 14000 5408 14006
rect 5276 13960 5356 13988
rect 5172 13728 5224 13734
rect 5172 13670 5224 13676
rect 5092 13518 5212 13546
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 4528 13320 4580 13326
rect 4528 13262 4580 13268
rect 4540 13190 4568 13262
rect 4528 13184 4580 13190
rect 4528 13126 4580 13132
rect 4632 12646 4660 13330
rect 4988 13184 5040 13190
rect 5040 13144 5120 13172
rect 4988 13126 5040 13132
rect 5092 12918 5120 13144
rect 5080 12912 5132 12918
rect 5080 12854 5132 12860
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 4988 12776 5040 12782
rect 4988 12718 5040 12724
rect 4620 12640 4672 12646
rect 4620 12582 4672 12588
rect 4528 11620 4580 11626
rect 4448 11580 4528 11608
rect 4344 11008 4396 11014
rect 4264 10968 4344 10996
rect 4344 10950 4396 10956
rect 4356 9625 4384 10950
rect 4342 9616 4398 9625
rect 4448 9586 4476 11580
rect 4528 11562 4580 11568
rect 4540 11354 4568 11562
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 4632 10470 4660 12582
rect 4712 11892 4764 11898
rect 4712 11834 4764 11840
rect 4724 11082 4752 11834
rect 4712 11076 4764 11082
rect 4712 11018 4764 11024
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 4528 10124 4580 10130
rect 4528 10066 4580 10072
rect 4342 9551 4398 9560
rect 4436 9580 4488 9586
rect 4436 9522 4488 9528
rect 4344 9444 4396 9450
rect 4344 9386 4396 9392
rect 4356 9178 4384 9386
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4160 8560 4212 8566
rect 4160 8502 4212 8508
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 4448 8362 4476 9522
rect 4540 8430 4568 10066
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4632 9722 4660 9998
rect 4620 9716 4672 9722
rect 4620 9658 4672 9664
rect 4712 9104 4764 9110
rect 4712 9046 4764 9052
rect 4724 8634 4752 9046
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 3884 8356 3936 8362
rect 3884 8298 3936 8304
rect 4436 8356 4488 8362
rect 4436 8298 4488 8304
rect 3792 7540 3844 7546
rect 3792 7482 3844 7488
rect 3896 7342 3924 8298
rect 4540 8090 4568 8366
rect 4528 8084 4580 8090
rect 4528 8026 4580 8032
rect 3884 7336 3936 7342
rect 3884 7278 3936 7284
rect 4620 7268 4672 7274
rect 4620 7210 4672 7216
rect 4632 6866 4660 7210
rect 4816 7002 4844 12718
rect 5000 12306 5028 12718
rect 4988 12300 5040 12306
rect 4988 12242 5040 12248
rect 4896 12096 4948 12102
rect 4896 12038 4948 12044
rect 4908 11830 4936 12038
rect 4896 11824 4948 11830
rect 4896 11766 4948 11772
rect 4908 11014 4936 11766
rect 5000 11354 5028 12242
rect 4988 11348 5040 11354
rect 4988 11290 5040 11296
rect 4896 11008 4948 11014
rect 4896 10950 4948 10956
rect 4908 7546 4936 10950
rect 5092 9110 5120 12854
rect 5184 11830 5212 13518
rect 5276 13394 5304 13960
rect 5356 13942 5408 13948
rect 5356 13796 5408 13802
rect 5460 13784 5488 14350
rect 5552 13870 5580 14418
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5540 13864 5592 13870
rect 5540 13806 5592 13812
rect 5408 13756 5488 13784
rect 5356 13738 5408 13744
rect 5460 13530 5488 13756
rect 5552 13705 5580 13806
rect 6012 13734 6040 14486
rect 6000 13728 6052 13734
rect 5538 13696 5594 13705
rect 6000 13670 6052 13676
rect 5538 13631 5594 13640
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 5264 13388 5316 13394
rect 5264 13330 5316 13336
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 5460 12918 5488 13330
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5448 12912 5500 12918
rect 5448 12854 5500 12860
rect 5816 12640 5868 12646
rect 5816 12582 5868 12588
rect 5828 12306 5856 12582
rect 6012 12374 6040 13670
rect 6000 12368 6052 12374
rect 6000 12310 6052 12316
rect 5816 12300 5868 12306
rect 5816 12242 5868 12248
rect 5264 12164 5316 12170
rect 5264 12106 5316 12112
rect 5172 11824 5224 11830
rect 5172 11766 5224 11772
rect 5172 11688 5224 11694
rect 5172 11630 5224 11636
rect 5184 11150 5212 11630
rect 5172 11144 5224 11150
rect 5172 11086 5224 11092
rect 5184 10742 5212 11086
rect 5172 10736 5224 10742
rect 5172 10678 5224 10684
rect 5184 10266 5212 10678
rect 5172 10260 5224 10266
rect 5172 10202 5224 10208
rect 5080 9104 5132 9110
rect 5080 9046 5132 9052
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 5000 8294 5028 8978
rect 5080 8968 5132 8974
rect 5080 8910 5132 8916
rect 4988 8288 5040 8294
rect 4988 8230 5040 8236
rect 5000 7954 5028 8230
rect 4988 7948 5040 7954
rect 4988 7890 5040 7896
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 5000 7274 5028 7890
rect 5092 7410 5120 8910
rect 5080 7404 5132 7410
rect 5080 7346 5132 7352
rect 4988 7268 5040 7274
rect 4988 7210 5040 7216
rect 4804 6996 4856 7002
rect 4804 6938 4856 6944
rect 4620 6860 4672 6866
rect 4620 6802 4672 6808
rect 4632 6118 4660 6802
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4632 1465 4660 6054
rect 5184 5778 5212 10202
rect 5276 8566 5304 12106
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5356 11620 5408 11626
rect 5356 11562 5408 11568
rect 5368 11218 5396 11562
rect 6012 11558 6040 12310
rect 6000 11552 6052 11558
rect 6000 11494 6052 11500
rect 5356 11212 5408 11218
rect 5356 11154 5408 11160
rect 5368 10130 5396 11154
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 5460 10470 5488 11086
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 5368 9926 5396 10066
rect 5552 10062 5580 10406
rect 6012 10130 6040 10950
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5448 9988 5500 9994
rect 5448 9930 5500 9936
rect 5356 9920 5408 9926
rect 5356 9862 5408 9868
rect 5368 9450 5396 9862
rect 5356 9444 5408 9450
rect 5356 9386 5408 9392
rect 5460 9382 5488 9930
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5460 8906 5488 9318
rect 5448 8900 5500 8906
rect 5448 8842 5500 8848
rect 5460 8634 5488 8842
rect 5552 8838 5580 9998
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5264 8560 5316 8566
rect 5264 8502 5316 8508
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 5368 7546 5396 8366
rect 5460 8090 5488 8570
rect 5552 8498 5580 8774
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5448 8084 5500 8090
rect 5448 8026 5500 8032
rect 5552 7818 5580 8434
rect 5632 8356 5684 8362
rect 5632 8298 5684 8304
rect 5644 7954 5672 8298
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5540 7812 5592 7818
rect 5540 7754 5592 7760
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5172 5772 5224 5778
rect 5172 5714 5224 5720
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 6012 5370 6040 5714
rect 6000 5364 6052 5370
rect 6000 5306 6052 5312
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 6104 2650 6132 19110
rect 6368 15632 6420 15638
rect 6368 15574 6420 15580
rect 6184 15496 6236 15502
rect 6184 15438 6236 15444
rect 6196 15026 6224 15438
rect 6276 15428 6328 15434
rect 6276 15370 6328 15376
rect 6288 15162 6316 15370
rect 6276 15156 6328 15162
rect 6276 15098 6328 15104
rect 6184 15020 6236 15026
rect 6184 14962 6236 14968
rect 6380 14822 6408 15574
rect 6368 14816 6420 14822
rect 6368 14758 6420 14764
rect 6380 14278 6408 14758
rect 6656 14618 6684 23462
rect 6748 22642 6776 24006
rect 6840 23118 6868 24006
rect 7748 23792 7800 23798
rect 7748 23734 7800 23740
rect 6920 23248 6972 23254
rect 6920 23190 6972 23196
rect 6828 23112 6880 23118
rect 6828 23054 6880 23060
rect 6932 22778 6960 23190
rect 7380 23044 7432 23050
rect 7380 22986 7432 22992
rect 6920 22772 6972 22778
rect 6920 22714 6972 22720
rect 6736 22636 6788 22642
rect 6736 22578 6788 22584
rect 6736 22432 6788 22438
rect 6736 22374 6788 22380
rect 6748 22098 6776 22374
rect 6932 22234 6960 22714
rect 7392 22642 7420 22986
rect 7760 22642 7788 23734
rect 8220 23730 8248 24210
rect 8956 23866 8984 27520
rect 10612 25786 10640 27520
rect 10612 25758 10732 25786
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10232 24064 10284 24070
rect 10232 24006 10284 24012
rect 8944 23860 8996 23866
rect 8944 23802 8996 23808
rect 10244 23730 10272 24006
rect 8208 23724 8260 23730
rect 8208 23666 8260 23672
rect 10232 23724 10284 23730
rect 10232 23666 10284 23672
rect 8220 23633 8248 23666
rect 8206 23624 8262 23633
rect 8206 23559 8262 23568
rect 9956 23520 10008 23526
rect 9956 23462 10008 23468
rect 9772 23248 9824 23254
rect 9772 23190 9824 23196
rect 7380 22636 7432 22642
rect 7380 22578 7432 22584
rect 7748 22636 7800 22642
rect 7748 22578 7800 22584
rect 8852 22636 8904 22642
rect 8852 22578 8904 22584
rect 9496 22636 9548 22642
rect 9496 22578 9548 22584
rect 6920 22228 6972 22234
rect 6920 22170 6972 22176
rect 6736 22092 6788 22098
rect 6736 22034 6788 22040
rect 6748 21350 6776 22034
rect 6736 21344 6788 21350
rect 6736 21286 6788 21292
rect 6748 16794 6776 21286
rect 7288 20936 7340 20942
rect 7288 20878 7340 20884
rect 7300 19990 7328 20878
rect 7288 19984 7340 19990
rect 7288 19926 7340 19932
rect 7196 18760 7248 18766
rect 7196 18702 7248 18708
rect 7012 18624 7064 18630
rect 7012 18566 7064 18572
rect 7024 18222 7052 18566
rect 6920 18216 6972 18222
rect 6920 18158 6972 18164
rect 7012 18216 7064 18222
rect 7012 18158 7064 18164
rect 6828 17672 6880 17678
rect 6828 17614 6880 17620
rect 6840 17338 6868 17614
rect 6828 17332 6880 17338
rect 6828 17274 6880 17280
rect 6736 16788 6788 16794
rect 6736 16730 6788 16736
rect 6932 16726 6960 18158
rect 7024 17746 7052 18158
rect 7208 17814 7236 18702
rect 7196 17808 7248 17814
rect 7196 17750 7248 17756
rect 7012 17740 7064 17746
rect 7012 17682 7064 17688
rect 7024 17134 7052 17682
rect 7392 17626 7420 22578
rect 8668 22432 8720 22438
rect 8668 22374 8720 22380
rect 8680 21554 8708 22374
rect 8864 22234 8892 22578
rect 9128 22432 9180 22438
rect 9128 22374 9180 22380
rect 8852 22228 8904 22234
rect 8852 22170 8904 22176
rect 8668 21548 8720 21554
rect 8668 21490 8720 21496
rect 9140 21486 9168 22374
rect 9128 21480 9180 21486
rect 9128 21422 9180 21428
rect 7564 21004 7616 21010
rect 7564 20946 7616 20952
rect 7576 20058 7604 20946
rect 8760 20528 8812 20534
rect 8760 20470 8812 20476
rect 7564 20052 7616 20058
rect 7564 19994 7616 20000
rect 7472 19236 7524 19242
rect 7472 19178 7524 19184
rect 7484 18970 7512 19178
rect 7576 19174 7604 19994
rect 8772 19990 8800 20470
rect 8208 19984 8260 19990
rect 8208 19926 8260 19932
rect 8760 19984 8812 19990
rect 8760 19926 8812 19932
rect 7840 19712 7892 19718
rect 7840 19654 7892 19660
rect 7852 19378 7880 19654
rect 8220 19514 8248 19926
rect 8484 19780 8536 19786
rect 8484 19722 8536 19728
rect 8208 19508 8260 19514
rect 8208 19450 8260 19456
rect 7840 19372 7892 19378
rect 7840 19314 7892 19320
rect 7564 19168 7616 19174
rect 7564 19110 7616 19116
rect 7472 18964 7524 18970
rect 7576 18952 7604 19110
rect 7656 18964 7708 18970
rect 7576 18924 7656 18952
rect 7472 18906 7524 18912
rect 7656 18906 7708 18912
rect 7484 18426 7512 18906
rect 7472 18420 7524 18426
rect 7472 18362 7524 18368
rect 7852 18290 7880 19314
rect 8496 18970 8524 19722
rect 8484 18964 8536 18970
rect 8484 18906 8536 18912
rect 8850 18728 8906 18737
rect 8850 18663 8906 18672
rect 8864 18630 8892 18663
rect 8852 18624 8904 18630
rect 8852 18566 8904 18572
rect 8864 18426 8892 18566
rect 8852 18420 8904 18426
rect 8852 18362 8904 18368
rect 7840 18284 7892 18290
rect 7840 18226 7892 18232
rect 8852 18284 8904 18290
rect 8852 18226 8904 18232
rect 8668 18148 8720 18154
rect 8668 18090 8720 18096
rect 7748 17808 7800 17814
rect 7748 17750 7800 17756
rect 7300 17598 7420 17626
rect 7012 17128 7064 17134
rect 7012 17070 7064 17076
rect 6920 16720 6972 16726
rect 6920 16662 6972 16668
rect 7104 15564 7156 15570
rect 7104 15506 7156 15512
rect 7116 14958 7144 15506
rect 7196 15360 7248 15366
rect 7196 15302 7248 15308
rect 7208 14958 7236 15302
rect 7300 15162 7328 17598
rect 7380 17536 7432 17542
rect 7380 17478 7432 17484
rect 7288 15156 7340 15162
rect 7288 15098 7340 15104
rect 7104 14952 7156 14958
rect 7104 14894 7156 14900
rect 7196 14952 7248 14958
rect 7196 14894 7248 14900
rect 6828 14884 6880 14890
rect 6828 14826 6880 14832
rect 6644 14612 6696 14618
rect 6644 14554 6696 14560
rect 6368 14272 6420 14278
rect 6368 14214 6420 14220
rect 6380 13938 6408 14214
rect 6368 13932 6420 13938
rect 6368 13874 6420 13880
rect 6656 13462 6684 14554
rect 6840 13870 6868 14826
rect 7116 14346 7144 14894
rect 7104 14340 7156 14346
rect 7104 14282 7156 14288
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 7196 13796 7248 13802
rect 7196 13738 7248 13744
rect 6736 13524 6788 13530
rect 6736 13466 6788 13472
rect 6644 13456 6696 13462
rect 6644 13398 6696 13404
rect 6552 13184 6604 13190
rect 6552 13126 6604 13132
rect 6564 12646 6592 13126
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 6564 12102 6592 12582
rect 6748 12442 6776 13466
rect 6736 12436 6788 12442
rect 6736 12378 6788 12384
rect 7104 12300 7156 12306
rect 7104 12242 7156 12248
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6564 11830 6592 12038
rect 6552 11824 6604 11830
rect 6552 11766 6604 11772
rect 6920 11824 6972 11830
rect 6920 11766 6972 11772
rect 6184 11552 6236 11558
rect 6184 11494 6236 11500
rect 6196 11150 6224 11494
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 6276 11076 6328 11082
rect 6276 11018 6328 11024
rect 6288 10742 6316 11018
rect 6276 10736 6328 10742
rect 6276 10678 6328 10684
rect 6644 10736 6696 10742
rect 6644 10678 6696 10684
rect 6288 9178 6316 10678
rect 6656 9926 6684 10678
rect 6840 10266 6868 11154
rect 6932 10742 6960 11766
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 7024 11558 7052 11698
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 6920 10736 6972 10742
rect 6920 10678 6972 10684
rect 7024 10674 7052 11494
rect 7116 11286 7144 12242
rect 7104 11280 7156 11286
rect 7104 11222 7156 11228
rect 7012 10668 7064 10674
rect 7012 10610 7064 10616
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 6736 9988 6788 9994
rect 6736 9930 6788 9936
rect 6368 9920 6420 9926
rect 6368 9862 6420 9868
rect 6644 9920 6696 9926
rect 6644 9862 6696 9868
rect 6276 9172 6328 9178
rect 6276 9114 6328 9120
rect 6276 8968 6328 8974
rect 6276 8910 6328 8916
rect 6184 7812 6236 7818
rect 6184 7754 6236 7760
rect 6196 6866 6224 7754
rect 6288 7750 6316 8910
rect 6380 8634 6408 9862
rect 6644 9648 6696 9654
rect 6644 9590 6696 9596
rect 6552 8832 6604 8838
rect 6656 8820 6684 9590
rect 6748 8838 6776 9930
rect 6840 9110 6868 10202
rect 6828 9104 6880 9110
rect 6828 9046 6880 9052
rect 6604 8792 6684 8820
rect 6552 8774 6604 8780
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 6656 8566 6684 8792
rect 6736 8832 6788 8838
rect 6736 8774 6788 8780
rect 6644 8560 6696 8566
rect 6644 8502 6696 8508
rect 6552 8288 6604 8294
rect 6748 8276 6776 8774
rect 6604 8248 6776 8276
rect 6552 8230 6604 8236
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 6196 6458 6224 6802
rect 6288 6730 6316 7686
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6472 7002 6500 7142
rect 6460 6996 6512 7002
rect 6460 6938 6512 6944
rect 6276 6724 6328 6730
rect 6276 6666 6328 6672
rect 6184 6452 6236 6458
rect 6184 6394 6236 6400
rect 6564 5370 6592 8230
rect 6840 7954 6868 9046
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6932 7410 6960 10474
rect 7024 10470 7052 10610
rect 7116 10606 7144 11222
rect 7208 11218 7236 13738
rect 7288 11620 7340 11626
rect 7288 11562 7340 11568
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 7196 11008 7248 11014
rect 7196 10950 7248 10956
rect 7208 10810 7236 10950
rect 7196 10804 7248 10810
rect 7196 10746 7248 10752
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 7024 9586 7052 10406
rect 7300 10198 7328 11562
rect 7288 10192 7340 10198
rect 7288 10134 7340 10140
rect 7102 10024 7158 10033
rect 7102 9959 7158 9968
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 7024 9382 7052 9522
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 6932 7002 6960 7346
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 7024 5914 7052 9318
rect 7116 8974 7144 9959
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 7208 9353 7236 9386
rect 7194 9344 7250 9353
rect 7194 9279 7250 9288
rect 7208 9110 7236 9279
rect 7300 9178 7328 10134
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7196 9104 7248 9110
rect 7196 9046 7248 9052
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 7116 8566 7144 8774
rect 7104 8560 7156 8566
rect 7104 8502 7156 8508
rect 7288 8424 7340 8430
rect 7288 8366 7340 8372
rect 7300 7954 7328 8366
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 7300 7342 7328 7890
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 7012 5908 7064 5914
rect 7012 5850 7064 5856
rect 6552 5364 6604 5370
rect 6552 5306 6604 5312
rect 7392 4154 7420 17478
rect 7760 16998 7788 17750
rect 8680 17270 8708 18090
rect 8864 17814 8892 18226
rect 8852 17808 8904 17814
rect 8852 17750 8904 17756
rect 8668 17264 8720 17270
rect 8668 17206 8720 17212
rect 8024 17128 8076 17134
rect 8024 17070 8076 17076
rect 8300 17128 8352 17134
rect 8300 17070 8352 17076
rect 7748 16992 7800 16998
rect 7748 16934 7800 16940
rect 7656 16652 7708 16658
rect 7656 16594 7708 16600
rect 7668 16250 7696 16594
rect 7760 16590 7788 16934
rect 7932 16652 7984 16658
rect 7932 16594 7984 16600
rect 7748 16584 7800 16590
rect 7748 16526 7800 16532
rect 7656 16244 7708 16250
rect 7656 16186 7708 16192
rect 7668 14482 7696 16186
rect 7944 15978 7972 16594
rect 7932 15972 7984 15978
rect 7932 15914 7984 15920
rect 7944 15570 7972 15914
rect 7932 15564 7984 15570
rect 7932 15506 7984 15512
rect 7840 15360 7892 15366
rect 7840 15302 7892 15308
rect 7852 15026 7880 15302
rect 7840 15020 7892 15026
rect 7840 14962 7892 14968
rect 7656 14476 7708 14482
rect 7656 14418 7708 14424
rect 7840 14476 7892 14482
rect 7840 14418 7892 14424
rect 7668 13734 7696 14418
rect 7656 13728 7708 13734
rect 7656 13670 7708 13676
rect 7564 13320 7616 13326
rect 7564 13262 7616 13268
rect 7472 12980 7524 12986
rect 7472 12922 7524 12928
rect 7484 12714 7512 12922
rect 7576 12850 7604 13262
rect 7852 13190 7880 14418
rect 7944 14278 7972 15506
rect 7932 14272 7984 14278
rect 7932 14214 7984 14220
rect 7840 13184 7892 13190
rect 7840 13126 7892 13132
rect 7564 12844 7616 12850
rect 7564 12786 7616 12792
rect 7472 12708 7524 12714
rect 7472 12650 7524 12656
rect 7656 12232 7708 12238
rect 7656 12174 7708 12180
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 7564 12096 7616 12102
rect 7564 12038 7616 12044
rect 7484 11830 7512 12038
rect 7576 11898 7604 12038
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7472 11824 7524 11830
rect 7472 11766 7524 11772
rect 7484 10742 7512 11766
rect 7668 11558 7696 12174
rect 7852 11898 7880 13126
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 7656 11552 7708 11558
rect 7656 11494 7708 11500
rect 7564 11076 7616 11082
rect 7564 11018 7616 11024
rect 7472 10736 7524 10742
rect 7472 10678 7524 10684
rect 7484 10266 7512 10678
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7484 9761 7512 9862
rect 7470 9752 7526 9761
rect 7576 9722 7604 11018
rect 7668 9994 7696 11494
rect 7944 11354 7972 14214
rect 8036 13814 8064 17070
rect 8116 16992 8168 16998
rect 8116 16934 8168 16940
rect 8128 15910 8156 16934
rect 8312 16454 8340 17070
rect 8300 16448 8352 16454
rect 8300 16390 8352 16396
rect 8208 16040 8260 16046
rect 8208 15982 8260 15988
rect 8116 15904 8168 15910
rect 8116 15846 8168 15852
rect 8128 15162 8156 15846
rect 8220 15366 8248 15982
rect 8312 15638 8340 16390
rect 9140 16250 9168 21422
rect 9220 21004 9272 21010
rect 9220 20946 9272 20952
rect 9232 20602 9260 20946
rect 9220 20596 9272 20602
rect 9220 20538 9272 20544
rect 9312 18080 9364 18086
rect 9312 18022 9364 18028
rect 9220 17604 9272 17610
rect 9220 17546 9272 17552
rect 9232 17338 9260 17546
rect 9220 17332 9272 17338
rect 9220 17274 9272 17280
rect 9128 16244 9180 16250
rect 9128 16186 9180 16192
rect 8300 15632 8352 15638
rect 8300 15574 8352 15580
rect 8392 15428 8444 15434
rect 8392 15370 8444 15376
rect 8208 15360 8260 15366
rect 8208 15302 8260 15308
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 8404 14958 8432 15370
rect 8116 14952 8168 14958
rect 8116 14894 8168 14900
rect 8392 14952 8444 14958
rect 8392 14894 8444 14900
rect 8128 14482 8156 14894
rect 8404 14550 8432 14894
rect 8392 14544 8444 14550
rect 8392 14486 8444 14492
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 8760 14272 8812 14278
rect 8760 14214 8812 14220
rect 8852 14272 8904 14278
rect 8852 14214 8904 14220
rect 8772 13938 8800 14214
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 8036 13786 8156 13814
rect 8024 12640 8076 12646
rect 8024 12582 8076 12588
rect 8036 12238 8064 12582
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 7932 11348 7984 11354
rect 7932 11290 7984 11296
rect 7932 11144 7984 11150
rect 8036 11132 8064 12174
rect 8128 11898 8156 13786
rect 8208 13728 8260 13734
rect 8208 13670 8260 13676
rect 8574 13696 8630 13705
rect 8116 11892 8168 11898
rect 8116 11834 8168 11840
rect 7984 11104 8064 11132
rect 7932 11086 7984 11092
rect 7748 10736 7800 10742
rect 7748 10678 7800 10684
rect 7656 9988 7708 9994
rect 7656 9930 7708 9936
rect 7470 9687 7526 9696
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 7668 9518 7696 9930
rect 7760 9654 7788 10678
rect 7840 10464 7892 10470
rect 7840 10406 7892 10412
rect 7748 9648 7800 9654
rect 7748 9590 7800 9596
rect 7656 9512 7708 9518
rect 7470 9480 7526 9489
rect 7656 9454 7708 9460
rect 7470 9415 7526 9424
rect 7484 7954 7512 9415
rect 7668 9382 7696 9454
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7472 7948 7524 7954
rect 7472 7890 7524 7896
rect 7484 7274 7512 7890
rect 7472 7268 7524 7274
rect 7472 7210 7524 7216
rect 7484 5778 7512 7210
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 7472 5772 7524 5778
rect 7472 5714 7524 5720
rect 7484 4826 7512 5714
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 7576 4282 7604 7142
rect 7668 5030 7696 9318
rect 7852 8430 7880 10406
rect 7944 10062 7972 11086
rect 7932 10056 7984 10062
rect 7930 10024 7932 10033
rect 7984 10024 7986 10033
rect 7930 9959 7986 9968
rect 7930 9752 7986 9761
rect 7930 9687 7986 9696
rect 7944 8498 7972 9687
rect 8220 9489 8248 13670
rect 8574 13631 8630 13640
rect 8588 13530 8616 13631
rect 8576 13524 8628 13530
rect 8576 13466 8628 13472
rect 8864 13433 8892 14214
rect 9128 13864 9180 13870
rect 9128 13806 9180 13812
rect 9140 13705 9168 13806
rect 9126 13696 9182 13705
rect 9126 13631 9182 13640
rect 9140 13530 9168 13631
rect 9128 13524 9180 13530
rect 9128 13466 9180 13472
rect 8850 13424 8906 13433
rect 8850 13359 8906 13368
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8588 12782 8616 13126
rect 8668 12912 8720 12918
rect 8668 12854 8720 12860
rect 8576 12776 8628 12782
rect 8576 12718 8628 12724
rect 8588 12170 8616 12718
rect 8680 12646 8708 12854
rect 8760 12708 8812 12714
rect 8864 12696 8892 13359
rect 8944 12776 8996 12782
rect 8944 12718 8996 12724
rect 8812 12668 8892 12696
rect 8760 12650 8812 12656
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 8850 12608 8906 12617
rect 8576 12164 8628 12170
rect 8576 12106 8628 12112
rect 8588 11626 8616 12106
rect 8680 11744 8708 12582
rect 8956 12594 8984 12718
rect 8906 12566 8984 12594
rect 8850 12543 8906 12552
rect 8864 12442 8892 12543
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 8864 11830 8892 12378
rect 8852 11824 8904 11830
rect 8852 11766 8904 11772
rect 8760 11756 8812 11762
rect 8680 11716 8760 11744
rect 8760 11698 8812 11704
rect 8576 11620 8628 11626
rect 8576 11562 8628 11568
rect 8300 9920 8352 9926
rect 8300 9862 8352 9868
rect 8206 9480 8262 9489
rect 8206 9415 8262 9424
rect 8312 9042 8340 9862
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8116 9036 8168 9042
rect 8116 8978 8168 8984
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 7840 8424 7892 8430
rect 7840 8366 7892 8372
rect 7852 7954 7880 8366
rect 8024 8356 8076 8362
rect 8024 8298 8076 8304
rect 7840 7948 7892 7954
rect 7840 7890 7892 7896
rect 7852 7002 7880 7890
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 7840 6996 7892 7002
rect 7840 6938 7892 6944
rect 7944 5778 7972 7278
rect 8036 6798 8064 8298
rect 8128 8294 8156 8978
rect 8208 8900 8260 8906
rect 8208 8842 8260 8848
rect 8116 8288 8168 8294
rect 8116 8230 8168 8236
rect 8128 7818 8156 8230
rect 8220 8090 8248 8842
rect 8312 8090 8340 8978
rect 8208 8084 8260 8090
rect 8208 8026 8260 8032
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8116 7812 8168 7818
rect 8116 7754 8168 7760
rect 8312 7546 8340 8026
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8208 6996 8260 7002
rect 8404 6984 8432 9318
rect 8588 9110 8616 11562
rect 8668 11212 8720 11218
rect 8668 11154 8720 11160
rect 8680 10606 8708 11154
rect 8772 11014 8800 11698
rect 8864 11354 8892 11766
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8760 11008 8812 11014
rect 8760 10950 8812 10956
rect 8772 10810 8800 10950
rect 8760 10804 8812 10810
rect 8760 10746 8812 10752
rect 8668 10600 8720 10606
rect 8668 10542 8720 10548
rect 8680 10198 8708 10542
rect 8772 10266 8800 10746
rect 8864 10742 8892 11290
rect 8852 10736 8904 10742
rect 8852 10678 8904 10684
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8668 10192 8720 10198
rect 8668 10134 8720 10140
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 8576 9104 8628 9110
rect 8576 9046 8628 9052
rect 8772 9042 8800 9454
rect 8760 9036 8812 9042
rect 8760 8978 8812 8984
rect 9140 8430 9168 13466
rect 9324 12986 9352 18022
rect 9404 17808 9456 17814
rect 9404 17750 9456 17756
rect 9416 16794 9444 17750
rect 9404 16788 9456 16794
rect 9404 16730 9456 16736
rect 9508 16250 9536 22578
rect 9784 22438 9812 23190
rect 9862 23080 9918 23089
rect 9862 23015 9918 23024
rect 9772 22432 9824 22438
rect 9772 22374 9824 22380
rect 9680 22092 9732 22098
rect 9680 22034 9732 22040
rect 9692 21690 9720 22034
rect 9876 21690 9904 23015
rect 9968 22574 9996 23462
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10140 23112 10192 23118
rect 10140 23054 10192 23060
rect 10232 23112 10284 23118
rect 10232 23054 10284 23060
rect 9956 22568 10008 22574
rect 9956 22510 10008 22516
rect 10152 22114 10180 23054
rect 10244 22642 10272 23054
rect 10232 22636 10284 22642
rect 10232 22578 10284 22584
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10704 22234 10732 25758
rect 11610 24848 11666 24857
rect 11610 24783 11666 24792
rect 11624 24274 11652 24783
rect 11612 24268 11664 24274
rect 11612 24210 11664 24216
rect 11336 24064 11388 24070
rect 11336 24006 11388 24012
rect 11348 23118 11376 24006
rect 11624 23866 11652 24210
rect 11612 23860 11664 23866
rect 11612 23802 11664 23808
rect 11612 23588 11664 23594
rect 11612 23530 11664 23536
rect 11428 23248 11480 23254
rect 11428 23190 11480 23196
rect 11336 23112 11388 23118
rect 11336 23054 11388 23060
rect 11348 22778 11376 23054
rect 11336 22772 11388 22778
rect 11336 22714 11388 22720
rect 11440 22642 11468 23190
rect 11624 23118 11652 23530
rect 11612 23112 11664 23118
rect 11612 23054 11664 23060
rect 11428 22636 11480 22642
rect 11428 22578 11480 22584
rect 10784 22568 10836 22574
rect 10784 22510 10836 22516
rect 10692 22228 10744 22234
rect 10692 22170 10744 22176
rect 10322 22128 10378 22137
rect 10152 22086 10322 22114
rect 10322 22063 10378 22072
rect 10336 22030 10364 22063
rect 10324 22024 10376 22030
rect 10324 21966 10376 21972
rect 9680 21684 9732 21690
rect 9680 21626 9732 21632
rect 9864 21684 9916 21690
rect 9864 21626 9916 21632
rect 9692 21146 9720 21626
rect 10796 21570 10824 22510
rect 10704 21542 10824 21570
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 9680 21140 9732 21146
rect 9680 21082 9732 21088
rect 9588 20392 9640 20398
rect 9588 20334 9640 20340
rect 9600 19514 9628 20334
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 9772 19984 9824 19990
rect 9772 19926 9824 19932
rect 9588 19508 9640 19514
rect 9588 19450 9640 19456
rect 9784 19174 9812 19926
rect 9864 19304 9916 19310
rect 9864 19246 9916 19252
rect 9772 19168 9824 19174
rect 9772 19110 9824 19116
rect 9876 17796 9904 19246
rect 10048 19168 10100 19174
rect 10048 19110 10100 19116
rect 9956 18760 10008 18766
rect 9956 18702 10008 18708
rect 9968 18290 9996 18702
rect 10060 18426 10088 19110
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10048 18420 10100 18426
rect 10048 18362 10100 18368
rect 9956 18284 10008 18290
rect 9956 18226 10008 18232
rect 10060 18136 10088 18362
rect 10140 18148 10192 18154
rect 10060 18108 10140 18136
rect 10140 18090 10192 18096
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 9956 17808 10008 17814
rect 9876 17768 9956 17796
rect 9876 17338 9904 17768
rect 9956 17750 10008 17756
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 9956 17128 10008 17134
rect 9956 17070 10008 17076
rect 9968 16726 9996 17070
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 9956 16720 10008 16726
rect 9956 16662 10008 16668
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 10140 16108 10192 16114
rect 10140 16050 10192 16056
rect 10152 15978 10180 16050
rect 10140 15972 10192 15978
rect 10140 15914 10192 15920
rect 9588 15904 9640 15910
rect 9588 15846 9640 15852
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 9508 14074 9536 14214
rect 9496 14068 9548 14074
rect 9496 14010 9548 14016
rect 9312 12980 9364 12986
rect 9312 12922 9364 12928
rect 9600 10810 9628 15846
rect 10152 15706 10180 15914
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 9956 15632 10008 15638
rect 9956 15574 10008 15580
rect 9968 15162 9996 15574
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 10152 15094 10180 15642
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 10336 15162 10364 15438
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 10140 15088 10192 15094
rect 10140 15030 10192 15036
rect 10048 15020 10100 15026
rect 10048 14962 10100 14968
rect 10060 14618 10088 14962
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10704 14618 10732 21542
rect 11060 21344 11112 21350
rect 11060 21286 11112 21292
rect 11072 20602 11100 21286
rect 11428 20936 11480 20942
rect 11428 20878 11480 20884
rect 11060 20596 11112 20602
rect 11060 20538 11112 20544
rect 11440 19990 11468 20878
rect 11428 19984 11480 19990
rect 11428 19926 11480 19932
rect 10876 19848 10928 19854
rect 10876 19790 10928 19796
rect 10888 19378 10916 19790
rect 11440 19514 11468 19926
rect 11428 19508 11480 19514
rect 11428 19450 11480 19456
rect 10876 19372 10928 19378
rect 10876 19314 10928 19320
rect 10784 19304 10836 19310
rect 10888 19281 10916 19314
rect 10784 19246 10836 19252
rect 10874 19272 10930 19281
rect 10796 18154 10824 19246
rect 10874 19207 10930 19216
rect 11152 18964 11204 18970
rect 11152 18906 11204 18912
rect 11164 18426 11192 18906
rect 11428 18760 11480 18766
rect 11428 18702 11480 18708
rect 11152 18420 11204 18426
rect 11152 18362 11204 18368
rect 10784 18148 10836 18154
rect 10784 18090 10836 18096
rect 10796 17814 10824 18090
rect 11164 17814 11192 18362
rect 11440 18086 11468 18702
rect 11428 18080 11480 18086
rect 11428 18022 11480 18028
rect 11520 18080 11572 18086
rect 11520 18022 11572 18028
rect 10784 17808 10836 17814
rect 10784 17750 10836 17756
rect 11152 17808 11204 17814
rect 11152 17750 11204 17756
rect 11336 17808 11388 17814
rect 11336 17750 11388 17756
rect 11152 17604 11204 17610
rect 11152 17546 11204 17552
rect 10876 17196 10928 17202
rect 10876 17138 10928 17144
rect 10888 16658 10916 17138
rect 10968 16720 11020 16726
rect 11020 16680 11100 16708
rect 10968 16662 11020 16668
rect 10876 16652 10928 16658
rect 10876 16594 10928 16600
rect 10784 15972 10836 15978
rect 10784 15914 10836 15920
rect 10796 15638 10824 15914
rect 10888 15910 10916 16594
rect 10968 16040 11020 16046
rect 10968 15982 11020 15988
rect 10876 15904 10928 15910
rect 10876 15846 10928 15852
rect 10784 15632 10836 15638
rect 10784 15574 10836 15580
rect 10980 15502 11008 15982
rect 11072 15910 11100 16680
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 10980 15026 11008 15438
rect 10968 15020 11020 15026
rect 10968 14962 11020 14968
rect 11072 14906 11100 15846
rect 10796 14878 11100 14906
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 10048 14612 10100 14618
rect 10048 14554 10100 14560
rect 10692 14612 10744 14618
rect 10692 14554 10744 14560
rect 9784 13734 9812 14554
rect 9772 13728 9824 13734
rect 9772 13670 9824 13676
rect 9956 13728 10008 13734
rect 9956 13670 10008 13676
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9692 12646 9720 13126
rect 9968 12714 9996 13670
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10140 13388 10192 13394
rect 10140 13330 10192 13336
rect 9956 12708 10008 12714
rect 9956 12650 10008 12656
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9692 12306 9720 12582
rect 10152 12442 10180 13330
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10140 12436 10192 12442
rect 10140 12378 10192 12384
rect 10704 12374 10732 12786
rect 10692 12368 10744 12374
rect 10692 12310 10744 12316
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 9588 10804 9640 10810
rect 9588 10746 9640 10752
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 9416 8906 9444 9998
rect 9404 8900 9456 8906
rect 9404 8842 9456 8848
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9140 8022 9168 8366
rect 9508 8090 9536 8366
rect 9692 8294 9720 12242
rect 10140 12096 10192 12102
rect 10140 12038 10192 12044
rect 10152 11898 10180 12038
rect 10796 11898 10824 14878
rect 10876 14272 10928 14278
rect 10876 14214 10928 14220
rect 10888 13870 10916 14214
rect 10876 13864 10928 13870
rect 10876 13806 10928 13812
rect 10968 13864 11020 13870
rect 10968 13806 11020 13812
rect 11164 13814 11192 17546
rect 11348 17338 11376 17750
rect 11336 17332 11388 17338
rect 11336 17274 11388 17280
rect 11348 17066 11376 17274
rect 11336 17060 11388 17066
rect 11336 17002 11388 17008
rect 11440 16726 11468 18022
rect 11428 16720 11480 16726
rect 11428 16662 11480 16668
rect 11244 14952 11296 14958
rect 11244 14894 11296 14900
rect 11256 14618 11284 14894
rect 11244 14612 11296 14618
rect 11244 14554 11296 14560
rect 11256 14006 11284 14554
rect 11244 14000 11296 14006
rect 11244 13942 11296 13948
rect 10980 13190 11008 13806
rect 11164 13786 11284 13814
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 11164 12850 11192 13126
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 10784 11892 10836 11898
rect 10784 11834 10836 11840
rect 10796 11694 10824 11834
rect 10784 11688 10836 11694
rect 10784 11630 10836 11636
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 9968 11082 9996 11494
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10048 11144 10100 11150
rect 10048 11086 10100 11092
rect 9956 11076 10008 11082
rect 9956 11018 10008 11024
rect 10060 10674 10088 11086
rect 10048 10668 10100 10674
rect 10048 10610 10100 10616
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 9956 10192 10008 10198
rect 9956 10134 10008 10140
rect 9968 9382 9996 10134
rect 10796 10130 10824 11630
rect 11256 11200 11284 13786
rect 11428 12368 11480 12374
rect 11428 12310 11480 12316
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 11348 11354 11376 12174
rect 11440 11898 11468 12310
rect 11428 11892 11480 11898
rect 11428 11834 11480 11840
rect 11336 11348 11388 11354
rect 11336 11290 11388 11296
rect 11428 11212 11480 11218
rect 11256 11172 11428 11200
rect 11428 11154 11480 11160
rect 11336 10600 11388 10606
rect 11336 10542 11388 10548
rect 10876 10464 10928 10470
rect 10876 10406 10928 10412
rect 10784 10124 10836 10130
rect 10784 10066 10836 10072
rect 10048 10056 10100 10062
rect 10048 9998 10100 10004
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 9784 9110 9812 9318
rect 9772 9104 9824 9110
rect 9824 9064 9904 9092
rect 9772 9046 9824 9052
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9784 8498 9812 8774
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9680 8288 9732 8294
rect 9680 8230 9732 8236
rect 9876 8090 9904 9064
rect 9496 8084 9548 8090
rect 9496 8026 9548 8032
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 8944 8016 8996 8022
rect 8944 7958 8996 7964
rect 9128 8016 9180 8022
rect 9128 7958 9180 7964
rect 8484 7880 8536 7886
rect 8956 7857 8984 7958
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 8484 7822 8536 7828
rect 8942 7848 8998 7857
rect 8260 6956 8432 6984
rect 8208 6938 8260 6944
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 8036 5778 8064 6734
rect 8220 6100 8248 6938
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 8312 6254 8340 6598
rect 8496 6254 8524 7822
rect 8942 7783 8998 7792
rect 9784 7546 9812 7890
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 8758 7440 8814 7449
rect 8758 7375 8814 7384
rect 8772 7274 8800 7375
rect 8760 7268 8812 7274
rect 8760 7210 8812 7216
rect 8852 7268 8904 7274
rect 8852 7210 8904 7216
rect 9404 7268 9456 7274
rect 9404 7210 9456 7216
rect 8772 7002 8800 7210
rect 8760 6996 8812 7002
rect 8760 6938 8812 6944
rect 8864 6662 8892 7210
rect 9312 7200 9364 7206
rect 9312 7142 9364 7148
rect 8852 6656 8904 6662
rect 8852 6598 8904 6604
rect 9324 6390 9352 7142
rect 9312 6384 9364 6390
rect 9312 6326 9364 6332
rect 9416 6372 9444 7210
rect 9876 6866 9904 8026
rect 9968 7002 9996 9318
rect 10060 8906 10088 9998
rect 10784 9920 10836 9926
rect 10784 9862 10836 9868
rect 10796 9722 10824 9862
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10048 8900 10100 8906
rect 10048 8842 10100 8848
rect 10704 8838 10732 9454
rect 10796 9110 10824 9658
rect 10784 9104 10836 9110
rect 10784 9046 10836 9052
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 10060 8362 10088 8570
rect 10048 8356 10100 8362
rect 10048 8298 10100 8304
rect 10060 7954 10088 8298
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10048 7948 10100 7954
rect 10048 7890 10100 7896
rect 10060 7546 10088 7890
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 10520 7410 10548 7822
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 10888 7342 10916 10406
rect 11348 10062 11376 10542
rect 11440 10470 11468 11154
rect 11428 10464 11480 10470
rect 11428 10406 11480 10412
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11428 9376 11480 9382
rect 11428 9318 11480 9324
rect 11244 8560 11296 8566
rect 11244 8502 11296 8508
rect 11256 7342 11284 8502
rect 11336 8356 11388 8362
rect 11336 8298 11388 8304
rect 11348 8090 11376 8298
rect 11336 8084 11388 8090
rect 11336 8026 11388 8032
rect 11440 7993 11468 9318
rect 11426 7984 11482 7993
rect 11426 7919 11482 7928
rect 10876 7336 10928 7342
rect 10876 7278 10928 7284
rect 11244 7336 11296 7342
rect 11244 7278 11296 7284
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 11256 7002 11284 7278
rect 9956 6996 10008 7002
rect 9956 6938 10008 6944
rect 11244 6996 11296 7002
rect 11244 6938 11296 6944
rect 9864 6860 9916 6866
rect 9784 6820 9864 6848
rect 9496 6384 9548 6390
rect 9416 6344 9496 6372
rect 8300 6248 8352 6254
rect 8300 6190 8352 6196
rect 8484 6248 8536 6254
rect 8484 6190 8536 6196
rect 8300 6112 8352 6118
rect 8220 6072 8300 6100
rect 8300 6054 8352 6060
rect 7932 5772 7984 5778
rect 7932 5714 7984 5720
rect 8024 5772 8076 5778
rect 8024 5714 8076 5720
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 7564 4276 7616 4282
rect 7564 4218 7616 4224
rect 7300 4126 7420 4154
rect 7300 2650 7328 4126
rect 6092 2644 6144 2650
rect 6092 2586 6144 2592
rect 7288 2644 7340 2650
rect 7288 2586 7340 2592
rect 7196 2508 7248 2514
rect 7196 2450 7248 2456
rect 5540 2304 5592 2310
rect 5540 2246 5592 2252
rect 4618 1456 4674 1465
rect 4618 1391 4674 1400
rect 3790 82 3846 480
rect 3712 54 3846 82
rect 754 0 810 54
rect 2226 0 2282 54
rect 3790 0 3846 54
rect 5354 82 5410 480
rect 5552 82 5580 2246
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 5354 54 5580 82
rect 6918 82 6974 480
rect 7208 82 7236 2450
rect 7668 105 7696 4966
rect 7944 4826 7972 5714
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8220 5234 8248 5646
rect 8208 5228 8260 5234
rect 8208 5170 8260 5176
rect 8220 4826 8248 5170
rect 8312 5030 8340 6054
rect 8496 5914 8524 6190
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 9416 5710 9444 6344
rect 9496 6326 9548 6332
rect 9784 6254 9812 6820
rect 9864 6802 9916 6808
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 9876 5846 9904 6394
rect 11152 6384 11204 6390
rect 11152 6326 11204 6332
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 9864 5840 9916 5846
rect 9864 5782 9916 5788
rect 10232 5840 10284 5846
rect 10232 5782 10284 5788
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 9876 5370 9904 5782
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 10244 5234 10272 5782
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 10520 5234 10548 5646
rect 10796 5574 10824 6258
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10796 5273 10824 5510
rect 11164 5370 11192 6326
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 10782 5264 10838 5273
rect 10232 5228 10284 5234
rect 10152 5188 10232 5216
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8312 4010 8340 4966
rect 8300 4004 8352 4010
rect 8300 3946 8352 3952
rect 9324 3942 9352 4966
rect 10152 4826 10180 5188
rect 10232 5170 10284 5176
rect 10508 5228 10560 5234
rect 10560 5188 10732 5216
rect 10782 5199 10838 5208
rect 10508 5170 10560 5176
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10704 4758 10732 5188
rect 11256 5098 11284 6734
rect 11348 6458 11376 6802
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 11244 5092 11296 5098
rect 11244 5034 11296 5040
rect 10692 4752 10744 4758
rect 10692 4694 10744 4700
rect 10704 4282 10732 4694
rect 11428 4684 11480 4690
rect 11428 4626 11480 4632
rect 11440 4282 11468 4626
rect 10692 4276 10744 4282
rect 10692 4218 10744 4224
rect 11428 4276 11480 4282
rect 11428 4218 11480 4224
rect 9864 4004 9916 4010
rect 9864 3946 9916 3952
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 9048 3602 9076 3878
rect 9876 3670 9904 3946
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 9864 3664 9916 3670
rect 9864 3606 9916 3612
rect 9036 3596 9088 3602
rect 9036 3538 9088 3544
rect 8024 3528 8076 3534
rect 8024 3470 8076 3476
rect 8036 3194 8064 3470
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 8036 2854 8064 3130
rect 9048 3058 9076 3538
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 9232 3194 9260 3470
rect 9876 3194 9904 3606
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9968 3126 9996 3878
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10416 3460 10468 3466
rect 10416 3402 10468 3408
rect 9956 3120 10008 3126
rect 9956 3062 10008 3068
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 8208 2916 8260 2922
rect 8208 2858 8260 2864
rect 8024 2848 8076 2854
rect 8024 2790 8076 2796
rect 8220 2650 8248 2858
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 9048 2582 9076 2994
rect 9968 2922 9996 3062
rect 10428 3058 10456 3402
rect 10416 3052 10468 3058
rect 10416 2994 10468 3000
rect 9956 2916 10008 2922
rect 9956 2858 10008 2864
rect 10140 2848 10192 2854
rect 10140 2790 10192 2796
rect 9036 2576 9088 2582
rect 9036 2518 9088 2524
rect 10152 2446 10180 2790
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 11532 2650 11560 18022
rect 11624 15638 11652 23054
rect 11796 20256 11848 20262
rect 11796 20198 11848 20204
rect 11808 19854 11836 20198
rect 11888 19984 11940 19990
rect 11888 19926 11940 19932
rect 11796 19848 11848 19854
rect 11796 19790 11848 19796
rect 11900 19446 11928 19926
rect 11888 19440 11940 19446
rect 11888 19382 11940 19388
rect 11796 17876 11848 17882
rect 12268 17864 12296 27520
rect 13728 23520 13780 23526
rect 13728 23462 13780 23468
rect 12348 20392 12400 20398
rect 12348 20334 12400 20340
rect 12360 19378 12388 20334
rect 12900 20256 12952 20262
rect 12900 20198 12952 20204
rect 12808 19848 12860 19854
rect 12808 19790 12860 19796
rect 12624 19712 12676 19718
rect 12624 19654 12676 19660
rect 12636 19378 12664 19654
rect 12820 19378 12848 19790
rect 12348 19372 12400 19378
rect 12348 19314 12400 19320
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 12808 19372 12860 19378
rect 12808 19314 12860 19320
rect 12532 19168 12584 19174
rect 12532 19110 12584 19116
rect 12544 18970 12572 19110
rect 12532 18964 12584 18970
rect 12532 18906 12584 18912
rect 12636 18698 12664 19314
rect 12912 18902 12940 20198
rect 13452 19916 13504 19922
rect 13452 19858 13504 19864
rect 13464 19514 13492 19858
rect 13452 19508 13504 19514
rect 13452 19450 13504 19456
rect 13464 19174 13492 19450
rect 13452 19168 13504 19174
rect 13452 19110 13504 19116
rect 12900 18896 12952 18902
rect 12900 18838 12952 18844
rect 12992 18896 13044 18902
rect 12992 18838 13044 18844
rect 12624 18692 12676 18698
rect 12624 18634 12676 18640
rect 12636 18290 12664 18634
rect 12624 18284 12676 18290
rect 12624 18226 12676 18232
rect 12624 18148 12676 18154
rect 12624 18090 12676 18096
rect 12268 17836 12388 17864
rect 11796 17818 11848 17824
rect 11808 17678 11836 17818
rect 12256 17740 12308 17746
rect 12256 17682 12308 17688
rect 11796 17672 11848 17678
rect 11796 17614 11848 17620
rect 11808 17338 11836 17614
rect 12268 17338 12296 17682
rect 11796 17332 11848 17338
rect 11796 17274 11848 17280
rect 12256 17332 12308 17338
rect 12256 17274 12308 17280
rect 11980 17264 12032 17270
rect 11980 17206 12032 17212
rect 11992 16658 12020 17206
rect 12268 17134 12296 17274
rect 12256 17128 12308 17134
rect 12256 17070 12308 17076
rect 11980 16652 12032 16658
rect 11980 16594 12032 16600
rect 11992 16250 12020 16594
rect 11980 16244 12032 16250
rect 11980 16186 12032 16192
rect 11612 15632 11664 15638
rect 11612 15574 11664 15580
rect 11624 14618 11652 15574
rect 12164 14816 12216 14822
rect 12164 14758 12216 14764
rect 11612 14612 11664 14618
rect 11612 14554 11664 14560
rect 12176 14550 12204 14758
rect 12164 14544 12216 14550
rect 12164 14486 12216 14492
rect 12176 13938 12204 14486
rect 12360 14006 12388 17836
rect 12636 17338 12664 18090
rect 12912 17814 12940 18838
rect 13004 18426 13032 18838
rect 12992 18420 13044 18426
rect 12992 18362 13044 18368
rect 12900 17808 12952 17814
rect 12900 17750 12952 17756
rect 13004 17746 13032 18362
rect 12992 17740 13044 17746
rect 12992 17682 13044 17688
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 13452 17672 13504 17678
rect 13452 17614 13504 17620
rect 13464 17338 13492 17614
rect 12624 17332 12676 17338
rect 12624 17274 12676 17280
rect 13452 17332 13504 17338
rect 13452 17274 13504 17280
rect 13556 17202 13584 17682
rect 13544 17196 13596 17202
rect 13544 17138 13596 17144
rect 12808 15632 12860 15638
rect 12808 15574 12860 15580
rect 12532 15496 12584 15502
rect 12532 15438 12584 15444
rect 12440 14884 12492 14890
rect 12440 14826 12492 14832
rect 12452 14550 12480 14826
rect 12440 14544 12492 14550
rect 12440 14486 12492 14492
rect 12452 14074 12480 14486
rect 12544 14414 12572 15438
rect 12820 15366 12848 15574
rect 13360 15496 13412 15502
rect 13360 15438 13412 15444
rect 12808 15360 12860 15366
rect 12808 15302 12860 15308
rect 12820 14958 12848 15302
rect 13372 15162 13400 15438
rect 13360 15156 13412 15162
rect 13360 15098 13412 15104
rect 12808 14952 12860 14958
rect 12808 14894 12860 14900
rect 13176 14476 13228 14482
rect 13176 14418 13228 14424
rect 12532 14408 12584 14414
rect 12532 14350 12584 14356
rect 13188 14074 13216 14418
rect 13636 14408 13688 14414
rect 13636 14350 13688 14356
rect 13648 14074 13676 14350
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 13636 14068 13688 14074
rect 13636 14010 13688 14016
rect 12348 14000 12400 14006
rect 12348 13942 12400 13948
rect 12164 13932 12216 13938
rect 12164 13874 12216 13880
rect 12532 13864 12584 13870
rect 12532 13806 12584 13812
rect 12544 13462 12572 13806
rect 13188 13462 13216 14010
rect 13648 13734 13676 14010
rect 13740 13938 13768 23462
rect 13924 20602 13952 27520
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15488 23866 15516 27520
rect 15476 23860 15528 23866
rect 15476 23802 15528 23808
rect 17144 23633 17172 27520
rect 18800 23866 18828 27520
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 20456 24857 20484 27520
rect 20442 24848 20498 24857
rect 20442 24783 20498 24792
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 20628 24064 20680 24070
rect 20628 24006 20680 24012
rect 18788 23860 18840 23866
rect 18788 23802 18840 23808
rect 17130 23624 17186 23633
rect 17130 23559 17186 23568
rect 15752 23520 15804 23526
rect 15752 23462 15804 23468
rect 19984 23520 20036 23526
rect 19984 23462 20036 23468
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15568 22432 15620 22438
rect 15568 22374 15620 22380
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 13912 20596 13964 20602
rect 13912 20538 13964 20544
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 15384 17740 15436 17746
rect 15384 17682 15436 17688
rect 14556 17536 14608 17542
rect 14556 17478 14608 17484
rect 13728 13932 13780 13938
rect 13728 13874 13780 13880
rect 14372 13796 14424 13802
rect 14372 13738 14424 13744
rect 13636 13728 13688 13734
rect 13636 13670 13688 13676
rect 14384 13462 14412 13738
rect 14464 13728 14516 13734
rect 14464 13670 14516 13676
rect 11980 13456 12032 13462
rect 11980 13398 12032 13404
rect 12532 13456 12584 13462
rect 12532 13398 12584 13404
rect 13176 13456 13228 13462
rect 13176 13398 13228 13404
rect 14372 13456 14424 13462
rect 14372 13398 14424 13404
rect 11886 13288 11942 13297
rect 11886 13223 11942 13232
rect 11900 12170 11928 13223
rect 11992 12646 12020 13398
rect 12256 13388 12308 13394
rect 12256 13330 12308 13336
rect 12268 13297 12296 13330
rect 12440 13320 12492 13326
rect 12254 13288 12310 13297
rect 12440 13262 12492 13268
rect 12254 13223 12310 13232
rect 12452 12850 12480 13262
rect 13188 12986 13216 13398
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13176 12980 13228 12986
rect 13176 12922 13228 12928
rect 12440 12844 12492 12850
rect 12440 12786 12492 12792
rect 11980 12640 12032 12646
rect 11980 12582 12032 12588
rect 12256 12640 12308 12646
rect 12256 12582 12308 12588
rect 11992 12306 12020 12582
rect 11980 12300 12032 12306
rect 11980 12242 12032 12248
rect 11888 12164 11940 12170
rect 11888 12106 11940 12112
rect 12164 11688 12216 11694
rect 12164 11630 12216 11636
rect 12176 11218 12204 11630
rect 12268 11558 12296 12582
rect 12452 12442 12480 12786
rect 13740 12442 13768 13262
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 14188 12708 14240 12714
rect 14188 12650 14240 12656
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 12820 11898 12848 12174
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 13832 11830 13860 12242
rect 13820 11824 13872 11830
rect 13820 11766 13872 11772
rect 12624 11688 12676 11694
rect 12624 11630 12676 11636
rect 12256 11552 12308 11558
rect 12256 11494 12308 11500
rect 12636 11286 12664 11630
rect 12808 11620 12860 11626
rect 12808 11562 12860 11568
rect 12624 11280 12676 11286
rect 12624 11222 12676 11228
rect 12820 11218 12848 11562
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13464 11286 13492 11494
rect 13452 11280 13504 11286
rect 13452 11222 13504 11228
rect 12164 11212 12216 11218
rect 12164 11154 12216 11160
rect 12808 11212 12860 11218
rect 12808 11154 12860 11160
rect 12176 10810 12204 11154
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12636 10130 12664 10474
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 11612 10124 11664 10130
rect 11612 10066 11664 10072
rect 12624 10124 12676 10130
rect 12624 10066 12676 10072
rect 11624 9722 11652 10066
rect 11612 9716 11664 9722
rect 11612 9658 11664 9664
rect 11624 9110 11652 9658
rect 12636 9654 12664 10066
rect 12728 9926 12756 10406
rect 12820 10266 12848 11154
rect 13084 11008 13136 11014
rect 13084 10950 13136 10956
rect 13096 10538 13124 10950
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 13084 10532 13136 10538
rect 13084 10474 13136 10480
rect 12808 10260 12860 10266
rect 12808 10202 12860 10208
rect 12992 10056 13044 10062
rect 12992 9998 13044 10004
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12624 9648 12676 9654
rect 12624 9590 12676 9596
rect 12728 9586 12756 9862
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 11980 9444 12032 9450
rect 11980 9386 12032 9392
rect 11612 9104 11664 9110
rect 11664 9064 11836 9092
rect 11612 9046 11664 9052
rect 11612 8968 11664 8974
rect 11664 8945 11744 8956
rect 11664 8936 11758 8945
rect 11664 8928 11702 8936
rect 11612 8910 11664 8916
rect 11702 8871 11758 8880
rect 11808 8634 11836 9064
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11900 8566 11928 8978
rect 11888 8560 11940 8566
rect 11888 8502 11940 8508
rect 11992 8022 12020 9386
rect 12452 9110 12480 9454
rect 12440 9104 12492 9110
rect 12440 9046 12492 9052
rect 13004 9042 13032 9998
rect 12992 9036 13044 9042
rect 12992 8978 13044 8984
rect 12716 8356 12768 8362
rect 12716 8298 12768 8304
rect 11980 8016 12032 8022
rect 11980 7958 12032 7964
rect 11992 7546 12020 7958
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 11992 7342 12020 7482
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 11980 7336 12032 7342
rect 11980 7278 12032 7284
rect 11992 5846 12020 7278
rect 12256 7268 12308 7274
rect 12256 7210 12308 7216
rect 11980 5840 12032 5846
rect 11980 5782 12032 5788
rect 12268 5778 12296 7210
rect 12452 7002 12480 7346
rect 12728 7002 12756 8298
rect 13004 8090 13032 8978
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 13096 8022 13124 10474
rect 13280 8566 13308 10610
rect 13464 10470 13492 11222
rect 14200 10810 14228 12650
rect 14292 11898 14320 12718
rect 14476 12102 14504 13670
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14280 11892 14332 11898
rect 14280 11834 14332 11840
rect 14292 11558 14320 11834
rect 14464 11756 14516 11762
rect 14464 11698 14516 11704
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 14476 11286 14504 11698
rect 14464 11280 14516 11286
rect 14464 11222 14516 11228
rect 14188 10804 14240 10810
rect 14188 10746 14240 10752
rect 14200 10470 14228 10746
rect 14372 10532 14424 10538
rect 14372 10474 14424 10480
rect 13452 10464 13504 10470
rect 13452 10406 13504 10412
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 13464 10198 13492 10406
rect 14384 10266 14412 10474
rect 14372 10260 14424 10266
rect 14372 10202 14424 10208
rect 13452 10192 13504 10198
rect 13452 10134 13504 10140
rect 13464 9450 13492 10134
rect 13728 9988 13780 9994
rect 13728 9930 13780 9936
rect 13544 9920 13596 9926
rect 13544 9862 13596 9868
rect 13452 9444 13504 9450
rect 13452 9386 13504 9392
rect 13360 9376 13412 9382
rect 13360 9318 13412 9324
rect 13268 8560 13320 8566
rect 13268 8502 13320 8508
rect 13372 8362 13400 9318
rect 13464 9110 13492 9386
rect 13452 9104 13504 9110
rect 13452 9046 13504 9052
rect 13464 8634 13492 9046
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13360 8356 13412 8362
rect 13360 8298 13412 8304
rect 13084 8016 13136 8022
rect 13084 7958 13136 7964
rect 13372 7954 13400 8298
rect 13360 7948 13412 7954
rect 13360 7890 13412 7896
rect 13176 7744 13228 7750
rect 13176 7686 13228 7692
rect 12440 6996 12492 7002
rect 12440 6938 12492 6944
rect 12716 6996 12768 7002
rect 12716 6938 12768 6944
rect 12256 5772 12308 5778
rect 12256 5714 12308 5720
rect 12268 5370 12296 5714
rect 12532 5704 12584 5710
rect 12532 5646 12584 5652
rect 12256 5364 12308 5370
rect 12256 5306 12308 5312
rect 12544 5234 12572 5646
rect 12728 5302 12756 6938
rect 13188 6458 13216 7686
rect 13372 7546 13400 7890
rect 13360 7540 13412 7546
rect 13360 7482 13412 7488
rect 13360 7200 13412 7206
rect 13360 7142 13412 7148
rect 13372 6934 13400 7142
rect 13360 6928 13412 6934
rect 13360 6870 13412 6876
rect 13452 6724 13504 6730
rect 13452 6666 13504 6672
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 13188 6186 13216 6394
rect 13464 6322 13492 6666
rect 13452 6316 13504 6322
rect 13452 6258 13504 6264
rect 13176 6180 13228 6186
rect 13176 6122 13228 6128
rect 12992 5840 13044 5846
rect 12992 5782 13044 5788
rect 13004 5370 13032 5782
rect 13176 5568 13228 5574
rect 13176 5510 13228 5516
rect 13188 5370 13216 5510
rect 12992 5364 13044 5370
rect 12992 5306 13044 5312
rect 13176 5364 13228 5370
rect 13176 5306 13228 5312
rect 12716 5296 12768 5302
rect 12716 5238 12768 5244
rect 12532 5228 12584 5234
rect 12532 5170 12584 5176
rect 12900 4480 12952 4486
rect 12900 4422 12952 4428
rect 11520 2644 11572 2650
rect 11520 2586 11572 2592
rect 11796 2508 11848 2514
rect 11796 2450 11848 2456
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 8576 2304 8628 2310
rect 8576 2246 8628 2252
rect 6918 54 7236 82
rect 7654 96 7710 105
rect 5354 0 5410 54
rect 6918 0 6974 54
rect 7654 31 7710 40
rect 8482 82 8538 480
rect 8588 82 8616 2246
rect 9876 1329 9904 2382
rect 9862 1320 9918 1329
rect 9862 1255 9918 1264
rect 8482 54 8616 82
rect 10046 82 10102 480
rect 10336 82 10364 2382
rect 11808 2310 11836 2450
rect 11796 2304 11848 2310
rect 11796 2246 11848 2252
rect 10046 54 10364 82
rect 11610 82 11666 480
rect 11808 82 11836 2246
rect 11610 54 11836 82
rect 12912 82 12940 4422
rect 13188 4282 13216 5306
rect 13176 4276 13228 4282
rect 13176 4218 13228 4224
rect 13188 4078 13216 4218
rect 13176 4072 13228 4078
rect 13176 4014 13228 4020
rect 13556 2650 13584 9862
rect 13740 9722 13768 9930
rect 14384 9926 14412 10202
rect 14372 9920 14424 9926
rect 14372 9862 14424 9868
rect 13728 9716 13780 9722
rect 13728 9658 13780 9664
rect 13912 9444 13964 9450
rect 13912 9386 13964 9392
rect 13924 9178 13952 9386
rect 13912 9172 13964 9178
rect 13912 9114 13964 9120
rect 14278 8936 14334 8945
rect 14278 8871 14334 8880
rect 14292 8838 14320 8871
rect 14280 8832 14332 8838
rect 14280 8774 14332 8780
rect 14372 8832 14424 8838
rect 14372 8774 14424 8780
rect 14280 8356 14332 8362
rect 14384 8344 14412 8774
rect 14332 8316 14412 8344
rect 14464 8356 14516 8362
rect 14280 8298 14332 8304
rect 14464 8298 14516 8304
rect 14292 7857 14320 8298
rect 14476 8022 14504 8298
rect 14568 8090 14596 17478
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15396 17202 15424 17682
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 15396 17105 15424 17138
rect 15382 17096 15438 17105
rect 15382 17031 15438 17040
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15292 14272 15344 14278
rect 15292 14214 15344 14220
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15304 13394 15332 14214
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15304 12986 15332 13330
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15384 12640 15436 12646
rect 15384 12582 15436 12588
rect 15292 12436 15344 12442
rect 15292 12378 15344 12384
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14832 11756 14884 11762
rect 14832 11698 14884 11704
rect 14844 10742 14872 11698
rect 15304 11558 15332 12378
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 15304 11354 15332 11494
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15396 11286 15424 12582
rect 15476 12232 15528 12238
rect 15476 12174 15528 12180
rect 15488 11762 15516 12174
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 15476 11620 15528 11626
rect 15476 11562 15528 11568
rect 15488 11286 15516 11562
rect 15384 11280 15436 11286
rect 15384 11222 15436 11228
rect 15476 11280 15528 11286
rect 15476 11222 15528 11228
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15396 10810 15424 11222
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15488 10742 15516 11222
rect 14832 10736 14884 10742
rect 14832 10678 14884 10684
rect 15476 10736 15528 10742
rect 15476 10678 15528 10684
rect 14832 10192 14884 10198
rect 14832 10134 14884 10140
rect 14844 9722 14872 10134
rect 15580 10062 15608 22374
rect 15764 16697 15792 23462
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 15844 22568 15896 22574
rect 15842 22536 15844 22545
rect 15896 22536 15898 22545
rect 15842 22471 15898 22480
rect 15856 22438 15884 22471
rect 15844 22432 15896 22438
rect 15844 22374 15896 22380
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 17132 20256 17184 20262
rect 17132 20198 17184 20204
rect 17144 19281 17172 20198
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 17130 19272 17186 19281
rect 17130 19207 17186 19216
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 15750 16688 15806 16697
rect 15750 16623 15806 16632
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19248 14816 19300 14822
rect 19248 14758 19300 14764
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 15672 14074 15700 14350
rect 15660 14068 15712 14074
rect 15660 14010 15712 14016
rect 15752 13252 15804 13258
rect 15752 13194 15804 13200
rect 15764 10810 15792 13194
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15752 10804 15804 10810
rect 15752 10746 15804 10752
rect 15568 10056 15620 10062
rect 15568 9998 15620 10004
rect 15292 9988 15344 9994
rect 15292 9930 15344 9936
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14832 9716 14884 9722
rect 14832 9658 14884 9664
rect 14556 8084 14608 8090
rect 14556 8026 14608 8032
rect 14464 8016 14516 8022
rect 14464 7958 14516 7964
rect 14278 7848 14334 7857
rect 14278 7783 14334 7792
rect 14568 7562 14596 8026
rect 14844 7954 14872 9658
rect 15304 9586 15332 9930
rect 15580 9722 15608 9998
rect 15568 9716 15620 9722
rect 15568 9658 15620 9664
rect 15292 9580 15344 9586
rect 15292 9522 15344 9528
rect 15304 9450 15332 9522
rect 15292 9444 15344 9450
rect 15292 9386 15344 9392
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15304 8498 15332 9386
rect 15660 9104 15712 9110
rect 15660 9046 15712 9052
rect 15672 8498 15700 9046
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 15660 8492 15712 8498
rect 15660 8434 15712 8440
rect 14832 7948 14884 7954
rect 14832 7890 14884 7896
rect 15384 7948 15436 7954
rect 15384 7890 15436 7896
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14384 7534 14596 7562
rect 15396 7546 15424 7890
rect 15384 7540 15436 7546
rect 14384 7410 14412 7534
rect 15384 7482 15436 7488
rect 14372 7404 14424 7410
rect 14372 7346 14424 7352
rect 14556 7404 14608 7410
rect 14556 7346 14608 7352
rect 14568 6934 14596 7346
rect 14648 7268 14700 7274
rect 14648 7210 14700 7216
rect 14660 6934 14688 7210
rect 13820 6928 13872 6934
rect 13820 6870 13872 6876
rect 14556 6928 14608 6934
rect 14556 6870 14608 6876
rect 14648 6928 14700 6934
rect 14648 6870 14700 6876
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13740 5914 13768 6734
rect 13832 6458 13860 6870
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 14648 6316 14700 6322
rect 14648 6258 14700 6264
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13740 5642 13768 5850
rect 14660 5778 14688 6258
rect 14740 6180 14792 6186
rect 14740 6122 14792 6128
rect 15016 6180 15068 6186
rect 15016 6122 15068 6128
rect 15108 6180 15160 6186
rect 15108 6122 15160 6128
rect 14752 5778 14780 6122
rect 14648 5772 14700 5778
rect 14648 5714 14700 5720
rect 14740 5772 14792 5778
rect 14740 5714 14792 5720
rect 13728 5636 13780 5642
rect 13728 5578 13780 5584
rect 14372 5568 14424 5574
rect 14372 5510 14424 5516
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 13912 5364 13964 5370
rect 13912 5306 13964 5312
rect 13832 5098 13860 5306
rect 13924 5273 13952 5306
rect 14004 5296 14056 5302
rect 13910 5264 13966 5273
rect 14004 5238 14056 5244
rect 13910 5199 13966 5208
rect 13820 5092 13872 5098
rect 13820 5034 13872 5040
rect 13820 4752 13872 4758
rect 13820 4694 13872 4700
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 13740 3738 13768 4558
rect 13832 4010 13860 4694
rect 14016 4622 14044 5238
rect 14384 4690 14412 5510
rect 14568 5137 14596 5510
rect 14660 5302 14688 5714
rect 15028 5710 15056 6122
rect 15120 5846 15148 6122
rect 15108 5840 15160 5846
rect 15108 5782 15160 5788
rect 15016 5704 15068 5710
rect 15016 5646 15068 5652
rect 15476 5636 15528 5642
rect 15476 5578 15528 5584
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15488 5302 15516 5578
rect 14648 5296 14700 5302
rect 14648 5238 14700 5244
rect 15476 5296 15528 5302
rect 15476 5238 15528 5244
rect 14554 5128 14610 5137
rect 14554 5063 14610 5072
rect 14568 5030 14596 5063
rect 14556 5024 14608 5030
rect 14556 4966 14608 4972
rect 14372 4684 14424 4690
rect 14372 4626 14424 4632
rect 15292 4684 15344 4690
rect 15292 4626 15344 4632
rect 14004 4616 14056 4622
rect 14004 4558 14056 4564
rect 14832 4480 14884 4486
rect 14832 4422 14884 4428
rect 13820 4004 13872 4010
rect 13820 3946 13872 3952
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 13740 3505 13768 3674
rect 13726 3496 13782 3505
rect 13726 3431 13782 3440
rect 13544 2644 13596 2650
rect 13544 2586 13596 2592
rect 13174 82 13230 480
rect 12912 54 13230 82
rect 8482 0 8538 54
rect 10046 0 10102 54
rect 11610 0 11666 54
rect 13174 0 13230 54
rect 14738 82 14794 480
rect 14844 82 14872 4422
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15304 4282 15332 4626
rect 15292 4276 15344 4282
rect 15292 4218 15344 4224
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14738 54 14872 82
rect 15856 82 15884 13126
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 16040 11286 16068 12174
rect 17224 12096 17276 12102
rect 17224 12038 17276 12044
rect 17236 11558 17264 12038
rect 17224 11552 17276 11558
rect 17224 11494 17276 11500
rect 16028 11280 16080 11286
rect 16028 11222 16080 11228
rect 16856 11212 16908 11218
rect 16856 11154 16908 11160
rect 16868 10810 16896 11154
rect 16856 10804 16908 10810
rect 16856 10746 16908 10752
rect 15936 9444 15988 9450
rect 15936 9386 15988 9392
rect 15948 9110 15976 9386
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 16764 9376 16816 9382
rect 16764 9318 16816 9324
rect 15936 9104 15988 9110
rect 15936 9046 15988 9052
rect 16316 8430 16344 9318
rect 16776 8974 16804 9318
rect 17132 9036 17184 9042
rect 17132 8978 17184 8984
rect 16764 8968 16816 8974
rect 16764 8910 16816 8916
rect 16776 8634 16804 8910
rect 17144 8634 17172 8978
rect 17316 8832 17368 8838
rect 17236 8809 17316 8820
rect 17222 8800 17316 8809
rect 17278 8792 17316 8800
rect 17316 8774 17368 8780
rect 17222 8735 17278 8744
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 16304 8424 16356 8430
rect 16304 8366 16356 8372
rect 16316 8090 16344 8366
rect 16304 8084 16356 8090
rect 16304 8026 16356 8032
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 15948 6458 15976 6802
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 16028 5772 16080 5778
rect 16028 5714 16080 5720
rect 16040 5302 16068 5714
rect 16028 5296 16080 5302
rect 16028 5238 16080 5244
rect 17500 5092 17552 5098
rect 17500 5034 17552 5040
rect 16210 82 16266 480
rect 15856 54 16266 82
rect 17512 82 17540 5034
rect 18788 2916 18840 2922
rect 18788 2858 18840 2864
rect 18800 2514 18828 2858
rect 19260 2582 19288 14758
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19996 11830 20024 23462
rect 20640 21457 20668 24006
rect 20626 21448 20682 21457
rect 20626 21383 20682 21392
rect 22112 20602 22140 27520
rect 22192 24132 22244 24138
rect 22192 24074 22244 24080
rect 22100 20596 22152 20602
rect 22100 20538 22152 20544
rect 22204 18737 22232 24074
rect 23768 23866 23796 27520
rect 25134 26208 25190 26217
rect 25134 26143 25190 26152
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 23940 24336 23992 24342
rect 23940 24278 23992 24284
rect 23952 23866 23980 24278
rect 25148 24274 25176 26143
rect 25424 24342 25452 27520
rect 25412 24336 25464 24342
rect 25412 24278 25464 24284
rect 25136 24268 25188 24274
rect 25136 24210 25188 24216
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 25148 23866 25176 24210
rect 27080 23866 27108 27520
rect 27618 24168 27674 24177
rect 27618 24103 27674 24112
rect 23756 23860 23808 23866
rect 23756 23802 23808 23808
rect 23940 23860 23992 23866
rect 23940 23802 23992 23808
rect 25136 23860 25188 23866
rect 25136 23802 25188 23808
rect 27068 23860 27120 23866
rect 27068 23802 27120 23808
rect 23940 23520 23992 23526
rect 23940 23462 23992 23468
rect 23952 22137 23980 23462
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 27632 22545 27660 24103
rect 27618 22536 27674 22545
rect 27618 22471 27674 22480
rect 23938 22128 23994 22137
rect 23938 22063 23994 22072
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 25134 21040 25190 21049
rect 25134 20975 25190 20984
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 25148 20602 25176 20975
rect 25136 20596 25188 20602
rect 25136 20538 25188 20544
rect 25148 20398 25176 20538
rect 25136 20392 25188 20398
rect 25136 20334 25188 20340
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 27618 19136 27674 19145
rect 27618 19071 27674 19080
rect 22190 18728 22246 18737
rect 22190 18663 22246 18672
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 27632 17105 27660 19071
rect 27618 17096 27674 17105
rect 27618 17031 27674 17040
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 25134 16008 25190 16017
rect 25134 15943 25190 15952
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 25148 15162 25176 15943
rect 25136 15156 25188 15162
rect 25136 15098 25188 15104
rect 25148 14958 25176 15098
rect 25136 14952 25188 14958
rect 25136 14894 25188 14900
rect 24216 14816 24268 14822
rect 24216 14758 24268 14764
rect 19984 11824 20036 11830
rect 19984 11766 20036 11772
rect 19432 11552 19484 11558
rect 19432 11494 19484 11500
rect 19248 2576 19300 2582
rect 19248 2518 19300 2524
rect 18788 2508 18840 2514
rect 18788 2450 18840 2456
rect 17774 82 17830 480
rect 17512 54 17830 82
rect 14738 0 14794 54
rect 16210 0 16266 54
rect 17774 0 17830 54
rect 19338 82 19394 480
rect 19444 82 19472 11494
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 20260 11008 20312 11014
rect 20260 10950 20312 10956
rect 20272 10849 20300 10950
rect 20258 10840 20314 10849
rect 20258 10775 20314 10784
rect 24122 10840 24178 10849
rect 24122 10775 24178 10784
rect 24136 10606 24164 10775
rect 24124 10600 24176 10606
rect 24124 10542 24176 10548
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 24228 10282 24256 14758
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24858 13696 24914 13705
rect 24858 13631 24914 13640
rect 24584 13524 24636 13530
rect 24584 13466 24636 13472
rect 24596 13433 24624 13466
rect 24582 13424 24638 13433
rect 24872 13394 24900 13631
rect 24582 13359 24638 13368
rect 24860 13388 24912 13394
rect 24860 13330 24912 13336
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24872 12986 24900 13330
rect 24860 12980 24912 12986
rect 24860 12922 24912 12928
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 25134 10976 25190 10985
rect 24289 10908 24585 10928
rect 25134 10911 25190 10920
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 25148 10810 25176 10911
rect 25136 10804 25188 10810
rect 25136 10746 25188 10752
rect 24228 10254 24348 10282
rect 24216 10192 24268 10198
rect 24216 10134 24268 10140
rect 24228 9586 24256 10134
rect 24320 10062 24348 10254
rect 24308 10056 24360 10062
rect 24308 9998 24360 10004
rect 25044 10056 25096 10062
rect 25044 9998 25096 10004
rect 24768 9988 24820 9994
rect 24768 9930 24820 9936
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24216 9580 24268 9586
rect 24216 9522 24268 9528
rect 24032 9376 24084 9382
rect 24032 9318 24084 9324
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 24044 9092 24072 9318
rect 24124 9104 24176 9110
rect 24044 9064 24124 9092
rect 24044 8294 24072 9064
rect 24124 9046 24176 9052
rect 24780 9042 24808 9930
rect 25056 9722 25084 9998
rect 25044 9716 25096 9722
rect 25044 9658 25096 9664
rect 24768 9036 24820 9042
rect 24768 8978 24820 8984
rect 24780 8945 24808 8978
rect 24860 8968 24912 8974
rect 24766 8936 24822 8945
rect 24860 8910 24912 8916
rect 24766 8871 24822 8880
rect 24122 8800 24178 8809
rect 24122 8735 24178 8744
rect 24136 8430 24164 8735
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24766 8664 24822 8673
rect 24766 8599 24822 8608
rect 24780 8566 24808 8599
rect 24768 8560 24820 8566
rect 24768 8502 24820 8508
rect 24124 8424 24176 8430
rect 24124 8366 24176 8372
rect 24872 8294 24900 8910
rect 24032 8288 24084 8294
rect 24032 8230 24084 8236
rect 24860 8288 24912 8294
rect 24860 8230 24912 8236
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 24044 7993 24072 8230
rect 24030 7984 24086 7993
rect 24030 7919 24086 7928
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24872 7546 24900 8230
rect 24860 7540 24912 7546
rect 24860 7482 24912 7488
rect 25136 7200 25188 7206
rect 25136 7142 25188 7148
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 25148 6905 25176 7142
rect 25134 6896 25190 6905
rect 25134 6831 25190 6840
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 23662 5128 23718 5137
rect 23662 5063 23718 5072
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 23676 4826 23704 5063
rect 23756 5024 23808 5030
rect 23756 4966 23808 4972
rect 23664 4820 23716 4826
rect 23664 4762 23716 4768
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 22560 2372 22612 2378
rect 22560 2314 22612 2320
rect 20628 2304 20680 2310
rect 20628 2246 20680 2252
rect 20720 2304 20772 2310
rect 20720 2246 20772 2252
rect 19338 54 19472 82
rect 20640 82 20668 2246
rect 20732 1329 20760 2246
rect 20718 1320 20774 1329
rect 20718 1255 20774 1264
rect 20902 82 20958 480
rect 20640 54 20958 82
rect 19338 0 19394 54
rect 20902 0 20958 54
rect 22466 82 22522 480
rect 22572 82 22600 2314
rect 22466 54 22600 82
rect 23768 82 23796 4966
rect 23940 4684 23992 4690
rect 23940 4626 23992 4632
rect 23952 3942 23980 4626
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 23940 3936 23992 3942
rect 23940 3878 23992 3884
rect 24032 3936 24084 3942
rect 24032 3878 24084 3884
rect 27620 3936 27672 3942
rect 27620 3878 27672 3884
rect 23952 2650 23980 3878
rect 24044 3505 24072 3878
rect 27632 3777 27660 3878
rect 27618 3768 27674 3777
rect 27618 3703 27674 3712
rect 24030 3496 24086 3505
rect 24030 3431 24086 3440
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 23940 2644 23992 2650
rect 23940 2586 23992 2592
rect 25228 2644 25280 2650
rect 25228 2586 25280 2592
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24030 82 24086 480
rect 23768 54 24086 82
rect 25240 82 25268 2586
rect 26884 2304 26936 2310
rect 26884 2246 26936 2252
rect 25594 82 25650 480
rect 25240 54 25650 82
rect 26896 82 26924 2246
rect 27618 1320 27674 1329
rect 27618 1255 27674 1264
rect 27158 82 27214 480
rect 27632 105 27660 1255
rect 26896 54 27214 82
rect 22466 0 22522 54
rect 24030 0 24086 54
rect 25594 0 25650 54
rect 27158 0 27214 54
rect 27618 96 27674 105
rect 27618 31 27674 40
<< via2 >>
rect 1490 26560 1546 26616
rect 1582 24792 1638 24848
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 1122 21256 1178 21312
rect 1306 19488 1362 19544
rect 110 18264 166 18320
rect 1490 15952 1546 16008
rect 1582 14456 1638 14512
rect 110 13096 166 13152
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5998 21392 6054 21448
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 2318 13232 2374 13288
rect 110 9560 166 9616
rect 110 7792 166 7848
rect 110 6024 166 6080
rect 1582 10784 1638 10840
rect 2134 12552 2190 12608
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 3146 9424 3202 9480
rect 3054 7384 3110 7440
rect 4158 16632 4214 16688
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 3790 9288 3846 9344
rect 2778 4800 2834 4856
rect 1766 2896 1822 2952
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 4342 9560 4398 9616
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5538 13640 5594 13696
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 8206 23568 8262 23624
rect 8850 18672 8906 18728
rect 7102 9968 7158 10024
rect 7194 9288 7250 9344
rect 7470 9696 7526 9752
rect 7470 9424 7526 9480
rect 7930 10004 7932 10024
rect 7932 10004 7984 10024
rect 7984 10004 7986 10024
rect 7930 9968 7986 10004
rect 7930 9696 7986 9752
rect 8574 13640 8630 13696
rect 9126 13640 9182 13696
rect 8850 13368 8906 13424
rect 8850 12552 8906 12608
rect 8206 9424 8262 9480
rect 9862 23024 9918 23080
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 11610 24792 11666 24848
rect 10322 22072 10378 22128
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10874 19216 10930 19272
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 8942 7792 8998 7848
rect 8758 7384 8814 7440
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 11426 7928 11482 7984
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 4618 1400 4674 1456
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10782 5208 10838 5264
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 20442 24792 20498 24848
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 17130 23568 17186 23624
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 11886 13232 11942 13288
rect 12254 13232 12310 13288
rect 11702 8880 11758 8936
rect 7654 40 7710 96
rect 9862 1264 9918 1320
rect 14278 8880 14334 8936
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 15382 17040 15438 17096
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 15842 22516 15844 22536
rect 15844 22516 15896 22536
rect 15896 22516 15898 22536
rect 15842 22480 15898 22516
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 17130 19216 17186 19272
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 15750 16632 15806 16688
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14278 7792 14334 7848
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 13910 5208 13966 5264
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14554 5072 14610 5128
rect 13726 3440 13782 3496
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 17222 8744 17278 8800
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 20626 21392 20682 21448
rect 25134 26152 25190 26208
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 27618 24112 27674 24168
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 27618 22480 27674 22536
rect 23938 22072 23994 22128
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 25134 20984 25190 21040
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 27618 19080 27674 19136
rect 22190 18672 22246 18728
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 27618 17040 27674 17096
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 25134 15952 25190 16008
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 20258 10784 20314 10840
rect 24122 10784 24178 10840
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24858 13640 24914 13696
rect 24582 13368 24638 13424
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 25134 10920 25190 10976
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 24766 8880 24822 8936
rect 24122 8744 24178 8800
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24766 8608 24822 8664
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 24030 7928 24086 7984
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 25134 6840 25190 6896
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 23662 5072 23718 5128
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 20718 1264 20774 1320
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 27618 3712 27674 3768
rect 24030 3440 24086 3496
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 27618 1264 27674 1320
rect 27618 40 27674 96
<< metal3 >>
rect 0 27072 480 27192
rect 62 26618 122 27072
rect 27520 26664 28000 26784
rect 1485 26618 1551 26621
rect 62 26616 1551 26618
rect 62 26560 1490 26616
rect 1546 26560 1551 26616
rect 62 26558 1551 26560
rect 1485 26555 1551 26558
rect 25129 26210 25195 26213
rect 27662 26210 27722 26664
rect 25129 26208 27722 26210
rect 25129 26152 25134 26208
rect 25190 26152 27722 26208
rect 25129 26150 27722 26152
rect 25129 26147 25195 26150
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 0 25304 480 25424
rect 62 24850 122 25304
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 1577 24850 1643 24853
rect 62 24848 1643 24850
rect 62 24792 1582 24848
rect 1638 24792 1643 24848
rect 62 24790 1643 24792
rect 1577 24787 1643 24790
rect 11605 24850 11671 24853
rect 20437 24850 20503 24853
rect 11605 24848 20503 24850
rect 11605 24792 11610 24848
rect 11666 24792 20442 24848
rect 20498 24792 20503 24848
rect 11605 24790 20503 24792
rect 11605 24787 11671 24790
rect 20437 24787 20503 24790
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 27520 24168 28000 24200
rect 27520 24112 27618 24168
rect 27674 24112 28000 24168
rect 27520 24080 28000 24112
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 0 23536 480 23656
rect 8201 23626 8267 23629
rect 17125 23626 17191 23629
rect 8201 23624 17191 23626
rect 8201 23568 8206 23624
rect 8262 23568 17130 23624
rect 17186 23568 17191 23624
rect 8201 23566 17191 23568
rect 8201 23563 8267 23566
rect 17125 23563 17191 23566
rect 62 23082 122 23536
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 9857 23082 9923 23085
rect 62 23080 9923 23082
rect 62 23024 9862 23080
rect 9918 23024 9923 23080
rect 62 23022 9923 23024
rect 9857 23019 9923 23022
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 15837 22538 15903 22541
rect 27613 22538 27679 22541
rect 15837 22536 27679 22538
rect 15837 22480 15842 22536
rect 15898 22480 27618 22536
rect 27674 22480 27679 22536
rect 15837 22478 27679 22480
rect 15837 22475 15903 22478
rect 27613 22475 27679 22478
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 10317 22130 10383 22133
rect 23933 22130 23999 22133
rect 10317 22128 23999 22130
rect 10317 22072 10322 22128
rect 10378 22072 23938 22128
rect 23994 22072 23999 22128
rect 10317 22070 23999 22072
rect 10317 22067 10383 22070
rect 23933 22067 23999 22070
rect 0 21768 480 21888
rect 5610 21792 5930 21793
rect 62 21314 122 21768
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 27520 21496 28000 21616
rect 5993 21450 6059 21453
rect 20621 21450 20687 21453
rect 5993 21448 20687 21450
rect 5993 21392 5998 21448
rect 6054 21392 20626 21448
rect 20682 21392 20687 21448
rect 5993 21390 20687 21392
rect 5993 21387 6059 21390
rect 20621 21387 20687 21390
rect 1117 21314 1183 21317
rect 62 21312 1183 21314
rect 62 21256 1122 21312
rect 1178 21256 1183 21312
rect 62 21254 1183 21256
rect 1117 21251 1183 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 25129 21042 25195 21045
rect 27662 21042 27722 21496
rect 25129 21040 27722 21042
rect 25129 20984 25134 21040
rect 25190 20984 27722 21040
rect 25129 20982 27722 20984
rect 25129 20979 25195 20982
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 10277 20160 10597 20161
rect 0 20000 480 20120
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 62 19546 122 20000
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 1301 19546 1367 19549
rect 62 19544 1367 19546
rect 62 19488 1306 19544
rect 1362 19488 1367 19544
rect 62 19486 1367 19488
rect 1301 19483 1367 19486
rect 10869 19274 10935 19277
rect 17125 19274 17191 19277
rect 10869 19272 17191 19274
rect 10869 19216 10874 19272
rect 10930 19216 17130 19272
rect 17186 19216 17191 19272
rect 10869 19214 17191 19216
rect 10869 19211 10935 19214
rect 17125 19211 17191 19214
rect 27520 19136 28000 19168
rect 27520 19080 27618 19136
rect 27674 19080 28000 19136
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 27520 19048 28000 19080
rect 19610 19007 19930 19008
rect 8845 18730 8911 18733
rect 22185 18730 22251 18733
rect 8845 18728 22251 18730
rect 8845 18672 8850 18728
rect 8906 18672 22190 18728
rect 22246 18672 22251 18728
rect 8845 18670 22251 18672
rect 8845 18667 8911 18670
rect 22185 18667 22251 18670
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 0 18320 480 18352
rect 0 18264 110 18320
rect 166 18264 480 18320
rect 0 18232 480 18264
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 15377 17098 15443 17101
rect 27613 17098 27679 17101
rect 15377 17096 27679 17098
rect 15377 17040 15382 17096
rect 15438 17040 27618 17096
rect 27674 17040 27679 17096
rect 15377 17038 27679 17040
rect 15377 17035 15443 17038
rect 27613 17035 27679 17038
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 4153 16690 4219 16693
rect 15745 16690 15811 16693
rect 4153 16688 15811 16690
rect 4153 16632 4158 16688
rect 4214 16632 15750 16688
rect 15806 16632 15811 16688
rect 4153 16630 15811 16632
rect 4153 16627 4219 16630
rect 15745 16627 15811 16630
rect 0 16464 480 16584
rect 27520 16464 28000 16584
rect 62 16010 122 16464
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 1485 16010 1551 16013
rect 62 16008 1551 16010
rect 62 15952 1490 16008
rect 1546 15952 1551 16008
rect 62 15950 1551 15952
rect 1485 15947 1551 15950
rect 25129 16010 25195 16013
rect 27662 16010 27722 16464
rect 25129 16008 27722 16010
rect 25129 15952 25134 16008
rect 25190 15952 27722 16008
rect 25129 15950 27722 15952
rect 25129 15947 25195 15950
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 0 14832 480 14952
rect 62 14514 122 14832
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 1577 14514 1643 14517
rect 62 14512 1643 14514
rect 62 14456 1582 14512
rect 1638 14456 1643 14512
rect 62 14454 1643 14456
rect 1577 14451 1643 14454
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 27520 13880 28000 14000
rect 5533 13698 5599 13701
rect 8569 13698 8635 13701
rect 9121 13698 9187 13701
rect 5533 13696 9187 13698
rect 5533 13640 5538 13696
rect 5594 13640 8574 13696
rect 8630 13640 9126 13696
rect 9182 13640 9187 13696
rect 5533 13638 9187 13640
rect 5533 13635 5599 13638
rect 8569 13635 8635 13638
rect 9121 13635 9187 13638
rect 24853 13698 24919 13701
rect 27662 13698 27722 13880
rect 24853 13696 27722 13698
rect 24853 13640 24858 13696
rect 24914 13640 27722 13696
rect 24853 13638 27722 13640
rect 24853 13635 24919 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 8845 13426 8911 13429
rect 24577 13426 24643 13429
rect 8845 13424 24643 13426
rect 8845 13368 8850 13424
rect 8906 13368 24582 13424
rect 24638 13368 24643 13424
rect 8845 13366 24643 13368
rect 8845 13363 8911 13366
rect 24577 13363 24643 13366
rect 2313 13290 2379 13293
rect 11881 13290 11947 13293
rect 12249 13290 12315 13293
rect 2313 13288 12315 13290
rect 2313 13232 2318 13288
rect 2374 13232 11886 13288
rect 11942 13232 12254 13288
rect 12310 13232 12315 13288
rect 2313 13230 12315 13232
rect 2313 13227 2379 13230
rect 11881 13227 11947 13230
rect 12249 13227 12315 13230
rect 0 13152 480 13184
rect 0 13096 110 13152
rect 166 13096 480 13152
rect 0 13064 480 13096
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 2129 12610 2195 12613
rect 8845 12610 8911 12613
rect 2129 12608 8911 12610
rect 2129 12552 2134 12608
rect 2190 12552 8850 12608
rect 8906 12552 8911 12608
rect 2129 12550 8911 12552
rect 2129 12547 2195 12550
rect 8845 12547 8911 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 10277 11456 10597 11457
rect 0 11296 480 11416
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 27520 11296 28000 11416
rect 62 10842 122 11296
rect 25129 10978 25195 10981
rect 27662 10978 27722 11296
rect 25129 10976 27722 10978
rect 25129 10920 25134 10976
rect 25190 10920 27722 10976
rect 25129 10918 27722 10920
rect 25129 10915 25195 10918
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 1577 10842 1643 10845
rect 62 10840 1643 10842
rect 62 10784 1582 10840
rect 1638 10784 1643 10840
rect 62 10782 1643 10784
rect 1577 10779 1643 10782
rect 20253 10842 20319 10845
rect 24117 10842 24183 10845
rect 20253 10840 24183 10842
rect 20253 10784 20258 10840
rect 20314 10784 24122 10840
rect 24178 10784 24183 10840
rect 20253 10782 24183 10784
rect 20253 10779 20319 10782
rect 24117 10779 24183 10782
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 7097 10026 7163 10029
rect 7925 10026 7991 10029
rect 7097 10024 7991 10026
rect 7097 9968 7102 10024
rect 7158 9968 7930 10024
rect 7986 9968 7991 10024
rect 7097 9966 7991 9968
rect 7097 9963 7163 9966
rect 7925 9963 7991 9966
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 7465 9754 7531 9757
rect 7925 9754 7991 9757
rect 7465 9752 7991 9754
rect 7465 9696 7470 9752
rect 7526 9696 7930 9752
rect 7986 9696 7991 9752
rect 7465 9694 7991 9696
rect 7465 9691 7531 9694
rect 7925 9691 7991 9694
rect 0 9616 480 9648
rect 4337 9618 4403 9621
rect 0 9560 110 9616
rect 166 9560 480 9616
rect 0 9528 480 9560
rect 4294 9616 4403 9618
rect 4294 9560 4342 9616
rect 4398 9560 4403 9616
rect 4294 9555 4403 9560
rect 3141 9482 3207 9485
rect 4294 9482 4354 9555
rect 7465 9482 7531 9485
rect 8201 9482 8267 9485
rect 3141 9480 8267 9482
rect 3141 9424 3146 9480
rect 3202 9424 7470 9480
rect 7526 9424 8206 9480
rect 8262 9424 8267 9480
rect 3141 9422 8267 9424
rect 3141 9419 3207 9422
rect 7465 9419 7531 9422
rect 8201 9419 8267 9422
rect 3785 9346 3851 9349
rect 7189 9346 7255 9349
rect 3785 9344 7255 9346
rect 3785 9288 3790 9344
rect 3846 9288 7194 9344
rect 7250 9288 7255 9344
rect 3785 9286 7255 9288
rect 3785 9283 3851 9286
rect 7189 9283 7255 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 11697 8938 11763 8941
rect 14273 8938 14339 8941
rect 24761 8938 24827 8941
rect 11697 8936 24827 8938
rect 11697 8880 11702 8936
rect 11758 8880 14278 8936
rect 14334 8880 24766 8936
rect 24822 8880 24827 8936
rect 11697 8878 24827 8880
rect 11697 8875 11763 8878
rect 14273 8875 14339 8878
rect 24761 8875 24827 8878
rect 27520 8848 28000 8968
rect 17217 8802 17283 8805
rect 24117 8802 24183 8805
rect 17217 8800 24183 8802
rect 17217 8744 17222 8800
rect 17278 8744 24122 8800
rect 24178 8744 24183 8800
rect 17217 8742 24183 8744
rect 17217 8739 17283 8742
rect 24117 8739 24183 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 24761 8666 24827 8669
rect 27662 8666 27722 8848
rect 24761 8664 27722 8666
rect 24761 8608 24766 8664
rect 24822 8608 27722 8664
rect 24761 8606 27722 8608
rect 24761 8603 24827 8606
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 11421 7986 11487 7989
rect 24025 7986 24091 7989
rect 11421 7984 24091 7986
rect 11421 7928 11426 7984
rect 11482 7928 24030 7984
rect 24086 7928 24091 7984
rect 11421 7926 24091 7928
rect 11421 7923 11487 7926
rect 24025 7923 24091 7926
rect 0 7848 480 7880
rect 0 7792 110 7848
rect 166 7792 480 7848
rect 0 7760 480 7792
rect 8937 7850 9003 7853
rect 14273 7850 14339 7853
rect 8937 7848 14339 7850
rect 8937 7792 8942 7848
rect 8998 7792 14278 7848
rect 14334 7792 14339 7848
rect 8937 7790 14339 7792
rect 8937 7787 9003 7790
rect 14273 7787 14339 7790
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 3049 7442 3115 7445
rect 8753 7442 8819 7445
rect 3049 7440 8819 7442
rect 3049 7384 3054 7440
rect 3110 7384 8758 7440
rect 8814 7384 8819 7440
rect 3049 7382 8819 7384
rect 3049 7379 3115 7382
rect 8753 7379 8819 7382
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 25129 6898 25195 6901
rect 25129 6896 27722 6898
rect 25129 6840 25134 6896
rect 25190 6840 27722 6896
rect 25129 6838 27722 6840
rect 25129 6835 25195 6838
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 27662 6384 27722 6838
rect 27520 6264 28000 6384
rect 0 6080 480 6112
rect 0 6024 110 6080
rect 166 6024 480 6080
rect 0 5992 480 6024
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 10777 5266 10843 5269
rect 13905 5266 13971 5269
rect 10777 5264 13971 5266
rect 10777 5208 10782 5264
rect 10838 5208 13910 5264
rect 13966 5208 13971 5264
rect 10777 5206 13971 5208
rect 10777 5203 10843 5206
rect 13905 5203 13971 5206
rect 14549 5130 14615 5133
rect 23657 5130 23723 5133
rect 14549 5128 23723 5130
rect 14549 5072 14554 5128
rect 14610 5072 23662 5128
rect 23718 5072 23723 5128
rect 14549 5070 23723 5072
rect 14549 5067 14615 5070
rect 23657 5067 23723 5070
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 2773 4858 2839 4861
rect 62 4856 2839 4858
rect 62 4800 2778 4856
rect 2834 4800 2839 4856
rect 62 4798 2839 4800
rect 62 4344 122 4798
rect 2773 4795 2839 4798
rect 5610 4384 5930 4385
rect 0 4224 480 4344
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 27520 3768 28000 3800
rect 27520 3712 27618 3768
rect 27674 3712 28000 3768
rect 27520 3680 28000 3712
rect 13721 3498 13787 3501
rect 24025 3498 24091 3501
rect 13721 3496 24091 3498
rect 13721 3440 13726 3496
rect 13782 3440 24030 3496
rect 24086 3440 24091 3496
rect 13721 3438 24091 3440
rect 13721 3435 13787 3438
rect 24025 3435 24091 3438
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 1761 2954 1827 2957
rect 62 2952 1827 2954
rect 62 2896 1766 2952
rect 1822 2896 1827 2952
rect 62 2894 1827 2896
rect 62 2576 122 2894
rect 1761 2891 1827 2894
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 0 2456 480 2576
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 4613 1458 4679 1461
rect 62 1456 4679 1458
rect 62 1400 4618 1456
rect 4674 1400 4679 1456
rect 62 1398 4679 1400
rect 62 944 122 1398
rect 4613 1395 4679 1398
rect 9857 1322 9923 1325
rect 20713 1322 20779 1325
rect 9857 1320 20779 1322
rect 9857 1264 9862 1320
rect 9918 1264 20718 1320
rect 20774 1264 20779 1320
rect 9857 1262 20779 1264
rect 9857 1259 9923 1262
rect 20713 1259 20779 1262
rect 27520 1320 28000 1352
rect 27520 1264 27618 1320
rect 27674 1264 28000 1320
rect 27520 1232 28000 1264
rect 0 824 480 944
rect 7649 98 7715 101
rect 27613 98 27679 101
rect 7649 96 27679 98
rect 7649 40 7654 96
rect 7710 40 27618 96
rect 27674 40 27679 96
rect 7649 38 27679 40
rect 7649 35 7715 38
rect 27613 35 27679 38
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_39
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5520 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5980 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_51 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_55 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6164 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_8  FILLER_1_51 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_59
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_61 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6716 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_68
timestamp 1586364061
transform 1 0 7360 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_66
timestamp 1586364061
transform 1 0 7176 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7176 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7360 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_12.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8096 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8372 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 7544 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_70
timestamp 1586364061
transform 1 0 7544 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_77
timestamp 1586364061
transform 1 0 8188 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_81
timestamp 1586364061
transform 1 0 8556 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_72
timestamp 1586364061
transform 1 0 7728 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_89
timestamp 1586364061
transform 1 0 9292 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_85
timestamp 1586364061
transform 1 0 8924 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9476 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_12.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_103
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_102
timestamp 1586364061
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_106
timestamp 1586364061
transform 1 0 10856 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_117
timestamp 1586364061
transform 1 0 11868 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_113
timestamp 1586364061
transform 1 0 11500 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_114
timestamp 1586364061
transform 1 0 11592 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11684 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_121
timestamp 1586364061
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_118
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12880 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13340 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_131
timestamp 1586364061
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_135
timestamp 1586364061
transform 1 0 13524 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _237_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 18768 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_4  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_191
timestamp 1586364061
transform 1 0 18676 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _235_
timestamp 1586364061
transform 1 0 19964 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__237__A
timestamp 1586364061
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_200
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_204
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__235__A
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_209
timestamp 1586364061
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_6  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_12.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_258
timestamp 1586364061
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_262
timestamp 1586364061
transform 1 0 25208 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_0_274
timestamp 1586364061
transform 1 0 26312 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 590 592
use scs8hd_inv_8  _185_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8004 0 -1 3808
box -38 -48 866 592
use scs8hd_fill_1  FILLER_2_74
timestamp 1586364061
transform 1 0 7912 0 -1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_103
timestamp 1586364061
transform 1 0 10580 0 -1 3808
box -38 -48 774 592
use scs8hd_conb_1  _219_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11316 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_114
timestamp 1586364061
transform 1 0 11592 0 -1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_126
timestamp 1586364061
transform 1 0 12696 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_2_134
timestamp 1586364061
transform 1 0 13432 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_138
timestamp 1586364061
transform 1 0 13800 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_2_150
timestamp 1586364061
transform 1 0 14904 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_12.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8096 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7544 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_72
timestamp 1586364061
transform 1 0 7728 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _184_
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_87
timestamp 1586364061
transform 1 0 9108 0 1 3808
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10856 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_104
timestamp 1586364061
transform 1 0 10672 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_108
timestamp 1586364061
transform 1 0 11040 0 1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__234__A
timestamp 1586364061
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 774 592
use scs8hd_decap_8  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 774 592
use scs8hd_inv_8  _183_
timestamp 1586364061
transform 1 0 13340 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 13156 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14352 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_142
timestamp 1586364061
transform 1 0 14168 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_146
timestamp 1586364061
transform 1 0 14536 0 1 3808
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__229__A
timestamp 1586364061
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_156
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_168
timestamp 1586364061
transform 1 0 16560 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_3_180
timestamp 1586364061
transform 1 0 17664 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_232
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_249
timestamp 1586364061
transform 1 0 24012 0 1 3808
box -38 -48 590 592
use scs8hd_inv_1  mux_top_track_10.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_258
timestamp 1586364061
transform 1 0 24840 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_262
timestamp 1586364061
transform 1 0 25208 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_3_274
timestamp 1586364061
transform 1 0 26312 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 7452 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8372 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_71
timestamp 1586364061
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_75
timestamp 1586364061
transform 1 0 8004 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_8  FILLER_4_81
timestamp 1586364061
transform 1 0 8556 0 -1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_89
timestamp 1586364061
transform 1 0 9292 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10396 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10120 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_97
timestamp 1586364061
transform 1 0 10028 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_100
timestamp 1586364061
transform 1 0 10304 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_104
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 774 592
use scs8hd_buf_2  _234_
timestamp 1586364061
transform 1 0 11408 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_116
timestamp 1586364061
transform 1 0 11776 0 -1 4896
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_4_128
timestamp 1586364061
transform 1 0 12880 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_8  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 774 592
use scs8hd_buf_2  _229_
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_158
timestamp 1586364061
transform 1 0 15640 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_170
timestamp 1586364061
transform 1 0 16744 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_182
timestamp 1586364061
transform 1 0 17848 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_194
timestamp 1586364061
transform 1 0 18952 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_4_206
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_10.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_6  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 590 592
use scs8hd_decap_12  FILLER_4_248
timestamp 1586364061
transform 1 0 23920 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_260
timestamp 1586364061
transform 1 0 25024 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_272
timestamp 1586364061
transform 1 0 26128 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_55
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 590 592
use scs8hd_buf_1  _098_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7084 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_68
timestamp 1586364061
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_12.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 7544 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_72
timestamp 1586364061
transform 1 0 7728 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_76
timestamp 1586364061
transform 1 0 8096 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9568 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_90
timestamp 1586364061
transform 1 0 9384 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_94
timestamp 1586364061
transform 1 0 9752 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_107
timestamp 1586364061
transform 1 0 10948 0 1 4896
box -38 -48 222 592
use scs8hd_conb_1  _209_
timestamp 1586364061
transform 1 0 12512 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_111
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_5_119
timestamp 1586364061
transform 1 0 12052 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12972 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_127
timestamp 1586364061
transform 1 0 12788 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_131
timestamp 1586364061
transform 1 0 13156 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_145
timestamp 1586364061
transform 1 0 14444 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_149
timestamp 1586364061
transform 1 0 14812 0 1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_11.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15180 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 16008 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_156
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_160
timestamp 1586364061
transform 1 0 15824 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_164
timestamp 1586364061
transform 1 0 16192 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_5_176
timestamp 1586364061
transform 1 0 17296 0 1 4896
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_182
timestamp 1586364061
transform 1 0 17848 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22080 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22540 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_231
timestamp 1586364061
transform 1 0 22356 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_235
timestamp 1586364061
transform 1 0 22724 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_243
timestamp 1586364061
transform 1 0 23460 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_6
timestamp 1586364061
transform 1 0 1656 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_10
timestamp 1586364061
transform 1 0 2024 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_7_14
timestamp 1586364061
transform 1 0 2392 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_26
timestamp 1586364061
transform 1 0 3496 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_40
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 406 592
use scs8hd_buf_1  _097_
timestamp 1586364061
transform 1 0 5980 0 -1 5984
box -38 -48 314 592
use scs8hd_buf_1  _106_
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 5612 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 6072 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_52
timestamp 1586364061
transform 1 0 5888 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_47
timestamp 1586364061
transform 1 0 5428 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 314 592
use scs8hd_nor2_4  _131_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7452 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_8  _191_
timestamp 1586364061
transform 1 0 6900 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_56
timestamp 1586364061
transform 1 0 6256 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8464 0 1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8280 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_78
timestamp 1586364061
transform 1 0 8280 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_82
timestamp 1586364061
transform 1 0 8648 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_72
timestamp 1586364061
transform 1 0 7728 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_76
timestamp 1586364061
transform 1 0 8096 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_86
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_91
timestamp 1586364061
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_95
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 222 592
use scs8hd_conb_1  _208_
timestamp 1586364061
transform 1 0 11224 0 -1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_102
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_106
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_108
timestamp 1586364061
transform 1 0 11040 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_10.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12236 0 -1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_113
timestamp 1586364061
transform 1 0 11500 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_8  FILLER_7_112
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_120
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13156 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_132
timestamp 1586364061
transform 1 0 13248 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_138
timestamp 1586364061
transform 1 0 13800 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_142
timestamp 1586364061
transform 1 0 14168 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_143
timestamp 1586364061
transform 1 0 14260 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14352 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_11.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_146
timestamp 1586364061
transform 1 0 14536 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_152
timestamp 1586364061
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_6_147
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14904 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14720 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14904 0 1 5984
box -38 -48 866 592
use scs8hd_inv_8  _200_
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 15916 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_159
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_163
timestamp 1586364061
transform 1 0 16100 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_175
timestamp 1586364061
transform 1 0 17204 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_187
timestamp 1586364061
transform 1 0 18308 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_199
timestamp 1586364061
transform 1 0 19412 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_6_211
timestamp 1586364061
transform 1 0 20516 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_220
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_232
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_263
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1748 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_10
timestamp 1586364061
transform 1 0 2024 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_8_22
timestamp 1586364061
transform 1 0 3128 0 -1 7072
box -38 -48 774 592
use scs8hd_buf_1  _132_
timestamp 1586364061
transform 1 0 4600 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_30
timestamp 1586364061
transform 1 0 3864 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_8_41
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 1142 592
use scs8hd_buf_1  _122_
timestamp 1586364061
transform 1 0 6072 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_53
timestamp 1586364061
transform 1 0 5980 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 7084 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_57
timestamp 1586364061
transform 1 0 6348 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_67
timestamp 1586364061
transform 1 0 7268 0 -1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_72
timestamp 1586364061
transform 1 0 7728 0 -1 7072
box -38 -48 130 592
use scs8hd_inv_8  _196_
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_88
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_8  _190_
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_107
timestamp 1586364061
transform 1 0 10948 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_119
timestamp 1586364061
transform 1 0 12052 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13340 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_125
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_135
timestamp 1586364061
transform 1 0 13524 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 774 592
use scs8hd_inv_8  _201_
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_163
timestamp 1586364061
transform 1 0 16100 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_175
timestamp 1586364061
transform 1 0 17204 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_187
timestamp 1586364061
transform 1 0 18308 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_199
timestamp 1586364061
transform 1 0 19412 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_211
timestamp 1586364061
transform 1 0 20516 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_263
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1656 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2116 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_9
timestamp 1586364061
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_13
timestamp 1586364061
transform 1 0 2300 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 2944 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_17
timestamp 1586364061
transform 1 0 2668 0 1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_9_22
timestamp 1586364061
transform 1 0 3128 0 1 7072
box -38 -48 774 592
use scs8hd_buf_1  _103_
timestamp 1586364061
transform 1 0 3864 0 1 7072
box -38 -48 314 592
use scs8hd_buf_1  _139_
timestamp 1586364061
transform 1 0 4876 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_33
timestamp 1586364061
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_37
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 5336 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 5704 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_44
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_48
timestamp 1586364061
transform 1 0 5520 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_52
timestamp 1586364061
transform 1 0 5888 0 1 7072
box -38 -48 590 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 7084 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_58
timestamp 1586364061
transform 1 0 6440 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8648 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 8096 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 8464 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_78
timestamp 1586364061
transform 1 0 8280 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_91
timestamp 1586364061
transform 1 0 9476 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_96
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_100
timestamp 1586364061
transform 1 0 10304 0 1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_11.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_134
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_138
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_151
timestamp 1586364061
transform 1 0 14996 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_156
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_168
timestamp 1586364061
transform 1 0 16560 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_9_180
timestamp 1586364061
transform 1 0 17664 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_196
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_208
timestamp 1586364061
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_220
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_232
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_253
timestamp 1586364061
transform 1 0 24380 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_258
timestamp 1586364061
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_262
timestamp 1586364061
transform 1 0 25208 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_9_274
timestamp 1586364061
transform 1 0 26312 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 1840 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_6
timestamp 1586364061
transform 1 0 1656 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_10
timestamp 1586364061
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 2944 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_6  FILLER_10_14
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_8  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 4784 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 4416 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_38
timestamp 1586364061
transform 1 0 4600 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_1  _155_
timestamp 1586364061
transform 1 0 4968 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__163__D
timestamp 1586364061
transform 1 0 5428 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 5796 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_45
timestamp 1586364061
transform 1 0 5244 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_49
timestamp 1586364061
transform 1 0 5612 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_53
timestamp 1586364061
transform 1 0 5980 0 -1 8160
box -38 -48 406 592
use scs8hd_conb_1  _215_
timestamp 1586364061
transform 1 0 6532 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__126__D
timestamp 1586364061
transform 1 0 6992 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 6348 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_62
timestamp 1586364061
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_66
timestamp 1586364061
transform 1 0 7176 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 7544 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 8556 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_79
timestamp 1586364061
transform 1 0 8372 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_83
timestamp 1586364061
transform 1 0 8740 0 -1 8160
box -38 -48 314 592
use scs8hd_nor2_4  _162_
timestamp 1586364061
transform 1 0 9752 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_88
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11132 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_103
timestamp 1586364061
transform 1 0 10580 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_107
timestamp 1586364061
transform 1 0 10948 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_11.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11316 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_10_122
timestamp 1586364061
transform 1 0 12328 0 -1 8160
box -38 -48 314 592
use scs8hd_inv_8  _182_
timestamp 1586364061
transform 1 0 13064 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_127
timestamp 1586364061
transform 1 0 12788 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_139
timestamp 1586364061
transform 1 0 13892 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_143
timestamp 1586364061
transform 1 0 14260 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_147
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 590 592
use scs8hd_inv_8  _177_
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_163
timestamp 1586364061
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_167
timestamp 1586364061
transform 1 0 16468 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_179
timestamp 1586364061
transform 1 0 17572 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_191
timestamp 1586364061
transform 1 0 18676 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_203
timestamp 1586364061
transform 1 0 19780 0 -1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_211
timestamp 1586364061
transform 1 0 20516 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_251
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_263
timestamp 1586364061
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_or2_4  _102_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1564 0 1 8160
box -38 -48 682 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_12
timestamp 1586364061
transform 1 0 2208 0 1 8160
box -38 -48 222 592
use scs8hd_buf_1  _114_
timestamp 1586364061
transform 1 0 3128 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 2392 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 2944 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_16
timestamp 1586364061
transform 1 0 2576 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_25
timestamp 1586364061
transform 1 0 3404 0 1 8160
box -38 -48 222 592
use scs8hd_buf_1  _152_
timestamp 1586364061
transform 1 0 4140 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 4876 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 3956 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_29
timestamp 1586364061
transform 1 0 3772 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_36
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_40
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 130 592
use scs8hd_or4_4  _163_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use scs8hd_fill_1  FILLER_11_43
timestamp 1586364061
transform 1 0 5060 0 1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _145_
timestamp 1586364061
transform 1 0 7268 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 6440 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__C
timestamp 1586364061
transform 1 0 6992 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_60
timestamp 1586364061
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_66
timestamp 1586364061
transform 1 0 7176 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__153__C
timestamp 1586364061
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 8648 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_76
timestamp 1586364061
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_80
timestamp 1586364061
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 866 592
use scs8hd_fill_2  FILLER_11_84
timestamp 1586364061
transform 1 0 8832 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_95
timestamp 1586364061
transform 1 0 9844 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _161_
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_99
timestamp 1586364061
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_112
timestamp 1586364061
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_116
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_120
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_134
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_138
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_151
timestamp 1586364061
transform 1 0 14996 0 1 8160
box -38 -48 406 592
use scs8hd_inv_8  _176_
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_155
timestamp 1586364061
transform 1 0 15364 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_158
timestamp 1586364061
transform 1 0 15640 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_168
timestamp 1586364061
transform 1 0 16560 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_172
timestamp 1586364061
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_176
timestamp 1586364061
transform 1 0 17296 0 1 8160
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_182
timestamp 1586364061
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_196
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_220
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_232
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24012 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 406 592
use scs8hd_buf_2  _241_
timestamp 1586364061
transform 1 0 24564 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24380 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__241__A
timestamp 1586364061
transform 1 0 25116 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_251
timestamp 1586364061
transform 1 0 24196 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_259
timestamp 1586364061
transform 1 0 24932 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_263
timestamp 1586364061
transform 1 0 25300 0 1 8160
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_11_275
timestamp 1586364061
transform 1 0 26404 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_inv_8  _101_
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_12_12
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 406 592
use scs8hd_buf_1  _129_
timestamp 1586364061
transform 1 0 2944 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 2576 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_18
timestamp 1586364061
transform 1 0 2760 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_8  _095_
timestamp 1586364061
transform 1 0 4876 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 4692 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 4232 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__231__A
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_36
timestamp 1586364061
transform 1 0 4416 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 5888 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_50
timestamp 1586364061
transform 1 0 5704 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_54
timestamp 1586364061
transform 1 0 6072 0 -1 9248
box -38 -48 222 592
use scs8hd_or4_4  _126_
timestamp 1586364061
transform 1 0 6440 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__153__D
timestamp 1586364061
transform 1 0 7452 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_67
timestamp 1586364061
transform 1 0 7268 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__115__D
timestamp 1586364061
transform 1 0 7820 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_71
timestamp 1586364061
transform 1 0 7636 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_88
timestamp 1586364061
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 11224 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 11040 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_102
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_106
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12236 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_119
timestamp 1586364061
transform 1 0 12052 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_123
timestamp 1586364061
transform 1 0 12420 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_127
timestamp 1586364061
transform 1 0 12788 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_140
timestamp 1586364061
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_144
timestamp 1586364061
transform 1 0 14352 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_148
timestamp 1586364061
transform 1 0 14720 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_152
timestamp 1586364061
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_165
timestamp 1586364061
transform 1 0 16284 0 -1 9248
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17020 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_176
timestamp 1586364061
transform 1 0 17296 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_188
timestamp 1586364061
transform 1 0 18400 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_200
timestamp 1586364061
transform 1 0 19504 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_212
timestamp 1586364061
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24012 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_12_239
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_247
timestamp 1586364061
transform 1 0 23828 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_258
timestamp 1586364061
transform 1 0 24840 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_270
timestamp 1586364061
transform 1 0 25944 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_274
timestamp 1586364061
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_nand2_4  _108_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 866 592
use scs8hd_buf_2  _231_
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 2024 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_12
timestamp 1586364061
transform 1 0 2208 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_7
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_12
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_20
timestamp 1586364061
transform 1 0 2944 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_16
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_24
timestamp 1586364061
transform 1 0 3312 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__130__D
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 3404 0 1 9248
box -38 -48 222 592
use scs8hd_inv_8  _137_
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 866 592
use scs8hd_or2_4  _099_
timestamp 1586364061
transform 1 0 2576 0 -1 10336
box -38 -48 682 592
use scs8hd_nand2_4  _138_
timestamp 1586364061
transform 1 0 4140 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_36
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_40
timestamp 1586364061
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_29
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_8  _113_
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 866 592
use scs8hd_or4_4  _160_
timestamp 1586364061
transform 1 0 5704 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__D
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__D
timestamp 1586364061
transform 1 0 5520 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_42
timestamp 1586364061
transform 1 0 4968 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_46
timestamp 1586364061
transform 1 0 5336 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_59
timestamp 1586364061
transform 1 0 6532 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__D
timestamp 1586364061
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__C
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_64
timestamp 1586364061
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 7176 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 6992 0 1 9248
box -38 -48 222 592
use scs8hd_or4_4  _153_
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 866 592
use scs8hd_or4_4  _115_
timestamp 1586364061
transform 1 0 7176 0 1 9248
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8740 0 1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 8740 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__D
timestamp 1586364061
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_75
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_79
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_77
timestamp 1586364061
transform 1 0 8188 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_81
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__D
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_94
timestamp 1586364061
transform 1 0 9752 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_85
timestamp 1586364061
transform 1 0 8924 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_89
timestamp 1586364061
transform 1 0 9292 0 -1 10336
box -38 -48 130 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10488 0 1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10304 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_98
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_102
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_107
timestamp 1586364061
transform 1 0 10948 0 -1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_10.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12236 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_113
timestamp 1586364061
transform 1 0 11500 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_117
timestamp 1586364061
transform 1 0 11868 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_119
timestamp 1586364061
transform 1 0 12052 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_123
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12788 0 -1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_134
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_138
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_138
timestamp 1586364061
transform 1 0 13800 0 -1 10336
box -38 -48 406 592
use scs8hd_conb_1  _218_
timestamp 1586364061
transform 1 0 14168 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14260 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_145
timestamp 1586364061
transform 1 0 14444 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_149
timestamp 1586364061
transform 1 0 14812 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_142
timestamp 1586364061
transform 1 0 14168 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15180 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16192 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_162
timestamp 1586364061
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_166
timestamp 1586364061
transform 1 0 16376 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_163
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 1142 592
use scs8hd_conb_1  _223_
timestamp 1586364061
transform 1 0 16744 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16560 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_173
timestamp 1586364061
transform 1 0 17020 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_175
timestamp 1586364061
transform 1 0 17204 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_181
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_187
timestamp 1586364061
transform 1 0 18308 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_196
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_199
timestamp 1586364061
transform 1 0 19412 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_220
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_14_211
timestamp 1586364061
transform 1 0 20516 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_8  _197_
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_240
timestamp 1586364061
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_14_247
timestamp 1586364061
transform 1 0 23828 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_254
timestamp 1586364061
transform 1 0 24472 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_258
timestamp 1586364061
transform 1 0 24840 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_262
timestamp 1586364061
transform 1 0 25208 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_259
timestamp 1586364061
transform 1 0 24932 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_13_274
timestamp 1586364061
transform 1 0 26312 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_271
timestamp 1586364061
transform 1 0 26036 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_or4_4  _166_
timestamp 1586364061
transform 1 0 2024 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 1840 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 130 592
use scs8hd_or4_4  _130_
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__C
timestamp 1586364061
transform 1 0 3404 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 3036 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_19
timestamp 1586364061
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_23
timestamp 1586364061
transform 1 0 3220 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 4876 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_36
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_40
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 130 592
use scs8hd_inv_8  _121_
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_43
timestamp 1586364061
transform 1 0 5060 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_or4_4  _143_
timestamp 1586364061
transform 1 0 7176 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 6992 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__C
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use scs8hd_or4_4  _110_
timestamp 1586364061
transform 1 0 8740 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 8556 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_75
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_79
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_92
timestamp 1586364061
transform 1 0 9568 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_96
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__C
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_100
timestamp 1586364061
transform 1 0 10304 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13708 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14076 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_139
timestamp 1586364061
transform 1 0 13892 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_152
timestamp 1586364061
transform 1 0 15088 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_10.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16284 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_156
timestamp 1586364061
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_163
timestamp 1586364061
transform 1 0 16100 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_167
timestamp 1586364061
transform 1 0 16468 0 1 10336
box -38 -48 406 592
use scs8hd_decap_8  FILLER_15_173
timestamp 1586364061
transform 1 0 17020 0 1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_181
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_220
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 774 592
use scs8hd_buf_2  _240_
timestamp 1586364061
transform 1 0 24564 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__240__A
timestamp 1586364061
transform 1 0 25116 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_253
timestamp 1586364061
transform 1 0 24380 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_259
timestamp 1586364061
transform 1 0 24932 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_263
timestamp 1586364061
transform 1 0 25300 0 1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_15_275
timestamp 1586364061
transform 1 0 26404 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_conb_1  _213_
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__166__C
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_6
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_12
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_8  _192_
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 406 592
use scs8hd_or4_4  _146_
timestamp 1586364061
transform 1 0 4876 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__149__D
timestamp 1586364061
transform 1 0 4692 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 4232 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_29
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_36
timestamp 1586364061
transform 1 0 4416 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__160__C
timestamp 1586364061
transform 1 0 5888 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_50
timestamp 1586364061
transform 1 0 5704 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_54
timestamp 1586364061
transform 1 0 6072 0 -1 11424
box -38 -48 314 592
use scs8hd_or4_4  _134_
timestamp 1586364061
transform 1 0 7268 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__143__D
timestamp 1586364061
transform 1 0 7084 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 6716 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 6348 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_59
timestamp 1586364061
transform 1 0 6532 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_63
timestamp 1586364061
transform 1 0 6900 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 8740 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__D
timestamp 1586364061
transform 1 0 8280 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_76
timestamp 1586364061
transform 1 0 8096 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 314 592
use scs8hd_or4_4  _118_
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__104__C
timestamp 1586364061
transform 1 0 9108 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_85
timestamp 1586364061
transform 1 0 8924 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_89
timestamp 1586364061
transform 1 0 9292 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_102
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_107
timestamp 1586364061
transform 1 0 10948 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 11316 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12328 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_120
timestamp 1586364061
transform 1 0 12144 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_124
timestamp 1586364061
transform 1 0 12512 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12880 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12696 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14352 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_139
timestamp 1586364061
transform 1 0 13892 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_143
timestamp 1586364061
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_146
timestamp 1586364061
transform 1 0 14536 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_152
timestamp 1586364061
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_163
timestamp 1586364061
transform 1 0 16100 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_174
timestamp 1586364061
transform 1 0 17112 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_186
timestamp 1586364061
transform 1 0 18216 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_198
timestamp 1586364061
transform 1 0 19320 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_210
timestamp 1586364061
transform 1 0 20424 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_buf_2  _233_
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__166__D
timestamp 1586364061
transform 1 0 2024 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_12
timestamp 1586364061
transform 1 0 2208 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_16
timestamp 1586364061
transform 1 0 2576 0 1 11424
box -38 -48 222 592
use scs8hd_or4_4  _149_
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 4508 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 4140 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_31
timestamp 1586364061
transform 1 0 3956 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_35
timestamp 1586364061
transform 1 0 4324 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_48
timestamp 1586364061
transform 1 0 5520 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_or4_4  _140_
timestamp 1586364061
transform 1 0 7176 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 6992 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__D
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use scs8hd_or4_4  _104_
timestamp 1586364061
transform 1 0 8740 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_75
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_79
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 9752 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_92
timestamp 1586364061
transform 1 0 9568 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_96
timestamp 1586364061
transform 1 0 9936 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__C
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_100
timestamp 1586364061
transform 1 0 10304 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12604 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_136
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14352 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14168 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_140
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 222 592
use scs8hd_inv_8  _178_
timestamp 1586364061
transform 1 0 15916 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15364 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_153
timestamp 1586364061
transform 1 0 15180 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_157
timestamp 1586364061
transform 1 0 15548 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17296 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16928 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_170
timestamp 1586364061
transform 1 0 16744 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_174
timestamp 1586364061
transform 1 0 17112 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_178
timestamp 1586364061
transform 1 0 17480 0 1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_17_182
timestamp 1586364061
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_buf_1  _167_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_6
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_10
timestamp 1586364061
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _147_
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_41
timestamp 1586364061
transform 1 0 4876 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5796 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__149__C
timestamp 1586364061
transform 1 0 5060 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__C
timestamp 1586364061
transform 1 0 5428 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_45
timestamp 1586364061
transform 1 0 5244 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_49
timestamp 1586364061
transform 1 0 5612 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 7176 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_62
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 222 592
use scs8hd_or4_4  _157_
timestamp 1586364061
transform 1 0 7544 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_4  FILLER_18_79
timestamp 1586364061
transform 1 0 8372 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_83
timestamp 1586364061
transform 1 0 8740 0 -1 12512
box -38 -48 130 592
use scs8hd_nor2_4  _158_
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__123__C
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__D
timestamp 1586364061
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_86
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_90
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 11040 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_106
timestamp 1586364061
transform 1 0 10856 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_119
timestamp 1586364061
transform 1 0 12052 0 -1 12512
box -38 -48 406 592
use scs8hd_inv_8  _198_
timestamp 1586364061
transform 1 0 12788 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_125
timestamp 1586364061
transform 1 0 12604 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_136
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_140
timestamp 1586364061
transform 1 0 13984 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_152
timestamp 1586364061
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_163
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17296 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_175
timestamp 1586364061
transform 1 0 17204 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_179
timestamp 1586364061
transform 1 0 17572 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_191
timestamp 1586364061
transform 1 0 18676 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_203
timestamp 1586364061
transform 1 0 19780 0 -1 12512
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_18_211
timestamp 1586364061
transform 1 0 20516 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_buf_2  _230_
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use scs8hd_buf_1  _100_
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_6
timestamp 1586364061
transform 1 0 1656 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__228__A
timestamp 1586364061
transform 1 0 1840 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 1932 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_10
timestamp 1586364061
transform 1 0 2024 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_11
timestamp 1586364061
transform 1 0 2116 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use scs8hd_inv_8  _193_
timestamp 1586364061
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2944 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2760 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_16
timestamp 1586364061
transform 1 0 2576 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_33
timestamp 1586364061
transform 1 0 4140 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_29
timestamp 1586364061
transform 1 0 3772 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 4232 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_40
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_36
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__C
timestamp 1586364061
transform 1 0 4416 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_nor3_4  _168_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4600 0 -1 13600
box -38 -48 1234 592
use scs8hd_nor2_4  _148_
timestamp 1586364061
transform 1 0 4876 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 5888 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5980 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_50
timestamp 1586364061
transform 1 0 5704 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_54
timestamp 1586364061
transform 1 0 6072 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_51
timestamp 1586364061
transform 1 0 5796 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_55
timestamp 1586364061
transform 1 0 6164 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_61
timestamp 1586364061
transform 1 0 6716 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_19_58
timestamp 1586364061
transform 1 0 6440 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__C
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__140__C
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 8648 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 8280 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 8096 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__C
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_76
timestamp 1586364061
transform 1 0 8096 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_80
timestamp 1586364061
transform 1 0 8464 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_74
timestamp 1586364061
transform 1 0 7912 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_78
timestamp 1586364061
transform 1 0 8280 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_82
timestamp 1586364061
transform 1 0 8648 0 -1 13600
box -38 -48 222 592
use scs8hd_or4_4  _123_
timestamp 1586364061
transform 1 0 8832 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 9752 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__123__D
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_93
timestamp 1586364061
transform 1 0 9660 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_86
timestamp 1586364061
transform 1 0 9016 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10396 0 1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__C
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11132 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_97
timestamp 1586364061
transform 1 0 10028 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_103
timestamp 1586364061
transform 1 0 10580 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_107
timestamp 1586364061
transform 1 0 10948 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_111
timestamp 1586364061
transform 1 0 11316 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_116
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_112
timestamp 1586364061
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_122
timestamp 1586364061
transform 1 0 12328 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12512 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11500 0 -1 13600
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__238__A
timestamp 1586364061
transform 1 0 12880 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_134
timestamp 1586364061
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_138
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_126
timestamp 1586364061
transform 1 0 12696 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_130
timestamp 1586364061
transform 1 0 13064 0 -1 13600
box -38 -48 590 592
use scs8hd_inv_8  _179_
timestamp 1586364061
transform 1 0 14168 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_151
timestamp 1586364061
transform 1 0 14996 0 1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 774 592
use scs8hd_conb_1  _224_
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 314 592
use scs8hd_buf_2  _226_
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__226__A
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_156
timestamp 1586364061
transform 1 0 15456 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_162
timestamp 1586364061
transform 1 0 16008 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_158
timestamp 1586364061
transform 1 0 15640 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_174
timestamp 1586364061
transform 1 0 17112 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_170
timestamp 1586364061
transform 1 0 16744 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_182
timestamp 1586364061
transform 1 0 17848 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_182
timestamp 1586364061
transform 1 0 17848 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_194
timestamp 1586364061
transform 1 0 18952 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_20_206
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_227
timestamp 1586364061
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_239
timestamp 1586364061
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_253
timestamp 1586364061
transform 1 0 24380 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_251
timestamp 1586364061
transform 1 0 24196 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_258
timestamp 1586364061
transform 1 0 24840 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use scs8hd_decap_4  FILLER_20_270
timestamp 1586364061
transform 1 0 25944 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_274
timestamp 1586364061
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_buf_2  _228_
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 2024 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_7
timestamp 1586364061
transform 1 0 1748 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_12
timestamp 1586364061
transform 1 0 2208 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _164_
timestamp 1586364061
transform 1 0 3036 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 2852 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_16
timestamp 1586364061
transform 1 0 2576 0 1 13600
box -38 -48 314 592
use scs8hd_nor3_4  _169_
timestamp 1586364061
transform 1 0 4600 0 1 13600
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_30
timestamp 1586364061
transform 1 0 3864 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_34
timestamp 1586364061
transform 1 0 4232 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_55
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 406 592
use scs8hd_inv_8  _202_
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_nor3_4  _171_
timestamp 1586364061
transform 1 0 8372 0 1 13600
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_71
timestamp 1586364061
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_75
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9752 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_92
timestamp 1586364061
transform 1 0 9568 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_96
timestamp 1586364061
transform 1 0 9936 0 1 13600
box -38 -48 222 592
use scs8hd_nor3_4  _170_
timestamp 1586364061
transform 1 0 10304 0 1 13600
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 10120 0 1 13600
box -38 -48 222 592
use scs8hd_buf_2  _238_
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12052 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_113
timestamp 1586364061
transform 1 0 11500 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_117
timestamp 1586364061
transform 1 0 11868 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_121
timestamp 1586364061
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 13064 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_127
timestamp 1586364061
transform 1 0 12788 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_132
timestamp 1586364061
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_145
timestamp 1586364061
transform 1 0 14444 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_149
timestamp 1586364061
transform 1 0 14812 0 1 13600
box -38 -48 406 592
use scs8hd_conb_1  _216_
timestamp 1586364061
transform 1 0 15180 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15640 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_156
timestamp 1586364061
transform 1 0 15456 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_160
timestamp 1586364061
transform 1 0 15824 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_172
timestamp 1586364061
transform 1 0 16928 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_21_180
timestamp 1586364061
transform 1 0 17664 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_196
timestamp 1586364061
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_220
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_232
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_257
timestamp 1586364061
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__233__A
timestamp 1586364061
transform 1 0 1840 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_6
timestamp 1586364061
transform 1 0 1656 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_10
timestamp 1586364061
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _165_
timestamp 1586364061
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use scs8hd_buf_1  _109_
timestamp 1586364061
transform 1 0 4416 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__169__C
timestamp 1586364061
transform 1 0 4876 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4232 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_39
timestamp 1586364061
transform 1 0 4692 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_13.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5428 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 5244 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_43
timestamp 1586364061
transform 1 0 5060 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 7084 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 7452 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6716 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_58
timestamp 1586364061
transform 1 0 6440 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_63
timestamp 1586364061
transform 1 0 6900 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_67
timestamp 1586364061
transform 1 0 7268 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 7636 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 8648 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_80
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_88
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 10856 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11224 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_104
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_108
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12052 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_112
timestamp 1586364061
transform 1 0 11408 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_118
timestamp 1586364061
transform 1 0 11960 0 -1 14688
box -38 -48 130 592
use scs8hd_inv_8  _199_
timestamp 1586364061
transform 1 0 13616 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_128
timestamp 1586364061
transform 1 0 12880 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_8  FILLER_22_145
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_157
timestamp 1586364061
transform 1 0 15548 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_169
timestamp 1586364061
transform 1 0 16652 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_181
timestamp 1586364061
transform 1 0 17756 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_193
timestamp 1586364061
transform 1 0 18860 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_22_205
timestamp 1586364061
transform 1 0 19964 0 -1 14688
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_213
timestamp 1586364061
transform 1 0 20700 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_239
timestamp 1586364061
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_251
timestamp 1586364061
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_263
timestamp 1586364061
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_buf_2  _227_
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__227__A
timestamp 1586364061
transform 1 0 1932 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_7
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_11
timestamp 1586364061
transform 1 0 2116 0 1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_15.LATCH_1_.latch
timestamp 1586364061
transform 1 0 3036 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2852 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 2392 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_16
timestamp 1586364061
transform 1 0 2576 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4232 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_32
timestamp 1586364061
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_36
timestamp 1586364061
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_40
timestamp 1586364061
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 7084 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8648 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8464 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 8096 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_74
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_78
timestamp 1586364061
transform 1 0 8280 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_93
timestamp 1586364061
transform 1 0 9660 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_97
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use scs8hd_inv_8  _206_
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_112
timestamp 1586364061
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_116
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_120
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_132
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 774 592
use scs8hd_conb_1  _212_
timestamp 1586364061
transform 1 0 13984 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_143
timestamp 1586364061
transform 1 0 14260 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_155
timestamp 1586364061
transform 1 0 15364 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_167
timestamp 1586364061
transform 1 0 16468 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_192
timestamp 1586364061
transform 1 0 18768 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18952 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19412 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_197
timestamp 1586364061
transform 1 0 19228 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_201
timestamp 1586364061
transform 1 0 19596 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_213
timestamp 1586364061
transform 1 0 20700 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_225
timestamp 1586364061
transform 1 0 21804 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_decap_6  FILLER_23_237
timestamp 1586364061
transform 1 0 22908 0 1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_23_243
timestamp 1586364061
transform 1 0 23460 0 1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_253
timestamp 1586364061
transform 1 0 24380 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_258
timestamp 1586364061
transform 1 0 24840 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_262
timestamp 1586364061
transform 1 0 25208 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_23_274
timestamp 1586364061
transform 1 0 26312 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_conb_1  _211_
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1840 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_6
timestamp 1586364061
transform 1 0 1656 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_10
timestamp 1586364061
transform 1 0 2024 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_8  _204_
timestamp 1586364061
transform 1 0 2392 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_15.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5980 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 5244 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__230__A
timestamp 1586364061
transform 1 0 5612 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_43
timestamp 1586364061
transform 1 0 5060 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_47
timestamp 1586364061
transform 1 0 5428 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_51
timestamp 1586364061
transform 1 0 5796 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 7084 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_62
timestamp 1586364061
transform 1 0 6808 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_67
timestamp 1586364061
transform 1 0 7268 0 -1 15776
box -38 -48 314 592
use scs8hd_nor2_4  _136_
timestamp 1586364061
transform 1 0 7544 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8556 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_79
timestamp 1586364061
transform 1 0 8372 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_83
timestamp 1586364061
transform 1 0 8740 0 -1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_87
timestamp 1586364061
transform 1 0 9108 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_91
timestamp 1586364061
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 -1 15776
box -38 -48 866 592
use scs8hd_fill_1  FILLER_24_98
timestamp 1586364061
transform 1 0 10120 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_108
timestamp 1586364061
transform 1 0 11040 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11776 0 -1 15776
box -38 -48 866 592
use scs8hd_conb_1  _221_
timestamp 1586364061
transform 1 0 13340 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 12788 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_125
timestamp 1586364061
transform 1 0 12604 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_129
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_136
timestamp 1586364061
transform 1 0 13616 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_24_148
timestamp 1586364061
transform 1 0 14720 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_152
timestamp 1586364061
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_166
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_178
timestamp 1586364061
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_190
timestamp 1586364061
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_202
timestamp 1586364061
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_239
timestamp 1586364061
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_251
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_263
timestamp 1586364061
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_12
timestamp 1586364061
transform 1 0 2208 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2944 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_16
timestamp 1586364061
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 4508 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_29
timestamp 1586364061
transform 1 0 3772 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_25_34
timestamp 1586364061
transform 1 0 4232 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_46
timestamp 1586364061
transform 1 0 5336 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_50
timestamp 1586364061
transform 1 0 5704 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_conb_1  _210_
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 7268 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_65
timestamp 1586364061
transform 1 0 7084 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_69
timestamp 1586364061
transform 1 0 7452 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8188 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_73
timestamp 1586364061
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 9752 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_88
timestamp 1586364061
transform 1 0 9200 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_92
timestamp 1586364061
transform 1 0 9568 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 10948 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_105
timestamp 1586364061
transform 1 0 10764 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_109
timestamp 1586364061
transform 1 0 11132 0 1 15776
box -38 -48 406 592
use scs8hd_inv_8  _188_
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 11868 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 11500 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_115
timestamp 1586364061
transform 1 0 11684 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_119
timestamp 1586364061
transform 1 0 12052 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_132
timestamp 1586364061
transform 1 0 13248 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_144
timestamp 1586364061
transform 1 0 14352 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_156
timestamp 1586364061
transform 1 0 15456 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_168
timestamp 1586364061
transform 1 0 16560 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_25_180
timestamp 1586364061
transform 1 0 17664 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_196
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_208
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_220
timestamp 1586364061
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_232
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_257
timestamp 1586364061
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_269
timestamp 1586364061
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_15.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_6
timestamp 1586364061
transform 1 0 1656 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1840 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_13.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_27_10
timestamp 1586364061
transform 1 0 2024 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_10
timestamp 1586364061
transform 1 0 2024 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 -1 16864
box -38 -48 222 592
use scs8hd_inv_8  _205_
timestamp 1586364061
transform 1 0 3036 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 2392 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 2760 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_16
timestamp 1586364061
transform 1 0 2576 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_20
timestamp 1586364061
transform 1 0 2944 0 1 16864
box -38 -48 130 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 4600 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 4416 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_41
timestamp 1586364061
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_30
timestamp 1586364061
transform 1 0 3864 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_34
timestamp 1586364061
transform 1 0 4232 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_13.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5796 0 -1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 5612 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_45
timestamp 1586364061
transform 1 0 5244 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_47
timestamp 1586364061
transform 1 0 5428 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 6440 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 6992 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_62
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_27_60
timestamp 1586364061
transform 1 0 6624 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_66
timestamp 1586364061
transform 1 0 7176 0 1 16864
box -38 -48 406 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 7636 0 -1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8188 0 1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8648 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_70
timestamp 1586364061
transform 1 0 7544 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_80
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_70
timestamp 1586364061
transform 1 0 7544 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_73
timestamp 1586364061
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_88
timestamp 1586364061
transform 1 0 9200 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_92
timestamp 1586364061
transform 1 0 9568 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9936 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9936 0 1 16864
box -38 -48 1050 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 10304 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_26_98
timestamp 1586364061
transform 1 0 10120 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_109
timestamp 1586364061
transform 1 0 11132 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_4  FILLER_27_107
timestamp 1586364061
transform 1 0 10948 0 1 16864
box -38 -48 406 592
use scs8hd_inv_8  _175_
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use scs8hd_inv_8  _187_
timestamp 1586364061
transform 1 0 11868 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11316 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11684 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_113
timestamp 1586364061
transform 1 0 11500 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_117
timestamp 1586364061
transform 1 0 11868 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 13432 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_126
timestamp 1586364061
transform 1 0 12696 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_138
timestamp 1586364061
transform 1 0 13800 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_136
timestamp 1586364061
transform 1 0 13616 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_150
timestamp 1586364061
transform 1 0 14904 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_27_140
timestamp 1586364061
transform 1 0 13984 0 1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_152
timestamp 1586364061
transform 1 0 15088 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_166
timestamp 1586364061
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_156
timestamp 1586364061
transform 1 0 15456 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_178
timestamp 1586364061
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_168
timestamp 1586364061
transform 1 0 16560 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_190
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_27_180
timestamp 1586364061
transform 1 0 17664 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_202
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_220
timestamp 1586364061
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_232
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_239
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_257
timestamp 1586364061
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_263
timestamp 1586364061
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_269
timestamp 1586364061
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_15.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2208 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_6
timestamp 1586364061
transform 1 0 1656 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_10
timestamp 1586364061
transform 1 0 2024 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_8  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5244 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5612 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_43
timestamp 1586364061
transform 1 0 5060 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_47
timestamp 1586364061
transform 1 0 5428 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_51
timestamp 1586364061
transform 1 0 5796 0 -1 17952
box -38 -48 590 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 6440 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7452 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_57
timestamp 1586364061
transform 1 0 6348 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_67
timestamp 1586364061
transform 1 0 7268 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_71
timestamp 1586364061
transform 1 0 7636 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_84
timestamp 1586364061
transform 1 0 8832 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_103
timestamp 1586364061
transform 1 0 10580 0 -1 17952
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11316 0 -1 17952
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_28_122
timestamp 1586364061
transform 1 0 12328 0 -1 17952
box -38 -48 406 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 13064 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_126
timestamp 1586364061
transform 1 0 12696 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_129
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_139
timestamp 1586364061
transform 1 0 13892 0 -1 17952
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_28_151
timestamp 1586364061
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_11.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_157
timestamp 1586364061
transform 1 0 15548 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_169
timestamp 1586364061
transform 1 0 16652 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_181
timestamp 1586364061
transform 1 0 17756 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_193
timestamp 1586364061
transform 1 0 18860 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_28_205
timestamp 1586364061
transform 1 0 19964 0 -1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_213
timestamp 1586364061
transform 1 0 20700 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_239
timestamp 1586364061
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_263
timestamp 1586364061
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 2300 0 1 17952
box -38 -48 1050 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_7
timestamp 1586364061
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 3496 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_24
timestamp 1586364061
transform 1 0 3312 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4416 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 3864 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_28
timestamp 1586364061
transform 1 0 3680 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_32
timestamp 1586364061
transform 1 0 4048 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_38
timestamp 1586364061
transform 1 0 4600 0 1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4968 0 1 17952
box -38 -48 1050 592
use scs8hd_decap_6  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 590 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 6900 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8464 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_72
timestamp 1586364061
transform 1 0 7728 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_76
timestamp 1586364061
transform 1 0 8096 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9476 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_89
timestamp 1586364061
transform 1 0 9292 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_93
timestamp 1586364061
transform 1 0 9660 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11040 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_106
timestamp 1586364061
transform 1 0 10856 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_110
timestamp 1586364061
transform 1 0 11224 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_132
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_136
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_148
timestamp 1586364061
transform 1 0 14720 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_160
timestamp 1586364061
transform 1 0 15824 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_172
timestamp 1586364061
transform 1 0 16928 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_29_180
timestamp 1586364061
transform 1 0 17664 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_220
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_232
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_6
timestamp 1586364061
transform 1 0 1656 0 -1 19040
box -38 -48 774 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 2392 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_8  FILLER_30_23
timestamp 1586364061
transform 1 0 3220 0 -1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4232 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_36
timestamp 1586364061
transform 1 0 4416 0 -1 19040
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4968 0 -1 19040
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_30_53
timestamp 1586364061
transform 1 0 5980 0 -1 19040
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7176 0 -1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 6900 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_61
timestamp 1586364061
transform 1 0 6716 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_65
timestamp 1586364061
transform 1 0 7084 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_77
timestamp 1586364061
transform 1 0 8188 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_81
timestamp 1586364061
transform 1 0 8556 0 -1 19040
box -38 -48 222 592
use scs8hd_conb_1  _220_
timestamp 1586364061
transform 1 0 9936 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_30_85
timestamp 1586364061
transform 1 0 8924 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_30_91
timestamp 1586364061
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11040 0 -1 19040
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_30_99
timestamp 1586364061
transform 1 0 10212 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_107
timestamp 1586364061
transform 1 0 10948 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_119
timestamp 1586364061
transform 1 0 12052 0 -1 19040
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 -1 19040
box -38 -48 866 592
use scs8hd_fill_2  FILLER_30_125
timestamp 1586364061
transform 1 0 12604 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_136
timestamp 1586364061
transform 1 0 13616 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_30_148
timestamp 1586364061
transform 1 0 14720 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_152
timestamp 1586364061
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_202
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 590 592
use scs8hd_decap_4  FILLER_31_11
timestamp 1586364061
transform 1 0 2116 0 1 19040
box -38 -48 406 592
use scs8hd_inv_8  _181_
timestamp 1586364061
transform 1 0 2668 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_26
timestamp 1586364061
transform 1 0 3496 0 1 19040
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4232 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5244 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6072 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_43
timestamp 1586364061
transform 1 0 5060 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_47
timestamp 1586364061
transform 1 0 5428 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7452 0 1 19040
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7268 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6440 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_56
timestamp 1586364061
transform 1 0 6256 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_60
timestamp 1586364061
transform 1 0 6624 0 1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_66
timestamp 1586364061
transform 1 0 7176 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8648 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_80
timestamp 1586364061
transform 1 0 8464 0 1 19040
box -38 -48 222 592
use scs8hd_inv_8  _186_
timestamp 1586364061
transform 1 0 9752 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9568 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 9200 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_84
timestamp 1586364061
transform 1 0 8832 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_90
timestamp 1586364061
transform 1 0 9384 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11132 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_103
timestamp 1586364061
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_107
timestamp 1586364061
transform 1 0 10948 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_114
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_132
timestamp 1586364061
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_136
timestamp 1586364061
transform 1 0 13616 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_148
timestamp 1586364061
transform 1 0 14720 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_160
timestamp 1586364061
transform 1 0 15824 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_172
timestamp 1586364061
transform 1 0 16928 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_decap_3  FILLER_31_180
timestamp 1586364061
transform 1 0 17664 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_inv_8  _195_
timestamp 1586364061
transform 1 0 1932 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1748 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_18
timestamp 1586364061
transform 1 0 2760 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_22
timestamp 1586364061
transform 1 0 3128 0 -1 20128
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4784 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4508 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_30
timestamp 1586364061
transform 1 0 3864 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_36
timestamp 1586364061
transform 1 0 4416 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_39
timestamp 1586364061
transform 1 0 4692 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_49
timestamp 1586364061
transform 1 0 5612 0 -1 20128
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6440 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 7452 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_57
timestamp 1586364061
transform 1 0 6348 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_67
timestamp 1586364061
transform 1 0 7268 0 -1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7820 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_71
timestamp 1586364061
transform 1 0 7636 0 -1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_84
timestamp 1586364061
transform 1 0 8832 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_32_102
timestamp 1586364061
transform 1 0 10488 0 -1 20128
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11592 0 -1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_32_123
timestamp 1586364061
transform 1 0 12420 0 -1 20128
box -38 -48 222 592
use scs8hd_inv_8  _174_
timestamp 1586364061
transform 1 0 13156 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12604 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_127
timestamp 1586364061
transform 1 0 12788 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_140
timestamp 1586364061
transform 1 0 13984 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_32_152
timestamp 1586364061
transform 1 0 15088 0 -1 20128
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 -1 21216
box -38 -48 866 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2208 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_6
timestamp 1586364061
transform 1 0 1656 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_10
timestamp 1586364061
transform 1 0 2024 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2852 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2668 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_14
timestamp 1586364061
transform 1 0 2392 0 1 20128
box -38 -48 314 592
use scs8hd_decap_6  FILLER_34_18
timestamp 1586364061
transform 1 0 2760 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_34_24
timestamp 1586364061
transform 1 0 3312 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_conb_1  _214_
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4508 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4324 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_28
timestamp 1586364061
transform 1 0 3680 0 1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_33_34
timestamp 1586364061
transform 1 0 4232 0 1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_34_35
timestamp 1586364061
transform 1 0 4324 0 -1 21216
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5520 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5888 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_46
timestamp 1586364061
transform 1 0 5336 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_50
timestamp 1586364061
transform 1 0 5704 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_54
timestamp 1586364061
transform 1 0 6072 0 1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_34_43
timestamp 1586364061
transform 1 0 5060 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_53
timestamp 1586364061
transform 1 0 5980 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_8  _173_
timestamp 1586364061
transform 1 0 7268 0 -1 21216
box -38 -48 866 592
use scs8hd_conb_1  _217_
timestamp 1586364061
transform 1 0 7084 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_33_60
timestamp 1586364061
transform 1 0 6624 0 1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_68
timestamp 1586364061
transform 1 0 7360 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_65
timestamp 1586364061
transform 1 0 7084 0 -1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8096 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7544 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_72
timestamp 1586364061
transform 1 0 7728 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_76
timestamp 1586364061
transform 1 0 8096 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_8  _172_
timestamp 1586364061
transform 1 0 9660 0 1 20128
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 9476 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9108 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_85
timestamp 1586364061
transform 1 0 8924 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_89
timestamp 1586364061
transform 1 0 9292 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_88
timestamp 1586364061
transform 1 0 9200 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_96
timestamp 1586364061
transform 1 0 9936 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_33_102
timestamp 1586364061
transform 1 0 10488 0 1 20128
box -38 -48 774 592
use scs8hd_decap_4  FILLER_34_108
timestamp 1586364061
transform 1 0 11040 0 -1 21216
box -38 -48 406 592
use scs8hd_conb_1  _222_
timestamp 1586364061
transform 1 0 11408 0 -1 21216
box -38 -48 314 592
use scs8hd_buf_2  _236_
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11684 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_113
timestamp 1586364061
transform 1 0 11500 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_117
timestamp 1586364061
transform 1 0 11868 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_121
timestamp 1586364061
transform 1 0 12236 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_115
timestamp 1586364061
transform 1 0 11684 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__236__A
timestamp 1586364061
transform 1 0 12972 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_127
timestamp 1586364061
transform 1 0 12788 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_131
timestamp 1586364061
transform 1 0 13156 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_138
timestamp 1586364061
transform 1 0 13800 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_127
timestamp 1586364061
transform 1 0 12788 0 -1 21216
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13984 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_142
timestamp 1586364061
transform 1 0 14168 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_139
timestamp 1586364061
transform 1 0 13892 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_34_151
timestamp 1586364061
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_154
timestamp 1586364061
transform 1 0 15272 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_166
timestamp 1586364061
transform 1 0 16376 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_33_178
timestamp 1586364061
transform 1 0 17480 0 1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_33_182
timestamp 1586364061
transform 1 0 17848 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_253
timestamp 1586364061
transform 1 0 24380 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_258
timestamp 1586364061
transform 1 0 24840 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_262
timestamp 1586364061
transform 1 0 25208 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  FILLER_33_274
timestamp 1586364061
transform 1 0 26312 0 1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1840 0 1 21216
box -38 -48 866 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_7
timestamp 1586364061
transform 1 0 1748 0 1 21216
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3404 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3220 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_17
timestamp 1586364061
transform 1 0 2668 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_21
timestamp 1586364061
transform 1 0 3036 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 4784 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4416 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_34
timestamp 1586364061
transform 1 0 4232 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_38
timestamp 1586364061
transform 1 0 4600 0 1 21216
box -38 -48 222 592
use scs8hd_inv_8  _180_
timestamp 1586364061
transform 1 0 4968 0 1 21216
box -38 -48 866 592
use scs8hd_decap_6  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 6348 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_inv_8  _189_
timestamp 1586364061
transform 1 0 8648 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 8464 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__243__A
timestamp 1586364061
transform 1 0 9660 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_91
timestamp 1586364061
transform 1 0 9476 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_95
timestamp 1586364061
transform 1 0 9844 0 1 21216
box -38 -48 590 592
use scs8hd_buf_2  _242_
timestamp 1586364061
transform 1 0 10396 0 1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__242__A
timestamp 1586364061
transform 1 0 10948 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_105
timestamp 1586364061
transform 1 0 10764 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_109
timestamp 1586364061
transform 1 0 11132 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_35_121
timestamp 1586364061
transform 1 0 12236 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_147
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_159
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_171
timestamp 1586364061
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1840 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_6
timestamp 1586364061
transform 1 0 1656 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_10
timestamp 1586364061
transform 1 0 2024 0 -1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_6  FILLER_36_14
timestamp 1586364061
transform 1 0 2392 0 -1 22304
box -38 -48 590 592
use scs8hd_decap_8  FILLER_36_23
timestamp 1586364061
transform 1 0 3220 0 -1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_35
timestamp 1586364061
transform 1 0 4324 0 -1 22304
box -38 -48 774 592
use scs8hd_conb_1  _225_
timestamp 1586364061
transform 1 0 5060 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_46
timestamp 1586364061
transform 1 0 5336 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_3  FILLER_36_54
timestamp 1586364061
transform 1 0 6072 0 -1 22304
box -38 -48 314 592
use scs8hd_inv_8  _203_
timestamp 1586364061
transform 1 0 6348 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_12  FILLER_36_66
timestamp 1586364061
transform 1 0 7176 0 -1 22304
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_78
timestamp 1586364061
transform 1 0 8280 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_82
timestamp 1586364061
transform 1 0 8648 0 -1 22304
box -38 -48 130 592
use scs8hd_buf_2  _243_
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_36_85
timestamp 1586364061
transform 1 0 8924 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_36_91
timestamp 1586364061
transform 1 0 9476 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_97
timestamp 1586364061
transform 1 0 10028 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_36_101
timestamp 1586364061
transform 1 0 10396 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_113
timestamp 1586364061
transform 1 0 11500 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_125
timestamp 1586364061
transform 1 0 12604 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_137
timestamp 1586364061
transform 1 0 13708 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_36_149
timestamp 1586364061
transform 1 0 14812 0 -1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_166
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_178
timestamp 1586364061
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_190
timestamp 1586364061
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_202
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__239__A
timestamp 1586364061
transform 1 0 1564 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_7
timestamp 1586364061
transform 1 0 1748 0 1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_37_13
timestamp 1586364061
transform 1 0 2300 0 1 22304
box -38 -48 130 592
use scs8hd_inv_8  _194_
timestamp 1586364061
transform 1 0 2944 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 2760 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__232__A
timestamp 1586364061
transform 1 0 2392 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_16
timestamp 1586364061
transform 1 0 2576 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_29
timestamp 1586364061
transform 1 0 3772 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_41
timestamp 1586364061
transform 1 0 4876 0 1 22304
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_49
timestamp 1586364061
transform 1 0 5612 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_53
timestamp 1586364061
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_57
timestamp 1586364061
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8740 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_71
timestamp 1586364061
transform 1 0 7636 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_75
timestamp 1586364061
transform 1 0 8004 0 1 22304
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_92
timestamp 1586364061
transform 1 0 9568 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_96
timestamp 1586364061
transform 1 0 9936 0 1 22304
box -38 -48 222 592
use scs8hd_inv_8  _207_
timestamp 1586364061
transform 1 0 10304 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_109
timestamp 1586364061
transform 1 0 11132 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11316 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_113
timestamp 1586364061
transform 1 0 11500 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_117
timestamp 1586364061
transform 1 0 11868 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_121
timestamp 1586364061
transform 1 0 12236 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_37_147
timestamp 1586364061
transform 1 0 14628 0 1 22304
box -38 -48 590 592
use scs8hd_inv_1  mux_top_track_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15732 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_153
timestamp 1586364061
transform 1 0 15180 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_157
timestamp 1586364061
transform 1 0 15548 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_161
timestamp 1586364061
transform 1 0 15916 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_173
timestamp 1586364061
transform 1 0 17020 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_181
timestamp 1586364061
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_196
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_208
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_220
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_232
timestamp 1586364061
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_buf_2  _239_
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_7
timestamp 1586364061
transform 1 0 1748 0 -1 23392
box -38 -48 1142 592
use scs8hd_buf_2  _232_
timestamp 1586364061
transform 1 0 2852 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_8  FILLER_38_23
timestamp 1586364061
transform 1 0 3220 0 -1 23392
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6716 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_4  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_60
timestamp 1586364061
transform 1 0 6624 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_70
timestamp 1586364061
transform 1 0 7544 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_38_82
timestamp 1586364061
transform 1 0 8648 0 -1 23392
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_90
timestamp 1586364061
transform 1 0 9384 0 -1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_8  FILLER_38_102
timestamp 1586364061
transform 1 0 10488 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_38_119
timestamp 1586364061
transform 1 0 12052 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_131
timestamp 1586364061
transform 1 0 13156 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_38_143
timestamp 1586364061
transform 1 0 14260 0 -1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_38_151
timestamp 1586364061
transform 1 0 14996 0 -1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_166
timestamp 1586364061
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_178
timestamp 1586364061
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_190
timestamp 1586364061
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_202
timestamp 1586364061
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_263
timestamp 1586364061
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2024 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_6  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_39_9
timestamp 1586364061
transform 1 0 1932 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_13
timestamp 1586364061
transform 1 0 2300 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_17
timestamp 1586364061
transform 1 0 2668 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_29
timestamp 1586364061
transform 1 0 3772 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_41
timestamp 1586364061
transform 1 0 4876 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_13.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6164 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_53
timestamp 1586364061
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_3  FILLER_40_52
timestamp 1586364061
transform 1 0 5888 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_13.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7268 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7268 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_57
timestamp 1586364061
transform 1 0 6348 0 1 23392
box -38 -48 406 592
use scs8hd_decap_4  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_66
timestamp 1586364061
transform 1 0 7176 0 1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_40_58
timestamp 1586364061
transform 1 0 6440 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_1  FILLER_40_66
timestamp 1586364061
transform 1 0 7176 0 -1 24480
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8740 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7728 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8096 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_70
timestamp 1586364061
transform 1 0 7544 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_78
timestamp 1586364061
transform 1 0 8280 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_82
timestamp 1586364061
transform 1 0 8648 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_70
timestamp 1586364061
transform 1 0 7544 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_82
timestamp 1586364061
transform 1 0 8648 0 -1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9200 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_90
timestamp 1586364061
transform 1 0 9384 0 1 23392
box -38 -48 590 592
use scs8hd_fill_2  FILLER_40_90
timestamp 1586364061
transform 1 0 9384 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10120 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_107
timestamp 1586364061
transform 1 0 10948 0 1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_40_97
timestamp 1586364061
transform 1 0 10028 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_100
timestamp 1586364061
transform 1 0 10304 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11500 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_115
timestamp 1586364061
transform 1 0 11684 0 1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_39_121
timestamp 1586364061
transform 1 0 12236 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_112
timestamp 1586364061
transform 1 0 11408 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_116
timestamp 1586364061
transform 1 0 11776 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13800 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_39_135
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_128
timestamp 1586364061
transform 1 0 12880 0 -1 24480
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14260 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_141
timestamp 1586364061
transform 1 0 14076 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_145
timestamp 1586364061
transform 1 0 14444 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_140
timestamp 1586364061
transform 1 0 13984 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_152
timestamp 1586364061
transform 1 0 15088 0 -1 24480
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_157
timestamp 1586364061
transform 1 0 15548 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_15.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17296 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_169
timestamp 1586364061
transform 1 0 16652 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_174
timestamp 1586364061
transform 1 0 17112 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_178
timestamp 1586364061
transform 1 0 17480 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_39_182
timestamp 1586364061
transform 1 0 17848 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_196
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_208
timestamp 1586364061
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_39_220
timestamp 1586364061
transform 1 0 21344 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21804 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22264 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_224
timestamp 1586364061
transform 1 0 21712 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_228
timestamp 1586364061
transform 1 0 22080 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_232
timestamp 1586364061
transform 1 0 22448 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23460 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_249
timestamp 1586364061
transform 1 0 24012 0 1 23392
box -38 -48 590 592
use scs8hd_decap_4  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_8  FILLER_40_246
timestamp 1586364061
transform 1 0 23736 0 -1 24480
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_258
timestamp 1586364061
transform 1 0 24840 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_262
timestamp 1586364061
transform 1 0 25208 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_254
timestamp 1586364061
transform 1 0 24472 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_258
timestamp 1586364061
transform 1 0 24840 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_266
timestamp 1586364061
transform 1 0 25576 0 1 23392
box -38 -48 774 592
use scs8hd_decap_3  FILLER_39_274
timestamp 1586364061
transform 1 0 26312 0 1 23392
box -38 -48 314 592
use scs8hd_decap_4  FILLER_40_270
timestamp 1586364061
transform 1 0 25944 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_274
timestamp 1586364061
transform 1 0 26312 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
<< labels >>
rlabel metal3 s 0 824 480 944 6 address[0]
port 0 nsew default input
rlabel metal3 s 0 2456 480 2576 6 address[1]
port 1 nsew default input
rlabel metal3 s 27520 1232 28000 1352 6 address[2]
port 2 nsew default input
rlabel metal2 s 754 27520 810 28000 6 address[3]
port 3 nsew default input
rlabel metal3 s 0 4224 480 4344 6 address[4]
port 4 nsew default input
rlabel metal2 s 3790 0 3846 480 6 address[5]
port 5 nsew default input
rlabel metal2 s 5354 0 5410 480 6 chanx_left_in[0]
port 6 nsew default input
rlabel metal2 s 2318 27520 2374 28000 6 chanx_left_in[1]
port 7 nsew default input
rlabel metal2 s 6918 0 6974 480 6 chanx_left_in[2]
port 8 nsew default input
rlabel metal2 s 8482 0 8538 480 6 chanx_left_in[3]
port 9 nsew default input
rlabel metal3 s 27520 3680 28000 3800 6 chanx_left_in[4]
port 10 nsew default input
rlabel metal3 s 0 5992 480 6112 6 chanx_left_in[5]
port 11 nsew default input
rlabel metal2 s 10046 0 10102 480 6 chanx_left_in[6]
port 12 nsew default input
rlabel metal3 s 0 7760 480 7880 6 chanx_left_in[7]
port 13 nsew default input
rlabel metal2 s 11610 0 11666 480 6 chanx_left_in[8]
port 14 nsew default input
rlabel metal2 s 13174 0 13230 480 6 chanx_left_out[0]
port 15 nsew default tristate
rlabel metal3 s 0 9528 480 9648 6 chanx_left_out[1]
port 16 nsew default tristate
rlabel metal2 s 3974 27520 4030 28000 6 chanx_left_out[2]
port 17 nsew default tristate
rlabel metal3 s 0 11296 480 11416 6 chanx_left_out[3]
port 18 nsew default tristate
rlabel metal3 s 0 13064 480 13184 6 chanx_left_out[4]
port 19 nsew default tristate
rlabel metal2 s 14738 0 14794 480 6 chanx_left_out[5]
port 20 nsew default tristate
rlabel metal3 s 0 14832 480 14952 6 chanx_left_out[6]
port 21 nsew default tristate
rlabel metal3 s 0 16464 480 16584 6 chanx_left_out[7]
port 22 nsew default tristate
rlabel metal2 s 16210 0 16266 480 6 chanx_left_out[8]
port 23 nsew default tristate
rlabel metal3 s 0 18232 480 18352 6 chany_top_in[0]
port 24 nsew default input
rlabel metal2 s 5630 27520 5686 28000 6 chany_top_in[1]
port 25 nsew default input
rlabel metal3 s 0 20000 480 20120 6 chany_top_in[2]
port 26 nsew default input
rlabel metal2 s 7286 27520 7342 28000 6 chany_top_in[3]
port 27 nsew default input
rlabel metal2 s 17774 0 17830 480 6 chany_top_in[4]
port 28 nsew default input
rlabel metal2 s 19338 0 19394 480 6 chany_top_in[5]
port 29 nsew default input
rlabel metal3 s 27520 6264 28000 6384 6 chany_top_in[6]
port 30 nsew default input
rlabel metal3 s 0 21768 480 21888 6 chany_top_in[7]
port 31 nsew default input
rlabel metal2 s 8942 27520 8998 28000 6 chany_top_in[8]
port 32 nsew default input
rlabel metal2 s 10598 27520 10654 28000 6 chany_top_out[0]
port 33 nsew default tristate
rlabel metal3 s 0 23536 480 23656 6 chany_top_out[1]
port 34 nsew default tristate
rlabel metal3 s 27520 8848 28000 8968 6 chany_top_out[2]
port 35 nsew default tristate
rlabel metal3 s 27520 11296 28000 11416 6 chany_top_out[3]
port 36 nsew default tristate
rlabel metal3 s 0 25304 480 25424 6 chany_top_out[4]
port 37 nsew default tristate
rlabel metal2 s 12254 27520 12310 28000 6 chany_top_out[5]
port 38 nsew default tristate
rlabel metal2 s 20902 0 20958 480 6 chany_top_out[6]
port 39 nsew default tristate
rlabel metal2 s 13910 27520 13966 28000 6 chany_top_out[7]
port 40 nsew default tristate
rlabel metal2 s 22466 0 22522 480 6 chany_top_out[8]
port 41 nsew default tristate
rlabel metal2 s 2226 0 2282 480 6 data_in
port 42 nsew default input
rlabel metal2 s 754 0 810 480 6 enable
port 43 nsew default input
rlabel metal2 s 17130 27520 17186 28000 6 left_bottom_grid_pin_11_
port 44 nsew default input
rlabel metal2 s 18786 27520 18842 28000 6 left_bottom_grid_pin_13_
port 45 nsew default input
rlabel metal2 s 20442 27520 20498 28000 6 left_bottom_grid_pin_15_
port 46 nsew default input
rlabel metal3 s 27520 13880 28000 14000 6 left_bottom_grid_pin_1_
port 47 nsew default input
rlabel metal3 s 0 27072 480 27192 6 left_bottom_grid_pin_3_
port 48 nsew default input
rlabel metal3 s 27520 16464 28000 16584 6 left_bottom_grid_pin_5_
port 49 nsew default input
rlabel metal2 s 15474 27520 15530 28000 6 left_bottom_grid_pin_7_
port 50 nsew default input
rlabel metal3 s 27520 19048 28000 19168 6 left_bottom_grid_pin_9_
port 51 nsew default input
rlabel metal2 s 24030 0 24086 480 6 left_top_grid_pin_10_
port 52 nsew default input
rlabel metal3 s 27520 21496 28000 21616 6 top_left_grid_pin_13_
port 53 nsew default input
rlabel metal2 s 27158 0 27214 480 6 top_right_grid_pin_11_
port 54 nsew default input
rlabel metal3 s 27520 26664 28000 26784 6 top_right_grid_pin_13_
port 55 nsew default input
rlabel metal2 s 27066 27520 27122 28000 6 top_right_grid_pin_15_
port 56 nsew default input
rlabel metal2 s 22098 27520 22154 28000 6 top_right_grid_pin_1_
port 57 nsew default input
rlabel metal3 s 27520 24080 28000 24200 6 top_right_grid_pin_3_
port 58 nsew default input
rlabel metal2 s 23754 27520 23810 28000 6 top_right_grid_pin_5_
port 59 nsew default input
rlabel metal2 s 25410 27520 25466 28000 6 top_right_grid_pin_7_
port 60 nsew default input
rlabel metal2 s 25594 0 25650 480 6 top_right_grid_pin_9_
port 61 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 62 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 63 nsew default input
<< end >>
