VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga_core
  CLASS BLOCK ;
  FOREIGN fpga_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 2310.000 BY 2486.000 ;
  PIN IO_ISOL_N
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.920 2.400 300.520 ;
    END
  END IO_ISOL_N
  PIN Test_en
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.560 2.400 129.160 ;
    END
  END Test_en
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2307.600 2330.400 2310.000 2331.000 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 2.400 43.480 ;
    END
  END ccff_tail
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 2.400 214.840 ;
    END
  END clk
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 42.870 2483.600 43.150 2486.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2307.600 465.840 2310.000 466.440 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[10]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2307.600 776.600 2310.000 777.200 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[11]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2307.600 1087.360 2310.000 1087.960 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[12]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2307.600 1398.120 2310.000 1398.720 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[13]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2307.600 1708.880 2310.000 1709.480 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[14]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2307.600 2019.640 2310.000 2020.240 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[15]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2026.390 0.000 2026.670 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[16]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2036.970 0.000 2037.250 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[17]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2047.550 0.000 2047.830 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[18]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2058.590 0.000 2058.870 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[19]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 128.430 2483.600 128.710 2486.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2069.170 0.000 2069.450 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[20]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2079.750 0.000 2080.030 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[21]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2090.330 0.000 2090.610 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[22]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2101.370 0.000 2101.650 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[23]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2111.950 0.000 2112.230 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[24]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1737.510 0.000 1737.790 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[25]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1748.090 0.000 1748.370 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[26]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1759.130 0.000 1759.410 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[27]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1769.710 0.000 1769.990 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[28]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1780.290 0.000 1780.570 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[29]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 213.990 2483.600 214.270 2486.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1790.870 0.000 1791.150 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[30]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1801.910 0.000 1802.190 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[31]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1812.490 0.000 1812.770 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[32]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1823.070 0.000 1823.350 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[33]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1448.630 0.000 1448.910 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[34]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1459.670 0.000 1459.950 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[35]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1470.250 0.000 1470.530 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[36]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1480.830 0.000 1481.110 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[37]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1491.410 0.000 1491.690 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[38]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1502.450 0.000 1502.730 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[39]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 299.550 2483.600 299.830 2486.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1513.030 0.000 1513.310 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[40]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1523.610 0.000 1523.890 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[41]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1534.190 0.000 1534.470 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[42]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1160.210 0.000 1160.490 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[43]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1170.790 0.000 1171.070 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[44]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1181.370 0.000 1181.650 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[45]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1191.950 0.000 1192.230 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[46]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1202.990 0.000 1203.270 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[47]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1213.570 0.000 1213.850 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[48]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1224.150 0.000 1224.430 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[49]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 385.110 2483.600 385.390 2486.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1234.730 0.000 1235.010 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[50]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1245.770 0.000 1246.050 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[51]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 871.330 0.000 871.610 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[52]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 881.910 0.000 882.190 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[53]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 892.490 0.000 892.770 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[54]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 903.530 0.000 903.810 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[55]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 914.110 0.000 914.390 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[56]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 924.690 0.000 924.970 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[57]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 935.270 0.000 935.550 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[58]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 946.310 0.000 946.590 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[59]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 470.670 2483.600 470.950 2486.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 956.890 0.000 957.170 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[60]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 582.450 0.000 582.730 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[61]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 593.030 0.000 593.310 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[62]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 604.070 0.000 604.350 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[63]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 614.650 0.000 614.930 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[64]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 625.230 0.000 625.510 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[65]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 635.810 0.000 636.090 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[66]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 646.850 0.000 647.130 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[67]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 657.430 0.000 657.710 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[68]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 668.010 0.000 668.290 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[69]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 556.230 2483.600 556.510 2486.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[70]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 304.610 0.000 304.890 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[71]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 315.190 0.000 315.470 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[72]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 325.770 0.000 326.050 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[73]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 336.350 0.000 336.630 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[74]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[75]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 357.970 0.000 358.250 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[76]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 368.550 0.000 368.830 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[77]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 379.130 0.000 379.410 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[78]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 5.150 0.000 5.430 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[79]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 641.790 2483.600 642.070 2486.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[80]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[81]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[82]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[83]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[84]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[85]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[86]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[87]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 385.600 2.400 386.200 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[88]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 642.640 2.400 643.240 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[89]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 727.350 2483.600 727.630 2486.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 899.680 2.400 900.280 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[90]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1156.720 2.400 1157.320 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[91]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1414.440 2.400 1415.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[92]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1671.480 2.400 1672.080 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[93]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1928.520 2.400 1929.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[94]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2185.560 2.400 2186.160 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[95]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2307.600 155.080 2310.000 155.680 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[9]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 812.910 2483.600 813.190 2486.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2307.600 569.200 2310.000 569.800 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[10]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2307.600 879.960 2310.000 880.560 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[11]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2307.600 1190.720 2310.000 1191.320 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[12]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2307.600 1501.480 2310.000 1502.080 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[13]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2307.600 1812.240 2310.000 1812.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[14]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2307.600 2123.000 2310.000 2123.600 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[15]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2122.530 0.000 2122.810 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[16]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2133.110 0.000 2133.390 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[17]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2144.150 0.000 2144.430 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[18]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2154.730 0.000 2155.010 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[19]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 898.470 2483.600 898.750 2486.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2165.310 0.000 2165.590 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[20]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2175.890 0.000 2176.170 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[21]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2186.930 0.000 2187.210 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[22]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2197.510 0.000 2197.790 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[23]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2208.090 0.000 2208.370 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[24]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1833.650 0.000 1833.930 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[25]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1844.690 0.000 1844.970 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[26]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1855.270 0.000 1855.550 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[27]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1865.850 0.000 1866.130 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[28]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1876.430 0.000 1876.710 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[29]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 984.030 2483.600 984.310 2486.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1887.470 0.000 1887.750 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[30]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1898.050 0.000 1898.330 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[31]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1908.630 0.000 1908.910 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[32]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1919.210 0.000 1919.490 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[33]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1545.230 0.000 1545.510 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[34]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1555.810 0.000 1556.090 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[35]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1566.390 0.000 1566.670 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[36]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1576.970 0.000 1577.250 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[37]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1588.010 0.000 1588.290 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[38]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1598.590 0.000 1598.870 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[39]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1069.590 2483.600 1069.870 2486.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1609.170 0.000 1609.450 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[40]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1619.750 0.000 1620.030 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[41]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1630.790 0.000 1631.070 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[42]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1256.350 0.000 1256.630 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[43]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1266.930 0.000 1267.210 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[44]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1277.510 0.000 1277.790 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[45]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1288.550 0.000 1288.830 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[46]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1299.130 0.000 1299.410 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[47]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1309.710 0.000 1309.990 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[48]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1320.290 0.000 1320.570 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[49]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1155.150 2483.600 1155.430 2486.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1331.330 0.000 1331.610 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[50]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1341.910 0.000 1342.190 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[51]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 967.470 0.000 967.750 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[52]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 978.050 0.000 978.330 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[53]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 989.090 0.000 989.370 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[54]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 999.670 0.000 999.950 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[55]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1010.250 0.000 1010.530 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[56]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1020.830 0.000 1021.110 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[57]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1031.870 0.000 1032.150 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[58]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1042.450 0.000 1042.730 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[59]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1240.710 2483.600 1240.990 2486.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1053.030 0.000 1053.310 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[60]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 678.590 0.000 678.870 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[61]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 689.630 0.000 689.910 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[62]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 700.210 0.000 700.490 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[63]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 710.790 0.000 711.070 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[64]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 721.370 0.000 721.650 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[65]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 732.410 0.000 732.690 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[66]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 742.990 0.000 743.270 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[67]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 753.570 0.000 753.850 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[68]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 764.150 0.000 764.430 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[69]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1326.270 2483.600 1326.550 2486.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 390.170 0.000 390.450 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[70]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 400.750 0.000 401.030 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[71]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 411.330 0.000 411.610 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[72]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[73]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 432.950 0.000 433.230 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[74]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 443.530 0.000 443.810 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[75]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[76]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 464.690 0.000 464.970 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[77]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 475.730 0.000 476.010 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[78]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[79]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1411.830 2483.600 1412.110 2486.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[80]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[81]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[82]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[83]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[84]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[85]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[86]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[87]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[88]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.280 2.400 471.880 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[88]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[89]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 728.320 2.400 728.920 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[89]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1497.390 2483.600 1497.670 2486.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[90]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 985.360 2.400 985.960 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[90]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[91]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1242.400 2.400 1243.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[91]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[92]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1500.120 2.400 1500.720 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[92]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[93]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1757.160 2.400 1757.760 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[93]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[94]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2014.200 2.400 2014.800 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[94]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[95]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2271.240 2.400 2271.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[95]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2307.600 258.440 2310.000 259.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[9]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1582.950 2483.600 1583.230 2486.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2307.600 673.240 2310.000 673.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[10]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2307.600 984.000 2310.000 984.600 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[11]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2307.600 1294.760 2310.000 1295.360 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[12]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2307.600 1605.520 2310.000 1606.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[13]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2307.600 1916.280 2310.000 1916.880 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[14]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2307.600 2227.040 2310.000 2227.640 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[15]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2218.670 0.000 2218.950 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[16]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2229.710 0.000 2229.990 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[17]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2240.290 0.000 2240.570 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[18]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2250.870 0.000 2251.150 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[19]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1668.510 2483.600 1668.790 2486.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2261.450 0.000 2261.730 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[20]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2272.490 0.000 2272.770 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[21]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2283.070 0.000 2283.350 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[22]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2293.650 0.000 2293.930 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[23]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2304.230 0.000 2304.510 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[24]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1930.250 0.000 1930.530 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[25]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1940.830 0.000 1941.110 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[26]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1951.410 0.000 1951.690 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[27]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1961.990 0.000 1962.270 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[28]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1973.030 0.000 1973.310 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[29]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1754.070 2483.600 1754.350 2486.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1983.610 0.000 1983.890 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[30]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1994.190 0.000 1994.470 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[31]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2004.770 0.000 2005.050 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[32]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2015.810 0.000 2016.090 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[33]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1641.370 0.000 1641.650 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[34]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1651.950 0.000 1652.230 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[35]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1662.530 0.000 1662.810 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[36]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1673.570 0.000 1673.850 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[37]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1684.150 0.000 1684.430 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[38]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1694.730 0.000 1695.010 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[39]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1839.630 2483.600 1839.910 2486.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1705.310 0.000 1705.590 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[40]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1716.350 0.000 1716.630 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[41]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1726.930 0.000 1727.210 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[42]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1352.490 0.000 1352.770 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[43]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1363.070 0.000 1363.350 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[44]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1374.110 0.000 1374.390 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[45]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1384.690 0.000 1384.970 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[46]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1395.270 0.000 1395.550 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[47]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1405.850 0.000 1406.130 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[48]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1416.890 0.000 1417.170 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[49]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1925.190 2483.600 1925.470 2486.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1427.470 0.000 1427.750 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[50]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1438.050 0.000 1438.330 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[51]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1063.610 0.000 1063.890 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[52]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1074.650 0.000 1074.930 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[53]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1085.230 0.000 1085.510 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[54]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1095.810 0.000 1096.090 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[55]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1106.390 0.000 1106.670 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[56]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1117.430 0.000 1117.710 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[57]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1128.010 0.000 1128.290 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[58]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1138.590 0.000 1138.870 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[59]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2010.750 2483.600 2011.030 2486.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1149.170 0.000 1149.450 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[60]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 775.190 0.000 775.470 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[61]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 785.770 0.000 786.050 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[62]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 796.350 0.000 796.630 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[63]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 806.930 0.000 807.210 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[64]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 817.970 0.000 818.250 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[65]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 828.550 0.000 828.830 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[66]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 839.130 0.000 839.410 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[67]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 849.710 0.000 849.990 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[68]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 860.750 0.000 861.030 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[69]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2096.310 2483.600 2096.590 2486.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 486.310 0.000 486.590 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[70]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 496.890 0.000 497.170 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[71]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 507.470 0.000 507.750 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[72]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 518.510 0.000 518.790 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[73]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 529.090 0.000 529.370 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[74]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 539.670 0.000 539.950 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[75]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 550.250 0.000 550.530 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[76]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 561.290 0.000 561.570 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[77]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 571.870 0.000 572.150 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[78]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[79]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2181.870 2483.600 2182.150 2486.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[80]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[81]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 229.630 0.000 229.910 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[82]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[83]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 250.790 0.000 251.070 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[84]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 261.830 0.000 262.110 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[85]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[86]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 282.990 0.000 283.270 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[87]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.960 2.400 557.560 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[88]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 814.000 2.400 814.600 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[89]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2267.430 2483.600 2267.710 2486.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1071.040 2.400 1071.640 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[90]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1328.760 2.400 1329.360 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[91]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1585.800 2.400 1586.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[92]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1842.840 2.400 1843.440 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[93]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2099.880 2.400 2100.480 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[94]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2356.920 2.400 2357.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[95]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2307.600 362.480 2310.000 363.080 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[9]
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2307.600 51.720 2310.000 52.320 ;
    END
  END prog_clk
  PIN sc_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2442.600 2.400 2443.200 ;
    END
  END sc_head
  PIN sc_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2307.600 2433.760 2310.000 2434.360 ;
    END
  END sc_tail
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 94.840 2304.140 96.440 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 124.840 2304.140 126.440 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2304.140 2472.565 ;
      LAYER met1 ;
        RECT 5.130 2.760 2304.530 2472.720 ;
      LAYER met2 ;
        RECT 5.160 2483.320 42.590 2483.600 ;
        RECT 43.430 2483.320 128.150 2483.600 ;
        RECT 128.990 2483.320 213.710 2483.600 ;
        RECT 214.550 2483.320 299.270 2483.600 ;
        RECT 300.110 2483.320 384.830 2483.600 ;
        RECT 385.670 2483.320 470.390 2483.600 ;
        RECT 471.230 2483.320 555.950 2483.600 ;
        RECT 556.790 2483.320 641.510 2483.600 ;
        RECT 642.350 2483.320 727.070 2483.600 ;
        RECT 727.910 2483.320 812.630 2483.600 ;
        RECT 813.470 2483.320 898.190 2483.600 ;
        RECT 899.030 2483.320 983.750 2483.600 ;
        RECT 984.590 2483.320 1069.310 2483.600 ;
        RECT 1070.150 2483.320 1154.870 2483.600 ;
        RECT 1155.710 2483.320 1240.430 2483.600 ;
        RECT 1241.270 2483.320 1325.990 2483.600 ;
        RECT 1326.830 2483.320 1411.550 2483.600 ;
        RECT 1412.390 2483.320 1497.110 2483.600 ;
        RECT 1497.950 2483.320 1582.670 2483.600 ;
        RECT 1583.510 2483.320 1668.230 2483.600 ;
        RECT 1669.070 2483.320 1753.790 2483.600 ;
        RECT 1754.630 2483.320 1839.350 2483.600 ;
        RECT 1840.190 2483.320 1924.910 2483.600 ;
        RECT 1925.750 2483.320 2010.470 2483.600 ;
        RECT 2011.310 2483.320 2096.030 2483.600 ;
        RECT 2096.870 2483.320 2181.590 2483.600 ;
        RECT 2182.430 2483.320 2267.150 2483.600 ;
        RECT 2267.990 2483.320 2304.500 2483.600 ;
        RECT 5.160 2.680 2304.500 2483.320 ;
        RECT 5.710 2.400 15.450 2.680 ;
        RECT 16.290 2.400 26.030 2.680 ;
        RECT 26.870 2.400 36.610 2.680 ;
        RECT 37.450 2.400 47.650 2.680 ;
        RECT 48.490 2.400 58.230 2.680 ;
        RECT 59.070 2.400 68.810 2.680 ;
        RECT 69.650 2.400 79.390 2.680 ;
        RECT 80.230 2.400 90.430 2.680 ;
        RECT 91.270 2.400 101.010 2.680 ;
        RECT 101.850 2.400 111.590 2.680 ;
        RECT 112.430 2.400 122.170 2.680 ;
        RECT 123.010 2.400 133.210 2.680 ;
        RECT 134.050 2.400 143.790 2.680 ;
        RECT 144.630 2.400 154.370 2.680 ;
        RECT 155.210 2.400 164.950 2.680 ;
        RECT 165.790 2.400 175.990 2.680 ;
        RECT 176.830 2.400 186.570 2.680 ;
        RECT 187.410 2.400 197.150 2.680 ;
        RECT 197.990 2.400 207.730 2.680 ;
        RECT 208.570 2.400 218.770 2.680 ;
        RECT 219.610 2.400 229.350 2.680 ;
        RECT 230.190 2.400 239.930 2.680 ;
        RECT 240.770 2.400 250.510 2.680 ;
        RECT 251.350 2.400 261.550 2.680 ;
        RECT 262.390 2.400 272.130 2.680 ;
        RECT 272.970 2.400 282.710 2.680 ;
        RECT 283.550 2.400 293.290 2.680 ;
        RECT 294.130 2.400 304.330 2.680 ;
        RECT 305.170 2.400 314.910 2.680 ;
        RECT 315.750 2.400 325.490 2.680 ;
        RECT 326.330 2.400 336.070 2.680 ;
        RECT 336.910 2.400 347.110 2.680 ;
        RECT 347.950 2.400 357.690 2.680 ;
        RECT 358.530 2.400 368.270 2.680 ;
        RECT 369.110 2.400 378.850 2.680 ;
        RECT 379.690 2.400 389.890 2.680 ;
        RECT 390.730 2.400 400.470 2.680 ;
        RECT 401.310 2.400 411.050 2.680 ;
        RECT 411.890 2.400 421.630 2.680 ;
        RECT 422.470 2.400 432.670 2.680 ;
        RECT 433.510 2.400 443.250 2.680 ;
        RECT 444.090 2.400 453.830 2.680 ;
        RECT 454.670 2.400 464.410 2.680 ;
        RECT 465.250 2.400 475.450 2.680 ;
        RECT 476.290 2.400 486.030 2.680 ;
        RECT 486.870 2.400 496.610 2.680 ;
        RECT 497.450 2.400 507.190 2.680 ;
        RECT 508.030 2.400 518.230 2.680 ;
        RECT 519.070 2.400 528.810 2.680 ;
        RECT 529.650 2.400 539.390 2.680 ;
        RECT 540.230 2.400 549.970 2.680 ;
        RECT 550.810 2.400 561.010 2.680 ;
        RECT 561.850 2.400 571.590 2.680 ;
        RECT 572.430 2.400 582.170 2.680 ;
        RECT 583.010 2.400 592.750 2.680 ;
        RECT 593.590 2.400 603.790 2.680 ;
        RECT 604.630 2.400 614.370 2.680 ;
        RECT 615.210 2.400 624.950 2.680 ;
        RECT 625.790 2.400 635.530 2.680 ;
        RECT 636.370 2.400 646.570 2.680 ;
        RECT 647.410 2.400 657.150 2.680 ;
        RECT 657.990 2.400 667.730 2.680 ;
        RECT 668.570 2.400 678.310 2.680 ;
        RECT 679.150 2.400 689.350 2.680 ;
        RECT 690.190 2.400 699.930 2.680 ;
        RECT 700.770 2.400 710.510 2.680 ;
        RECT 711.350 2.400 721.090 2.680 ;
        RECT 721.930 2.400 732.130 2.680 ;
        RECT 732.970 2.400 742.710 2.680 ;
        RECT 743.550 2.400 753.290 2.680 ;
        RECT 754.130 2.400 763.870 2.680 ;
        RECT 764.710 2.400 774.910 2.680 ;
        RECT 775.750 2.400 785.490 2.680 ;
        RECT 786.330 2.400 796.070 2.680 ;
        RECT 796.910 2.400 806.650 2.680 ;
        RECT 807.490 2.400 817.690 2.680 ;
        RECT 818.530 2.400 828.270 2.680 ;
        RECT 829.110 2.400 838.850 2.680 ;
        RECT 839.690 2.400 849.430 2.680 ;
        RECT 850.270 2.400 860.470 2.680 ;
        RECT 861.310 2.400 871.050 2.680 ;
        RECT 871.890 2.400 881.630 2.680 ;
        RECT 882.470 2.400 892.210 2.680 ;
        RECT 893.050 2.400 903.250 2.680 ;
        RECT 904.090 2.400 913.830 2.680 ;
        RECT 914.670 2.400 924.410 2.680 ;
        RECT 925.250 2.400 934.990 2.680 ;
        RECT 935.830 2.400 946.030 2.680 ;
        RECT 946.870 2.400 956.610 2.680 ;
        RECT 957.450 2.400 967.190 2.680 ;
        RECT 968.030 2.400 977.770 2.680 ;
        RECT 978.610 2.400 988.810 2.680 ;
        RECT 989.650 2.400 999.390 2.680 ;
        RECT 1000.230 2.400 1009.970 2.680 ;
        RECT 1010.810 2.400 1020.550 2.680 ;
        RECT 1021.390 2.400 1031.590 2.680 ;
        RECT 1032.430 2.400 1042.170 2.680 ;
        RECT 1043.010 2.400 1052.750 2.680 ;
        RECT 1053.590 2.400 1063.330 2.680 ;
        RECT 1064.170 2.400 1074.370 2.680 ;
        RECT 1075.210 2.400 1084.950 2.680 ;
        RECT 1085.790 2.400 1095.530 2.680 ;
        RECT 1096.370 2.400 1106.110 2.680 ;
        RECT 1106.950 2.400 1117.150 2.680 ;
        RECT 1117.990 2.400 1127.730 2.680 ;
        RECT 1128.570 2.400 1138.310 2.680 ;
        RECT 1139.150 2.400 1148.890 2.680 ;
        RECT 1149.730 2.400 1159.930 2.680 ;
        RECT 1160.770 2.400 1170.510 2.680 ;
        RECT 1171.350 2.400 1181.090 2.680 ;
        RECT 1181.930 2.400 1191.670 2.680 ;
        RECT 1192.510 2.400 1202.710 2.680 ;
        RECT 1203.550 2.400 1213.290 2.680 ;
        RECT 1214.130 2.400 1223.870 2.680 ;
        RECT 1224.710 2.400 1234.450 2.680 ;
        RECT 1235.290 2.400 1245.490 2.680 ;
        RECT 1246.330 2.400 1256.070 2.680 ;
        RECT 1256.910 2.400 1266.650 2.680 ;
        RECT 1267.490 2.400 1277.230 2.680 ;
        RECT 1278.070 2.400 1288.270 2.680 ;
        RECT 1289.110 2.400 1298.850 2.680 ;
        RECT 1299.690 2.400 1309.430 2.680 ;
        RECT 1310.270 2.400 1320.010 2.680 ;
        RECT 1320.850 2.400 1331.050 2.680 ;
        RECT 1331.890 2.400 1341.630 2.680 ;
        RECT 1342.470 2.400 1352.210 2.680 ;
        RECT 1353.050 2.400 1362.790 2.680 ;
        RECT 1363.630 2.400 1373.830 2.680 ;
        RECT 1374.670 2.400 1384.410 2.680 ;
        RECT 1385.250 2.400 1394.990 2.680 ;
        RECT 1395.830 2.400 1405.570 2.680 ;
        RECT 1406.410 2.400 1416.610 2.680 ;
        RECT 1417.450 2.400 1427.190 2.680 ;
        RECT 1428.030 2.400 1437.770 2.680 ;
        RECT 1438.610 2.400 1448.350 2.680 ;
        RECT 1449.190 2.400 1459.390 2.680 ;
        RECT 1460.230 2.400 1469.970 2.680 ;
        RECT 1470.810 2.400 1480.550 2.680 ;
        RECT 1481.390 2.400 1491.130 2.680 ;
        RECT 1491.970 2.400 1502.170 2.680 ;
        RECT 1503.010 2.400 1512.750 2.680 ;
        RECT 1513.590 2.400 1523.330 2.680 ;
        RECT 1524.170 2.400 1533.910 2.680 ;
        RECT 1534.750 2.400 1544.950 2.680 ;
        RECT 1545.790 2.400 1555.530 2.680 ;
        RECT 1556.370 2.400 1566.110 2.680 ;
        RECT 1566.950 2.400 1576.690 2.680 ;
        RECT 1577.530 2.400 1587.730 2.680 ;
        RECT 1588.570 2.400 1598.310 2.680 ;
        RECT 1599.150 2.400 1608.890 2.680 ;
        RECT 1609.730 2.400 1619.470 2.680 ;
        RECT 1620.310 2.400 1630.510 2.680 ;
        RECT 1631.350 2.400 1641.090 2.680 ;
        RECT 1641.930 2.400 1651.670 2.680 ;
        RECT 1652.510 2.400 1662.250 2.680 ;
        RECT 1663.090 2.400 1673.290 2.680 ;
        RECT 1674.130 2.400 1683.870 2.680 ;
        RECT 1684.710 2.400 1694.450 2.680 ;
        RECT 1695.290 2.400 1705.030 2.680 ;
        RECT 1705.870 2.400 1716.070 2.680 ;
        RECT 1716.910 2.400 1726.650 2.680 ;
        RECT 1727.490 2.400 1737.230 2.680 ;
        RECT 1738.070 2.400 1747.810 2.680 ;
        RECT 1748.650 2.400 1758.850 2.680 ;
        RECT 1759.690 2.400 1769.430 2.680 ;
        RECT 1770.270 2.400 1780.010 2.680 ;
        RECT 1780.850 2.400 1790.590 2.680 ;
        RECT 1791.430 2.400 1801.630 2.680 ;
        RECT 1802.470 2.400 1812.210 2.680 ;
        RECT 1813.050 2.400 1822.790 2.680 ;
        RECT 1823.630 2.400 1833.370 2.680 ;
        RECT 1834.210 2.400 1844.410 2.680 ;
        RECT 1845.250 2.400 1854.990 2.680 ;
        RECT 1855.830 2.400 1865.570 2.680 ;
        RECT 1866.410 2.400 1876.150 2.680 ;
        RECT 1876.990 2.400 1887.190 2.680 ;
        RECT 1888.030 2.400 1897.770 2.680 ;
        RECT 1898.610 2.400 1908.350 2.680 ;
        RECT 1909.190 2.400 1918.930 2.680 ;
        RECT 1919.770 2.400 1929.970 2.680 ;
        RECT 1930.810 2.400 1940.550 2.680 ;
        RECT 1941.390 2.400 1951.130 2.680 ;
        RECT 1951.970 2.400 1961.710 2.680 ;
        RECT 1962.550 2.400 1972.750 2.680 ;
        RECT 1973.590 2.400 1983.330 2.680 ;
        RECT 1984.170 2.400 1993.910 2.680 ;
        RECT 1994.750 2.400 2004.490 2.680 ;
        RECT 2005.330 2.400 2015.530 2.680 ;
        RECT 2016.370 2.400 2026.110 2.680 ;
        RECT 2026.950 2.400 2036.690 2.680 ;
        RECT 2037.530 2.400 2047.270 2.680 ;
        RECT 2048.110 2.400 2058.310 2.680 ;
        RECT 2059.150 2.400 2068.890 2.680 ;
        RECT 2069.730 2.400 2079.470 2.680 ;
        RECT 2080.310 2.400 2090.050 2.680 ;
        RECT 2090.890 2.400 2101.090 2.680 ;
        RECT 2101.930 2.400 2111.670 2.680 ;
        RECT 2112.510 2.400 2122.250 2.680 ;
        RECT 2123.090 2.400 2132.830 2.680 ;
        RECT 2133.670 2.400 2143.870 2.680 ;
        RECT 2144.710 2.400 2154.450 2.680 ;
        RECT 2155.290 2.400 2165.030 2.680 ;
        RECT 2165.870 2.400 2175.610 2.680 ;
        RECT 2176.450 2.400 2186.650 2.680 ;
        RECT 2187.490 2.400 2197.230 2.680 ;
        RECT 2198.070 2.400 2207.810 2.680 ;
        RECT 2208.650 2.400 2218.390 2.680 ;
        RECT 2219.230 2.400 2229.430 2.680 ;
        RECT 2230.270 2.400 2240.010 2.680 ;
        RECT 2240.850 2.400 2250.590 2.680 ;
        RECT 2251.430 2.400 2261.170 2.680 ;
        RECT 2262.010 2.400 2272.210 2.680 ;
        RECT 2273.050 2.400 2282.790 2.680 ;
        RECT 2283.630 2.400 2293.370 2.680 ;
        RECT 2294.210 2.400 2303.950 2.680 ;
      LAYER met3 ;
        RECT 2.400 2443.600 2307.600 2472.645 ;
        RECT 2.800 2442.200 2307.600 2443.600 ;
        RECT 2.400 2434.760 2307.600 2442.200 ;
        RECT 2.400 2433.360 2307.200 2434.760 ;
        RECT 2.400 2357.920 2307.600 2433.360 ;
        RECT 2.800 2356.520 2307.600 2357.920 ;
        RECT 2.400 2331.400 2307.600 2356.520 ;
        RECT 2.400 2330.000 2307.200 2331.400 ;
        RECT 2.400 2272.240 2307.600 2330.000 ;
        RECT 2.800 2270.840 2307.600 2272.240 ;
        RECT 2.400 2228.040 2307.600 2270.840 ;
        RECT 2.400 2226.640 2307.200 2228.040 ;
        RECT 2.400 2186.560 2307.600 2226.640 ;
        RECT 2.800 2185.160 2307.600 2186.560 ;
        RECT 2.400 2124.000 2307.600 2185.160 ;
        RECT 2.400 2122.600 2307.200 2124.000 ;
        RECT 2.400 2100.880 2307.600 2122.600 ;
        RECT 2.800 2099.480 2307.600 2100.880 ;
        RECT 2.400 2020.640 2307.600 2099.480 ;
        RECT 2.400 2019.240 2307.200 2020.640 ;
        RECT 2.400 2015.200 2307.600 2019.240 ;
        RECT 2.800 2013.800 2307.600 2015.200 ;
        RECT 2.400 1929.520 2307.600 2013.800 ;
        RECT 2.800 1928.120 2307.600 1929.520 ;
        RECT 2.400 1917.280 2307.600 1928.120 ;
        RECT 2.400 1915.880 2307.200 1917.280 ;
        RECT 2.400 1843.840 2307.600 1915.880 ;
        RECT 2.800 1842.440 2307.600 1843.840 ;
        RECT 2.400 1813.240 2307.600 1842.440 ;
        RECT 2.400 1811.840 2307.200 1813.240 ;
        RECT 2.400 1758.160 2307.600 1811.840 ;
        RECT 2.800 1756.760 2307.600 1758.160 ;
        RECT 2.400 1709.880 2307.600 1756.760 ;
        RECT 2.400 1708.480 2307.200 1709.880 ;
        RECT 2.400 1672.480 2307.600 1708.480 ;
        RECT 2.800 1671.080 2307.600 1672.480 ;
        RECT 2.400 1606.520 2307.600 1671.080 ;
        RECT 2.400 1605.120 2307.200 1606.520 ;
        RECT 2.400 1586.800 2307.600 1605.120 ;
        RECT 2.800 1585.400 2307.600 1586.800 ;
        RECT 2.400 1502.480 2307.600 1585.400 ;
        RECT 2.400 1501.120 2307.200 1502.480 ;
        RECT 2.800 1501.080 2307.200 1501.120 ;
        RECT 2.800 1499.720 2307.600 1501.080 ;
        RECT 2.400 1415.440 2307.600 1499.720 ;
        RECT 2.800 1414.040 2307.600 1415.440 ;
        RECT 2.400 1399.120 2307.600 1414.040 ;
        RECT 2.400 1397.720 2307.200 1399.120 ;
        RECT 2.400 1329.760 2307.600 1397.720 ;
        RECT 2.800 1328.360 2307.600 1329.760 ;
        RECT 2.400 1295.760 2307.600 1328.360 ;
        RECT 2.400 1294.360 2307.200 1295.760 ;
        RECT 2.400 1243.400 2307.600 1294.360 ;
        RECT 2.800 1242.000 2307.600 1243.400 ;
        RECT 2.400 1191.720 2307.600 1242.000 ;
        RECT 2.400 1190.320 2307.200 1191.720 ;
        RECT 2.400 1157.720 2307.600 1190.320 ;
        RECT 2.800 1156.320 2307.600 1157.720 ;
        RECT 2.400 1088.360 2307.600 1156.320 ;
        RECT 2.400 1086.960 2307.200 1088.360 ;
        RECT 2.400 1072.040 2307.600 1086.960 ;
        RECT 2.800 1070.640 2307.600 1072.040 ;
        RECT 2.400 986.360 2307.600 1070.640 ;
        RECT 2.800 985.000 2307.600 986.360 ;
        RECT 2.800 984.960 2307.200 985.000 ;
        RECT 2.400 983.600 2307.200 984.960 ;
        RECT 2.400 900.680 2307.600 983.600 ;
        RECT 2.800 899.280 2307.600 900.680 ;
        RECT 2.400 880.960 2307.600 899.280 ;
        RECT 2.400 879.560 2307.200 880.960 ;
        RECT 2.400 815.000 2307.600 879.560 ;
        RECT 2.800 813.600 2307.600 815.000 ;
        RECT 2.400 777.600 2307.600 813.600 ;
        RECT 2.400 776.200 2307.200 777.600 ;
        RECT 2.400 729.320 2307.600 776.200 ;
        RECT 2.800 727.920 2307.600 729.320 ;
        RECT 2.400 674.240 2307.600 727.920 ;
        RECT 2.400 672.840 2307.200 674.240 ;
        RECT 2.400 643.640 2307.600 672.840 ;
        RECT 2.800 642.240 2307.600 643.640 ;
        RECT 2.400 570.200 2307.600 642.240 ;
        RECT 2.400 568.800 2307.200 570.200 ;
        RECT 2.400 557.960 2307.600 568.800 ;
        RECT 2.800 556.560 2307.600 557.960 ;
        RECT 2.400 472.280 2307.600 556.560 ;
        RECT 2.800 470.880 2307.600 472.280 ;
        RECT 2.400 466.840 2307.600 470.880 ;
        RECT 2.400 465.440 2307.200 466.840 ;
        RECT 2.400 386.600 2307.600 465.440 ;
        RECT 2.800 385.200 2307.600 386.600 ;
        RECT 2.400 363.480 2307.600 385.200 ;
        RECT 2.400 362.080 2307.200 363.480 ;
        RECT 2.400 300.920 2307.600 362.080 ;
        RECT 2.800 299.520 2307.600 300.920 ;
        RECT 2.400 259.440 2307.600 299.520 ;
        RECT 2.400 258.040 2307.200 259.440 ;
        RECT 2.400 215.240 2307.600 258.040 ;
        RECT 2.800 213.840 2307.600 215.240 ;
        RECT 2.400 156.080 2307.600 213.840 ;
        RECT 2.400 154.680 2307.200 156.080 ;
        RECT 2.400 129.560 2307.600 154.680 ;
        RECT 2.800 128.160 2307.600 129.560 ;
        RECT 2.400 52.720 2307.600 128.160 ;
        RECT 2.400 51.320 2307.200 52.720 ;
        RECT 2.400 43.880 2307.600 51.320 ;
        RECT 2.800 42.480 2307.600 43.880 ;
        RECT 2.400 10.715 2307.600 42.480 ;
      LAYER met4 ;
        RECT 21.040 10.640 2297.640 2472.720 ;
      LAYER met5 ;
        RECT 5.520 154.840 2304.140 2466.440 ;
  END
END fpga_core
END LIBRARY

