magic
tech sky130A
magscale 1 2
timestamp 1609016931
<< locali >>
rect 9413 18675 9447 18777
rect 7573 18131 7607 18233
rect 14289 17927 14323 18097
rect 8953 16839 8987 17077
rect 8861 11467 8895 11705
rect 22017 11535 22051 12113
rect 11713 9223 11747 9325
rect 22017 8271 22051 8849
<< viali >>
rect 20177 20409 20211 20443
rect 20729 20409 20763 20443
rect 19993 20205 20027 20239
rect 20545 20205 20579 20239
rect 14381 19865 14415 19899
rect 16497 19865 16531 19899
rect 18245 19865 18279 19899
rect 19349 19865 19383 19899
rect 21005 19865 21039 19899
rect 20085 19797 20119 19831
rect 4813 19729 4847 19763
rect 5080 19729 5114 19763
rect 6837 19729 6871 19763
rect 8033 19729 8067 19763
rect 8300 19729 8334 19763
rect 14749 19729 14783 19763
rect 15393 19729 15427 19763
rect 16405 19729 16439 19763
rect 17049 19729 17083 19763
rect 18061 19729 18095 19763
rect 19809 19729 19843 19763
rect 20821 19729 20855 19763
rect 7113 19661 7147 19695
rect 9689 19661 9723 19695
rect 14841 19661 14875 19695
rect 14933 19661 14967 19695
rect 16589 19661 16623 19695
rect 6193 19525 6227 19559
rect 9413 19525 9447 19559
rect 14013 19525 14047 19559
rect 16037 19525 16071 19559
rect 20453 19321 20487 19355
rect 21097 19321 21131 19355
rect 9689 19253 9723 19287
rect 12449 19253 12483 19287
rect 8953 19185 8987 19219
rect 10241 19185 10275 19219
rect 4077 19117 4111 19151
rect 6193 19117 6227 19151
rect 6449 19117 6483 19151
rect 8861 19117 8895 19151
rect 10057 19117 10091 19151
rect 11069 19117 11103 19151
rect 12725 19117 12759 19151
rect 12981 19117 13015 19151
rect 15301 19117 15335 19151
rect 17049 19117 17083 19151
rect 17325 19117 17359 19151
rect 18245 19117 18279 19151
rect 19533 19117 19567 19151
rect 19809 19117 19843 19151
rect 20269 19117 20303 19151
rect 20913 19117 20947 19151
rect 4322 19049 4356 19083
rect 11336 19049 11370 19083
rect 15546 19049 15580 19083
rect 19073 19049 19107 19083
rect 5457 18981 5491 19015
rect 7573 18981 7607 19015
rect 8401 18981 8435 19015
rect 8769 18981 8803 19015
rect 10149 18981 10183 19015
rect 14105 18981 14139 19015
rect 16681 18981 16715 19015
rect 4537 18777 4571 18811
rect 5089 18777 5123 18811
rect 6837 18777 6871 18811
rect 9229 18777 9263 18811
rect 9413 18777 9447 18811
rect 9689 18777 9723 18811
rect 11621 18777 11655 18811
rect 14933 18777 14967 18811
rect 16497 18777 16531 18811
rect 18521 18777 18555 18811
rect 21005 18777 21039 18811
rect 13820 18709 13854 18743
rect 18429 18709 18463 18743
rect 19441 18709 19475 18743
rect 20177 18709 20211 18743
rect 2688 18641 2722 18675
rect 4445 18641 4479 18675
rect 6285 18641 6319 18675
rect 7205 18641 7239 18675
rect 9413 18641 9447 18675
rect 10508 18641 10542 18675
rect 12817 18641 12851 18675
rect 16865 18641 16899 18675
rect 17509 18641 17543 18675
rect 19165 18641 19199 18675
rect 19901 18641 19935 18675
rect 20821 18641 20855 18675
rect 2421 18573 2455 18607
rect 4629 18573 4663 18607
rect 7297 18573 7331 18607
rect 7389 18573 7423 18607
rect 10241 18573 10275 18607
rect 12909 18573 12943 18607
rect 13001 18573 13035 18607
rect 13553 18573 13587 18607
rect 16957 18573 16991 18607
rect 17049 18573 17083 18607
rect 18613 18573 18647 18607
rect 3801 18505 3835 18539
rect 18061 18505 18095 18539
rect 4077 18437 4111 18471
rect 5549 18437 5583 18471
rect 11989 18437 12023 18471
rect 12449 18437 12483 18471
rect 16129 18437 16163 18471
rect 6653 18233 6687 18267
rect 7573 18233 7607 18267
rect 7757 18233 7791 18267
rect 11069 18233 11103 18267
rect 16957 18233 16991 18267
rect 11345 18165 11379 18199
rect 7113 18097 7147 18131
rect 7205 18097 7239 18131
rect 7573 18097 7607 18131
rect 11897 18097 11931 18131
rect 13921 18097 13955 18131
rect 14105 18097 14139 18131
rect 14289 18097 14323 18131
rect 18889 18097 18923 18131
rect 9689 18029 9723 18063
rect 9956 18029 9990 18063
rect 11713 17961 11747 17995
rect 12357 17961 12391 17995
rect 13829 17961 13863 17995
rect 15577 18029 15611 18063
rect 15844 18029 15878 18063
rect 17233 18029 17267 18063
rect 17489 18029 17523 18063
rect 20913 18029 20947 18063
rect 14473 17961 14507 17995
rect 7021 17893 7055 17927
rect 8033 17893 8067 17927
rect 11805 17893 11839 17927
rect 13093 17893 13127 17927
rect 13461 17893 13495 17927
rect 14289 17893 14323 17927
rect 18613 17893 18647 17927
rect 19349 17893 19383 17927
rect 21097 17893 21131 17927
rect 4721 17689 4755 17723
rect 9505 17689 9539 17723
rect 9873 17689 9907 17723
rect 19533 17689 19567 17723
rect 10333 17621 10367 17655
rect 4629 17553 4663 17587
rect 8033 17553 8067 17587
rect 10241 17553 10275 17587
rect 10885 17553 10919 17587
rect 19349 17553 19383 17587
rect 20269 17553 20303 17587
rect 20821 17553 20855 17587
rect 4905 17485 4939 17519
rect 10517 17485 10551 17519
rect 20453 17417 20487 17451
rect 4261 17349 4295 17383
rect 21005 17349 21039 17383
rect 3157 17145 3191 17179
rect 6745 17145 6779 17179
rect 6193 17077 6227 17111
rect 7113 17077 7147 17111
rect 8953 17077 8987 17111
rect 10333 17077 10367 17111
rect 11437 17077 11471 17111
rect 4353 17009 4387 17043
rect 7665 17009 7699 17043
rect 8677 17009 8711 17043
rect 1777 16941 1811 16975
rect 4813 16941 4847 16975
rect 5080 16941 5114 16975
rect 7573 16941 7607 16975
rect 2044 16873 2078 16907
rect 7481 16873 7515 16907
rect 8493 16873 8527 16907
rect 12081 17009 12115 17043
rect 18889 17009 18923 17043
rect 20085 17009 20119 17043
rect 11161 16941 11195 16975
rect 15761 16941 15795 16975
rect 18613 16941 18647 16975
rect 19809 16941 19843 16975
rect 20913 16941 20947 16975
rect 9137 16873 9171 16907
rect 11897 16873 11931 16907
rect 3433 16805 3467 16839
rect 8125 16805 8159 16839
rect 8585 16805 8619 16839
rect 8953 16805 8987 16839
rect 11805 16805 11839 16839
rect 21097 16805 21131 16839
rect 3617 16601 3651 16635
rect 4169 16601 4203 16635
rect 8217 16601 8251 16635
rect 10517 16601 10551 16635
rect 10885 16601 10919 16635
rect 10977 16601 11011 16635
rect 11805 16601 11839 16635
rect 13001 16601 13035 16635
rect 14841 16601 14875 16635
rect 15945 16601 15979 16635
rect 18061 16601 18095 16635
rect 7082 16533 7116 16567
rect 9014 16533 9048 16567
rect 12725 16533 12759 16567
rect 13461 16533 13495 16567
rect 16405 16533 16439 16567
rect 16957 16533 16991 16567
rect 18429 16533 18463 16567
rect 19993 16533 20027 16567
rect 3525 16465 3559 16499
rect 4721 16465 4755 16499
rect 4997 16465 5031 16499
rect 13369 16465 13403 16499
rect 14013 16465 14047 16499
rect 14749 16465 14783 16499
rect 15393 16465 15427 16499
rect 16313 16465 16347 16499
rect 18521 16465 18555 16499
rect 19717 16465 19751 16499
rect 20453 16465 20487 16499
rect 20729 16465 20763 16499
rect 3709 16397 3743 16431
rect 6837 16397 6871 16431
rect 8769 16397 8803 16431
rect 11069 16397 11103 16431
rect 13553 16397 13587 16431
rect 14933 16397 14967 16431
rect 16589 16397 16623 16431
rect 18705 16397 18739 16431
rect 14381 16329 14415 16363
rect 3157 16261 3191 16295
rect 10149 16261 10183 16295
rect 2789 16057 2823 16091
rect 6561 16057 6595 16091
rect 7665 16057 7699 16091
rect 13277 16057 13311 16091
rect 14933 16057 14967 16091
rect 16681 16057 16715 16091
rect 18337 16057 18371 16091
rect 21097 16057 21131 16091
rect 3249 15921 3283 15955
rect 3341 15921 3375 15955
rect 5181 15921 5215 15955
rect 8953 15921 8987 15955
rect 10241 15921 10275 15955
rect 18613 15921 18647 15955
rect 4261 15853 4295 15887
rect 7849 15853 7883 15887
rect 8677 15853 8711 15887
rect 10497 15853 10531 15887
rect 11897 15853 11931 15887
rect 13553 15853 13587 15887
rect 13809 15853 13843 15887
rect 15301 15853 15335 15887
rect 15557 15853 15591 15887
rect 16957 15853 16991 15887
rect 17213 15853 17247 15887
rect 20913 15853 20947 15887
rect 3157 15785 3191 15819
rect 5448 15785 5482 15819
rect 12164 15785 12198 15819
rect 11621 15717 11655 15751
rect 3157 15513 3191 15547
rect 7205 15513 7239 15547
rect 8309 15445 8343 15479
rect 18328 15445 18362 15479
rect 20085 15445 20119 15479
rect 1777 15377 1811 15411
rect 2044 15377 2078 15411
rect 7573 15377 7607 15411
rect 18061 15377 18095 15411
rect 19809 15377 19843 15411
rect 20821 15377 20855 15411
rect 7665 15309 7699 15343
rect 7757 15309 7791 15343
rect 19441 15173 19475 15207
rect 21005 15173 21039 15207
rect 7113 14969 7147 15003
rect 4169 14901 4203 14935
rect 4721 14833 4755 14867
rect 7665 14833 7699 14867
rect 8125 14833 8159 14867
rect 7573 14765 7607 14799
rect 8769 14765 8803 14799
rect 19901 14765 19935 14799
rect 20913 14765 20947 14799
rect 4537 14697 4571 14731
rect 5181 14697 5215 14731
rect 7481 14697 7515 14731
rect 20177 14697 20211 14731
rect 4629 14629 4663 14663
rect 8585 14629 8619 14663
rect 13369 14629 13403 14663
rect 21097 14629 21131 14663
rect 4445 14425 4479 14459
rect 4721 14425 4755 14459
rect 5089 14425 5123 14459
rect 11989 14425 12023 14459
rect 12909 14425 12943 14459
rect 17601 14425 17635 14459
rect 18521 14425 18555 14459
rect 21005 14425 21039 14459
rect 3332 14357 3366 14391
rect 7104 14357 7138 14391
rect 8585 14357 8619 14391
rect 10149 14357 10183 14391
rect 12817 14357 12851 14391
rect 19073 14357 19107 14391
rect 5825 14289 5859 14323
rect 9229 14289 9263 14323
rect 9873 14289 9907 14323
rect 13737 14289 13771 14323
rect 14280 14289 14314 14323
rect 16037 14289 16071 14323
rect 18429 14289 18463 14323
rect 19993 14289 20027 14323
rect 20821 14289 20855 14323
rect 3065 14221 3099 14255
rect 5181 14221 5215 14255
rect 5273 14221 5307 14255
rect 6837 14221 6871 14255
rect 9321 14221 9355 14255
rect 9505 14221 9539 14255
rect 13093 14221 13127 14255
rect 14013 14221 14047 14255
rect 16129 14221 16163 14255
rect 16221 14221 16255 14255
rect 18705 14221 18739 14255
rect 20269 14221 20303 14255
rect 8217 14153 8251 14187
rect 8861 14153 8895 14187
rect 12449 14153 12483 14187
rect 13553 14085 13587 14119
rect 15393 14085 15427 14119
rect 15669 14085 15703 14119
rect 18061 14085 18095 14119
rect 19717 14085 19751 14119
rect 4537 13881 4571 13915
rect 7205 13881 7239 13915
rect 8033 13881 8067 13915
rect 8401 13881 8435 13915
rect 15301 13881 15335 13915
rect 18705 13881 18739 13915
rect 18981 13881 19015 13915
rect 20453 13881 20487 13915
rect 21097 13881 21131 13915
rect 13645 13813 13679 13847
rect 13921 13813 13955 13847
rect 8861 13745 8895 13779
rect 9045 13745 9079 13779
rect 9965 13745 9999 13779
rect 12265 13745 12299 13779
rect 14381 13745 14415 13779
rect 14565 13745 14599 13779
rect 15853 13745 15887 13779
rect 16589 13745 16623 13779
rect 17325 13745 17359 13779
rect 19441 13745 19475 13779
rect 19533 13745 19567 13779
rect 5825 13677 5859 13711
rect 6092 13677 6126 13711
rect 10232 13677 10266 13711
rect 15669 13677 15703 13711
rect 16313 13677 16347 13711
rect 17592 13677 17626 13711
rect 20269 13677 20303 13711
rect 20913 13677 20947 13711
rect 12510 13609 12544 13643
rect 15761 13609 15795 13643
rect 8769 13541 8803 13575
rect 11345 13541 11379 13575
rect 14289 13541 14323 13575
rect 19349 13541 19383 13575
rect 5181 13337 5215 13371
rect 9413 13337 9447 13371
rect 11529 13337 11563 13371
rect 12541 13337 12575 13371
rect 15485 13337 15519 13371
rect 16221 13337 16255 13371
rect 18429 13337 18463 13371
rect 20545 13337 20579 13371
rect 21097 13337 21131 13371
rect 8024 13269 8058 13303
rect 10241 13269 10275 13303
rect 13001 13269 13035 13303
rect 13921 13269 13955 13303
rect 3801 13201 3835 13235
rect 4068 13201 4102 13235
rect 12909 13201 12943 13235
rect 18797 13201 18831 13235
rect 19441 13201 19475 13235
rect 20361 13201 20395 13235
rect 20913 13201 20947 13235
rect 7757 13133 7791 13167
rect 13093 13133 13127 13167
rect 18889 13133 18923 13167
rect 19073 13133 19107 13167
rect 20085 13133 20119 13167
rect 9137 13065 9171 13099
rect 13645 12997 13679 13031
rect 7757 12793 7791 12827
rect 9965 12793 9999 12827
rect 12357 12793 12391 12827
rect 13093 12793 13127 12827
rect 18981 12793 19015 12827
rect 19901 12793 19935 12827
rect 20453 12793 20487 12827
rect 21097 12793 21131 12827
rect 15669 12725 15703 12759
rect 17049 12725 17083 12759
rect 10609 12657 10643 12691
rect 16221 12657 16255 12691
rect 17601 12657 17635 12691
rect 7941 12589 7975 12623
rect 10333 12589 10367 12623
rect 10977 12589 11011 12623
rect 13277 12589 13311 12623
rect 17509 12589 17543 12623
rect 19441 12589 19475 12623
rect 19717 12589 19751 12623
rect 20269 12589 20303 12623
rect 20913 12589 20947 12623
rect 11222 12521 11256 12555
rect 12633 12521 12667 12555
rect 16037 12521 16071 12555
rect 18153 12521 18187 12555
rect 10425 12453 10459 12487
rect 14197 12453 14231 12487
rect 16129 12453 16163 12487
rect 16773 12453 16807 12487
rect 17417 12453 17451 12487
rect 18429 12453 18463 12487
rect 10333 12249 10367 12283
rect 13645 12249 13679 12283
rect 15669 12249 15703 12283
rect 16681 12249 16715 12283
rect 21005 12249 21039 12283
rect 11713 12181 11747 12215
rect 16037 12181 16071 12215
rect 17141 12181 17175 12215
rect 18429 12181 18463 12215
rect 20177 12181 20211 12215
rect 10701 12113 10735 12147
rect 11437 12113 11471 12147
rect 14289 12113 14323 12147
rect 17049 12113 17083 12147
rect 18521 12113 18555 12147
rect 19901 12113 19935 12147
rect 20821 12113 20855 12147
rect 22017 12113 22051 12147
rect 10793 12045 10827 12079
rect 10977 12045 11011 12079
rect 12909 12045 12943 12079
rect 13737 12045 13771 12079
rect 13921 12045 13955 12079
rect 14565 12045 14599 12079
rect 15393 12045 15427 12079
rect 16129 12045 16163 12079
rect 16313 12045 16347 12079
rect 17325 12045 17359 12079
rect 18613 12045 18647 12079
rect 19625 12045 19659 12079
rect 13277 11909 13311 11943
rect 18061 11909 18095 11943
rect 19165 11909 19199 11943
rect 7665 11705 7699 11739
rect 8861 11705 8895 11739
rect 9137 11705 9171 11739
rect 11069 11705 11103 11739
rect 11345 11705 11379 11739
rect 14473 11705 14507 11739
rect 18153 11705 18187 11739
rect 19349 11705 19383 11739
rect 21097 11705 21131 11739
rect 8493 11569 8527 11603
rect 8677 11569 8711 11603
rect 13093 11569 13127 11603
rect 17693 11569 17727 11603
rect 18797 11569 18831 11603
rect 9689 11501 9723 11535
rect 15301 11501 15335 11535
rect 15568 11501 15602 11535
rect 19165 11501 19199 11535
rect 20545 11501 20579 11535
rect 20913 11501 20947 11535
rect 22017 11501 22051 11535
rect 8401 11433 8435 11467
rect 8861 11433 8895 11467
rect 9956 11433 9990 11467
rect 13360 11433 13394 11467
rect 18521 11433 18555 11467
rect 8033 11365 8067 11399
rect 16681 11365 16715 11399
rect 18613 11365 18647 11399
rect 19717 11365 19751 11399
rect 8585 11161 8619 11195
rect 9137 11161 9171 11195
rect 10517 11161 10551 11195
rect 13553 11161 13587 11195
rect 21005 11161 21039 11195
rect 19441 11093 19475 11127
rect 8493 11025 8527 11059
rect 9597 11025 9631 11059
rect 10885 11025 10919 11059
rect 10977 11025 11011 11059
rect 13737 11025 13771 11059
rect 19165 11025 19199 11059
rect 20177 11025 20211 11059
rect 20821 11025 20855 11059
rect 8769 10957 8803 10991
rect 11069 10957 11103 10991
rect 8125 10889 8159 10923
rect 20545 10889 20579 10923
rect 8033 10617 8067 10651
rect 11161 10617 11195 10651
rect 12541 10617 12575 10651
rect 19257 10617 19291 10651
rect 21097 10617 21131 10651
rect 12265 10549 12299 10583
rect 8493 10481 8527 10515
rect 8677 10481 8711 10515
rect 10701 10481 10735 10515
rect 11621 10481 11655 10515
rect 11713 10481 11747 10515
rect 14197 10481 14231 10515
rect 19901 10481 19935 10515
rect 8401 10413 8435 10447
rect 11529 10413 11563 10447
rect 15301 10413 15335 10447
rect 20913 10413 20947 10447
rect 13921 10345 13955 10379
rect 19625 10345 19659 10379
rect 20269 10345 20303 10379
rect 13553 10277 13587 10311
rect 14013 10277 14047 10311
rect 14565 10277 14599 10311
rect 18981 10277 19015 10311
rect 19717 10277 19751 10311
rect 9321 10073 9355 10107
rect 13461 10073 13495 10107
rect 13553 10073 13587 10107
rect 17601 10073 17635 10107
rect 19441 10073 19475 10107
rect 19717 10073 19751 10107
rect 20085 10073 20119 10107
rect 21005 10073 21039 10107
rect 14442 10005 14476 10039
rect 16488 10005 16522 10039
rect 20177 10005 20211 10039
rect 7941 9937 7975 9971
rect 8208 9937 8242 9971
rect 14197 9937 14231 9971
rect 16221 9937 16255 9971
rect 18061 9937 18095 9971
rect 18328 9937 18362 9971
rect 20821 9937 20855 9971
rect 13645 9869 13679 9903
rect 20269 9869 20303 9903
rect 13093 9733 13127 9767
rect 15577 9733 15611 9767
rect 11529 9529 11563 9563
rect 20085 9529 20119 9563
rect 13185 9461 13219 9495
rect 21097 9461 21131 9495
rect 13921 9393 13955 9427
rect 14013 9393 14047 9427
rect 15853 9393 15887 9427
rect 18705 9393 18739 9427
rect 10149 9325 10183 9359
rect 11713 9325 11747 9359
rect 11805 9325 11839 9359
rect 12072 9325 12106 9359
rect 18972 9325 19006 9359
rect 20545 9325 20579 9359
rect 20913 9325 20947 9359
rect 10416 9257 10450 9291
rect 13829 9257 13863 9291
rect 11713 9189 11747 9223
rect 13461 9189 13495 9223
rect 15301 9189 15335 9223
rect 15669 9189 15703 9223
rect 15761 9189 15795 9223
rect 16405 9189 16439 9223
rect 11897 8985 11931 9019
rect 13461 8985 13495 9019
rect 15393 8985 15427 9019
rect 16221 8985 16255 9019
rect 20085 8985 20119 9019
rect 20545 8985 20579 9019
rect 11713 8849 11747 8883
rect 13277 8849 13311 8883
rect 16037 8849 16071 8883
rect 19809 8849 19843 8883
rect 20821 8849 20855 8883
rect 22017 8849 22051 8883
rect 21005 8713 21039 8747
rect 21097 8441 21131 8475
rect 11345 8305 11379 8339
rect 13645 8305 13679 8339
rect 16589 8305 16623 8339
rect 11069 8237 11103 8271
rect 13461 8237 13495 8271
rect 16405 8237 16439 8271
rect 20545 8237 20579 8271
rect 20913 8237 20947 8271
rect 22017 8237 22051 8271
rect 11161 7897 11195 7931
rect 16957 7897 16991 7931
rect 19625 7897 19659 7931
rect 21005 7897 21039 7931
rect 17325 7829 17359 7863
rect 10701 7761 10735 7795
rect 11529 7761 11563 7795
rect 13645 7761 13679 7795
rect 13912 7761 13946 7795
rect 18501 7761 18535 7795
rect 20545 7761 20579 7795
rect 20821 7761 20855 7795
rect 11621 7693 11655 7727
rect 11713 7693 11747 7727
rect 15301 7693 15335 7727
rect 17417 7693 17451 7727
rect 17601 7693 17635 7727
rect 18245 7693 18279 7727
rect 15025 7557 15059 7591
rect 11253 7353 11287 7387
rect 18429 7353 18463 7387
rect 18705 7353 18739 7387
rect 21097 7353 21131 7387
rect 13277 7285 13311 7319
rect 9873 7217 9907 7251
rect 14749 7217 14783 7251
rect 15393 7217 15427 7251
rect 19165 7217 19199 7251
rect 19257 7217 19291 7251
rect 11897 7149 11931 7183
rect 12153 7149 12187 7183
rect 14565 7149 14599 7183
rect 17049 7149 17083 7183
rect 17316 7149 17350 7183
rect 20545 7149 20579 7183
rect 20913 7149 20947 7183
rect 10140 7081 10174 7115
rect 13921 7081 13955 7115
rect 15638 7081 15672 7115
rect 19073 7081 19107 7115
rect 14197 7013 14231 7047
rect 14657 7013 14691 7047
rect 16773 7013 16807 7047
rect 19717 7013 19751 7047
rect 11345 6809 11379 6843
rect 11805 6809 11839 6843
rect 14657 6809 14691 6843
rect 18613 6809 18647 6843
rect 11713 6741 11747 6775
rect 14565 6741 14599 6775
rect 8657 6673 8691 6707
rect 11069 6673 11103 6707
rect 18061 6673 18095 6707
rect 8401 6605 8435 6639
rect 11897 6605 11931 6639
rect 14749 6605 14783 6639
rect 9781 6537 9815 6571
rect 14197 6537 14231 6571
rect 8033 6469 8067 6503
rect 12541 6469 12575 6503
rect 15301 6469 15335 6503
rect 21373 6469 21407 6503
rect 21097 6265 21131 6299
rect 20913 6061 20947 6095
rect 21005 5721 21039 5755
rect 20821 5585 20855 5619
rect 21281 5109 21315 5143
rect 21005 4633 21039 4667
rect 20821 4497 20855 4531
rect 21281 4089 21315 4123
<< metal1 >>
rect 1104 20554 21896 20576
rect 1104 20502 4447 20554
rect 4499 20502 4511 20554
rect 4563 20502 4575 20554
rect 4627 20502 4639 20554
rect 4691 20502 11378 20554
rect 11430 20502 11442 20554
rect 11494 20502 11506 20554
rect 11558 20502 11570 20554
rect 11622 20502 18308 20554
rect 18360 20502 18372 20554
rect 18424 20502 18436 20554
rect 18488 20502 18500 20554
rect 18552 20502 21896 20554
rect 1104 20480 21896 20502
rect 20162 20440 20168 20452
rect 20123 20412 20168 20440
rect 20162 20400 20168 20412
rect 20220 20400 20226 20452
rect 20530 20400 20536 20452
rect 20588 20440 20594 20452
rect 20717 20443 20775 20449
rect 20717 20440 20729 20443
rect 20588 20412 20729 20440
rect 20588 20400 20594 20412
rect 20717 20409 20729 20412
rect 20763 20409 20775 20443
rect 20717 20403 20775 20409
rect 19978 20236 19984 20248
rect 19939 20208 19984 20236
rect 19978 20196 19984 20208
rect 20036 20196 20042 20248
rect 20070 20196 20076 20248
rect 20128 20236 20134 20248
rect 20533 20239 20591 20245
rect 20533 20236 20545 20239
rect 20128 20208 20545 20236
rect 20128 20196 20134 20208
rect 20533 20205 20545 20208
rect 20579 20205 20591 20239
rect 20533 20199 20591 20205
rect 1104 20010 21896 20032
rect 1104 19958 7912 20010
rect 7964 19958 7976 20010
rect 8028 19958 8040 20010
rect 8092 19958 8104 20010
rect 8156 19958 14843 20010
rect 14895 19958 14907 20010
rect 14959 19958 14971 20010
rect 15023 19958 15035 20010
rect 15087 19958 21896 20010
rect 1104 19936 21896 19958
rect 14369 19899 14427 19905
rect 14369 19865 14381 19899
rect 14415 19896 14427 19899
rect 16485 19899 16543 19905
rect 16485 19896 16497 19899
rect 14415 19868 16497 19896
rect 14415 19865 14427 19868
rect 14369 19859 14427 19865
rect 16485 19865 16497 19868
rect 16531 19865 16543 19899
rect 16485 19859 16543 19865
rect 18233 19899 18291 19905
rect 18233 19865 18245 19899
rect 18279 19896 18291 19899
rect 18598 19896 18604 19908
rect 18279 19868 18604 19896
rect 18279 19865 18291 19868
rect 18233 19859 18291 19865
rect 18598 19856 18604 19868
rect 18656 19856 18662 19908
rect 19242 19856 19248 19908
rect 19300 19896 19306 19908
rect 19337 19899 19395 19905
rect 19337 19896 19349 19899
rect 19300 19868 19349 19896
rect 19300 19856 19306 19868
rect 19337 19865 19349 19868
rect 19383 19865 19395 19899
rect 19337 19859 19395 19865
rect 20622 19856 20628 19908
rect 20680 19896 20686 19908
rect 20993 19899 21051 19905
rect 20993 19896 21005 19899
rect 20680 19868 21005 19896
rect 20680 19856 20686 19868
rect 20993 19865 21005 19868
rect 21039 19865 21051 19899
rect 20993 19859 21051 19865
rect 20070 19828 20076 19840
rect 4908 19800 8064 19828
rect 20031 19800 20076 19828
rect 4908 19772 4936 19800
rect 4801 19763 4859 19769
rect 4801 19729 4813 19763
rect 4847 19760 4859 19763
rect 4890 19760 4896 19772
rect 4847 19732 4896 19760
rect 4847 19729 4859 19732
rect 4801 19723 4859 19729
rect 4890 19720 4896 19732
rect 4948 19720 4954 19772
rect 5068 19763 5126 19769
rect 5068 19729 5080 19763
rect 5114 19760 5126 19763
rect 6546 19760 6552 19772
rect 5114 19732 6552 19760
rect 5114 19729 5126 19732
rect 5068 19723 5126 19729
rect 6546 19720 6552 19732
rect 6604 19720 6610 19772
rect 6822 19760 6828 19772
rect 6783 19732 6828 19760
rect 6822 19720 6828 19732
rect 6880 19720 6886 19772
rect 8036 19769 8064 19800
rect 20070 19788 20076 19800
rect 20128 19788 20134 19840
rect 8294 19769 8300 19772
rect 8021 19763 8079 19769
rect 8021 19729 8033 19763
rect 8067 19729 8079 19763
rect 8288 19760 8300 19769
rect 8255 19732 8300 19760
rect 8021 19723 8079 19729
rect 8288 19723 8300 19732
rect 8294 19720 8300 19723
rect 8352 19720 8358 19772
rect 14182 19720 14188 19772
rect 14240 19760 14246 19772
rect 14737 19763 14795 19769
rect 14737 19760 14749 19763
rect 14240 19732 14749 19760
rect 14240 19720 14246 19732
rect 14737 19729 14749 19732
rect 14783 19760 14795 19763
rect 15381 19763 15439 19769
rect 15381 19760 15393 19763
rect 14783 19732 15393 19760
rect 14783 19729 14795 19732
rect 14737 19723 14795 19729
rect 15381 19729 15393 19732
rect 15427 19729 15439 19763
rect 15381 19723 15439 19729
rect 16393 19763 16451 19769
rect 16393 19729 16405 19763
rect 16439 19760 16451 19763
rect 17037 19763 17095 19769
rect 17037 19760 17049 19763
rect 16439 19732 17049 19760
rect 16439 19729 16451 19732
rect 16393 19723 16451 19729
rect 17037 19729 17049 19732
rect 17083 19729 17095 19763
rect 18046 19760 18052 19772
rect 18007 19732 18052 19760
rect 17037 19723 17095 19729
rect 18046 19720 18052 19732
rect 18104 19720 18110 19772
rect 18138 19720 18144 19772
rect 18196 19760 18202 19772
rect 19797 19763 19855 19769
rect 19797 19760 19809 19763
rect 18196 19732 19809 19760
rect 18196 19720 18202 19732
rect 19797 19729 19809 19732
rect 19843 19729 19855 19763
rect 19797 19723 19855 19729
rect 20162 19720 20168 19772
rect 20220 19760 20226 19772
rect 20809 19763 20867 19769
rect 20809 19760 20821 19763
rect 20220 19732 20821 19760
rect 20220 19720 20226 19732
rect 20809 19729 20821 19732
rect 20855 19729 20867 19763
rect 20809 19723 20867 19729
rect 7101 19695 7159 19701
rect 7101 19661 7113 19695
rect 7147 19692 7159 19695
rect 7742 19692 7748 19704
rect 7147 19664 7748 19692
rect 7147 19661 7159 19664
rect 7101 19655 7159 19661
rect 7742 19652 7748 19664
rect 7800 19652 7806 19704
rect 9674 19692 9680 19704
rect 9635 19664 9680 19692
rect 9674 19652 9680 19664
rect 9732 19652 9738 19704
rect 14829 19695 14887 19701
rect 14829 19692 14841 19695
rect 14016 19664 14841 19692
rect 14016 19568 14044 19664
rect 14829 19661 14841 19664
rect 14875 19661 14887 19695
rect 14829 19655 14887 19661
rect 14921 19695 14979 19701
rect 14921 19661 14933 19695
rect 14967 19661 14979 19695
rect 16577 19695 16635 19701
rect 16577 19692 16589 19695
rect 14921 19655 14979 19661
rect 16408 19664 16589 19692
rect 14734 19584 14740 19636
rect 14792 19624 14798 19636
rect 14936 19624 14964 19655
rect 16408 19636 16436 19664
rect 16577 19661 16589 19664
rect 16623 19661 16635 19695
rect 16577 19655 16635 19661
rect 14792 19596 14964 19624
rect 14792 19584 14798 19596
rect 16390 19584 16396 19636
rect 16448 19584 16454 19636
rect 6181 19559 6239 19565
rect 6181 19525 6193 19559
rect 6227 19556 6239 19559
rect 6270 19556 6276 19568
rect 6227 19528 6276 19556
rect 6227 19525 6239 19528
rect 6181 19519 6239 19525
rect 6270 19516 6276 19528
rect 6328 19516 6334 19568
rect 9401 19559 9459 19565
rect 9401 19525 9413 19559
rect 9447 19556 9459 19559
rect 10226 19556 10232 19568
rect 9447 19528 10232 19556
rect 9447 19525 9459 19528
rect 9401 19519 9459 19525
rect 10226 19516 10232 19528
rect 10284 19516 10290 19568
rect 13998 19556 14004 19568
rect 13959 19528 14004 19556
rect 13998 19516 14004 19528
rect 14056 19516 14062 19568
rect 16025 19559 16083 19565
rect 16025 19525 16037 19559
rect 16071 19556 16083 19559
rect 17034 19556 17040 19568
rect 16071 19528 17040 19556
rect 16071 19525 16083 19528
rect 16025 19519 16083 19525
rect 17034 19516 17040 19528
rect 17092 19516 17098 19568
rect 1104 19466 21896 19488
rect 1104 19414 4447 19466
rect 4499 19414 4511 19466
rect 4563 19414 4575 19466
rect 4627 19414 4639 19466
rect 4691 19414 11378 19466
rect 11430 19414 11442 19466
rect 11494 19414 11506 19466
rect 11558 19414 11570 19466
rect 11622 19414 18308 19466
rect 18360 19414 18372 19466
rect 18424 19414 18436 19466
rect 18488 19414 18500 19466
rect 18552 19414 21896 19466
rect 1104 19392 21896 19414
rect 20438 19352 20444 19364
rect 20399 19324 20444 19352
rect 20438 19312 20444 19324
rect 20496 19312 20502 19364
rect 21082 19352 21088 19364
rect 21043 19324 21088 19352
rect 21082 19312 21088 19324
rect 21140 19312 21146 19364
rect 9677 19287 9735 19293
rect 9677 19284 9689 19287
rect 9600 19256 9689 19284
rect 8294 19176 8300 19228
rect 8352 19216 8358 19228
rect 8941 19219 8999 19225
rect 8941 19216 8953 19219
rect 8352 19188 8953 19216
rect 8352 19176 8358 19188
rect 8941 19185 8953 19188
rect 8987 19185 8999 19219
rect 8941 19179 8999 19185
rect 1946 19108 1952 19160
rect 2004 19148 2010 19160
rect 3878 19148 3884 19160
rect 2004 19120 3884 19148
rect 2004 19108 2010 19120
rect 3878 19108 3884 19120
rect 3936 19108 3942 19160
rect 4065 19151 4123 19157
rect 4065 19117 4077 19151
rect 4111 19148 4123 19151
rect 4890 19148 4896 19160
rect 4111 19120 4896 19148
rect 4111 19117 4123 19120
rect 4065 19111 4123 19117
rect 2498 19040 2504 19092
rect 2556 19080 2562 19092
rect 3970 19080 3976 19092
rect 2556 19052 3976 19080
rect 2556 19040 2562 19052
rect 3970 19040 3976 19052
rect 4028 19040 4034 19092
rect 2406 18972 2412 19024
rect 2464 19012 2470 19024
rect 4080 19012 4108 19111
rect 4890 19108 4896 19120
rect 4948 19148 4954 19160
rect 6181 19151 6239 19157
rect 6181 19148 6193 19151
rect 4948 19120 6193 19148
rect 4948 19108 4954 19120
rect 6181 19117 6193 19120
rect 6227 19117 6239 19151
rect 6181 19111 6239 19117
rect 6270 19108 6276 19160
rect 6328 19148 6334 19160
rect 6437 19151 6495 19157
rect 6437 19148 6449 19151
rect 6328 19120 6449 19148
rect 6328 19108 6334 19120
rect 6437 19117 6449 19120
rect 6483 19117 6495 19151
rect 6437 19111 6495 19117
rect 8662 19108 8668 19160
rect 8720 19148 8726 19160
rect 8849 19151 8907 19157
rect 8849 19148 8861 19151
rect 8720 19120 8861 19148
rect 8720 19108 8726 19120
rect 8849 19117 8861 19120
rect 8895 19117 8907 19151
rect 8849 19111 8907 19117
rect 4246 19040 4252 19092
rect 4304 19089 4310 19092
rect 4304 19083 4368 19089
rect 4304 19049 4322 19083
rect 4356 19049 4368 19083
rect 9600 19080 9628 19256
rect 9677 19253 9689 19256
rect 9723 19253 9735 19287
rect 9677 19247 9735 19253
rect 12437 19287 12495 19293
rect 12437 19253 12449 19287
rect 12483 19253 12495 19287
rect 12437 19247 12495 19253
rect 9950 19176 9956 19228
rect 10008 19216 10014 19228
rect 10226 19216 10232 19228
rect 10008 19188 10232 19216
rect 10008 19176 10014 19188
rect 10226 19176 10232 19188
rect 10284 19176 10290 19228
rect 12452 19216 12480 19247
rect 19242 19216 19248 19228
rect 10888 19188 11192 19216
rect 12452 19188 12848 19216
rect 9674 19108 9680 19160
rect 9732 19148 9738 19160
rect 10045 19151 10103 19157
rect 10045 19148 10057 19151
rect 9732 19120 10057 19148
rect 9732 19108 9738 19120
rect 10045 19117 10057 19120
rect 10091 19117 10103 19151
rect 10045 19111 10103 19117
rect 10134 19108 10140 19160
rect 10192 19148 10198 19160
rect 10888 19148 10916 19188
rect 11054 19148 11060 19160
rect 10192 19120 10916 19148
rect 11015 19120 11060 19148
rect 10192 19108 10198 19120
rect 11054 19108 11060 19120
rect 11112 19108 11118 19160
rect 11164 19148 11192 19188
rect 12526 19148 12532 19160
rect 11164 19120 12532 19148
rect 12526 19108 12532 19120
rect 12584 19108 12590 19160
rect 12713 19151 12771 19157
rect 12713 19117 12725 19151
rect 12759 19117 12771 19151
rect 12820 19148 12848 19188
rect 18248 19188 19248 19216
rect 12986 19157 12992 19160
rect 12969 19151 12992 19157
rect 12969 19148 12981 19151
rect 12820 19120 12981 19148
rect 12713 19111 12771 19117
rect 12969 19117 12981 19120
rect 13044 19148 13050 19160
rect 15289 19151 15347 19157
rect 15289 19148 15301 19151
rect 13044 19120 13117 19148
rect 13556 19120 15301 19148
rect 12969 19111 12992 19117
rect 11146 19080 11152 19092
rect 4304 19043 4368 19049
rect 8404 19052 9352 19080
rect 9600 19052 11152 19080
rect 4304 19040 4310 19043
rect 5442 19012 5448 19024
rect 2464 18984 4108 19012
rect 5403 18984 5448 19012
rect 2464 18972 2470 18984
rect 5442 18972 5448 18984
rect 5500 18972 5506 19024
rect 7561 19015 7619 19021
rect 7561 18981 7573 19015
rect 7607 19012 7619 19015
rect 8294 19012 8300 19024
rect 7607 18984 8300 19012
rect 7607 18981 7619 18984
rect 7561 18975 7619 18981
rect 8294 18972 8300 18984
rect 8352 18972 8358 19024
rect 8404 19021 8432 19052
rect 8389 19015 8447 19021
rect 8389 18981 8401 19015
rect 8435 18981 8447 19015
rect 8754 19012 8760 19024
rect 8715 18984 8760 19012
rect 8389 18975 8447 18981
rect 8754 18972 8760 18984
rect 8812 18972 8818 19024
rect 9324 19012 9352 19052
rect 11146 19040 11152 19052
rect 11204 19040 11210 19092
rect 11324 19083 11382 19089
rect 11324 19049 11336 19083
rect 11370 19080 11382 19083
rect 11606 19080 11612 19092
rect 11370 19052 11612 19080
rect 11370 19049 11382 19052
rect 11324 19043 11382 19049
rect 11606 19040 11612 19052
rect 11664 19040 11670 19092
rect 12728 19080 12756 19111
rect 12986 19108 12992 19111
rect 13044 19108 13050 19120
rect 13556 19092 13584 19120
rect 15289 19117 15301 19120
rect 15335 19117 15347 19151
rect 17034 19148 17040 19160
rect 16995 19120 17040 19148
rect 15289 19111 15347 19117
rect 17034 19108 17040 19120
rect 17092 19108 17098 19160
rect 17313 19151 17371 19157
rect 17313 19117 17325 19151
rect 17359 19148 17371 19151
rect 18046 19148 18052 19160
rect 17359 19120 18052 19148
rect 17359 19117 17371 19120
rect 17313 19111 17371 19117
rect 18046 19108 18052 19120
rect 18104 19108 18110 19160
rect 18248 19157 18276 19188
rect 19242 19176 19248 19188
rect 19300 19176 19306 19228
rect 18233 19151 18291 19157
rect 18233 19117 18245 19151
rect 18279 19117 18291 19151
rect 18233 19111 18291 19117
rect 18322 19108 18328 19160
rect 18380 19148 18386 19160
rect 19521 19151 19579 19157
rect 19521 19148 19533 19151
rect 18380 19120 19533 19148
rect 18380 19108 18386 19120
rect 19521 19117 19533 19120
rect 19567 19117 19579 19151
rect 19521 19111 19579 19117
rect 19797 19151 19855 19157
rect 19797 19117 19809 19151
rect 19843 19148 19855 19151
rect 20257 19151 20315 19157
rect 20257 19148 20269 19151
rect 19843 19120 20269 19148
rect 19843 19117 19855 19120
rect 19797 19111 19855 19117
rect 20257 19117 20269 19120
rect 20303 19117 20315 19151
rect 20257 19111 20315 19117
rect 20901 19151 20959 19157
rect 20901 19117 20913 19151
rect 20947 19117 20959 19151
rect 20901 19111 20959 19117
rect 13538 19080 13544 19092
rect 12728 19052 13544 19080
rect 13538 19040 13544 19052
rect 13596 19040 13602 19092
rect 14734 19040 14740 19092
rect 14792 19080 14798 19092
rect 15534 19083 15592 19089
rect 15534 19080 15546 19083
rect 14792 19052 15546 19080
rect 14792 19040 14798 19052
rect 15534 19049 15546 19052
rect 15580 19049 15592 19083
rect 19058 19080 19064 19092
rect 19019 19052 19064 19080
rect 15534 19043 15592 19049
rect 19058 19040 19064 19052
rect 19116 19040 19122 19092
rect 10137 19015 10195 19021
rect 10137 19012 10149 19015
rect 9324 18984 10149 19012
rect 10137 18981 10149 18984
rect 10183 18981 10195 19015
rect 10137 18975 10195 18981
rect 10410 18972 10416 19024
rect 10468 19012 10474 19024
rect 10962 19012 10968 19024
rect 10468 18984 10968 19012
rect 10468 18972 10474 18984
rect 10962 18972 10968 18984
rect 11020 18972 11026 19024
rect 12526 18972 12532 19024
rect 12584 19012 12590 19024
rect 12894 19012 12900 19024
rect 12584 18984 12900 19012
rect 12584 18972 12590 18984
rect 12894 18972 12900 18984
rect 12952 18972 12958 19024
rect 14090 19012 14096 19024
rect 14051 18984 14096 19012
rect 14090 18972 14096 18984
rect 14148 18972 14154 19024
rect 16390 18972 16396 19024
rect 16448 19012 16454 19024
rect 16669 19015 16727 19021
rect 16669 19012 16681 19015
rect 16448 18984 16681 19012
rect 16448 18972 16454 18984
rect 16669 18981 16681 18984
rect 16715 18981 16727 19015
rect 16669 18975 16727 18981
rect 16758 18972 16764 19024
rect 16816 19012 16822 19024
rect 20916 19012 20944 19111
rect 16816 18984 20944 19012
rect 16816 18972 16822 18984
rect 1104 18922 21896 18944
rect 1104 18870 7912 18922
rect 7964 18870 7976 18922
rect 8028 18870 8040 18922
rect 8092 18870 8104 18922
rect 8156 18870 14843 18922
rect 14895 18870 14907 18922
rect 14959 18870 14971 18922
rect 15023 18870 15035 18922
rect 15087 18870 21896 18922
rect 1104 18848 21896 18870
rect 4154 18768 4160 18820
rect 4212 18808 4218 18820
rect 4525 18811 4583 18817
rect 4525 18808 4537 18811
rect 4212 18780 4537 18808
rect 4212 18768 4218 18780
rect 4525 18777 4537 18780
rect 4571 18808 4583 18811
rect 5077 18811 5135 18817
rect 5077 18808 5089 18811
rect 4571 18780 5089 18808
rect 4571 18777 4583 18780
rect 4525 18771 4583 18777
rect 5077 18777 5089 18780
rect 5123 18777 5135 18811
rect 6822 18808 6828 18820
rect 6783 18780 6828 18808
rect 5077 18771 5135 18777
rect 6822 18768 6828 18780
rect 6880 18768 6886 18820
rect 8570 18808 8576 18820
rect 6932 18780 8576 18808
rect 5810 18700 5816 18752
rect 5868 18740 5874 18752
rect 6932 18740 6960 18780
rect 8570 18768 8576 18780
rect 8628 18768 8634 18820
rect 8662 18768 8668 18820
rect 8720 18808 8726 18820
rect 9217 18811 9275 18817
rect 9217 18808 9229 18811
rect 8720 18780 9229 18808
rect 8720 18768 8726 18780
rect 9217 18777 9229 18780
rect 9263 18777 9275 18811
rect 9217 18771 9275 18777
rect 9401 18811 9459 18817
rect 9401 18777 9413 18811
rect 9447 18808 9459 18811
rect 9677 18811 9735 18817
rect 9677 18808 9689 18811
rect 9447 18780 9689 18808
rect 9447 18777 9459 18780
rect 9401 18771 9459 18777
rect 9677 18777 9689 18780
rect 9723 18808 9735 18811
rect 10134 18808 10140 18820
rect 9723 18780 10140 18808
rect 9723 18777 9735 18780
rect 9677 18771 9735 18777
rect 10134 18768 10140 18780
rect 10192 18768 10198 18820
rect 11422 18808 11428 18820
rect 10244 18780 11428 18808
rect 5868 18712 6960 18740
rect 5868 18700 5874 18712
rect 7006 18700 7012 18752
rect 7064 18740 7070 18752
rect 10244 18740 10272 18780
rect 11422 18768 11428 18780
rect 11480 18768 11486 18820
rect 11606 18808 11612 18820
rect 11567 18780 11612 18808
rect 11606 18768 11612 18780
rect 11664 18768 11670 18820
rect 14734 18768 14740 18820
rect 14792 18808 14798 18820
rect 14921 18811 14979 18817
rect 14921 18808 14933 18811
rect 14792 18780 14933 18808
rect 14792 18768 14798 18780
rect 14921 18777 14933 18780
rect 14967 18777 14979 18811
rect 14921 18771 14979 18777
rect 16485 18811 16543 18817
rect 16485 18777 16497 18811
rect 16531 18808 16543 18811
rect 18509 18811 18567 18817
rect 18509 18808 18521 18811
rect 16531 18780 18521 18808
rect 16531 18777 16543 18780
rect 16485 18771 16543 18777
rect 18509 18777 18521 18780
rect 18555 18777 18567 18811
rect 20990 18808 20996 18820
rect 18509 18771 18567 18777
rect 18616 18780 20852 18808
rect 20951 18780 20996 18808
rect 13808 18743 13866 18749
rect 7064 18712 10272 18740
rect 12544 18712 12940 18740
rect 7064 18700 7070 18712
rect 2676 18675 2734 18681
rect 2676 18641 2688 18675
rect 2722 18672 2734 18675
rect 3142 18672 3148 18684
rect 2722 18644 3148 18672
rect 2722 18641 2734 18644
rect 2676 18635 2734 18641
rect 3142 18632 3148 18644
rect 3200 18632 3206 18684
rect 4433 18675 4491 18681
rect 4433 18641 4445 18675
rect 4479 18672 4491 18675
rect 6273 18675 6331 18681
rect 4479 18644 5580 18672
rect 4479 18641 4491 18644
rect 4433 18635 4491 18641
rect 1762 18564 1768 18616
rect 1820 18604 1826 18616
rect 2406 18604 2412 18616
rect 1820 18576 2412 18604
rect 1820 18564 1826 18576
rect 2406 18564 2412 18576
rect 2464 18564 2470 18616
rect 4617 18607 4675 18613
rect 4617 18573 4629 18607
rect 4663 18573 4675 18607
rect 4617 18567 4675 18573
rect 3789 18539 3847 18545
rect 3789 18505 3801 18539
rect 3835 18536 3847 18539
rect 4246 18536 4252 18548
rect 3835 18508 4252 18536
rect 3835 18505 3847 18508
rect 3789 18499 3847 18505
rect 4246 18496 4252 18508
rect 4304 18536 4310 18548
rect 4632 18536 4660 18567
rect 4304 18508 4660 18536
rect 4304 18496 4310 18508
rect 4065 18471 4123 18477
rect 4065 18437 4077 18471
rect 4111 18468 4123 18471
rect 4338 18468 4344 18480
rect 4111 18440 4344 18468
rect 4111 18437 4123 18440
rect 4065 18431 4123 18437
rect 4338 18428 4344 18440
rect 4396 18428 4402 18480
rect 5552 18477 5580 18644
rect 6273 18641 6285 18675
rect 6319 18672 6331 18675
rect 7193 18675 7251 18681
rect 7193 18672 7205 18675
rect 6319 18644 7205 18672
rect 6319 18641 6331 18644
rect 6273 18635 6331 18641
rect 7193 18641 7205 18644
rect 7239 18641 7251 18675
rect 7193 18635 7251 18641
rect 8754 18632 8760 18684
rect 8812 18672 8818 18684
rect 9401 18675 9459 18681
rect 9401 18672 9413 18675
rect 8812 18644 9413 18672
rect 8812 18632 8818 18644
rect 9401 18641 9413 18644
rect 9447 18641 9459 18675
rect 9401 18635 9459 18641
rect 10496 18675 10554 18681
rect 10496 18641 10508 18675
rect 10542 18672 10554 18675
rect 10962 18672 10968 18684
rect 10542 18644 10968 18672
rect 10542 18641 10554 18644
rect 10496 18635 10554 18641
rect 10962 18632 10968 18644
rect 11020 18632 11026 18684
rect 12434 18632 12440 18684
rect 12492 18672 12498 18684
rect 12544 18672 12572 18712
rect 12492 18644 12572 18672
rect 12492 18632 12498 18644
rect 12710 18632 12716 18684
rect 12768 18672 12774 18684
rect 12805 18675 12863 18681
rect 12805 18672 12817 18675
rect 12768 18644 12817 18672
rect 12768 18632 12774 18644
rect 12805 18641 12817 18644
rect 12851 18641 12863 18675
rect 12912 18672 12940 18712
rect 13808 18709 13820 18743
rect 13854 18740 13866 18743
rect 14090 18740 14096 18752
rect 13854 18712 14096 18740
rect 13854 18709 13866 18712
rect 13808 18703 13866 18709
rect 14090 18700 14096 18712
rect 14148 18700 14154 18752
rect 16758 18740 16764 18752
rect 14200 18712 16764 18740
rect 14200 18672 14228 18712
rect 16758 18700 16764 18712
rect 16816 18700 16822 18752
rect 17126 18700 17132 18752
rect 17184 18740 17190 18752
rect 18414 18740 18420 18752
rect 17184 18712 18276 18740
rect 18375 18712 18420 18740
rect 17184 18700 17190 18712
rect 12912 18644 14228 18672
rect 12805 18635 12863 18641
rect 14274 18632 14280 18684
rect 14332 18672 14338 18684
rect 15654 18672 15660 18684
rect 14332 18644 15660 18672
rect 14332 18632 14338 18644
rect 15654 18632 15660 18644
rect 15712 18632 15718 18684
rect 16850 18672 16856 18684
rect 16763 18644 16856 18672
rect 16850 18632 16856 18644
rect 16908 18672 16914 18684
rect 17497 18675 17555 18681
rect 17497 18672 17509 18675
rect 16908 18644 17509 18672
rect 16908 18632 16914 18644
rect 17497 18641 17509 18644
rect 17543 18641 17555 18675
rect 18248 18672 18276 18712
rect 18414 18700 18420 18712
rect 18472 18700 18478 18752
rect 18616 18672 18644 18780
rect 19429 18743 19487 18749
rect 19429 18709 19441 18743
rect 19475 18740 19487 18743
rect 19978 18740 19984 18752
rect 19475 18712 19984 18740
rect 19475 18709 19487 18712
rect 19429 18703 19487 18709
rect 19978 18700 19984 18712
rect 20036 18700 20042 18752
rect 20162 18740 20168 18752
rect 20123 18712 20168 18740
rect 20162 18700 20168 18712
rect 20220 18700 20226 18752
rect 20824 18740 20852 18780
rect 20990 18768 20996 18780
rect 21048 18768 21054 18820
rect 21726 18740 21732 18752
rect 20824 18712 21732 18740
rect 21726 18700 21732 18712
rect 21784 18700 21790 18752
rect 19153 18675 19211 18681
rect 19153 18672 19165 18675
rect 18248 18644 18644 18672
rect 18708 18644 19165 18672
rect 17497 18635 17555 18641
rect 6638 18564 6644 18616
rect 6696 18604 6702 18616
rect 7285 18607 7343 18613
rect 7285 18604 7297 18607
rect 6696 18576 7297 18604
rect 6696 18564 6702 18576
rect 7285 18573 7297 18576
rect 7331 18573 7343 18607
rect 7285 18567 7343 18573
rect 7377 18607 7435 18613
rect 7377 18573 7389 18607
rect 7423 18573 7435 18607
rect 7377 18567 7435 18573
rect 6270 18496 6276 18548
rect 6328 18536 6334 18548
rect 7392 18536 7420 18567
rect 6328 18508 7420 18536
rect 6328 18496 6334 18508
rect 5537 18471 5595 18477
rect 5537 18437 5549 18471
rect 5583 18468 5595 18471
rect 8772 18468 8800 18632
rect 9674 18564 9680 18616
rect 9732 18604 9738 18616
rect 10134 18604 10140 18616
rect 9732 18576 10140 18604
rect 9732 18564 9738 18576
rect 10134 18564 10140 18576
rect 10192 18604 10198 18616
rect 10229 18607 10287 18613
rect 10229 18604 10241 18607
rect 10192 18576 10241 18604
rect 10192 18564 10198 18576
rect 10229 18573 10241 18576
rect 10275 18573 10287 18607
rect 12897 18607 12955 18613
rect 12897 18604 12909 18607
rect 10229 18567 10287 18573
rect 11992 18576 12909 18604
rect 5583 18440 8800 18468
rect 5583 18437 5595 18440
rect 5537 18431 5595 18437
rect 9766 18428 9772 18480
rect 9824 18468 9830 18480
rect 11992 18477 12020 18576
rect 12897 18573 12909 18576
rect 12943 18573 12955 18607
rect 12897 18567 12955 18573
rect 12986 18564 12992 18616
rect 13044 18604 13050 18616
rect 13538 18604 13544 18616
rect 13044 18576 13089 18604
rect 13499 18576 13544 18604
rect 13044 18564 13050 18576
rect 13538 18564 13544 18576
rect 13596 18564 13602 18616
rect 16945 18607 17003 18613
rect 16945 18604 16957 18607
rect 16132 18576 16957 18604
rect 11977 18471 12035 18477
rect 11977 18468 11989 18471
rect 9824 18440 11989 18468
rect 9824 18428 9830 18440
rect 11977 18437 11989 18440
rect 12023 18437 12035 18471
rect 11977 18431 12035 18437
rect 12437 18471 12495 18477
rect 12437 18437 12449 18471
rect 12483 18468 12495 18471
rect 13906 18468 13912 18480
rect 12483 18440 13912 18468
rect 12483 18437 12495 18440
rect 12437 18431 12495 18437
rect 13906 18428 13912 18440
rect 13964 18428 13970 18480
rect 15470 18428 15476 18480
rect 15528 18468 15534 18480
rect 16132 18477 16160 18576
rect 16945 18573 16957 18576
rect 16991 18573 17003 18607
rect 16945 18567 17003 18573
rect 17034 18564 17040 18616
rect 17092 18604 17098 18616
rect 18598 18604 18604 18616
rect 17092 18576 17137 18604
rect 18559 18576 18604 18604
rect 17092 18564 17098 18576
rect 18598 18564 18604 18576
rect 18656 18564 18662 18616
rect 16206 18496 16212 18548
rect 16264 18536 16270 18548
rect 18049 18539 18107 18545
rect 16264 18508 17632 18536
rect 16264 18496 16270 18508
rect 16117 18471 16175 18477
rect 16117 18468 16129 18471
rect 15528 18440 16129 18468
rect 15528 18428 15534 18440
rect 16117 18437 16129 18440
rect 16163 18437 16175 18471
rect 17604 18468 17632 18508
rect 18049 18505 18061 18539
rect 18095 18536 18107 18539
rect 18708 18536 18736 18644
rect 19153 18641 19165 18644
rect 19199 18641 19211 18675
rect 19153 18635 19211 18641
rect 19889 18675 19947 18681
rect 19889 18641 19901 18675
rect 19935 18641 19947 18675
rect 20806 18672 20812 18684
rect 20767 18644 20812 18672
rect 19889 18635 19947 18641
rect 18095 18508 18736 18536
rect 18095 18505 18107 18508
rect 18049 18499 18107 18505
rect 19904 18468 19932 18635
rect 20806 18632 20812 18644
rect 20864 18632 20870 18684
rect 17604 18440 19932 18468
rect 16117 18431 16175 18437
rect 1104 18378 21896 18400
rect 1104 18326 4447 18378
rect 4499 18326 4511 18378
rect 4563 18326 4575 18378
rect 4627 18326 4639 18378
rect 4691 18326 11378 18378
rect 11430 18326 11442 18378
rect 11494 18326 11506 18378
rect 11558 18326 11570 18378
rect 11622 18326 18308 18378
rect 18360 18326 18372 18378
rect 18424 18326 18436 18378
rect 18488 18326 18500 18378
rect 18552 18326 21896 18378
rect 1104 18304 21896 18326
rect 6362 18264 6368 18276
rect 5184 18236 6368 18264
rect 290 18156 296 18208
rect 348 18196 354 18208
rect 5184 18196 5212 18236
rect 6362 18224 6368 18236
rect 6420 18224 6426 18276
rect 6638 18264 6644 18276
rect 6599 18236 6644 18264
rect 6638 18224 6644 18236
rect 6696 18224 6702 18276
rect 7561 18267 7619 18273
rect 7561 18264 7573 18267
rect 7024 18236 7573 18264
rect 348 18168 5212 18196
rect 348 18156 354 18168
rect 5258 18156 5264 18208
rect 5316 18196 5322 18208
rect 7024 18196 7052 18236
rect 7561 18233 7573 18236
rect 7607 18233 7619 18267
rect 7561 18227 7619 18233
rect 7745 18267 7803 18273
rect 7745 18233 7757 18267
rect 7791 18264 7803 18267
rect 8202 18264 8208 18276
rect 7791 18236 8208 18264
rect 7791 18233 7803 18236
rect 7745 18227 7803 18233
rect 7760 18196 7788 18227
rect 8202 18224 8208 18236
rect 8260 18224 8266 18276
rect 9692 18236 10916 18264
rect 5316 18168 7052 18196
rect 7116 18168 7788 18196
rect 5316 18156 5322 18168
rect 1394 18088 1400 18140
rect 1452 18128 1458 18140
rect 6638 18128 6644 18140
rect 1452 18100 6644 18128
rect 1452 18088 1458 18100
rect 6638 18088 6644 18100
rect 6696 18088 6702 18140
rect 7116 18137 7144 18168
rect 7926 18156 7932 18208
rect 7984 18196 7990 18208
rect 9692 18196 9720 18236
rect 7984 18168 9720 18196
rect 10888 18196 10916 18236
rect 10962 18224 10968 18276
rect 11020 18264 11026 18276
rect 11057 18267 11115 18273
rect 11057 18264 11069 18267
rect 11020 18236 11069 18264
rect 11020 18224 11026 18236
rect 11057 18233 11069 18236
rect 11103 18233 11115 18267
rect 12434 18264 12440 18276
rect 11057 18227 11115 18233
rect 11164 18236 12440 18264
rect 11164 18196 11192 18236
rect 12434 18224 12440 18236
rect 12492 18224 12498 18276
rect 12526 18224 12532 18276
rect 12584 18264 12590 18276
rect 15286 18264 15292 18276
rect 12584 18236 15292 18264
rect 12584 18224 12590 18236
rect 15286 18224 15292 18236
rect 15344 18224 15350 18276
rect 16206 18264 16212 18276
rect 15580 18236 16212 18264
rect 10888 18168 11192 18196
rect 11333 18199 11391 18205
rect 7984 18156 7990 18168
rect 11333 18165 11345 18199
rect 11379 18196 11391 18199
rect 15580 18196 15608 18236
rect 16206 18224 16212 18236
rect 16264 18224 16270 18276
rect 16945 18267 17003 18273
rect 16945 18233 16957 18267
rect 16991 18264 17003 18267
rect 17034 18264 17040 18276
rect 16991 18236 17040 18264
rect 16991 18233 17003 18236
rect 16945 18227 17003 18233
rect 17034 18224 17040 18236
rect 17092 18224 17098 18276
rect 17862 18224 17868 18276
rect 17920 18264 17926 18276
rect 21634 18264 21640 18276
rect 17920 18236 21640 18264
rect 17920 18224 17926 18236
rect 21634 18224 21640 18236
rect 21692 18224 21698 18276
rect 11379 18168 15608 18196
rect 11379 18165 11391 18168
rect 11333 18159 11391 18165
rect 7101 18131 7159 18137
rect 7101 18097 7113 18131
rect 7147 18097 7159 18131
rect 7101 18091 7159 18097
rect 7193 18131 7251 18137
rect 7193 18097 7205 18131
rect 7239 18097 7251 18131
rect 7193 18091 7251 18097
rect 7561 18131 7619 18137
rect 7561 18097 7573 18131
rect 7607 18128 7619 18131
rect 7607 18100 9812 18128
rect 7607 18097 7619 18100
rect 7561 18091 7619 18097
rect 6546 18020 6552 18072
rect 6604 18060 6610 18072
rect 7208 18060 7236 18091
rect 9784 18072 9812 18100
rect 11698 18088 11704 18140
rect 11756 18128 11762 18140
rect 11885 18131 11943 18137
rect 11885 18128 11897 18131
rect 11756 18100 11897 18128
rect 11756 18088 11762 18100
rect 11885 18097 11897 18100
rect 11931 18097 11943 18131
rect 13906 18128 13912 18140
rect 13867 18100 13912 18128
rect 11885 18091 11943 18097
rect 13906 18088 13912 18100
rect 13964 18088 13970 18140
rect 14090 18128 14096 18140
rect 14051 18100 14096 18128
rect 14090 18088 14096 18100
rect 14148 18088 14154 18140
rect 14277 18131 14335 18137
rect 14277 18097 14289 18131
rect 14323 18128 14335 18131
rect 17052 18128 17080 18224
rect 18690 18156 18696 18208
rect 18748 18196 18754 18208
rect 21450 18196 21456 18208
rect 18748 18168 21456 18196
rect 18748 18156 18754 18168
rect 21450 18156 21456 18168
rect 21508 18156 21514 18208
rect 18874 18128 18880 18140
rect 14323 18100 15700 18128
rect 17052 18100 17356 18128
rect 18835 18100 18880 18128
rect 14323 18097 14335 18100
rect 14277 18091 14335 18097
rect 9674 18060 9680 18072
rect 6604 18032 7236 18060
rect 9635 18032 9680 18060
rect 6604 18020 6610 18032
rect 9674 18020 9680 18032
rect 9732 18020 9738 18072
rect 9766 18020 9772 18072
rect 9824 18020 9830 18072
rect 9950 18069 9956 18072
rect 9944 18060 9956 18069
rect 9911 18032 9956 18060
rect 9944 18023 9956 18032
rect 9950 18020 9956 18023
rect 10008 18020 10014 18072
rect 10870 18020 10876 18072
rect 10928 18060 10934 18072
rect 15470 18060 15476 18072
rect 10928 18032 15476 18060
rect 10928 18020 10934 18032
rect 15470 18020 15476 18032
rect 15528 18020 15534 18072
rect 15565 18063 15623 18069
rect 15565 18029 15577 18063
rect 15611 18029 15623 18063
rect 15565 18023 15623 18029
rect 6454 17952 6460 18004
rect 6512 17992 6518 18004
rect 11238 17992 11244 18004
rect 6512 17964 11244 17992
rect 6512 17952 6518 17964
rect 11238 17952 11244 17964
rect 11296 17952 11302 18004
rect 11701 17995 11759 18001
rect 11701 17961 11713 17995
rect 11747 17992 11759 17995
rect 12345 17995 12403 18001
rect 12345 17992 12357 17995
rect 11747 17964 12357 17992
rect 11747 17961 11759 17964
rect 11701 17955 11759 17961
rect 12345 17961 12357 17964
rect 12391 17961 12403 17995
rect 12345 17955 12403 17961
rect 12894 17952 12900 18004
rect 12952 17992 12958 18004
rect 13722 17992 13728 18004
rect 12952 17964 13728 17992
rect 12952 17952 12958 17964
rect 13722 17952 13728 17964
rect 13780 17952 13786 18004
rect 13817 17995 13875 18001
rect 13817 17961 13829 17995
rect 13863 17992 13875 17995
rect 14461 17995 14519 18001
rect 14461 17992 14473 17995
rect 13863 17964 14473 17992
rect 13863 17961 13875 17964
rect 13817 17955 13875 17961
rect 14461 17961 14473 17964
rect 14507 17961 14519 17995
rect 14461 17955 14519 17961
rect 14734 17952 14740 18004
rect 14792 17992 14798 18004
rect 15580 17992 15608 18023
rect 14792 17964 15608 17992
rect 15672 17992 15700 18100
rect 15832 18063 15890 18069
rect 15832 18029 15844 18063
rect 15878 18060 15890 18063
rect 16390 18060 16396 18072
rect 15878 18032 16396 18060
rect 15878 18029 15890 18032
rect 15832 18023 15890 18029
rect 16390 18020 16396 18032
rect 16448 18020 16454 18072
rect 17218 18060 17224 18072
rect 17179 18032 17224 18060
rect 17218 18020 17224 18032
rect 17276 18020 17282 18072
rect 17328 18060 17356 18100
rect 18874 18088 18880 18100
rect 18932 18088 18938 18140
rect 20162 18088 20168 18140
rect 20220 18128 20226 18140
rect 21542 18128 21548 18140
rect 20220 18100 21548 18128
rect 20220 18088 20226 18100
rect 21542 18088 21548 18100
rect 21600 18088 21606 18140
rect 17477 18063 17535 18069
rect 17477 18060 17489 18063
rect 17328 18032 17489 18060
rect 17477 18029 17489 18032
rect 17523 18029 17535 18063
rect 17477 18023 17535 18029
rect 20070 18020 20076 18072
rect 20128 18060 20134 18072
rect 20901 18063 20959 18069
rect 20901 18060 20913 18063
rect 20128 18032 20913 18060
rect 20128 18020 20134 18032
rect 20901 18029 20913 18032
rect 20947 18029 20959 18063
rect 20901 18023 20959 18029
rect 18138 17992 18144 18004
rect 15672 17964 18144 17992
rect 14792 17952 14798 17964
rect 18138 17952 18144 17964
rect 18196 17952 18202 18004
rect 18782 17952 18788 18004
rect 18840 17992 18846 18004
rect 19610 17992 19616 18004
rect 18840 17964 19616 17992
rect 18840 17952 18846 17964
rect 19610 17952 19616 17964
rect 19668 17952 19674 18004
rect 20530 17952 20536 18004
rect 20588 17992 20594 18004
rect 22094 17992 22100 18004
rect 20588 17964 22100 17992
rect 20588 17952 20594 17964
rect 22094 17952 22100 17964
rect 22152 17952 22158 18004
rect 3050 17884 3056 17936
rect 3108 17924 3114 17936
rect 4154 17924 4160 17936
rect 3108 17896 4160 17924
rect 3108 17884 3114 17896
rect 4154 17884 4160 17896
rect 4212 17884 4218 17936
rect 4798 17884 4804 17936
rect 4856 17924 4862 17936
rect 6730 17924 6736 17936
rect 4856 17896 6736 17924
rect 4856 17884 4862 17896
rect 6730 17884 6736 17896
rect 6788 17884 6794 17936
rect 7009 17927 7067 17933
rect 7009 17893 7021 17927
rect 7055 17924 7067 17927
rect 7466 17924 7472 17936
rect 7055 17896 7472 17924
rect 7055 17893 7067 17896
rect 7009 17887 7067 17893
rect 7466 17884 7472 17896
rect 7524 17924 7530 17936
rect 8021 17927 8079 17933
rect 8021 17924 8033 17927
rect 7524 17896 8033 17924
rect 7524 17884 7530 17896
rect 8021 17893 8033 17896
rect 8067 17893 8079 17927
rect 8021 17887 8079 17893
rect 8570 17884 8576 17936
rect 8628 17924 8634 17936
rect 11146 17924 11152 17936
rect 8628 17896 11152 17924
rect 8628 17884 8634 17896
rect 11146 17884 11152 17896
rect 11204 17884 11210 17936
rect 11790 17924 11796 17936
rect 11751 17896 11796 17924
rect 11790 17884 11796 17896
rect 11848 17884 11854 17936
rect 11882 17884 11888 17936
rect 11940 17924 11946 17936
rect 12526 17924 12532 17936
rect 11940 17896 12532 17924
rect 11940 17884 11946 17896
rect 12526 17884 12532 17896
rect 12584 17884 12590 17936
rect 12710 17884 12716 17936
rect 12768 17924 12774 17936
rect 13081 17927 13139 17933
rect 13081 17924 13093 17927
rect 12768 17896 13093 17924
rect 12768 17884 12774 17896
rect 13081 17893 13093 17896
rect 13127 17893 13139 17927
rect 13081 17887 13139 17893
rect 13449 17927 13507 17933
rect 13449 17893 13461 17927
rect 13495 17924 13507 17927
rect 14277 17927 14335 17933
rect 14277 17924 14289 17927
rect 13495 17896 14289 17924
rect 13495 17893 13507 17896
rect 13449 17887 13507 17893
rect 14277 17893 14289 17896
rect 14323 17893 14335 17927
rect 14277 17887 14335 17893
rect 15378 17884 15384 17936
rect 15436 17924 15442 17936
rect 15838 17924 15844 17936
rect 15436 17896 15844 17924
rect 15436 17884 15442 17896
rect 15838 17884 15844 17896
rect 15896 17884 15902 17936
rect 18598 17924 18604 17936
rect 18559 17896 18604 17924
rect 18598 17884 18604 17896
rect 18656 17924 18662 17936
rect 19337 17927 19395 17933
rect 19337 17924 19349 17927
rect 18656 17896 19349 17924
rect 18656 17884 18662 17896
rect 19337 17893 19349 17896
rect 19383 17893 19395 17927
rect 19337 17887 19395 17893
rect 19794 17884 19800 17936
rect 19852 17924 19858 17936
rect 20346 17924 20352 17936
rect 19852 17896 20352 17924
rect 19852 17884 19858 17896
rect 20346 17884 20352 17896
rect 20404 17884 20410 17936
rect 21082 17924 21088 17936
rect 21043 17896 21088 17924
rect 21082 17884 21088 17896
rect 21140 17884 21146 17936
rect 21174 17884 21180 17936
rect 21232 17924 21238 17936
rect 22646 17924 22652 17936
rect 21232 17896 22652 17924
rect 21232 17884 21238 17896
rect 22646 17884 22652 17896
rect 22704 17884 22710 17936
rect 1104 17834 21896 17856
rect 1104 17782 7912 17834
rect 7964 17782 7976 17834
rect 8028 17782 8040 17834
rect 8092 17782 8104 17834
rect 8156 17782 14843 17834
rect 14895 17782 14907 17834
rect 14959 17782 14971 17834
rect 15023 17782 15035 17834
rect 15087 17782 21896 17834
rect 1104 17760 21896 17782
rect 4338 17680 4344 17732
rect 4396 17720 4402 17732
rect 4709 17723 4767 17729
rect 4709 17720 4721 17723
rect 4396 17692 4721 17720
rect 4396 17680 4402 17692
rect 4709 17689 4721 17692
rect 4755 17689 4767 17723
rect 4709 17683 4767 17689
rect 9214 17680 9220 17732
rect 9272 17720 9278 17732
rect 9493 17723 9551 17729
rect 9493 17720 9505 17723
rect 9272 17692 9505 17720
rect 9272 17680 9278 17692
rect 9493 17689 9505 17692
rect 9539 17689 9551 17723
rect 9493 17683 9551 17689
rect 9861 17723 9919 17729
rect 9861 17689 9873 17723
rect 9907 17720 9919 17723
rect 11790 17720 11796 17732
rect 9907 17692 11796 17720
rect 9907 17689 9919 17692
rect 9861 17683 9919 17689
rect 9508 17652 9536 17683
rect 11790 17680 11796 17692
rect 11848 17680 11854 17732
rect 12526 17680 12532 17732
rect 12584 17720 12590 17732
rect 15194 17720 15200 17732
rect 12584 17692 15200 17720
rect 12584 17680 12590 17692
rect 15194 17680 15200 17692
rect 15252 17680 15258 17732
rect 19518 17720 19524 17732
rect 19479 17692 19524 17720
rect 19518 17680 19524 17692
rect 19576 17680 19582 17732
rect 10321 17655 10379 17661
rect 10321 17652 10333 17655
rect 9508 17624 10333 17652
rect 10321 17621 10333 17624
rect 10367 17621 10379 17655
rect 10321 17615 10379 17621
rect 4338 17544 4344 17596
rect 4396 17584 4402 17596
rect 4617 17587 4675 17593
rect 4617 17584 4629 17587
rect 4396 17556 4629 17584
rect 4396 17544 4402 17556
rect 4617 17553 4629 17556
rect 4663 17553 4675 17587
rect 4617 17547 4675 17553
rect 8021 17587 8079 17593
rect 8021 17553 8033 17587
rect 8067 17584 8079 17587
rect 9858 17584 9864 17596
rect 8067 17556 9864 17584
rect 8067 17553 8079 17556
rect 8021 17547 8079 17553
rect 9858 17544 9864 17556
rect 9916 17584 9922 17596
rect 10229 17587 10287 17593
rect 10229 17584 10241 17587
rect 9916 17556 10241 17584
rect 9916 17544 9922 17556
rect 10229 17553 10241 17556
rect 10275 17584 10287 17587
rect 10873 17587 10931 17593
rect 10873 17584 10885 17587
rect 10275 17556 10885 17584
rect 10275 17553 10287 17556
rect 10229 17547 10287 17553
rect 10873 17553 10885 17556
rect 10919 17553 10931 17587
rect 18598 17584 18604 17596
rect 10873 17547 10931 17553
rect 13372 17556 18604 17584
rect 4893 17519 4951 17525
rect 4893 17485 4905 17519
rect 4939 17516 4951 17519
rect 5442 17516 5448 17528
rect 4939 17488 5448 17516
rect 4939 17485 4951 17488
rect 4893 17479 4951 17485
rect 5442 17476 5448 17488
rect 5500 17476 5506 17528
rect 10505 17519 10563 17525
rect 10505 17485 10517 17519
rect 10551 17516 10563 17519
rect 10962 17516 10968 17528
rect 10551 17488 10968 17516
rect 10551 17485 10563 17488
rect 10505 17479 10563 17485
rect 10962 17476 10968 17488
rect 11020 17476 11026 17528
rect 13372 17516 13400 17556
rect 18598 17544 18604 17556
rect 18656 17544 18662 17596
rect 18874 17544 18880 17596
rect 18932 17584 18938 17596
rect 19337 17587 19395 17593
rect 19337 17584 19349 17587
rect 18932 17556 19349 17584
rect 18932 17544 18938 17556
rect 19337 17553 19349 17556
rect 19383 17553 19395 17587
rect 19337 17547 19395 17553
rect 20257 17587 20315 17593
rect 20257 17553 20269 17587
rect 20303 17584 20315 17587
rect 20714 17584 20720 17596
rect 20303 17556 20720 17584
rect 20303 17553 20315 17556
rect 20257 17547 20315 17553
rect 20714 17544 20720 17556
rect 20772 17544 20778 17596
rect 20809 17587 20867 17593
rect 20809 17553 20821 17587
rect 20855 17553 20867 17587
rect 20809 17547 20867 17553
rect 20824 17516 20852 17547
rect 12360 17488 13400 17516
rect 13464 17488 20852 17516
rect 4798 17408 4804 17460
rect 4856 17448 4862 17460
rect 12360 17448 12388 17488
rect 4856 17420 12388 17448
rect 4856 17408 4862 17420
rect 4246 17380 4252 17392
rect 4207 17352 4252 17380
rect 4246 17340 4252 17352
rect 4304 17340 4310 17392
rect 8938 17340 8944 17392
rect 8996 17380 9002 17392
rect 13464 17380 13492 17488
rect 20438 17448 20444 17460
rect 20399 17420 20444 17448
rect 20438 17408 20444 17420
rect 20496 17408 20502 17460
rect 20990 17380 20996 17392
rect 8996 17352 13492 17380
rect 20951 17352 20996 17380
rect 8996 17340 9002 17352
rect 20990 17340 20996 17352
rect 21048 17340 21054 17392
rect 1104 17290 21896 17312
rect 1104 17238 4447 17290
rect 4499 17238 4511 17290
rect 4563 17238 4575 17290
rect 4627 17238 4639 17290
rect 4691 17238 11378 17290
rect 11430 17238 11442 17290
rect 11494 17238 11506 17290
rect 11558 17238 11570 17290
rect 11622 17238 18308 17290
rect 18360 17238 18372 17290
rect 18424 17238 18436 17290
rect 18488 17238 18500 17290
rect 18552 17238 21896 17290
rect 1104 17216 21896 17238
rect 3142 17176 3148 17188
rect 3103 17148 3148 17176
rect 3142 17136 3148 17148
rect 3200 17176 3206 17188
rect 3326 17176 3332 17188
rect 3200 17148 3332 17176
rect 3200 17136 3206 17148
rect 3326 17136 3332 17148
rect 3384 17136 3390 17188
rect 3510 17136 3516 17188
rect 3568 17176 3574 17188
rect 6730 17176 6736 17188
rect 3568 17148 6316 17176
rect 6691 17148 6736 17176
rect 3568 17136 3574 17148
rect 6181 17111 6239 17117
rect 6181 17077 6193 17111
rect 6227 17077 6239 17111
rect 6288 17108 6316 17148
rect 6730 17136 6736 17148
rect 6788 17136 6794 17188
rect 19702 17176 19708 17188
rect 6840 17148 19708 17176
rect 6840 17108 6868 17148
rect 19702 17136 19708 17148
rect 19760 17136 19766 17188
rect 6288 17080 6868 17108
rect 7101 17111 7159 17117
rect 6181 17071 6239 17077
rect 7101 17077 7113 17111
rect 7147 17108 7159 17111
rect 8941 17111 8999 17117
rect 8941 17108 8953 17111
rect 7147 17080 8953 17108
rect 7147 17077 7159 17080
rect 7101 17071 7159 17077
rect 8941 17077 8953 17080
rect 8987 17077 8999 17111
rect 8941 17071 8999 17077
rect 4338 17040 4344 17052
rect 4299 17012 4344 17040
rect 4338 17000 4344 17012
rect 4396 17000 4402 17052
rect 6196 17040 6224 17071
rect 9766 17068 9772 17120
rect 9824 17108 9830 17120
rect 10321 17111 10379 17117
rect 10321 17108 10333 17111
rect 9824 17080 10333 17108
rect 9824 17068 9830 17080
rect 10321 17077 10333 17080
rect 10367 17108 10379 17111
rect 10962 17108 10968 17120
rect 10367 17080 10968 17108
rect 10367 17077 10379 17080
rect 10321 17071 10379 17077
rect 10962 17068 10968 17080
rect 11020 17068 11026 17120
rect 11425 17111 11483 17117
rect 11425 17077 11437 17111
rect 11471 17108 11483 17111
rect 20438 17108 20444 17120
rect 11471 17080 20444 17108
rect 11471 17077 11483 17080
rect 11425 17071 11483 17077
rect 20438 17068 20444 17080
rect 20496 17068 20502 17120
rect 7006 17040 7012 17052
rect 6196 17012 7012 17040
rect 7006 17000 7012 17012
rect 7064 17040 7070 17052
rect 7653 17043 7711 17049
rect 7653 17040 7665 17043
rect 7064 17012 7665 17040
rect 7064 17000 7070 17012
rect 7653 17009 7665 17012
rect 7699 17009 7711 17043
rect 8662 17040 8668 17052
rect 8623 17012 8668 17040
rect 7653 17003 7711 17009
rect 8662 17000 8668 17012
rect 8720 17000 8726 17052
rect 12069 17043 12127 17049
rect 12069 17009 12081 17043
rect 12115 17040 12127 17043
rect 12158 17040 12164 17052
rect 12115 17012 12164 17040
rect 12115 17009 12127 17012
rect 12069 17003 12127 17009
rect 12158 17000 12164 17012
rect 12216 17000 12222 17052
rect 14366 17000 14372 17052
rect 14424 17040 14430 17052
rect 18874 17040 18880 17052
rect 14424 17012 18736 17040
rect 18835 17012 18880 17040
rect 14424 17000 14430 17012
rect 1762 16972 1768 16984
rect 1723 16944 1768 16972
rect 1762 16932 1768 16944
rect 1820 16932 1826 16984
rect 4801 16975 4859 16981
rect 4801 16941 4813 16975
rect 4847 16972 4859 16975
rect 4890 16972 4896 16984
rect 4847 16944 4896 16972
rect 4847 16941 4859 16944
rect 4801 16935 4859 16941
rect 4890 16932 4896 16944
rect 4948 16932 4954 16984
rect 5068 16975 5126 16981
rect 5068 16941 5080 16975
rect 5114 16972 5126 16975
rect 5442 16972 5448 16984
rect 5114 16944 5448 16972
rect 5114 16941 5126 16944
rect 5068 16935 5126 16941
rect 5442 16932 5448 16944
rect 5500 16932 5506 16984
rect 6730 16932 6736 16984
rect 6788 16972 6794 16984
rect 7561 16975 7619 16981
rect 7561 16972 7573 16975
rect 6788 16944 7573 16972
rect 6788 16932 6794 16944
rect 7561 16941 7573 16944
rect 7607 16941 7619 16975
rect 9858 16972 9864 16984
rect 7561 16935 7619 16941
rect 8404 16944 9864 16972
rect 2032 16907 2090 16913
rect 2032 16873 2044 16907
rect 2078 16904 2090 16907
rect 3694 16904 3700 16916
rect 2078 16876 3700 16904
rect 2078 16873 2090 16876
rect 2032 16867 2090 16873
rect 3694 16864 3700 16876
rect 3752 16864 3758 16916
rect 7469 16907 7527 16913
rect 7469 16873 7481 16907
rect 7515 16904 7527 16907
rect 8404 16904 8432 16944
rect 9858 16932 9864 16944
rect 9916 16932 9922 16984
rect 10870 16932 10876 16984
rect 10928 16972 10934 16984
rect 11149 16975 11207 16981
rect 11149 16972 11161 16975
rect 10928 16944 11161 16972
rect 10928 16932 10934 16944
rect 11149 16941 11161 16944
rect 11195 16972 11207 16975
rect 12710 16972 12716 16984
rect 11195 16944 12716 16972
rect 11195 16941 11207 16944
rect 11149 16935 11207 16941
rect 12710 16932 12716 16944
rect 12768 16932 12774 16984
rect 15286 16932 15292 16984
rect 15344 16972 15350 16984
rect 15746 16972 15752 16984
rect 15344 16944 15752 16972
rect 15344 16932 15350 16944
rect 15746 16932 15752 16944
rect 15804 16932 15810 16984
rect 18046 16932 18052 16984
rect 18104 16972 18110 16984
rect 18601 16975 18659 16981
rect 18601 16972 18613 16975
rect 18104 16944 18613 16972
rect 18104 16932 18110 16944
rect 18601 16941 18613 16944
rect 18647 16941 18659 16975
rect 18708 16972 18736 17012
rect 18874 17000 18880 17012
rect 18932 17000 18938 17052
rect 20070 17040 20076 17052
rect 20031 17012 20076 17040
rect 20070 17000 20076 17012
rect 20128 17000 20134 17052
rect 19797 16975 19855 16981
rect 19797 16972 19809 16975
rect 18708 16944 19809 16972
rect 18601 16935 18659 16941
rect 19797 16941 19809 16944
rect 19843 16941 19855 16975
rect 19797 16935 19855 16941
rect 20901 16975 20959 16981
rect 20901 16941 20913 16975
rect 20947 16941 20959 16975
rect 20901 16935 20959 16941
rect 7515 16876 8432 16904
rect 8481 16907 8539 16913
rect 7515 16873 7527 16876
rect 7469 16867 7527 16873
rect 8481 16873 8493 16907
rect 8527 16904 8539 16907
rect 9125 16907 9183 16913
rect 9125 16904 9137 16907
rect 8527 16876 9137 16904
rect 8527 16873 8539 16876
rect 8481 16867 8539 16873
rect 9125 16873 9137 16876
rect 9171 16873 9183 16907
rect 9125 16867 9183 16873
rect 10502 16864 10508 16916
rect 10560 16904 10566 16916
rect 11885 16907 11943 16913
rect 11885 16904 11897 16907
rect 10560 16876 11897 16904
rect 10560 16864 10566 16876
rect 11885 16873 11897 16876
rect 11931 16873 11943 16907
rect 11885 16867 11943 16873
rect 12526 16864 12532 16916
rect 12584 16904 12590 16916
rect 20916 16904 20944 16935
rect 12584 16876 20944 16904
rect 12584 16864 12590 16876
rect 3418 16836 3424 16848
rect 3379 16808 3424 16836
rect 3418 16796 3424 16808
rect 3476 16796 3482 16848
rect 8113 16839 8171 16845
rect 8113 16805 8125 16839
rect 8159 16836 8171 16839
rect 8386 16836 8392 16848
rect 8159 16808 8392 16836
rect 8159 16805 8171 16808
rect 8113 16799 8171 16805
rect 8386 16796 8392 16808
rect 8444 16796 8450 16848
rect 8573 16839 8631 16845
rect 8573 16805 8585 16839
rect 8619 16836 8631 16839
rect 8941 16839 8999 16845
rect 8941 16836 8953 16839
rect 8619 16808 8953 16836
rect 8619 16805 8631 16808
rect 8573 16799 8631 16805
rect 8941 16805 8953 16808
rect 8987 16805 8999 16839
rect 11790 16836 11796 16848
rect 11751 16808 11796 16836
rect 8941 16799 8999 16805
rect 11790 16796 11796 16808
rect 11848 16796 11854 16848
rect 19334 16796 19340 16848
rect 19392 16836 19398 16848
rect 19978 16836 19984 16848
rect 19392 16808 19984 16836
rect 19392 16796 19398 16808
rect 19978 16796 19984 16808
rect 20036 16796 20042 16848
rect 21082 16836 21088 16848
rect 21043 16808 21088 16836
rect 21082 16796 21088 16808
rect 21140 16796 21146 16848
rect 1104 16746 21896 16768
rect 1104 16694 7912 16746
rect 7964 16694 7976 16746
rect 8028 16694 8040 16746
rect 8092 16694 8104 16746
rect 8156 16694 14843 16746
rect 14895 16694 14907 16746
rect 14959 16694 14971 16746
rect 15023 16694 15035 16746
rect 15087 16694 21896 16746
rect 1104 16672 21896 16694
rect 3602 16632 3608 16644
rect 3563 16604 3608 16632
rect 3602 16592 3608 16604
rect 3660 16632 3666 16644
rect 4157 16635 4215 16641
rect 4157 16632 4169 16635
rect 3660 16604 4169 16632
rect 3660 16592 3666 16604
rect 4157 16601 4169 16604
rect 4203 16601 4215 16635
rect 4157 16595 4215 16601
rect 8205 16635 8263 16641
rect 8205 16601 8217 16635
rect 8251 16601 8263 16635
rect 10502 16632 10508 16644
rect 10463 16604 10508 16632
rect 8205 16595 8263 16601
rect 7006 16524 7012 16576
rect 7064 16573 7070 16576
rect 7064 16567 7128 16573
rect 7064 16533 7082 16567
rect 7116 16533 7128 16567
rect 8220 16564 8248 16595
rect 10502 16592 10508 16604
rect 10560 16592 10566 16644
rect 10870 16632 10876 16644
rect 10831 16604 10876 16632
rect 10870 16592 10876 16604
rect 10928 16592 10934 16644
rect 10962 16592 10968 16644
rect 11020 16632 11026 16644
rect 11790 16632 11796 16644
rect 11020 16604 11065 16632
rect 11751 16604 11796 16632
rect 11020 16592 11026 16604
rect 11790 16592 11796 16604
rect 11848 16592 11854 16644
rect 12989 16635 13047 16641
rect 12989 16601 13001 16635
rect 13035 16632 13047 16635
rect 14829 16635 14887 16641
rect 14829 16632 14841 16635
rect 13035 16604 14841 16632
rect 13035 16601 13047 16604
rect 12989 16595 13047 16601
rect 14829 16601 14841 16604
rect 14875 16601 14887 16635
rect 14829 16595 14887 16601
rect 15933 16635 15991 16641
rect 15933 16601 15945 16635
rect 15979 16632 15991 16635
rect 18046 16632 18052 16644
rect 15979 16604 17264 16632
rect 18007 16604 18052 16632
rect 15979 16601 15991 16604
rect 15933 16595 15991 16601
rect 8662 16564 8668 16576
rect 8220 16536 8668 16564
rect 7064 16527 7128 16533
rect 7064 16524 7070 16527
rect 8662 16524 8668 16536
rect 8720 16564 8726 16576
rect 9002 16567 9060 16573
rect 9002 16564 9014 16567
rect 8720 16536 9014 16564
rect 8720 16524 8726 16536
rect 9002 16533 9014 16536
rect 9048 16533 9060 16567
rect 12526 16564 12532 16576
rect 9002 16527 9060 16533
rect 9140 16536 12532 16564
rect 3513 16499 3571 16505
rect 3513 16465 3525 16499
rect 3559 16496 3571 16499
rect 4062 16496 4068 16508
rect 3559 16468 4068 16496
rect 3559 16465 3571 16468
rect 3513 16459 3571 16465
rect 4062 16456 4068 16468
rect 4120 16456 4126 16508
rect 4246 16456 4252 16508
rect 4304 16496 4310 16508
rect 4709 16499 4767 16505
rect 4709 16496 4721 16499
rect 4304 16468 4721 16496
rect 4304 16456 4310 16468
rect 4709 16465 4721 16468
rect 4755 16465 4767 16499
rect 4709 16459 4767 16465
rect 4985 16499 5043 16505
rect 4985 16465 4997 16499
rect 5031 16496 5043 16499
rect 9140 16496 9168 16536
rect 12526 16524 12532 16536
rect 12584 16524 12590 16576
rect 12713 16567 12771 16573
rect 12713 16533 12725 16567
rect 12759 16564 12771 16567
rect 13449 16567 13507 16573
rect 13449 16564 13461 16567
rect 12759 16536 13461 16564
rect 12759 16533 12771 16536
rect 12713 16527 12771 16533
rect 13449 16533 13461 16536
rect 13495 16533 13507 16567
rect 13449 16527 13507 16533
rect 5031 16468 9168 16496
rect 5031 16465 5043 16468
rect 4985 16459 5043 16465
rect 11146 16456 11152 16508
rect 11204 16496 11210 16508
rect 12728 16496 12756 16527
rect 15746 16524 15752 16576
rect 15804 16564 15810 16576
rect 16393 16567 16451 16573
rect 16393 16564 16405 16567
rect 15804 16536 16405 16564
rect 15804 16524 15810 16536
rect 16393 16533 16405 16536
rect 16439 16533 16451 16567
rect 16393 16527 16451 16533
rect 16850 16524 16856 16576
rect 16908 16564 16914 16576
rect 16945 16567 17003 16573
rect 16945 16564 16957 16567
rect 16908 16536 16957 16564
rect 16908 16524 16914 16536
rect 16945 16533 16957 16536
rect 16991 16533 17003 16567
rect 16945 16527 17003 16533
rect 11204 16468 12756 16496
rect 13357 16499 13415 16505
rect 11204 16456 11210 16468
rect 13357 16465 13369 16499
rect 13403 16496 13415 16499
rect 13998 16496 14004 16508
rect 13403 16468 14004 16496
rect 13403 16465 13415 16468
rect 13357 16459 13415 16465
rect 13998 16456 14004 16468
rect 14056 16456 14062 16508
rect 14366 16456 14372 16508
rect 14424 16456 14430 16508
rect 14737 16499 14795 16505
rect 14737 16465 14749 16499
rect 14783 16496 14795 16499
rect 15381 16499 15439 16505
rect 15381 16496 15393 16499
rect 14783 16468 15393 16496
rect 14783 16465 14795 16468
rect 14737 16459 14795 16465
rect 15381 16465 15393 16468
rect 15427 16465 15439 16499
rect 15381 16459 15439 16465
rect 16301 16499 16359 16505
rect 16301 16465 16313 16499
rect 16347 16496 16359 16499
rect 16482 16496 16488 16508
rect 16347 16468 16488 16496
rect 16347 16465 16359 16468
rect 16301 16459 16359 16465
rect 16482 16456 16488 16468
rect 16540 16496 16546 16508
rect 16868 16496 16896 16524
rect 16540 16468 16896 16496
rect 17236 16496 17264 16604
rect 18046 16592 18052 16604
rect 18104 16592 18110 16644
rect 18417 16567 18475 16573
rect 18417 16533 18429 16567
rect 18463 16564 18475 16567
rect 18598 16564 18604 16576
rect 18463 16536 18604 16564
rect 18463 16533 18475 16536
rect 18417 16527 18475 16533
rect 18598 16524 18604 16536
rect 18656 16524 18662 16576
rect 19981 16567 20039 16573
rect 19981 16533 19993 16567
rect 20027 16564 20039 16567
rect 20898 16564 20904 16576
rect 20027 16536 20904 16564
rect 20027 16533 20039 16536
rect 19981 16527 20039 16533
rect 20898 16524 20904 16536
rect 20956 16524 20962 16576
rect 18509 16499 18567 16505
rect 18509 16496 18521 16499
rect 17236 16468 18521 16496
rect 16540 16456 16546 16468
rect 18509 16465 18521 16468
rect 18555 16465 18567 16499
rect 19702 16496 19708 16508
rect 19663 16468 19708 16496
rect 18509 16459 18567 16465
rect 19702 16456 19708 16468
rect 19760 16456 19766 16508
rect 20438 16496 20444 16508
rect 20399 16468 20444 16496
rect 20438 16456 20444 16468
rect 20496 16456 20502 16508
rect 20714 16496 20720 16508
rect 20675 16468 20720 16496
rect 20714 16456 20720 16468
rect 20772 16456 20778 16508
rect 3694 16428 3700 16440
rect 3655 16400 3700 16428
rect 3694 16388 3700 16400
rect 3752 16388 3758 16440
rect 4890 16388 4896 16440
rect 4948 16428 4954 16440
rect 6822 16428 6828 16440
rect 4948 16400 6828 16428
rect 4948 16388 4954 16400
rect 6822 16388 6828 16400
rect 6880 16388 6886 16440
rect 8757 16431 8815 16437
rect 8757 16428 8769 16431
rect 7852 16400 8769 16428
rect 3142 16292 3148 16304
rect 3103 16264 3148 16292
rect 3142 16252 3148 16264
rect 3200 16252 3206 16304
rect 6822 16252 6828 16304
rect 6880 16292 6886 16304
rect 7852 16292 7880 16400
rect 8757 16397 8769 16400
rect 8803 16397 8815 16431
rect 8757 16391 8815 16397
rect 11057 16431 11115 16437
rect 11057 16397 11069 16431
rect 11103 16397 11115 16431
rect 11057 16391 11115 16397
rect 6880 16264 7880 16292
rect 8772 16292 8800 16391
rect 11072 16360 11100 16391
rect 13262 16388 13268 16440
rect 13320 16428 13326 16440
rect 13541 16431 13599 16437
rect 13541 16428 13553 16431
rect 13320 16400 13553 16428
rect 13320 16388 13326 16400
rect 13541 16397 13553 16400
rect 13587 16397 13599 16431
rect 13541 16391 13599 16397
rect 14384 16369 14412 16456
rect 14918 16428 14924 16440
rect 14879 16400 14924 16428
rect 14918 16388 14924 16400
rect 14976 16388 14982 16440
rect 16577 16431 16635 16437
rect 16577 16397 16589 16431
rect 16623 16428 16635 16431
rect 16666 16428 16672 16440
rect 16623 16400 16672 16428
rect 16623 16397 16635 16400
rect 16577 16391 16635 16397
rect 16666 16388 16672 16400
rect 16724 16388 16730 16440
rect 18690 16428 18696 16440
rect 18651 16400 18696 16428
rect 18690 16388 18696 16400
rect 18748 16388 18754 16440
rect 10336 16332 11100 16360
rect 14369 16363 14427 16369
rect 10336 16304 10364 16332
rect 14369 16329 14381 16363
rect 14415 16329 14427 16363
rect 14369 16323 14427 16329
rect 9674 16292 9680 16304
rect 8772 16264 9680 16292
rect 6880 16252 6886 16264
rect 9674 16252 9680 16264
rect 9732 16252 9738 16304
rect 10137 16295 10195 16301
rect 10137 16261 10149 16295
rect 10183 16292 10195 16295
rect 10318 16292 10324 16304
rect 10183 16264 10324 16292
rect 10183 16261 10195 16264
rect 10137 16255 10195 16261
rect 10318 16252 10324 16264
rect 10376 16252 10382 16304
rect 1104 16202 21896 16224
rect 1104 16150 4447 16202
rect 4499 16150 4511 16202
rect 4563 16150 4575 16202
rect 4627 16150 4639 16202
rect 4691 16150 11378 16202
rect 11430 16150 11442 16202
rect 11494 16150 11506 16202
rect 11558 16150 11570 16202
rect 11622 16150 18308 16202
rect 18360 16150 18372 16202
rect 18424 16150 18436 16202
rect 18488 16150 18500 16202
rect 18552 16150 21896 16202
rect 1104 16128 21896 16150
rect 2777 16091 2835 16097
rect 2777 16057 2789 16091
rect 2823 16088 2835 16091
rect 3510 16088 3516 16100
rect 2823 16060 3516 16088
rect 2823 16057 2835 16060
rect 2777 16051 2835 16057
rect 3510 16048 3516 16060
rect 3568 16048 3574 16100
rect 6546 16088 6552 16100
rect 6507 16060 6552 16088
rect 6546 16048 6552 16060
rect 6604 16048 6610 16100
rect 6822 16048 6828 16100
rect 6880 16088 6886 16100
rect 7653 16091 7711 16097
rect 7653 16088 7665 16091
rect 6880 16060 7665 16088
rect 6880 16048 6886 16060
rect 7653 16057 7665 16060
rect 7699 16057 7711 16091
rect 13262 16088 13268 16100
rect 13223 16060 13268 16088
rect 7653 16051 7711 16057
rect 13262 16048 13268 16060
rect 13320 16048 13326 16100
rect 14918 16088 14924 16100
rect 14879 16060 14924 16088
rect 14918 16048 14924 16060
rect 14976 16048 14982 16100
rect 16666 16088 16672 16100
rect 16627 16060 16672 16088
rect 16666 16048 16672 16060
rect 16724 16048 16730 16100
rect 18325 16091 18383 16097
rect 18325 16057 18337 16091
rect 18371 16088 18383 16091
rect 18690 16088 18696 16100
rect 18371 16060 18696 16088
rect 18371 16057 18383 16060
rect 18325 16051 18383 16057
rect 18690 16048 18696 16060
rect 18748 16048 18754 16100
rect 21082 16088 21088 16100
rect 21043 16060 21088 16088
rect 21082 16048 21088 16060
rect 21140 16048 21146 16100
rect 3142 15912 3148 15964
rect 3200 15952 3206 15964
rect 3237 15955 3295 15961
rect 3237 15952 3249 15955
rect 3200 15924 3249 15952
rect 3200 15912 3206 15924
rect 3237 15921 3249 15924
rect 3283 15921 3295 15955
rect 3237 15915 3295 15921
rect 3326 15912 3332 15964
rect 3384 15952 3390 15964
rect 3384 15924 3429 15952
rect 3384 15912 3390 15924
rect 4890 15912 4896 15964
rect 4948 15952 4954 15964
rect 5169 15955 5227 15961
rect 5169 15952 5181 15955
rect 4948 15924 5181 15952
rect 4948 15912 4954 15924
rect 5169 15921 5181 15924
rect 5215 15921 5227 15955
rect 5169 15915 5227 15921
rect 7466 15912 7472 15964
rect 7524 15912 7530 15964
rect 8938 15952 8944 15964
rect 8899 15924 8944 15952
rect 8938 15912 8944 15924
rect 8996 15912 9002 15964
rect 9674 15912 9680 15964
rect 9732 15952 9738 15964
rect 10229 15955 10287 15961
rect 10229 15952 10241 15955
rect 9732 15924 10241 15952
rect 9732 15912 9738 15924
rect 10229 15921 10241 15924
rect 10275 15921 10287 15955
rect 13280 15952 13308 16048
rect 14936 15952 14964 16048
rect 16684 15952 16712 16048
rect 18598 15952 18604 15964
rect 13280 15924 13676 15952
rect 14936 15924 15424 15952
rect 16684 15924 17080 15952
rect 18559 15924 18604 15952
rect 10229 15915 10287 15921
rect 4062 15844 4068 15896
rect 4120 15884 4126 15896
rect 4249 15887 4307 15893
rect 4249 15884 4261 15887
rect 4120 15856 4261 15884
rect 4120 15844 4126 15856
rect 4249 15853 4261 15856
rect 4295 15884 4307 15887
rect 7484 15884 7512 15912
rect 4295 15856 7512 15884
rect 7837 15887 7895 15893
rect 4295 15853 4307 15856
rect 4249 15847 4307 15853
rect 7837 15853 7849 15887
rect 7883 15884 7895 15887
rect 8202 15884 8208 15896
rect 7883 15856 8208 15884
rect 7883 15853 7895 15856
rect 7837 15847 7895 15853
rect 8202 15844 8208 15856
rect 8260 15844 8266 15896
rect 8386 15844 8392 15896
rect 8444 15884 8450 15896
rect 8665 15887 8723 15893
rect 8665 15884 8677 15887
rect 8444 15856 8677 15884
rect 8444 15844 8450 15856
rect 8665 15853 8677 15856
rect 8711 15853 8723 15887
rect 8665 15847 8723 15853
rect 10318 15844 10324 15896
rect 10376 15884 10382 15896
rect 10485 15887 10543 15893
rect 10485 15884 10497 15887
rect 10376 15856 10497 15884
rect 10376 15844 10382 15856
rect 10485 15853 10497 15856
rect 10531 15853 10543 15887
rect 10485 15847 10543 15853
rect 11885 15887 11943 15893
rect 11885 15853 11897 15887
rect 11931 15884 11943 15887
rect 13538 15884 13544 15896
rect 11931 15856 13544 15884
rect 11931 15853 11943 15856
rect 11885 15847 11943 15853
rect 13538 15844 13544 15856
rect 13596 15844 13602 15896
rect 13648 15884 13676 15924
rect 13797 15887 13855 15893
rect 13797 15884 13809 15887
rect 13648 15856 13809 15884
rect 13797 15853 13809 15856
rect 13843 15853 13855 15887
rect 13797 15847 13855 15853
rect 15289 15887 15347 15893
rect 15289 15853 15301 15887
rect 15335 15853 15347 15887
rect 15396 15884 15424 15924
rect 15545 15887 15603 15893
rect 15545 15884 15557 15887
rect 15396 15856 15557 15884
rect 15289 15847 15347 15853
rect 15545 15853 15557 15856
rect 15591 15853 15603 15887
rect 15545 15847 15603 15853
rect 16945 15887 17003 15893
rect 16945 15853 16957 15887
rect 16991 15853 17003 15887
rect 17052 15884 17080 15924
rect 18598 15912 18604 15924
rect 18656 15912 18662 15964
rect 17201 15887 17259 15893
rect 17201 15884 17213 15887
rect 17052 15856 17213 15884
rect 16945 15847 17003 15853
rect 17201 15853 17213 15856
rect 17247 15853 17259 15887
rect 20898 15884 20904 15896
rect 20859 15856 20904 15884
rect 17201 15847 17259 15853
rect 3145 15819 3203 15825
rect 3145 15785 3157 15819
rect 3191 15816 3203 15819
rect 3418 15816 3424 15828
rect 3191 15788 3424 15816
rect 3191 15785 3203 15788
rect 3145 15779 3203 15785
rect 3418 15776 3424 15788
rect 3476 15776 3482 15828
rect 5436 15819 5494 15825
rect 5436 15785 5448 15819
rect 5482 15816 5494 15819
rect 7742 15816 7748 15828
rect 5482 15788 7748 15816
rect 5482 15785 5494 15788
rect 5436 15779 5494 15785
rect 7742 15776 7748 15788
rect 7800 15776 7806 15828
rect 12158 15825 12164 15828
rect 12152 15816 12164 15825
rect 11624 15788 12164 15816
rect 11624 15757 11652 15788
rect 12152 15779 12164 15788
rect 12158 15776 12164 15779
rect 12216 15776 12222 15828
rect 13556 15816 13584 15844
rect 14734 15816 14740 15828
rect 13556 15788 14740 15816
rect 14734 15776 14740 15788
rect 14792 15816 14798 15828
rect 15304 15816 15332 15847
rect 16960 15816 16988 15847
rect 20898 15844 20904 15856
rect 20956 15844 20962 15896
rect 17310 15816 17316 15828
rect 14792 15788 17316 15816
rect 14792 15776 14798 15788
rect 17310 15776 17316 15788
rect 17368 15776 17374 15828
rect 11609 15751 11667 15757
rect 11609 15717 11621 15751
rect 11655 15717 11667 15751
rect 11609 15711 11667 15717
rect 1104 15658 21896 15680
rect 1104 15606 7912 15658
rect 7964 15606 7976 15658
rect 8028 15606 8040 15658
rect 8092 15606 8104 15658
rect 8156 15606 14843 15658
rect 14895 15606 14907 15658
rect 14959 15606 14971 15658
rect 15023 15606 15035 15658
rect 15087 15606 21896 15658
rect 1104 15584 21896 15606
rect 3145 15547 3203 15553
rect 3145 15513 3157 15547
rect 3191 15544 3203 15547
rect 3694 15544 3700 15556
rect 3191 15516 3700 15544
rect 3191 15513 3203 15516
rect 3145 15507 3203 15513
rect 3694 15504 3700 15516
rect 3752 15504 3758 15556
rect 7193 15547 7251 15553
rect 7193 15513 7205 15547
rect 7239 15544 7251 15547
rect 20806 15544 20812 15556
rect 7239 15516 19840 15544
rect 7239 15513 7251 15516
rect 7193 15507 7251 15513
rect 7650 15436 7656 15488
rect 7708 15476 7714 15488
rect 8297 15479 8355 15485
rect 8297 15476 8309 15479
rect 7708 15448 8309 15476
rect 7708 15436 7714 15448
rect 8297 15445 8309 15448
rect 8343 15445 8355 15479
rect 8297 15439 8355 15445
rect 18316 15479 18374 15485
rect 18316 15445 18328 15479
rect 18362 15476 18374 15479
rect 18690 15476 18696 15488
rect 18362 15448 18696 15476
rect 18362 15445 18374 15448
rect 18316 15439 18374 15445
rect 18690 15436 18696 15448
rect 18748 15436 18754 15488
rect 1762 15408 1768 15420
rect 1723 15380 1768 15408
rect 1762 15368 1768 15380
rect 1820 15368 1826 15420
rect 2032 15411 2090 15417
rect 2032 15377 2044 15411
rect 2078 15408 2090 15411
rect 4338 15408 4344 15420
rect 2078 15380 4344 15408
rect 2078 15377 2090 15380
rect 2032 15371 2090 15377
rect 4338 15368 4344 15380
rect 4396 15368 4402 15420
rect 7561 15411 7619 15417
rect 7561 15377 7573 15411
rect 7607 15408 7619 15411
rect 8110 15408 8116 15420
rect 7607 15380 8116 15408
rect 7607 15377 7619 15380
rect 7561 15371 7619 15377
rect 8110 15368 8116 15380
rect 8168 15368 8174 15420
rect 17310 15368 17316 15420
rect 17368 15408 17374 15420
rect 19812 15417 19840 15516
rect 20088 15516 20812 15544
rect 20088 15485 20116 15516
rect 20806 15504 20812 15516
rect 20864 15504 20870 15556
rect 20073 15479 20131 15485
rect 20073 15445 20085 15479
rect 20119 15445 20131 15479
rect 20073 15439 20131 15445
rect 18049 15411 18107 15417
rect 18049 15408 18061 15411
rect 17368 15380 18061 15408
rect 17368 15368 17374 15380
rect 18049 15377 18061 15380
rect 18095 15377 18107 15411
rect 18049 15371 18107 15377
rect 19797 15411 19855 15417
rect 19797 15377 19809 15411
rect 19843 15377 19855 15411
rect 20806 15408 20812 15420
rect 20767 15380 20812 15408
rect 19797 15371 19855 15377
rect 20806 15368 20812 15380
rect 20864 15368 20870 15420
rect 7650 15340 7656 15352
rect 7611 15312 7656 15340
rect 7650 15300 7656 15312
rect 7708 15300 7714 15352
rect 7742 15300 7748 15352
rect 7800 15340 7806 15352
rect 7800 15312 7845 15340
rect 7800 15300 7806 15312
rect 19426 15204 19432 15216
rect 19387 15176 19432 15204
rect 19426 15164 19432 15176
rect 19484 15164 19490 15216
rect 20990 15204 20996 15216
rect 20951 15176 20996 15204
rect 20990 15164 20996 15176
rect 21048 15164 21054 15216
rect 1104 15114 21896 15136
rect 1104 15062 4447 15114
rect 4499 15062 4511 15114
rect 4563 15062 4575 15114
rect 4627 15062 4639 15114
rect 4691 15062 11378 15114
rect 11430 15062 11442 15114
rect 11494 15062 11506 15114
rect 11558 15062 11570 15114
rect 11622 15062 18308 15114
rect 18360 15062 18372 15114
rect 18424 15062 18436 15114
rect 18488 15062 18500 15114
rect 18552 15062 21896 15114
rect 1104 15040 21896 15062
rect 7101 15003 7159 15009
rect 7101 14969 7113 15003
rect 7147 15000 7159 15003
rect 7650 15000 7656 15012
rect 7147 14972 7656 15000
rect 7147 14969 7159 14972
rect 7101 14963 7159 14969
rect 7650 14960 7656 14972
rect 7708 14960 7714 15012
rect 4157 14935 4215 14941
rect 4157 14901 4169 14935
rect 4203 14932 4215 14935
rect 4203 14904 8892 14932
rect 4203 14901 4215 14904
rect 4157 14895 4215 14901
rect 4338 14824 4344 14876
rect 4396 14864 4402 14876
rect 4709 14867 4767 14873
rect 4709 14864 4721 14867
rect 4396 14836 4721 14864
rect 4396 14824 4402 14836
rect 4709 14833 4721 14836
rect 4755 14833 4767 14867
rect 7650 14864 7656 14876
rect 7611 14836 7656 14864
rect 4709 14827 4767 14833
rect 7650 14824 7656 14836
rect 7708 14824 7714 14876
rect 8110 14864 8116 14876
rect 8071 14836 8116 14864
rect 8110 14824 8116 14836
rect 8168 14824 8174 14876
rect 3878 14756 3884 14808
rect 3936 14796 3942 14808
rect 7374 14796 7380 14808
rect 3936 14768 7380 14796
rect 3936 14756 3942 14768
rect 7374 14756 7380 14768
rect 7432 14756 7438 14808
rect 7558 14796 7564 14808
rect 7519 14768 7564 14796
rect 7558 14756 7564 14768
rect 7616 14756 7622 14808
rect 8757 14799 8815 14805
rect 8757 14765 8769 14799
rect 8803 14765 8815 14799
rect 8864 14796 8892 14904
rect 10134 14824 10140 14876
rect 10192 14864 10198 14876
rect 20806 14864 20812 14876
rect 10192 14836 20812 14864
rect 10192 14824 10198 14836
rect 20806 14824 20812 14836
rect 20864 14824 20870 14876
rect 19889 14799 19947 14805
rect 19889 14796 19901 14799
rect 8864 14768 19901 14796
rect 8757 14759 8815 14765
rect 19889 14765 19901 14768
rect 19935 14765 19947 14799
rect 20901 14799 20959 14805
rect 20901 14796 20913 14799
rect 19889 14759 19947 14765
rect 19996 14768 20913 14796
rect 4525 14731 4583 14737
rect 4525 14697 4537 14731
rect 4571 14728 4583 14731
rect 5169 14731 5227 14737
rect 5169 14728 5181 14731
rect 4571 14700 5181 14728
rect 4571 14697 4583 14700
rect 4525 14691 4583 14697
rect 5169 14697 5181 14700
rect 5215 14697 5227 14731
rect 5169 14691 5227 14697
rect 7469 14731 7527 14737
rect 7469 14697 7481 14731
rect 7515 14728 7527 14731
rect 8386 14728 8392 14740
rect 7515 14700 8392 14728
rect 7515 14697 7527 14700
rect 7469 14691 7527 14697
rect 8386 14688 8392 14700
rect 8444 14688 8450 14740
rect 8772 14728 8800 14759
rect 10962 14728 10968 14740
rect 8772 14700 10968 14728
rect 10962 14688 10968 14700
rect 11020 14688 11026 14740
rect 16574 14688 16580 14740
rect 16632 14728 16638 14740
rect 19996 14728 20024 14768
rect 20901 14765 20913 14768
rect 20947 14765 20959 14799
rect 20901 14759 20959 14765
rect 16632 14700 20024 14728
rect 20165 14731 20223 14737
rect 16632 14688 16638 14700
rect 20165 14697 20177 14731
rect 20211 14728 20223 14731
rect 20806 14728 20812 14740
rect 20211 14700 20812 14728
rect 20211 14697 20223 14700
rect 20165 14691 20223 14697
rect 20806 14688 20812 14700
rect 20864 14688 20870 14740
rect 4617 14663 4675 14669
rect 4617 14629 4629 14663
rect 4663 14660 4675 14663
rect 4706 14660 4712 14672
rect 4663 14632 4712 14660
rect 4663 14629 4675 14632
rect 4617 14623 4675 14629
rect 4706 14620 4712 14632
rect 4764 14620 4770 14672
rect 8202 14620 8208 14672
rect 8260 14660 8266 14672
rect 8573 14663 8631 14669
rect 8573 14660 8585 14663
rect 8260 14632 8585 14660
rect 8260 14620 8266 14632
rect 8573 14629 8585 14632
rect 8619 14629 8631 14663
rect 8573 14623 8631 14629
rect 12802 14620 12808 14672
rect 12860 14660 12866 14672
rect 13357 14663 13415 14669
rect 13357 14660 13369 14663
rect 12860 14632 13369 14660
rect 12860 14620 12866 14632
rect 13357 14629 13369 14632
rect 13403 14660 13415 14663
rect 14550 14660 14556 14672
rect 13403 14632 14556 14660
rect 13403 14629 13415 14632
rect 13357 14623 13415 14629
rect 14550 14620 14556 14632
rect 14608 14620 14614 14672
rect 21082 14660 21088 14672
rect 21043 14632 21088 14660
rect 21082 14620 21088 14632
rect 21140 14620 21146 14672
rect 1104 14570 21896 14592
rect 1104 14518 7912 14570
rect 7964 14518 7976 14570
rect 8028 14518 8040 14570
rect 8092 14518 8104 14570
rect 8156 14518 14843 14570
rect 14895 14518 14907 14570
rect 14959 14518 14971 14570
rect 15023 14518 15035 14570
rect 15087 14518 21896 14570
rect 1104 14496 21896 14518
rect 4338 14416 4344 14468
rect 4396 14456 4402 14468
rect 4433 14459 4491 14465
rect 4433 14456 4445 14459
rect 4396 14428 4445 14456
rect 4396 14416 4402 14428
rect 4433 14425 4445 14428
rect 4479 14425 4491 14459
rect 4706 14456 4712 14468
rect 4667 14428 4712 14456
rect 4433 14419 4491 14425
rect 4706 14416 4712 14428
rect 4764 14416 4770 14468
rect 5077 14459 5135 14465
rect 5077 14425 5089 14459
rect 5123 14456 5135 14459
rect 5123 14428 5856 14456
rect 5123 14425 5135 14428
rect 5077 14419 5135 14425
rect 3320 14391 3378 14397
rect 3320 14357 3332 14391
rect 3366 14388 3378 14391
rect 3366 14360 5212 14388
rect 3366 14357 3378 14360
rect 3320 14351 3378 14357
rect 5184 14320 5212 14360
rect 5828 14329 5856 14428
rect 7374 14416 7380 14468
rect 7432 14456 7438 14468
rect 11977 14459 12035 14465
rect 11977 14456 11989 14459
rect 7432 14428 7788 14456
rect 7432 14416 7438 14428
rect 7092 14391 7150 14397
rect 7092 14357 7104 14391
rect 7138 14388 7150 14391
rect 7190 14388 7196 14400
rect 7138 14360 7196 14388
rect 7138 14357 7150 14360
rect 7092 14351 7150 14357
rect 7190 14348 7196 14360
rect 7248 14388 7254 14400
rect 7650 14388 7656 14400
rect 7248 14360 7656 14388
rect 7248 14348 7254 14360
rect 7650 14348 7656 14360
rect 7708 14348 7714 14400
rect 7760 14388 7788 14428
rect 8312 14428 11989 14456
rect 8312 14388 8340 14428
rect 11977 14425 11989 14428
rect 12023 14456 12035 14459
rect 12897 14459 12955 14465
rect 12897 14456 12909 14459
rect 12023 14428 12909 14456
rect 12023 14425 12035 14428
rect 11977 14419 12035 14425
rect 12897 14425 12909 14428
rect 12943 14425 12955 14459
rect 12897 14419 12955 14425
rect 15562 14416 15568 14468
rect 15620 14456 15626 14468
rect 17589 14459 17647 14465
rect 17589 14456 17601 14459
rect 15620 14428 17601 14456
rect 15620 14416 15626 14428
rect 17589 14425 17601 14428
rect 17635 14456 17647 14459
rect 18509 14459 18567 14465
rect 18509 14456 18521 14459
rect 17635 14428 18521 14456
rect 17635 14425 17647 14428
rect 17589 14419 17647 14425
rect 18509 14425 18521 14428
rect 18555 14425 18567 14459
rect 18509 14419 18567 14425
rect 20993 14459 21051 14465
rect 20993 14425 21005 14459
rect 21039 14456 21051 14459
rect 21174 14456 21180 14468
rect 21039 14428 21180 14456
rect 21039 14425 21051 14428
rect 20993 14419 21051 14425
rect 21174 14416 21180 14428
rect 21232 14416 21238 14468
rect 7760 14360 8340 14388
rect 8386 14348 8392 14400
rect 8444 14388 8450 14400
rect 8573 14391 8631 14397
rect 8573 14388 8585 14391
rect 8444 14360 8585 14388
rect 8444 14348 8450 14360
rect 8573 14357 8585 14360
rect 8619 14388 8631 14391
rect 10134 14388 10140 14400
rect 8619 14360 9996 14388
rect 10095 14360 10140 14388
rect 8619 14357 8631 14360
rect 8573 14351 8631 14357
rect 5813 14323 5871 14329
rect 5184 14292 5304 14320
rect 5276 14264 5304 14292
rect 5813 14289 5825 14323
rect 5859 14320 5871 14323
rect 8404 14320 8432 14348
rect 5859 14292 8432 14320
rect 9217 14323 9275 14329
rect 5859 14289 5871 14292
rect 5813 14283 5871 14289
rect 9217 14289 9229 14323
rect 9263 14320 9275 14323
rect 9674 14320 9680 14332
rect 9263 14292 9680 14320
rect 9263 14289 9275 14292
rect 9217 14283 9275 14289
rect 9674 14280 9680 14292
rect 9732 14280 9738 14332
rect 9861 14323 9919 14329
rect 9861 14320 9873 14323
rect 9784 14292 9873 14320
rect 3050 14252 3056 14264
rect 3011 14224 3056 14252
rect 3050 14212 3056 14224
rect 3108 14212 3114 14264
rect 4154 14212 4160 14264
rect 4212 14252 4218 14264
rect 5169 14255 5227 14261
rect 5169 14252 5181 14255
rect 4212 14224 5181 14252
rect 4212 14212 4218 14224
rect 5169 14221 5181 14224
rect 5215 14221 5227 14255
rect 5169 14215 5227 14221
rect 5258 14212 5264 14264
rect 5316 14252 5322 14264
rect 6822 14252 6828 14264
rect 5316 14224 5409 14252
rect 6783 14224 6828 14252
rect 5316 14212 5322 14224
rect 6822 14212 6828 14224
rect 6880 14212 6886 14264
rect 8386 14212 8392 14264
rect 8444 14252 8450 14264
rect 9309 14255 9367 14261
rect 9309 14252 9321 14255
rect 8444 14224 9321 14252
rect 8444 14212 8450 14224
rect 9309 14221 9321 14224
rect 9355 14221 9367 14255
rect 9490 14252 9496 14264
rect 9451 14224 9496 14252
rect 9309 14215 9367 14221
rect 9490 14212 9496 14224
rect 9548 14212 9554 14264
rect 7834 14144 7840 14196
rect 7892 14184 7898 14196
rect 8205 14187 8263 14193
rect 8205 14184 8217 14187
rect 7892 14156 8217 14184
rect 7892 14144 7898 14156
rect 8205 14153 8217 14156
rect 8251 14153 8263 14187
rect 8205 14147 8263 14153
rect 8849 14187 8907 14193
rect 8849 14153 8861 14187
rect 8895 14184 8907 14187
rect 9784 14184 9812 14292
rect 9861 14289 9873 14292
rect 9907 14289 9919 14323
rect 9968 14320 9996 14360
rect 10134 14348 10140 14360
rect 10192 14348 10198 14400
rect 12802 14388 12808 14400
rect 12452 14360 12808 14388
rect 12452 14320 12480 14360
rect 12802 14348 12808 14360
rect 12860 14388 12866 14400
rect 18046 14388 18052 14400
rect 12860 14360 12905 14388
rect 13556 14360 18052 14388
rect 12860 14348 12866 14360
rect 13556 14320 13584 14360
rect 18046 14348 18052 14360
rect 18104 14348 18110 14400
rect 19061 14391 19119 14397
rect 19061 14388 19073 14391
rect 18432 14360 19073 14388
rect 13722 14320 13728 14332
rect 9968 14292 12480 14320
rect 12544 14292 13584 14320
rect 13683 14292 13728 14320
rect 9861 14283 9919 14289
rect 12544 14252 12572 14292
rect 13722 14280 13728 14292
rect 13780 14280 13786 14332
rect 14274 14329 14280 14332
rect 14268 14320 14280 14329
rect 14235 14292 14280 14320
rect 14268 14283 14280 14292
rect 14274 14280 14280 14283
rect 14332 14280 14338 14332
rect 15286 14280 15292 14332
rect 15344 14320 15350 14332
rect 16025 14323 16083 14329
rect 16025 14320 16037 14323
rect 15344 14292 16037 14320
rect 15344 14280 15350 14292
rect 16025 14289 16037 14292
rect 16071 14289 16083 14323
rect 16025 14283 16083 14289
rect 18138 14280 18144 14332
rect 18196 14320 18202 14332
rect 18432 14329 18460 14360
rect 19061 14357 19073 14360
rect 19107 14357 19119 14391
rect 19061 14351 19119 14357
rect 18417 14323 18475 14329
rect 18417 14320 18429 14323
rect 18196 14292 18429 14320
rect 18196 14280 18202 14292
rect 18417 14289 18429 14292
rect 18463 14289 18475 14323
rect 18417 14283 18475 14289
rect 18966 14280 18972 14332
rect 19024 14320 19030 14332
rect 19981 14323 20039 14329
rect 19981 14320 19993 14323
rect 19024 14292 19993 14320
rect 19024 14280 19030 14292
rect 19981 14289 19993 14292
rect 20027 14289 20039 14323
rect 20806 14320 20812 14332
rect 20767 14292 20812 14320
rect 19981 14283 20039 14289
rect 20806 14280 20812 14292
rect 20864 14280 20870 14332
rect 13078 14252 13084 14264
rect 8895 14156 9812 14184
rect 9876 14224 12572 14252
rect 13039 14224 13084 14252
rect 8895 14153 8907 14156
rect 8849 14147 8907 14153
rect 3970 14076 3976 14128
rect 4028 14116 4034 14128
rect 8018 14116 8024 14128
rect 4028 14088 8024 14116
rect 4028 14076 4034 14088
rect 8018 14076 8024 14088
rect 8076 14076 8082 14128
rect 9214 14076 9220 14128
rect 9272 14116 9278 14128
rect 9876 14116 9904 14224
rect 13078 14212 13084 14224
rect 13136 14212 13142 14264
rect 14001 14255 14059 14261
rect 14001 14221 14013 14255
rect 14047 14221 14059 14255
rect 16114 14252 16120 14264
rect 16075 14224 16120 14252
rect 14001 14215 14059 14221
rect 12437 14187 12495 14193
rect 12437 14153 12449 14187
rect 12483 14184 12495 14187
rect 13814 14184 13820 14196
rect 12483 14156 13820 14184
rect 12483 14153 12495 14156
rect 12437 14147 12495 14153
rect 13814 14144 13820 14156
rect 13872 14144 13878 14196
rect 9272 14088 9904 14116
rect 9272 14076 9278 14088
rect 12250 14076 12256 14128
rect 12308 14116 12314 14128
rect 13538 14116 13544 14128
rect 12308 14088 13544 14116
rect 12308 14076 12314 14088
rect 13538 14076 13544 14088
rect 13596 14116 13602 14128
rect 14016 14116 14044 14215
rect 16114 14212 16120 14224
rect 16172 14212 16178 14264
rect 16209 14255 16267 14261
rect 16209 14221 16221 14255
rect 16255 14221 16267 14255
rect 16209 14215 16267 14221
rect 18693 14255 18751 14261
rect 18693 14221 18705 14255
rect 18739 14252 18751 14255
rect 19426 14252 19432 14264
rect 18739 14224 19432 14252
rect 18739 14221 18751 14224
rect 18693 14215 18751 14221
rect 16224 14184 16252 14215
rect 19426 14212 19432 14224
rect 19484 14212 19490 14264
rect 20257 14255 20315 14261
rect 20257 14221 20269 14255
rect 20303 14252 20315 14255
rect 20898 14252 20904 14264
rect 20303 14224 20904 14252
rect 20303 14221 20315 14224
rect 20257 14215 20315 14221
rect 20898 14212 20904 14224
rect 20956 14212 20962 14264
rect 15396 14156 16252 14184
rect 13596 14088 14044 14116
rect 13596 14076 13602 14088
rect 15102 14076 15108 14128
rect 15160 14116 15166 14128
rect 15396 14125 15424 14156
rect 15381 14119 15439 14125
rect 15381 14116 15393 14119
rect 15160 14088 15393 14116
rect 15160 14076 15166 14088
rect 15381 14085 15393 14088
rect 15427 14085 15439 14119
rect 15381 14079 15439 14085
rect 15657 14119 15715 14125
rect 15657 14085 15669 14119
rect 15703 14116 15715 14119
rect 16298 14116 16304 14128
rect 15703 14088 16304 14116
rect 15703 14085 15715 14088
rect 15657 14079 15715 14085
rect 16298 14076 16304 14088
rect 16356 14076 16362 14128
rect 18049 14119 18107 14125
rect 18049 14085 18061 14119
rect 18095 14116 18107 14119
rect 18690 14116 18696 14128
rect 18095 14088 18696 14116
rect 18095 14085 18107 14088
rect 18049 14079 18107 14085
rect 18690 14076 18696 14088
rect 18748 14076 18754 14128
rect 19705 14119 19763 14125
rect 19705 14085 19717 14119
rect 19751 14116 19763 14119
rect 20254 14116 20260 14128
rect 19751 14088 20260 14116
rect 19751 14085 19763 14088
rect 19705 14079 19763 14085
rect 20254 14076 20260 14088
rect 20312 14076 20318 14128
rect 1104 14026 21896 14048
rect 1104 13974 4447 14026
rect 4499 13974 4511 14026
rect 4563 13974 4575 14026
rect 4627 13974 4639 14026
rect 4691 13974 11378 14026
rect 11430 13974 11442 14026
rect 11494 13974 11506 14026
rect 11558 13974 11570 14026
rect 11622 13974 18308 14026
rect 18360 13974 18372 14026
rect 18424 13974 18436 14026
rect 18488 13974 18500 14026
rect 18552 13974 21896 14026
rect 1104 13952 21896 13974
rect 4154 13872 4160 13924
rect 4212 13912 4218 13924
rect 4525 13915 4583 13921
rect 4525 13912 4537 13915
rect 4212 13884 4537 13912
rect 4212 13872 4218 13884
rect 4525 13881 4537 13884
rect 4571 13881 4583 13915
rect 6914 13912 6920 13924
rect 4525 13875 4583 13881
rect 5828 13884 6920 13912
rect 3050 13668 3056 13720
rect 3108 13708 3114 13720
rect 5828 13717 5856 13884
rect 6914 13872 6920 13884
rect 6972 13872 6978 13924
rect 7190 13912 7196 13924
rect 7151 13884 7196 13912
rect 7190 13872 7196 13884
rect 7248 13872 7254 13924
rect 8018 13912 8024 13924
rect 7979 13884 8024 13912
rect 8018 13872 8024 13884
rect 8076 13872 8082 13924
rect 8386 13912 8392 13924
rect 8347 13884 8392 13912
rect 8386 13872 8392 13884
rect 8444 13872 8450 13924
rect 15102 13912 15108 13924
rect 11256 13884 15108 13912
rect 6932 13844 6960 13872
rect 6932 13816 9996 13844
rect 8018 13736 8024 13788
rect 8076 13776 8082 13788
rect 8849 13779 8907 13785
rect 8849 13776 8861 13779
rect 8076 13748 8861 13776
rect 8076 13736 8082 13748
rect 8849 13745 8861 13748
rect 8895 13745 8907 13779
rect 9030 13776 9036 13788
rect 8943 13748 9036 13776
rect 8849 13739 8907 13745
rect 9030 13736 9036 13748
rect 9088 13776 9094 13788
rect 9968 13785 9996 13816
rect 9953 13779 10011 13785
rect 9088 13748 9720 13776
rect 9088 13736 9094 13748
rect 5813 13711 5871 13717
rect 5813 13708 5825 13711
rect 3108 13680 5825 13708
rect 3108 13668 3114 13680
rect 5813 13677 5825 13680
rect 5859 13677 5871 13711
rect 5813 13671 5871 13677
rect 6080 13711 6138 13717
rect 6080 13677 6092 13711
rect 6126 13708 6138 13711
rect 9214 13708 9220 13720
rect 6126 13680 9220 13708
rect 6126 13677 6138 13680
rect 6080 13671 6138 13677
rect 9214 13668 9220 13680
rect 9272 13668 9278 13720
rect 9692 13640 9720 13748
rect 9953 13745 9965 13779
rect 9999 13745 10011 13779
rect 9953 13739 10011 13745
rect 10220 13711 10278 13717
rect 10220 13677 10232 13711
rect 10266 13708 10278 13711
rect 11256 13708 11284 13884
rect 15102 13872 15108 13884
rect 15160 13872 15166 13924
rect 15286 13912 15292 13924
rect 15247 13884 15292 13912
rect 15286 13872 15292 13884
rect 15344 13872 15350 13924
rect 18046 13872 18052 13924
rect 18104 13912 18110 13924
rect 18693 13915 18751 13921
rect 18693 13912 18705 13915
rect 18104 13884 18705 13912
rect 18104 13872 18110 13884
rect 18693 13881 18705 13884
rect 18739 13881 18751 13915
rect 18966 13912 18972 13924
rect 18927 13884 18972 13912
rect 18693 13875 18751 13881
rect 13633 13847 13691 13853
rect 13633 13813 13645 13847
rect 13679 13813 13691 13847
rect 13633 13807 13691 13813
rect 13909 13847 13967 13853
rect 13909 13813 13921 13847
rect 13955 13844 13967 13847
rect 16114 13844 16120 13856
rect 13955 13816 16120 13844
rect 13955 13813 13967 13816
rect 13909 13807 13967 13813
rect 12250 13776 12256 13788
rect 12211 13748 12256 13776
rect 12250 13736 12256 13748
rect 12308 13736 12314 13788
rect 10266 13680 11284 13708
rect 13648 13708 13676 13807
rect 16114 13804 16120 13816
rect 16172 13804 16178 13856
rect 18708 13844 18736 13875
rect 18966 13872 18972 13884
rect 19024 13872 19030 13924
rect 20438 13912 20444 13924
rect 20399 13884 20444 13912
rect 20438 13872 20444 13884
rect 20496 13872 20502 13924
rect 20622 13872 20628 13924
rect 20680 13912 20686 13924
rect 21085 13915 21143 13921
rect 21085 13912 21097 13915
rect 20680 13884 21097 13912
rect 20680 13872 20686 13884
rect 21085 13881 21097 13884
rect 21131 13881 21143 13915
rect 21085 13875 21143 13881
rect 18708 13816 19564 13844
rect 13814 13736 13820 13788
rect 13872 13776 13878 13788
rect 14369 13779 14427 13785
rect 14369 13776 14381 13779
rect 13872 13748 14381 13776
rect 13872 13736 13878 13748
rect 14369 13745 14381 13748
rect 14415 13745 14427 13779
rect 14369 13739 14427 13745
rect 14553 13779 14611 13785
rect 14553 13745 14565 13779
rect 14599 13776 14611 13779
rect 15841 13779 15899 13785
rect 15841 13776 15853 13779
rect 14599 13748 15853 13776
rect 14599 13745 14611 13748
rect 14553 13739 14611 13745
rect 15841 13745 15853 13748
rect 15887 13745 15899 13779
rect 16574 13776 16580 13788
rect 16535 13748 16580 13776
rect 15841 13739 15899 13745
rect 14274 13708 14280 13720
rect 13648 13680 14280 13708
rect 10266 13677 10278 13680
rect 10220 13671 10278 13677
rect 14274 13668 14280 13680
rect 14332 13708 14338 13720
rect 14568 13708 14596 13739
rect 16574 13736 16580 13748
rect 16632 13736 16638 13788
rect 17310 13776 17316 13788
rect 17271 13748 17316 13776
rect 17310 13736 17316 13748
rect 17368 13736 17374 13788
rect 18690 13736 18696 13788
rect 18748 13776 18754 13788
rect 19536 13785 19564 13816
rect 19429 13779 19487 13785
rect 19429 13776 19441 13779
rect 18748 13748 19441 13776
rect 18748 13736 18754 13748
rect 19429 13745 19441 13748
rect 19475 13745 19487 13779
rect 19429 13739 19487 13745
rect 19521 13779 19579 13785
rect 19521 13745 19533 13779
rect 19567 13745 19579 13779
rect 19521 13739 19579 13745
rect 14332 13680 14596 13708
rect 14332 13668 14338 13680
rect 15470 13668 15476 13720
rect 15528 13708 15534 13720
rect 15657 13711 15715 13717
rect 15657 13708 15669 13711
rect 15528 13680 15669 13708
rect 15528 13668 15534 13680
rect 15657 13677 15669 13680
rect 15703 13677 15715 13711
rect 16298 13708 16304 13720
rect 16259 13680 16304 13708
rect 15657 13671 15715 13677
rect 16298 13668 16304 13680
rect 16356 13668 16362 13720
rect 17580 13711 17638 13717
rect 17580 13677 17592 13711
rect 17626 13708 17638 13711
rect 19334 13708 19340 13720
rect 17626 13680 19340 13708
rect 17626 13677 17638 13680
rect 17580 13671 17638 13677
rect 19334 13668 19340 13680
rect 19392 13668 19398 13720
rect 20254 13708 20260 13720
rect 20215 13680 20260 13708
rect 20254 13668 20260 13680
rect 20312 13668 20318 13720
rect 20898 13708 20904 13720
rect 20859 13680 20904 13708
rect 20898 13668 20904 13680
rect 20956 13668 20962 13720
rect 9692 13612 10640 13640
rect 10612 13584 10640 13612
rect 12434 13600 12440 13652
rect 12492 13649 12498 13652
rect 12492 13643 12556 13649
rect 12492 13609 12510 13643
rect 12544 13609 12556 13643
rect 12492 13603 12556 13609
rect 12492 13600 12498 13603
rect 12802 13600 12808 13652
rect 12860 13640 12866 13652
rect 15749 13643 15807 13649
rect 12860 13612 15700 13640
rect 12860 13600 12866 13612
rect 8754 13572 8760 13584
rect 8715 13544 8760 13572
rect 8754 13532 8760 13544
rect 8812 13532 8818 13584
rect 10594 13532 10600 13584
rect 10652 13572 10658 13584
rect 11333 13575 11391 13581
rect 11333 13572 11345 13575
rect 10652 13544 11345 13572
rect 10652 13532 10658 13544
rect 11333 13541 11345 13544
rect 11379 13541 11391 13575
rect 14274 13572 14280 13584
rect 14235 13544 14280 13572
rect 11333 13535 11391 13541
rect 14274 13532 14280 13544
rect 14332 13532 14338 13584
rect 15672 13572 15700 13612
rect 15749 13609 15761 13643
rect 15795 13640 15807 13643
rect 16482 13640 16488 13652
rect 15795 13612 16488 13640
rect 15795 13609 15807 13612
rect 15749 13603 15807 13609
rect 16482 13600 16488 13612
rect 16540 13600 16546 13652
rect 19058 13572 19064 13584
rect 15672 13544 19064 13572
rect 19058 13532 19064 13544
rect 19116 13532 19122 13584
rect 19334 13572 19340 13584
rect 19295 13544 19340 13572
rect 19334 13532 19340 13544
rect 19392 13532 19398 13584
rect 1104 13482 21896 13504
rect 1104 13430 7912 13482
rect 7964 13430 7976 13482
rect 8028 13430 8040 13482
rect 8092 13430 8104 13482
rect 8156 13430 14843 13482
rect 14895 13430 14907 13482
rect 14959 13430 14971 13482
rect 15023 13430 15035 13482
rect 15087 13430 21896 13482
rect 1104 13408 21896 13430
rect 5169 13371 5227 13377
rect 5169 13337 5181 13371
rect 5215 13368 5227 13371
rect 5258 13368 5264 13380
rect 5215 13340 5264 13368
rect 5215 13337 5227 13340
rect 5169 13331 5227 13337
rect 5258 13328 5264 13340
rect 5316 13328 5322 13380
rect 8754 13328 8760 13380
rect 8812 13368 8818 13380
rect 9401 13371 9459 13377
rect 9401 13368 9413 13371
rect 8812 13340 9413 13368
rect 8812 13328 8818 13340
rect 9401 13337 9413 13340
rect 9447 13368 9459 13371
rect 9490 13368 9496 13380
rect 9447 13340 9496 13368
rect 9447 13337 9459 13340
rect 9401 13331 9459 13337
rect 9490 13328 9496 13340
rect 9548 13328 9554 13380
rect 10962 13328 10968 13380
rect 11020 13368 11026 13380
rect 11517 13371 11575 13377
rect 11517 13368 11529 13371
rect 11020 13340 11529 13368
rect 11020 13328 11026 13340
rect 11517 13337 11529 13340
rect 11563 13337 11575 13371
rect 11517 13331 11575 13337
rect 12529 13371 12587 13377
rect 12529 13337 12541 13371
rect 12575 13368 12587 13371
rect 14274 13368 14280 13380
rect 12575 13340 14280 13368
rect 12575 13337 12587 13340
rect 12529 13331 12587 13337
rect 14274 13328 14280 13340
rect 14332 13328 14338 13380
rect 15470 13368 15476 13380
rect 15431 13340 15476 13368
rect 15470 13328 15476 13340
rect 15528 13328 15534 13380
rect 16209 13371 16267 13377
rect 16209 13337 16221 13371
rect 16255 13368 16267 13371
rect 16482 13368 16488 13380
rect 16255 13340 16488 13368
rect 16255 13337 16267 13340
rect 16209 13331 16267 13337
rect 16482 13328 16488 13340
rect 16540 13328 16546 13380
rect 18417 13371 18475 13377
rect 18417 13337 18429 13371
rect 18463 13368 18475 13371
rect 19334 13368 19340 13380
rect 18463 13340 19340 13368
rect 18463 13337 18475 13340
rect 18417 13331 18475 13337
rect 19334 13328 19340 13340
rect 19392 13328 19398 13380
rect 20530 13368 20536 13380
rect 20491 13340 20536 13368
rect 20530 13328 20536 13340
rect 20588 13328 20594 13380
rect 21085 13371 21143 13377
rect 21085 13337 21097 13371
rect 21131 13368 21143 13371
rect 21266 13368 21272 13380
rect 21131 13340 21272 13368
rect 21131 13337 21143 13340
rect 21085 13331 21143 13337
rect 21266 13328 21272 13340
rect 21324 13328 21330 13380
rect 8012 13303 8070 13309
rect 8012 13269 8024 13303
rect 8058 13300 8070 13303
rect 9030 13300 9036 13312
rect 8058 13272 9036 13300
rect 8058 13269 8070 13272
rect 8012 13263 8070 13269
rect 9030 13260 9036 13272
rect 9088 13260 9094 13312
rect 10229 13303 10287 13309
rect 10229 13269 10241 13303
rect 10275 13300 10287 13303
rect 12802 13300 12808 13312
rect 10275 13272 12808 13300
rect 10275 13269 10287 13272
rect 10229 13263 10287 13269
rect 12802 13260 12808 13272
rect 12860 13260 12866 13312
rect 12986 13300 12992 13312
rect 12947 13272 12992 13300
rect 12986 13260 12992 13272
rect 13044 13300 13050 13312
rect 13906 13300 13912 13312
rect 13044 13272 13912 13300
rect 13044 13260 13050 13272
rect 13906 13260 13912 13272
rect 13964 13260 13970 13312
rect 15286 13260 15292 13312
rect 15344 13300 15350 13312
rect 15344 13272 20392 13300
rect 15344 13260 15350 13272
rect 3050 13192 3056 13244
rect 3108 13232 3114 13244
rect 3789 13235 3847 13241
rect 3789 13232 3801 13235
rect 3108 13204 3801 13232
rect 3108 13192 3114 13204
rect 3789 13201 3801 13204
rect 3835 13201 3847 13235
rect 3789 13195 3847 13201
rect 4056 13235 4114 13241
rect 4056 13201 4068 13235
rect 4102 13232 4114 13235
rect 9398 13232 9404 13244
rect 4102 13204 9404 13232
rect 4102 13201 4114 13204
rect 4056 13195 4114 13201
rect 6914 13124 6920 13176
rect 6972 13164 6978 13176
rect 7742 13164 7748 13176
rect 6972 13136 7748 13164
rect 6972 13124 6978 13136
rect 7742 13124 7748 13136
rect 7800 13124 7806 13176
rect 9140 13105 9168 13204
rect 9398 13192 9404 13204
rect 9456 13192 9462 13244
rect 12710 13192 12716 13244
rect 12768 13232 12774 13244
rect 20364 13241 20392 13272
rect 12897 13235 12955 13241
rect 12897 13232 12909 13235
rect 12768 13204 12909 13232
rect 12768 13192 12774 13204
rect 12897 13201 12909 13204
rect 12943 13232 12955 13235
rect 18785 13235 18843 13241
rect 12943 13204 13676 13232
rect 12943 13201 12955 13204
rect 12897 13195 12955 13201
rect 12434 13124 12440 13176
rect 12492 13164 12498 13176
rect 13078 13164 13084 13176
rect 12492 13136 13084 13164
rect 12492 13124 12498 13136
rect 13078 13124 13084 13136
rect 13136 13124 13142 13176
rect 9125 13099 9183 13105
rect 9125 13065 9137 13099
rect 9171 13065 9183 13099
rect 9125 13059 9183 13065
rect 13648 13037 13676 13204
rect 18785 13201 18797 13235
rect 18831 13232 18843 13235
rect 19429 13235 19487 13241
rect 19429 13232 19441 13235
rect 18831 13204 19441 13232
rect 18831 13201 18843 13204
rect 18785 13195 18843 13201
rect 19429 13201 19441 13204
rect 19475 13201 19487 13235
rect 19429 13195 19487 13201
rect 20349 13235 20407 13241
rect 20349 13201 20361 13235
rect 20395 13201 20407 13235
rect 20349 13195 20407 13201
rect 20901 13235 20959 13241
rect 20901 13201 20913 13235
rect 20947 13201 20959 13235
rect 20901 13195 20959 13201
rect 18874 13164 18880 13176
rect 18835 13136 18880 13164
rect 18874 13124 18880 13136
rect 18932 13124 18938 13176
rect 19061 13167 19119 13173
rect 19061 13133 19073 13167
rect 19107 13164 19119 13167
rect 19334 13164 19340 13176
rect 19107 13136 19340 13164
rect 19107 13133 19119 13136
rect 19061 13127 19119 13133
rect 19334 13124 19340 13136
rect 19392 13124 19398 13176
rect 20073 13167 20131 13173
rect 20073 13133 20085 13167
rect 20119 13164 20131 13167
rect 20622 13164 20628 13176
rect 20119 13136 20628 13164
rect 20119 13133 20131 13136
rect 20073 13127 20131 13133
rect 20622 13124 20628 13136
rect 20680 13164 20686 13176
rect 20916 13164 20944 13195
rect 20680 13136 20944 13164
rect 20680 13124 20686 13136
rect 13633 13031 13691 13037
rect 13633 12997 13645 13031
rect 13679 13028 13691 13031
rect 13814 13028 13820 13040
rect 13679 13000 13820 13028
rect 13679 12997 13691 13000
rect 13633 12991 13691 12997
rect 13814 12988 13820 13000
rect 13872 12988 13878 13040
rect 1104 12938 21896 12960
rect 1104 12886 4447 12938
rect 4499 12886 4511 12938
rect 4563 12886 4575 12938
rect 4627 12886 4639 12938
rect 4691 12886 11378 12938
rect 11430 12886 11442 12938
rect 11494 12886 11506 12938
rect 11558 12886 11570 12938
rect 11622 12886 18308 12938
rect 18360 12886 18372 12938
rect 18424 12886 18436 12938
rect 18488 12886 18500 12938
rect 18552 12886 21896 12938
rect 1104 12864 21896 12886
rect 7742 12824 7748 12836
rect 7703 12796 7748 12824
rect 7742 12784 7748 12796
rect 7800 12784 7806 12836
rect 9674 12784 9680 12836
rect 9732 12824 9738 12836
rect 9953 12827 10011 12833
rect 9953 12824 9965 12827
rect 9732 12796 9965 12824
rect 9732 12784 9738 12796
rect 9953 12793 9965 12796
rect 9999 12793 10011 12827
rect 9953 12787 10011 12793
rect 10962 12784 10968 12836
rect 11020 12824 11026 12836
rect 12345 12827 12403 12833
rect 11020 12796 12020 12824
rect 11020 12784 11026 12796
rect 10594 12688 10600 12700
rect 10555 12660 10600 12688
rect 10594 12648 10600 12660
rect 10652 12648 10658 12700
rect 10796 12660 11100 12688
rect 7929 12623 7987 12629
rect 7929 12589 7941 12623
rect 7975 12620 7987 12623
rect 8202 12620 8208 12632
rect 7975 12592 8208 12620
rect 7975 12589 7987 12592
rect 7929 12583 7987 12589
rect 8202 12580 8208 12592
rect 8260 12580 8266 12632
rect 10321 12623 10379 12629
rect 10321 12589 10333 12623
rect 10367 12620 10379 12623
rect 10796 12620 10824 12660
rect 10962 12620 10968 12632
rect 10367 12592 10824 12620
rect 10923 12592 10968 12620
rect 10367 12589 10379 12592
rect 10321 12583 10379 12589
rect 10962 12580 10968 12592
rect 11020 12580 11026 12632
rect 11072 12620 11100 12660
rect 11992 12620 12020 12796
rect 12345 12793 12357 12827
rect 12391 12824 12403 12827
rect 12434 12824 12440 12836
rect 12391 12796 12440 12824
rect 12391 12793 12403 12796
rect 12345 12787 12403 12793
rect 12434 12784 12440 12796
rect 12492 12784 12498 12836
rect 13081 12827 13139 12833
rect 13081 12793 13093 12827
rect 13127 12824 13139 12827
rect 13722 12824 13728 12836
rect 13127 12796 13728 12824
rect 13127 12793 13139 12796
rect 13081 12787 13139 12793
rect 13722 12784 13728 12796
rect 13780 12784 13786 12836
rect 18874 12784 18880 12836
rect 18932 12824 18938 12836
rect 18969 12827 19027 12833
rect 18969 12824 18981 12827
rect 18932 12796 18981 12824
rect 18932 12784 18938 12796
rect 18969 12793 18981 12796
rect 19015 12824 19027 12827
rect 19058 12824 19064 12836
rect 19015 12796 19064 12824
rect 19015 12793 19027 12796
rect 18969 12787 19027 12793
rect 19058 12784 19064 12796
rect 19116 12784 19122 12836
rect 19889 12827 19947 12833
rect 19889 12793 19901 12827
rect 19935 12824 19947 12827
rect 20162 12824 20168 12836
rect 19935 12796 20168 12824
rect 19935 12793 19947 12796
rect 19889 12787 19947 12793
rect 20162 12784 20168 12796
rect 20220 12784 20226 12836
rect 20438 12824 20444 12836
rect 20399 12796 20444 12824
rect 20438 12784 20444 12796
rect 20496 12784 20502 12836
rect 21082 12824 21088 12836
rect 21043 12796 21088 12824
rect 21082 12784 21088 12796
rect 21140 12784 21146 12836
rect 15657 12759 15715 12765
rect 15657 12725 15669 12759
rect 15703 12725 15715 12759
rect 15657 12719 15715 12725
rect 17037 12759 17095 12765
rect 17037 12725 17049 12759
rect 17083 12756 17095 12759
rect 19242 12756 19248 12768
rect 17083 12728 19248 12756
rect 17083 12725 17095 12728
rect 17037 12719 17095 12725
rect 13265 12623 13323 12629
rect 13265 12620 13277 12623
rect 11072 12592 11376 12620
rect 11992 12592 13277 12620
rect 11054 12512 11060 12564
rect 11112 12552 11118 12564
rect 11210 12555 11268 12561
rect 11210 12552 11222 12555
rect 11112 12524 11222 12552
rect 11112 12512 11118 12524
rect 11210 12521 11222 12524
rect 11256 12521 11268 12555
rect 11348 12552 11376 12592
rect 13265 12589 13277 12592
rect 13311 12589 13323 12623
rect 15672 12620 15700 12719
rect 19242 12716 19248 12728
rect 19300 12716 19306 12768
rect 16206 12688 16212 12700
rect 16167 12660 16212 12688
rect 16206 12648 16212 12660
rect 16264 12648 16270 12700
rect 17586 12688 17592 12700
rect 17547 12660 17592 12688
rect 17586 12648 17592 12660
rect 17644 12648 17650 12700
rect 17770 12648 17776 12700
rect 17828 12688 17834 12700
rect 17828 12660 20300 12688
rect 17828 12648 17834 12660
rect 17497 12623 17555 12629
rect 17497 12620 17509 12623
rect 15672 12592 17509 12620
rect 13265 12583 13323 12589
rect 17497 12589 17509 12592
rect 17543 12589 17555 12623
rect 17497 12583 17555 12589
rect 19429 12623 19487 12629
rect 19429 12589 19441 12623
rect 19475 12620 19487 12623
rect 19702 12620 19708 12632
rect 19475 12592 19708 12620
rect 19475 12589 19487 12592
rect 19429 12583 19487 12589
rect 19702 12580 19708 12592
rect 19760 12580 19766 12632
rect 20272 12629 20300 12660
rect 20257 12623 20315 12629
rect 20257 12589 20269 12623
rect 20303 12589 20315 12623
rect 20257 12583 20315 12589
rect 20346 12580 20352 12632
rect 20404 12620 20410 12632
rect 20901 12623 20959 12629
rect 20901 12620 20913 12623
rect 20404 12592 20913 12620
rect 20404 12580 20410 12592
rect 20901 12589 20913 12592
rect 20947 12589 20959 12623
rect 20901 12583 20959 12589
rect 12621 12555 12679 12561
rect 12621 12552 12633 12555
rect 11348 12524 12633 12552
rect 11210 12515 11268 12521
rect 12621 12521 12633 12524
rect 12667 12521 12679 12555
rect 12621 12515 12679 12521
rect 16025 12555 16083 12561
rect 16025 12521 16037 12555
rect 16071 12552 16083 12555
rect 16574 12552 16580 12564
rect 16071 12524 16580 12552
rect 16071 12521 16083 12524
rect 16025 12515 16083 12521
rect 16574 12512 16580 12524
rect 16632 12512 16638 12564
rect 17126 12512 17132 12564
rect 17184 12552 17190 12564
rect 18141 12555 18199 12561
rect 18141 12552 18153 12555
rect 17184 12524 18153 12552
rect 17184 12512 17190 12524
rect 18141 12521 18153 12524
rect 18187 12521 18199 12555
rect 18141 12515 18199 12521
rect 7742 12444 7748 12496
rect 7800 12484 7806 12496
rect 8202 12484 8208 12496
rect 7800 12456 8208 12484
rect 7800 12444 7806 12456
rect 8202 12444 8208 12456
rect 8260 12444 8266 12496
rect 10413 12487 10471 12493
rect 10413 12453 10425 12487
rect 10459 12484 10471 12487
rect 11330 12484 11336 12496
rect 10459 12456 11336 12484
rect 10459 12453 10471 12456
rect 10413 12447 10471 12453
rect 11330 12444 11336 12456
rect 11388 12444 11394 12496
rect 14185 12487 14243 12493
rect 14185 12453 14197 12487
rect 14231 12484 14243 12487
rect 14550 12484 14556 12496
rect 14231 12456 14556 12484
rect 14231 12453 14243 12456
rect 14185 12447 14243 12453
rect 14550 12444 14556 12456
rect 14608 12444 14614 12496
rect 16114 12444 16120 12496
rect 16172 12484 16178 12496
rect 16758 12484 16764 12496
rect 16172 12456 16217 12484
rect 16719 12456 16764 12484
rect 16172 12444 16178 12456
rect 16758 12444 16764 12456
rect 16816 12444 16822 12496
rect 17402 12484 17408 12496
rect 17363 12456 17408 12484
rect 17402 12444 17408 12456
rect 17460 12444 17466 12496
rect 18046 12444 18052 12496
rect 18104 12484 18110 12496
rect 18417 12487 18475 12493
rect 18417 12484 18429 12487
rect 18104 12456 18429 12484
rect 18104 12444 18110 12456
rect 18417 12453 18429 12456
rect 18463 12484 18475 12487
rect 18966 12484 18972 12496
rect 18463 12456 18972 12484
rect 18463 12453 18475 12456
rect 18417 12447 18475 12453
rect 18966 12444 18972 12456
rect 19024 12444 19030 12496
rect 1104 12394 21896 12416
rect 1104 12342 7912 12394
rect 7964 12342 7976 12394
rect 8028 12342 8040 12394
rect 8092 12342 8104 12394
rect 8156 12342 14843 12394
rect 14895 12342 14907 12394
rect 14959 12342 14971 12394
rect 15023 12342 15035 12394
rect 15087 12342 21896 12394
rect 1104 12320 21896 12342
rect 10321 12283 10379 12289
rect 10321 12249 10333 12283
rect 10367 12249 10379 12283
rect 10321 12243 10379 12249
rect 10336 12212 10364 12243
rect 10962 12240 10968 12292
rect 11020 12280 11026 12292
rect 13078 12280 13084 12292
rect 11020 12252 13084 12280
rect 11020 12240 11026 12252
rect 13078 12240 13084 12252
rect 13136 12240 13142 12292
rect 13633 12283 13691 12289
rect 13633 12249 13645 12283
rect 13679 12280 13691 12283
rect 14550 12280 14556 12292
rect 13679 12252 14556 12280
rect 13679 12249 13691 12252
rect 13633 12243 13691 12249
rect 14550 12240 14556 12252
rect 14608 12240 14614 12292
rect 15657 12283 15715 12289
rect 15657 12249 15669 12283
rect 15703 12280 15715 12283
rect 16114 12280 16120 12292
rect 15703 12252 16120 12280
rect 15703 12249 15715 12252
rect 15657 12243 15715 12249
rect 16114 12240 16120 12252
rect 16172 12240 16178 12292
rect 16574 12240 16580 12292
rect 16632 12280 16638 12292
rect 16669 12283 16727 12289
rect 16669 12280 16681 12283
rect 16632 12252 16681 12280
rect 16632 12240 16638 12252
rect 16669 12249 16681 12252
rect 16715 12249 16727 12283
rect 16669 12243 16727 12249
rect 16758 12240 16764 12292
rect 16816 12280 16822 12292
rect 18230 12280 18236 12292
rect 16816 12252 18236 12280
rect 16816 12240 16822 12252
rect 18230 12240 18236 12252
rect 18288 12280 18294 12292
rect 18874 12280 18880 12292
rect 18288 12252 18880 12280
rect 18288 12240 18294 12252
rect 18874 12240 18880 12252
rect 18932 12240 18938 12292
rect 19794 12240 19800 12292
rect 19852 12280 19858 12292
rect 20993 12283 21051 12289
rect 20993 12280 21005 12283
rect 19852 12252 21005 12280
rect 19852 12240 19858 12252
rect 20993 12249 21005 12252
rect 21039 12249 21051 12283
rect 20993 12243 21051 12249
rect 11701 12215 11759 12221
rect 10336 12184 11468 12212
rect 10502 12104 10508 12156
rect 10560 12144 10566 12156
rect 11440 12153 11468 12184
rect 11701 12181 11713 12215
rect 11747 12212 11759 12215
rect 15286 12212 15292 12224
rect 11747 12184 15292 12212
rect 11747 12181 11759 12184
rect 11701 12175 11759 12181
rect 15286 12172 15292 12184
rect 15344 12172 15350 12224
rect 16025 12215 16083 12221
rect 16025 12181 16037 12215
rect 16071 12212 16083 12215
rect 16776 12212 16804 12240
rect 17126 12212 17132 12224
rect 16071 12184 16804 12212
rect 17087 12184 17132 12212
rect 16071 12181 16083 12184
rect 16025 12175 16083 12181
rect 10689 12147 10747 12153
rect 10689 12144 10701 12147
rect 10560 12116 10701 12144
rect 10560 12104 10566 12116
rect 10689 12113 10701 12116
rect 10735 12113 10747 12147
rect 10689 12107 10747 12113
rect 11425 12147 11483 12153
rect 11425 12113 11437 12147
rect 11471 12113 11483 12147
rect 14277 12147 14335 12153
rect 14277 12144 14289 12147
rect 11425 12107 11483 12113
rect 13832 12116 14289 12144
rect 8478 12036 8484 12088
rect 8536 12076 8542 12088
rect 10781 12079 10839 12085
rect 10781 12076 10793 12079
rect 8536 12048 10793 12076
rect 8536 12036 8542 12048
rect 10781 12045 10793 12048
rect 10827 12045 10839 12079
rect 10781 12039 10839 12045
rect 10965 12079 11023 12085
rect 10965 12045 10977 12079
rect 11011 12076 11023 12079
rect 11054 12076 11060 12088
rect 11011 12048 11060 12076
rect 11011 12045 11023 12048
rect 10965 12039 11023 12045
rect 11054 12036 11060 12048
rect 11112 12036 11118 12088
rect 12897 12079 12955 12085
rect 12897 12076 12909 12079
rect 12084 12048 12909 12076
rect 842 11968 848 12020
rect 900 12008 906 12020
rect 12084 12008 12112 12048
rect 12897 12045 12909 12048
rect 12943 12076 12955 12079
rect 13725 12079 13783 12085
rect 13725 12076 13737 12079
rect 12943 12048 13737 12076
rect 12943 12045 12955 12048
rect 12897 12039 12955 12045
rect 13725 12045 13737 12048
rect 13771 12045 13783 12079
rect 13725 12039 13783 12045
rect 900 11980 12112 12008
rect 900 11968 906 11980
rect 13630 11968 13636 12020
rect 13688 12008 13694 12020
rect 13832 12008 13860 12116
rect 14277 12113 14289 12116
rect 14323 12113 14335 12147
rect 16040 12144 16068 12175
rect 17126 12172 17132 12184
rect 17184 12172 17190 12224
rect 17678 12172 17684 12224
rect 17736 12212 17742 12224
rect 18417 12215 18475 12221
rect 18417 12212 18429 12215
rect 17736 12184 18429 12212
rect 17736 12172 17742 12184
rect 18417 12181 18429 12184
rect 18463 12181 18475 12215
rect 18417 12175 18475 12181
rect 20165 12215 20223 12221
rect 20165 12181 20177 12215
rect 20211 12212 20223 12215
rect 20346 12212 20352 12224
rect 20211 12184 20352 12212
rect 20211 12181 20223 12184
rect 20165 12175 20223 12181
rect 20346 12172 20352 12184
rect 20404 12172 20410 12224
rect 14277 12107 14335 12113
rect 14476 12116 16068 12144
rect 17037 12147 17095 12153
rect 13909 12079 13967 12085
rect 13909 12045 13921 12079
rect 13955 12076 13967 12079
rect 14366 12076 14372 12088
rect 13955 12048 14372 12076
rect 13955 12045 13967 12048
rect 13909 12039 13967 12045
rect 14366 12036 14372 12048
rect 14424 12036 14430 12088
rect 13688 11980 13860 12008
rect 13688 11968 13694 11980
rect 14274 11968 14280 12020
rect 14332 12008 14338 12020
rect 14476 12008 14504 12116
rect 17037 12113 17049 12147
rect 17083 12144 17095 12147
rect 18046 12144 18052 12156
rect 17083 12116 18052 12144
rect 17083 12113 17095 12116
rect 17037 12107 17095 12113
rect 18046 12104 18052 12116
rect 18104 12104 18110 12156
rect 18138 12104 18144 12156
rect 18196 12144 18202 12156
rect 18509 12147 18567 12153
rect 18509 12144 18521 12147
rect 18196 12116 18521 12144
rect 18196 12104 18202 12116
rect 18509 12113 18521 12116
rect 18555 12113 18567 12147
rect 18509 12107 18567 12113
rect 19242 12104 19248 12156
rect 19300 12144 19306 12156
rect 19889 12147 19947 12153
rect 19889 12144 19901 12147
rect 19300 12116 19901 12144
rect 19300 12104 19306 12116
rect 19889 12113 19901 12116
rect 19935 12113 19947 12147
rect 19889 12107 19947 12113
rect 20809 12147 20867 12153
rect 20809 12113 20821 12147
rect 20855 12144 20867 12147
rect 22005 12147 22063 12153
rect 22005 12144 22017 12147
rect 20855 12116 22017 12144
rect 20855 12113 20867 12116
rect 20809 12107 20867 12113
rect 22005 12113 22017 12116
rect 22051 12113 22063 12147
rect 22005 12107 22063 12113
rect 14553 12079 14611 12085
rect 14553 12045 14565 12079
rect 14599 12045 14611 12079
rect 14553 12039 14611 12045
rect 14332 11980 14504 12008
rect 14568 12008 14596 12039
rect 15194 12036 15200 12088
rect 15252 12076 15258 12088
rect 15381 12079 15439 12085
rect 15381 12076 15393 12079
rect 15252 12048 15393 12076
rect 15252 12036 15258 12048
rect 15381 12045 15393 12048
rect 15427 12076 15439 12079
rect 16117 12079 16175 12085
rect 16117 12076 16129 12079
rect 15427 12048 16129 12076
rect 15427 12045 15439 12048
rect 15381 12039 15439 12045
rect 16117 12045 16129 12048
rect 16163 12045 16175 12079
rect 16117 12039 16175 12045
rect 16301 12079 16359 12085
rect 16301 12045 16313 12079
rect 16347 12076 16359 12079
rect 17313 12079 17371 12085
rect 17313 12076 17325 12079
rect 16347 12048 17325 12076
rect 16347 12045 16359 12048
rect 16301 12039 16359 12045
rect 17313 12045 17325 12048
rect 17359 12076 17371 12079
rect 17862 12076 17868 12088
rect 17359 12048 17868 12076
rect 17359 12045 17371 12048
rect 17313 12039 17371 12045
rect 17862 12036 17868 12048
rect 17920 12036 17926 12088
rect 18598 12076 18604 12088
rect 18559 12048 18604 12076
rect 18598 12036 18604 12048
rect 18656 12036 18662 12088
rect 19613 12079 19671 12085
rect 19613 12045 19625 12079
rect 19659 12076 19671 12079
rect 20824 12076 20852 12107
rect 19659 12048 20852 12076
rect 19659 12045 19671 12048
rect 19613 12039 19671 12045
rect 17770 12008 17776 12020
rect 14568 11980 17776 12008
rect 14332 11968 14338 11980
rect 17770 11968 17776 11980
rect 17828 11968 17834 12020
rect 13265 11943 13323 11949
rect 13265 11909 13277 11943
rect 13311 11940 13323 11943
rect 13538 11940 13544 11952
rect 13311 11912 13544 11940
rect 13311 11909 13323 11912
rect 13265 11903 13323 11909
rect 13538 11900 13544 11912
rect 13596 11900 13602 11952
rect 17402 11900 17408 11952
rect 17460 11940 17466 11952
rect 18049 11943 18107 11949
rect 18049 11940 18061 11943
rect 17460 11912 18061 11940
rect 17460 11900 17466 11912
rect 18049 11909 18061 11912
rect 18095 11909 18107 11943
rect 18049 11903 18107 11909
rect 19058 11900 19064 11952
rect 19116 11940 19122 11952
rect 19153 11943 19211 11949
rect 19153 11940 19165 11943
rect 19116 11912 19165 11940
rect 19116 11900 19122 11912
rect 19153 11909 19165 11912
rect 19199 11909 19211 11943
rect 19153 11903 19211 11909
rect 1104 11850 21896 11872
rect 1104 11798 4447 11850
rect 4499 11798 4511 11850
rect 4563 11798 4575 11850
rect 4627 11798 4639 11850
rect 4691 11798 11378 11850
rect 11430 11798 11442 11850
rect 11494 11798 11506 11850
rect 11558 11798 11570 11850
rect 11622 11798 18308 11850
rect 18360 11798 18372 11850
rect 18424 11798 18436 11850
rect 18488 11798 18500 11850
rect 18552 11798 21896 11850
rect 1104 11776 21896 11798
rect 6638 11696 6644 11748
rect 6696 11736 6702 11748
rect 7653 11739 7711 11745
rect 7653 11736 7665 11739
rect 6696 11708 7665 11736
rect 6696 11696 6702 11708
rect 7653 11705 7665 11708
rect 7699 11736 7711 11739
rect 8849 11739 8907 11745
rect 7699 11708 8524 11736
rect 7699 11705 7711 11708
rect 7653 11699 7711 11705
rect 8294 11560 8300 11612
rect 8352 11560 8358 11612
rect 8496 11609 8524 11708
rect 8849 11705 8861 11739
rect 8895 11736 8907 11739
rect 9125 11739 9183 11745
rect 9125 11736 9137 11739
rect 8895 11708 9137 11736
rect 8895 11705 8907 11708
rect 8849 11699 8907 11705
rect 9125 11705 9137 11708
rect 9171 11736 9183 11739
rect 9490 11736 9496 11748
rect 9171 11708 9496 11736
rect 9171 11705 9183 11708
rect 9125 11699 9183 11705
rect 9490 11696 9496 11708
rect 9548 11736 9554 11748
rect 11054 11736 11060 11748
rect 9548 11708 10732 11736
rect 11015 11708 11060 11736
rect 9548 11696 9554 11708
rect 10704 11668 10732 11708
rect 11054 11696 11060 11708
rect 11112 11696 11118 11748
rect 11238 11696 11244 11748
rect 11296 11736 11302 11748
rect 11333 11739 11391 11745
rect 11333 11736 11345 11739
rect 11296 11708 11345 11736
rect 11296 11696 11302 11708
rect 11333 11705 11345 11708
rect 11379 11705 11391 11739
rect 14274 11736 14280 11748
rect 11333 11699 11391 11705
rect 11440 11708 14280 11736
rect 11440 11668 11468 11708
rect 14274 11696 14280 11708
rect 14332 11696 14338 11748
rect 14366 11696 14372 11748
rect 14424 11736 14430 11748
rect 14461 11739 14519 11745
rect 14461 11736 14473 11739
rect 14424 11708 14473 11736
rect 14424 11696 14430 11708
rect 14461 11705 14473 11708
rect 14507 11705 14519 11739
rect 14461 11699 14519 11705
rect 16206 11696 16212 11748
rect 16264 11696 16270 11748
rect 18138 11736 18144 11748
rect 18099 11708 18144 11736
rect 18138 11696 18144 11708
rect 18196 11696 18202 11748
rect 19337 11739 19395 11745
rect 19337 11705 19349 11739
rect 19383 11736 19395 11739
rect 19610 11736 19616 11748
rect 19383 11708 19616 11736
rect 19383 11705 19395 11708
rect 19337 11699 19395 11705
rect 19610 11696 19616 11708
rect 19668 11696 19674 11748
rect 20070 11696 20076 11748
rect 20128 11736 20134 11748
rect 21085 11739 21143 11745
rect 21085 11736 21097 11739
rect 20128 11708 21097 11736
rect 20128 11696 20134 11708
rect 21085 11705 21097 11708
rect 21131 11705 21143 11739
rect 21085 11699 21143 11705
rect 10704 11640 11468 11668
rect 16224 11668 16252 11696
rect 17770 11668 17776 11680
rect 16224 11640 17776 11668
rect 8481 11603 8539 11609
rect 8481 11569 8493 11603
rect 8527 11569 8539 11603
rect 8481 11563 8539 11569
rect 8665 11603 8723 11609
rect 8665 11569 8677 11603
rect 8711 11600 8723 11603
rect 8754 11600 8760 11612
rect 8711 11572 8760 11600
rect 8711 11569 8723 11572
rect 8665 11563 8723 11569
rect 8754 11560 8760 11572
rect 8812 11560 8818 11612
rect 13078 11600 13084 11612
rect 13039 11572 13084 11600
rect 13078 11560 13084 11572
rect 13136 11560 13142 11612
rect 8312 11532 8340 11560
rect 9677 11535 9735 11541
rect 9677 11532 9689 11535
rect 8312 11504 9689 11532
rect 9677 11501 9689 11504
rect 9723 11501 9735 11535
rect 13096 11532 13124 11560
rect 15194 11532 15200 11544
rect 13096 11504 15200 11532
rect 9677 11495 9735 11501
rect 15194 11492 15200 11504
rect 15252 11532 15258 11544
rect 15289 11535 15347 11541
rect 15289 11532 15301 11535
rect 15252 11504 15301 11532
rect 15252 11492 15258 11504
rect 15289 11501 15301 11504
rect 15335 11501 15347 11535
rect 15289 11495 15347 11501
rect 15556 11535 15614 11541
rect 15556 11501 15568 11535
rect 15602 11532 15614 11535
rect 16316 11532 16344 11640
rect 17770 11628 17776 11640
rect 17828 11668 17834 11680
rect 18598 11668 18604 11680
rect 17828 11640 18604 11668
rect 17828 11628 17834 11640
rect 18598 11628 18604 11640
rect 18656 11628 18662 11680
rect 17678 11600 17684 11612
rect 17639 11572 17684 11600
rect 17678 11560 17684 11572
rect 17736 11560 17742 11612
rect 17862 11560 17868 11612
rect 17920 11600 17926 11612
rect 18782 11600 18788 11612
rect 17920 11572 18788 11600
rect 17920 11560 17926 11572
rect 18782 11560 18788 11572
rect 18840 11560 18846 11612
rect 15602 11504 16344 11532
rect 19153 11535 19211 11541
rect 15602 11501 15614 11504
rect 15556 11495 15614 11501
rect 19153 11501 19165 11535
rect 19199 11532 19211 11535
rect 19426 11532 19432 11544
rect 19199 11504 19432 11532
rect 19199 11501 19211 11504
rect 19153 11495 19211 11501
rect 19426 11492 19432 11504
rect 19484 11492 19490 11544
rect 20533 11535 20591 11541
rect 20533 11501 20545 11535
rect 20579 11532 20591 11535
rect 20898 11532 20904 11544
rect 20579 11504 20904 11532
rect 20579 11501 20591 11504
rect 20533 11495 20591 11501
rect 20898 11492 20904 11504
rect 20956 11492 20962 11544
rect 22002 11532 22008 11544
rect 21963 11504 22008 11532
rect 22002 11492 22008 11504
rect 22060 11492 22066 11544
rect 9950 11473 9956 11476
rect 8389 11467 8447 11473
rect 8389 11433 8401 11467
rect 8435 11464 8447 11467
rect 8849 11467 8907 11473
rect 8849 11464 8861 11467
rect 8435 11436 8861 11464
rect 8435 11433 8447 11436
rect 8389 11427 8447 11433
rect 8849 11433 8861 11436
rect 8895 11433 8907 11467
rect 9944 11464 9956 11473
rect 9911 11436 9956 11464
rect 8849 11427 8907 11433
rect 9944 11427 9956 11436
rect 9950 11424 9956 11427
rect 10008 11424 10014 11476
rect 13348 11467 13406 11473
rect 13348 11433 13360 11467
rect 13394 11464 13406 11467
rect 18506 11464 18512 11476
rect 13394 11436 15608 11464
rect 18419 11436 18512 11464
rect 13394 11433 13406 11436
rect 13348 11427 13406 11433
rect 8021 11399 8079 11405
rect 8021 11365 8033 11399
rect 8067 11396 8079 11399
rect 8294 11396 8300 11408
rect 8067 11368 8300 11396
rect 8067 11365 8079 11368
rect 8021 11359 8079 11365
rect 8294 11356 8300 11368
rect 8352 11356 8358 11408
rect 11238 11356 11244 11408
rect 11296 11396 11302 11408
rect 12342 11396 12348 11408
rect 11296 11368 12348 11396
rect 11296 11356 11302 11368
rect 12342 11356 12348 11368
rect 12400 11396 12406 11408
rect 15470 11396 15476 11408
rect 12400 11368 15476 11396
rect 12400 11356 12406 11368
rect 15470 11356 15476 11368
rect 15528 11356 15534 11408
rect 15580 11396 15608 11436
rect 18506 11424 18512 11436
rect 18564 11464 18570 11476
rect 19242 11464 19248 11476
rect 18564 11436 19248 11464
rect 18564 11424 18570 11436
rect 19242 11424 19248 11436
rect 19300 11424 19306 11476
rect 16669 11399 16727 11405
rect 16669 11396 16681 11399
rect 15580 11368 16681 11396
rect 16669 11365 16681 11368
rect 16715 11396 16727 11399
rect 17586 11396 17592 11408
rect 16715 11368 17592 11396
rect 16715 11365 16727 11368
rect 16669 11359 16727 11365
rect 17586 11356 17592 11368
rect 17644 11356 17650 11408
rect 18598 11396 18604 11408
rect 18511 11368 18604 11396
rect 18598 11356 18604 11368
rect 18656 11396 18662 11408
rect 19334 11396 19340 11408
rect 18656 11368 19340 11396
rect 18656 11356 18662 11368
rect 19334 11356 19340 11368
rect 19392 11396 19398 11408
rect 19705 11399 19763 11405
rect 19705 11396 19717 11399
rect 19392 11368 19717 11396
rect 19392 11356 19398 11368
rect 19705 11365 19717 11368
rect 19751 11365 19763 11399
rect 19705 11359 19763 11365
rect 1104 11306 21896 11328
rect 1104 11254 7912 11306
rect 7964 11254 7976 11306
rect 8028 11254 8040 11306
rect 8092 11254 8104 11306
rect 8156 11254 14843 11306
rect 14895 11254 14907 11306
rect 14959 11254 14971 11306
rect 15023 11254 15035 11306
rect 15087 11254 21896 11306
rect 1104 11232 21896 11254
rect 7466 11152 7472 11204
rect 7524 11192 7530 11204
rect 8573 11195 8631 11201
rect 8573 11192 8585 11195
rect 7524 11164 8585 11192
rect 7524 11152 7530 11164
rect 8573 11161 8585 11164
rect 8619 11192 8631 11195
rect 9125 11195 9183 11201
rect 9125 11192 9137 11195
rect 8619 11164 9137 11192
rect 8619 11161 8631 11164
rect 8573 11155 8631 11161
rect 9125 11161 9137 11164
rect 9171 11161 9183 11195
rect 10502 11192 10508 11204
rect 10463 11164 10508 11192
rect 9125 11155 9183 11161
rect 9140 11124 9168 11155
rect 10502 11152 10508 11164
rect 10560 11152 10566 11204
rect 13078 11152 13084 11204
rect 13136 11192 13142 11204
rect 13541 11195 13599 11201
rect 13541 11192 13553 11195
rect 13136 11164 13553 11192
rect 13136 11152 13142 11164
rect 13541 11161 13553 11164
rect 13587 11161 13599 11195
rect 13541 11155 13599 11161
rect 15470 11152 15476 11204
rect 15528 11192 15534 11204
rect 18506 11192 18512 11204
rect 15528 11164 18512 11192
rect 15528 11152 15534 11164
rect 18506 11152 18512 11164
rect 18564 11152 18570 11204
rect 19978 11152 19984 11204
rect 20036 11192 20042 11204
rect 20993 11195 21051 11201
rect 20993 11192 21005 11195
rect 20036 11164 21005 11192
rect 20036 11152 20042 11164
rect 20993 11161 21005 11164
rect 21039 11161 21051 11195
rect 20993 11155 21051 11161
rect 17126 11124 17132 11136
rect 9140 11096 17132 11124
rect 17126 11084 17132 11096
rect 17184 11124 17190 11136
rect 19058 11124 19064 11136
rect 17184 11096 19064 11124
rect 17184 11084 17190 11096
rect 19058 11084 19064 11096
rect 19116 11084 19122 11136
rect 19426 11124 19432 11136
rect 19387 11096 19432 11124
rect 19426 11084 19432 11096
rect 19484 11084 19490 11136
rect 8481 11059 8539 11065
rect 8481 11025 8493 11059
rect 8527 11056 8539 11059
rect 9585 11059 9643 11065
rect 9585 11056 9597 11059
rect 8527 11028 9597 11056
rect 8527 11025 8539 11028
rect 8481 11019 8539 11025
rect 9585 11025 9597 11028
rect 9631 11056 9643 11059
rect 9858 11056 9864 11068
rect 9631 11028 9864 11056
rect 9631 11025 9643 11028
rect 9585 11019 9643 11025
rect 9858 11016 9864 11028
rect 9916 11016 9922 11068
rect 10870 11056 10876 11068
rect 10831 11028 10876 11056
rect 10870 11016 10876 11028
rect 10928 11016 10934 11068
rect 10965 11059 11023 11065
rect 10965 11025 10977 11059
rect 11011 11056 11023 11059
rect 11146 11056 11152 11068
rect 11011 11028 11152 11056
rect 11011 11025 11023 11028
rect 10965 11019 11023 11025
rect 11146 11016 11152 11028
rect 11204 11016 11210 11068
rect 13722 11056 13728 11068
rect 13683 11028 13728 11056
rect 13722 11016 13728 11028
rect 13780 11016 13786 11068
rect 19150 11056 19156 11068
rect 19111 11028 19156 11056
rect 19150 11016 19156 11028
rect 19208 11016 19214 11068
rect 20165 11059 20223 11065
rect 20165 11025 20177 11059
rect 20211 11056 20223 11059
rect 20622 11056 20628 11068
rect 20211 11028 20628 11056
rect 20211 11025 20223 11028
rect 20165 11019 20223 11025
rect 20622 11016 20628 11028
rect 20680 11056 20686 11068
rect 20809 11059 20867 11065
rect 20809 11056 20821 11059
rect 20680 11028 20821 11056
rect 20680 11016 20686 11028
rect 20809 11025 20821 11028
rect 20855 11025 20867 11059
rect 20809 11019 20867 11025
rect 8754 10988 8760 11000
rect 8667 10960 8760 10988
rect 8754 10948 8760 10960
rect 8812 10988 8818 11000
rect 8812 10960 9628 10988
rect 8812 10948 8818 10960
rect 8113 10923 8171 10929
rect 8113 10889 8125 10923
rect 8159 10920 8171 10923
rect 8386 10920 8392 10932
rect 8159 10892 8392 10920
rect 8159 10889 8171 10892
rect 8113 10883 8171 10889
rect 8386 10880 8392 10892
rect 8444 10880 8450 10932
rect 9600 10852 9628 10960
rect 9876 10920 9904 11016
rect 9950 10948 9956 11000
rect 10008 10988 10014 11000
rect 11057 10991 11115 10997
rect 11057 10988 11069 10991
rect 10008 10960 11069 10988
rect 10008 10948 10014 10960
rect 11057 10957 11069 10960
rect 11103 10957 11115 10991
rect 11057 10951 11115 10957
rect 18690 10920 18696 10932
rect 9876 10892 18696 10920
rect 18690 10880 18696 10892
rect 18748 10920 18754 10932
rect 18966 10920 18972 10932
rect 18748 10892 18972 10920
rect 18748 10880 18754 10892
rect 18966 10880 18972 10892
rect 19024 10880 19030 10932
rect 20530 10920 20536 10932
rect 20491 10892 20536 10920
rect 20530 10880 20536 10892
rect 20588 10880 20594 10932
rect 11698 10852 11704 10864
rect 9600 10824 11704 10852
rect 11698 10812 11704 10824
rect 11756 10812 11762 10864
rect 13998 10812 14004 10864
rect 14056 10852 14062 10864
rect 18598 10852 18604 10864
rect 14056 10824 18604 10852
rect 14056 10812 14062 10824
rect 18598 10812 18604 10824
rect 18656 10812 18662 10864
rect 1104 10762 21896 10784
rect 1104 10710 4447 10762
rect 4499 10710 4511 10762
rect 4563 10710 4575 10762
rect 4627 10710 4639 10762
rect 4691 10710 11378 10762
rect 11430 10710 11442 10762
rect 11494 10710 11506 10762
rect 11558 10710 11570 10762
rect 11622 10710 18308 10762
rect 18360 10710 18372 10762
rect 18424 10710 18436 10762
rect 18488 10710 18500 10762
rect 18552 10710 21896 10762
rect 1104 10688 21896 10710
rect 8021 10651 8079 10657
rect 8021 10617 8033 10651
rect 8067 10648 8079 10651
rect 8478 10648 8484 10660
rect 8067 10620 8484 10648
rect 8067 10617 8079 10620
rect 8021 10611 8079 10617
rect 8478 10608 8484 10620
rect 8536 10608 8542 10660
rect 11146 10648 11152 10660
rect 11107 10620 11152 10648
rect 11146 10608 11152 10620
rect 11204 10608 11210 10660
rect 12342 10608 12348 10660
rect 12400 10648 12406 10660
rect 12529 10651 12587 10657
rect 12529 10648 12541 10651
rect 12400 10620 12541 10648
rect 12400 10608 12406 10620
rect 12529 10617 12541 10620
rect 12575 10617 12587 10651
rect 12529 10611 12587 10617
rect 19150 10608 19156 10660
rect 19208 10648 19214 10660
rect 19245 10651 19303 10657
rect 19245 10648 19257 10651
rect 19208 10620 19257 10648
rect 19208 10608 19214 10620
rect 19245 10617 19257 10620
rect 19291 10617 19303 10651
rect 19245 10611 19303 10617
rect 21085 10651 21143 10657
rect 21085 10617 21097 10651
rect 21131 10648 21143 10651
rect 21450 10648 21456 10660
rect 21131 10620 21456 10648
rect 21131 10617 21143 10620
rect 21085 10611 21143 10617
rect 21450 10608 21456 10620
rect 21508 10608 21514 10660
rect 12253 10583 12311 10589
rect 12253 10580 12265 10583
rect 11624 10552 12265 10580
rect 8294 10472 8300 10524
rect 8352 10512 8358 10524
rect 8481 10515 8539 10521
rect 8481 10512 8493 10515
rect 8352 10484 8493 10512
rect 8352 10472 8358 10484
rect 8481 10481 8493 10484
rect 8527 10481 8539 10515
rect 8481 10475 8539 10481
rect 8665 10515 8723 10521
rect 8665 10481 8677 10515
rect 8711 10512 8723 10515
rect 9950 10512 9956 10524
rect 8711 10484 9956 10512
rect 8711 10481 8723 10484
rect 8665 10475 8723 10481
rect 9950 10472 9956 10484
rect 10008 10472 10014 10524
rect 10689 10515 10747 10521
rect 10689 10481 10701 10515
rect 10735 10512 10747 10515
rect 10870 10512 10876 10524
rect 10735 10484 10876 10512
rect 10735 10481 10747 10484
rect 10689 10475 10747 10481
rect 10870 10472 10876 10484
rect 10928 10472 10934 10524
rect 11624 10521 11652 10552
rect 12253 10549 12265 10552
rect 12299 10580 12311 10583
rect 13998 10580 14004 10592
rect 12299 10552 14004 10580
rect 12299 10549 12311 10552
rect 12253 10543 12311 10549
rect 13998 10540 14004 10552
rect 14056 10540 14062 10592
rect 11609 10515 11667 10521
rect 11609 10481 11621 10515
rect 11655 10481 11667 10515
rect 11609 10475 11667 10481
rect 11698 10472 11704 10524
rect 11756 10512 11762 10524
rect 14185 10515 14243 10521
rect 11756 10484 11801 10512
rect 11756 10472 11762 10484
rect 14185 10481 14197 10515
rect 14231 10512 14243 10515
rect 14366 10512 14372 10524
rect 14231 10484 14372 10512
rect 14231 10481 14243 10484
rect 14185 10475 14243 10481
rect 14366 10472 14372 10484
rect 14424 10472 14430 10524
rect 19886 10512 19892 10524
rect 19847 10484 19892 10512
rect 19886 10472 19892 10484
rect 19944 10472 19950 10524
rect 8386 10444 8392 10456
rect 8347 10416 8392 10444
rect 8386 10404 8392 10416
rect 8444 10404 8450 10456
rect 11517 10447 11575 10453
rect 11517 10413 11529 10447
rect 11563 10444 11575 10447
rect 12342 10444 12348 10456
rect 11563 10416 12348 10444
rect 11563 10413 11575 10416
rect 11517 10407 11575 10413
rect 12342 10404 12348 10416
rect 12400 10404 12406 10456
rect 13998 10404 14004 10456
rect 14056 10444 14062 10456
rect 15289 10447 15347 10453
rect 15289 10444 15301 10447
rect 14056 10416 15301 10444
rect 14056 10404 14062 10416
rect 15289 10413 15301 10416
rect 15335 10413 15347 10447
rect 15289 10407 15347 10413
rect 20622 10404 20628 10456
rect 20680 10444 20686 10456
rect 20901 10447 20959 10453
rect 20901 10444 20913 10447
rect 20680 10416 20913 10444
rect 20680 10404 20686 10416
rect 20901 10413 20913 10416
rect 20947 10413 20959 10447
rect 20901 10407 20959 10413
rect 13814 10336 13820 10388
rect 13872 10376 13878 10388
rect 13909 10379 13967 10385
rect 13909 10376 13921 10379
rect 13872 10348 13921 10376
rect 13872 10336 13878 10348
rect 13909 10345 13921 10348
rect 13955 10376 13967 10379
rect 19613 10379 19671 10385
rect 13955 10348 14320 10376
rect 13955 10345 13967 10348
rect 13909 10339 13967 10345
rect 14292 10320 14320 10348
rect 19613 10345 19625 10379
rect 19659 10376 19671 10379
rect 20257 10379 20315 10385
rect 20257 10376 20269 10379
rect 19659 10348 20269 10376
rect 19659 10345 19671 10348
rect 19613 10339 19671 10345
rect 20257 10345 20269 10348
rect 20303 10345 20315 10379
rect 20257 10339 20315 10345
rect 13446 10268 13452 10320
rect 13504 10308 13510 10320
rect 13541 10311 13599 10317
rect 13541 10308 13553 10311
rect 13504 10280 13553 10308
rect 13504 10268 13510 10280
rect 13541 10277 13553 10280
rect 13587 10277 13599 10311
rect 13998 10308 14004 10320
rect 13959 10280 14004 10308
rect 13541 10271 13599 10277
rect 13998 10268 14004 10280
rect 14056 10268 14062 10320
rect 14274 10268 14280 10320
rect 14332 10308 14338 10320
rect 14553 10311 14611 10317
rect 14553 10308 14565 10311
rect 14332 10280 14565 10308
rect 14332 10268 14338 10280
rect 14553 10277 14565 10280
rect 14599 10277 14611 10311
rect 18966 10308 18972 10320
rect 18927 10280 18972 10308
rect 14553 10271 14611 10277
rect 18966 10268 18972 10280
rect 19024 10268 19030 10320
rect 19702 10308 19708 10320
rect 19663 10280 19708 10308
rect 19702 10268 19708 10280
rect 19760 10268 19766 10320
rect 1104 10218 21896 10240
rect 1104 10166 7912 10218
rect 7964 10166 7976 10218
rect 8028 10166 8040 10218
rect 8092 10166 8104 10218
rect 8156 10166 14843 10218
rect 14895 10166 14907 10218
rect 14959 10166 14971 10218
rect 15023 10166 15035 10218
rect 15087 10166 21896 10218
rect 1104 10144 21896 10166
rect 8202 10104 8208 10116
rect 7944 10076 8208 10104
rect 7944 9977 7972 10076
rect 8202 10064 8208 10076
rect 8260 10064 8266 10116
rect 9309 10107 9367 10113
rect 9309 10073 9321 10107
rect 9355 10104 9367 10107
rect 9950 10104 9956 10116
rect 9355 10076 9956 10104
rect 9355 10073 9367 10076
rect 9309 10067 9367 10073
rect 9950 10064 9956 10076
rect 10008 10064 10014 10116
rect 13446 10104 13452 10116
rect 13407 10076 13452 10104
rect 13446 10064 13452 10076
rect 13504 10064 13510 10116
rect 13538 10064 13544 10116
rect 13596 10104 13602 10116
rect 17589 10107 17647 10113
rect 13596 10076 13641 10104
rect 13596 10064 13602 10076
rect 17589 10073 17601 10107
rect 17635 10104 17647 10107
rect 17770 10104 17776 10116
rect 17635 10076 17776 10104
rect 17635 10073 17647 10076
rect 17589 10067 17647 10073
rect 17770 10064 17776 10076
rect 17828 10064 17834 10116
rect 18782 10064 18788 10116
rect 18840 10104 18846 10116
rect 19429 10107 19487 10113
rect 19429 10104 19441 10107
rect 18840 10076 19441 10104
rect 18840 10064 18846 10076
rect 19429 10073 19441 10076
rect 19475 10073 19487 10107
rect 19702 10104 19708 10116
rect 19663 10076 19708 10104
rect 19429 10067 19487 10073
rect 19702 10064 19708 10076
rect 19760 10064 19766 10116
rect 20070 10104 20076 10116
rect 20031 10076 20076 10104
rect 20070 10064 20076 10076
rect 20128 10064 20134 10116
rect 20993 10107 21051 10113
rect 20993 10073 21005 10107
rect 21039 10104 21051 10107
rect 21634 10104 21640 10116
rect 21039 10076 21640 10104
rect 21039 10073 21051 10076
rect 20993 10067 21051 10073
rect 21634 10064 21640 10076
rect 21692 10064 21698 10116
rect 14366 9996 14372 10048
rect 14424 10045 14430 10048
rect 14424 10039 14488 10045
rect 14424 10005 14442 10039
rect 14476 10005 14488 10039
rect 14424 9999 14488 10005
rect 16476 10039 16534 10045
rect 16476 10005 16488 10039
rect 16522 10036 16534 10039
rect 18800 10036 18828 10064
rect 16522 10008 18828 10036
rect 16522 10005 16534 10008
rect 16476 9999 16534 10005
rect 14424 9996 14430 9999
rect 18966 9996 18972 10048
rect 19024 10036 19030 10048
rect 20165 10039 20223 10045
rect 20165 10036 20177 10039
rect 19024 10008 20177 10036
rect 19024 9996 19030 10008
rect 20165 10005 20177 10008
rect 20211 10005 20223 10039
rect 20165 9999 20223 10005
rect 7929 9971 7987 9977
rect 7929 9937 7941 9971
rect 7975 9937 7987 9971
rect 7929 9931 7987 9937
rect 8196 9971 8254 9977
rect 8196 9937 8208 9971
rect 8242 9968 8254 9971
rect 8754 9968 8760 9980
rect 8242 9940 8760 9968
rect 8242 9937 8254 9940
rect 8196 9931 8254 9937
rect 8754 9928 8760 9940
rect 8812 9928 8818 9980
rect 14185 9971 14243 9977
rect 14185 9937 14197 9971
rect 14231 9968 14243 9971
rect 15194 9968 15200 9980
rect 14231 9940 15200 9968
rect 14231 9937 14243 9940
rect 14185 9931 14243 9937
rect 15194 9928 15200 9940
rect 15252 9968 15258 9980
rect 16209 9971 16267 9977
rect 16209 9968 16221 9971
rect 15252 9940 16221 9968
rect 15252 9928 15258 9940
rect 16209 9937 16221 9940
rect 16255 9968 16267 9971
rect 18046 9968 18052 9980
rect 16255 9940 18052 9968
rect 16255 9937 16267 9940
rect 16209 9931 16267 9937
rect 18046 9928 18052 9940
rect 18104 9928 18110 9980
rect 18316 9971 18374 9977
rect 18316 9937 18328 9971
rect 18362 9968 18374 9971
rect 19886 9968 19892 9980
rect 18362 9940 19892 9968
rect 18362 9937 18374 9940
rect 18316 9931 18374 9937
rect 19886 9928 19892 9940
rect 19944 9928 19950 9980
rect 20530 9928 20536 9980
rect 20588 9968 20594 9980
rect 20809 9971 20867 9977
rect 20809 9968 20821 9971
rect 20588 9940 20821 9968
rect 20588 9928 20594 9940
rect 20809 9937 20821 9940
rect 20855 9937 20867 9971
rect 20809 9931 20867 9937
rect 13078 9860 13084 9912
rect 13136 9900 13142 9912
rect 13633 9903 13691 9909
rect 13633 9900 13645 9903
rect 13136 9872 13645 9900
rect 13136 9860 13142 9872
rect 13633 9869 13645 9872
rect 13679 9869 13691 9903
rect 20254 9900 20260 9912
rect 20215 9872 20260 9900
rect 13633 9863 13691 9869
rect 13648 9832 13676 9863
rect 20254 9860 20260 9872
rect 20312 9860 20318 9912
rect 13648 9804 14136 9832
rect 13081 9767 13139 9773
rect 13081 9733 13093 9767
rect 13127 9764 13139 9767
rect 13906 9764 13912 9776
rect 13127 9736 13912 9764
rect 13127 9733 13139 9736
rect 13081 9727 13139 9733
rect 13906 9724 13912 9736
rect 13964 9724 13970 9776
rect 14108 9764 14136 9804
rect 15565 9767 15623 9773
rect 15565 9764 15577 9767
rect 14108 9736 15577 9764
rect 15565 9733 15577 9736
rect 15611 9764 15623 9767
rect 15838 9764 15844 9776
rect 15611 9736 15844 9764
rect 15611 9733 15623 9736
rect 15565 9727 15623 9733
rect 15838 9724 15844 9736
rect 15896 9724 15902 9776
rect 1104 9674 21896 9696
rect 1104 9622 4447 9674
rect 4499 9622 4511 9674
rect 4563 9622 4575 9674
rect 4627 9622 4639 9674
rect 4691 9622 11378 9674
rect 11430 9622 11442 9674
rect 11494 9622 11506 9674
rect 11558 9622 11570 9674
rect 11622 9622 18308 9674
rect 18360 9622 18372 9674
rect 18424 9622 18436 9674
rect 18488 9622 18500 9674
rect 18552 9622 21896 9674
rect 1104 9600 21896 9622
rect 11517 9563 11575 9569
rect 11517 9529 11529 9563
rect 11563 9560 11575 9563
rect 11698 9560 11704 9572
rect 11563 9532 11704 9560
rect 11563 9529 11575 9532
rect 11517 9523 11575 9529
rect 11698 9520 11704 9532
rect 11756 9520 11762 9572
rect 19886 9520 19892 9572
rect 19944 9560 19950 9572
rect 20073 9563 20131 9569
rect 20073 9560 20085 9563
rect 19944 9532 20085 9560
rect 19944 9520 19950 9532
rect 20073 9529 20085 9532
rect 20119 9529 20131 9563
rect 20073 9523 20131 9529
rect 13173 9495 13231 9501
rect 13173 9461 13185 9495
rect 13219 9492 13231 9495
rect 21085 9495 21143 9501
rect 13219 9464 14044 9492
rect 13219 9461 13231 9464
rect 13173 9455 13231 9461
rect 10137 9359 10195 9365
rect 10137 9325 10149 9359
rect 10183 9356 10195 9359
rect 11701 9359 11759 9365
rect 11701 9356 11713 9359
rect 10183 9328 11713 9356
rect 10183 9325 10195 9328
rect 10137 9319 10195 9325
rect 11701 9325 11713 9328
rect 11747 9356 11759 9359
rect 11793 9359 11851 9365
rect 11793 9356 11805 9359
rect 11747 9328 11805 9356
rect 11747 9325 11759 9328
rect 11701 9319 11759 9325
rect 11793 9325 11805 9328
rect 11839 9325 11851 9359
rect 11793 9319 11851 9325
rect 12060 9359 12118 9365
rect 12060 9325 12072 9359
rect 12106 9356 12118 9359
rect 13078 9356 13084 9368
rect 12106 9328 13084 9356
rect 12106 9325 12118 9328
rect 12060 9319 12118 9325
rect 13078 9316 13084 9328
rect 13136 9316 13142 9368
rect 10404 9291 10462 9297
rect 10404 9257 10416 9291
rect 10450 9288 10462 9291
rect 13188 9288 13216 9455
rect 13906 9424 13912 9436
rect 13867 9396 13912 9424
rect 13906 9384 13912 9396
rect 13964 9384 13970 9436
rect 14016 9433 14044 9464
rect 21085 9461 21097 9495
rect 21131 9492 21143 9495
rect 21726 9492 21732 9504
rect 21131 9464 21732 9492
rect 21131 9461 21143 9464
rect 21085 9455 21143 9461
rect 21726 9452 21732 9464
rect 21784 9452 21790 9504
rect 14001 9427 14059 9433
rect 14001 9393 14013 9427
rect 14047 9393 14059 9427
rect 15838 9424 15844 9436
rect 15799 9396 15844 9424
rect 14001 9387 14059 9393
rect 15838 9384 15844 9396
rect 15896 9384 15902 9436
rect 18046 9384 18052 9436
rect 18104 9424 18110 9436
rect 18693 9427 18751 9433
rect 18693 9424 18705 9427
rect 18104 9396 18705 9424
rect 18104 9384 18110 9396
rect 18693 9393 18705 9396
rect 18739 9393 18751 9427
rect 18693 9387 18751 9393
rect 18960 9359 19018 9365
rect 18960 9325 18972 9359
rect 19006 9356 19018 9359
rect 19702 9356 19708 9368
rect 19006 9328 19708 9356
rect 19006 9325 19018 9328
rect 18960 9319 19018 9325
rect 19702 9316 19708 9328
rect 19760 9356 19766 9368
rect 20254 9356 20260 9368
rect 19760 9328 20260 9356
rect 19760 9316 19766 9328
rect 20254 9316 20260 9328
rect 20312 9316 20318 9368
rect 20533 9359 20591 9365
rect 20533 9325 20545 9359
rect 20579 9356 20591 9359
rect 20898 9356 20904 9368
rect 20579 9328 20904 9356
rect 20579 9325 20591 9328
rect 20533 9319 20591 9325
rect 20898 9316 20904 9328
rect 20956 9316 20962 9368
rect 10450 9260 13216 9288
rect 13817 9291 13875 9297
rect 10450 9257 10462 9260
rect 10404 9251 10462 9257
rect 13817 9257 13829 9291
rect 13863 9288 13875 9291
rect 13863 9260 15332 9288
rect 13863 9257 13875 9260
rect 13817 9251 13875 9257
rect 11701 9223 11759 9229
rect 11701 9189 11713 9223
rect 11747 9220 11759 9223
rect 12986 9220 12992 9232
rect 11747 9192 12992 9220
rect 11747 9189 11759 9192
rect 11701 9183 11759 9189
rect 12986 9180 12992 9192
rect 13044 9180 13050 9232
rect 13449 9223 13507 9229
rect 13449 9189 13461 9223
rect 13495 9220 13507 9223
rect 13630 9220 13636 9232
rect 13495 9192 13636 9220
rect 13495 9189 13507 9192
rect 13449 9183 13507 9189
rect 13630 9180 13636 9192
rect 13688 9180 13694 9232
rect 15304 9229 15332 9260
rect 15289 9223 15347 9229
rect 15289 9189 15301 9223
rect 15335 9189 15347 9223
rect 15289 9183 15347 9189
rect 15378 9180 15384 9232
rect 15436 9220 15442 9232
rect 15657 9223 15715 9229
rect 15657 9220 15669 9223
rect 15436 9192 15669 9220
rect 15436 9180 15442 9192
rect 15657 9189 15669 9192
rect 15703 9189 15715 9223
rect 15657 9183 15715 9189
rect 15749 9223 15807 9229
rect 15749 9189 15761 9223
rect 15795 9220 15807 9223
rect 16393 9223 16451 9229
rect 16393 9220 16405 9223
rect 15795 9192 16405 9220
rect 15795 9189 15807 9192
rect 15749 9183 15807 9189
rect 16393 9189 16405 9192
rect 16439 9220 16451 9223
rect 16482 9220 16488 9232
rect 16439 9192 16488 9220
rect 16439 9189 16451 9192
rect 16393 9183 16451 9189
rect 16482 9180 16488 9192
rect 16540 9180 16546 9232
rect 1104 9130 21896 9152
rect 1104 9078 7912 9130
rect 7964 9078 7976 9130
rect 8028 9078 8040 9130
rect 8092 9078 8104 9130
rect 8156 9078 14843 9130
rect 14895 9078 14907 9130
rect 14959 9078 14971 9130
rect 15023 9078 15035 9130
rect 15087 9078 21896 9130
rect 1104 9056 21896 9078
rect 11885 9019 11943 9025
rect 11885 8985 11897 9019
rect 11931 9016 11943 9019
rect 12066 9016 12072 9028
rect 11931 8988 12072 9016
rect 11931 8985 11943 8988
rect 11885 8979 11943 8985
rect 12066 8976 12072 8988
rect 12124 8976 12130 9028
rect 13170 8976 13176 9028
rect 13228 9016 13234 9028
rect 13449 9019 13507 9025
rect 13449 9016 13461 9019
rect 13228 8988 13461 9016
rect 13228 8976 13234 8988
rect 13449 8985 13461 8988
rect 13495 8985 13507 9019
rect 15378 9016 15384 9028
rect 15339 8988 15384 9016
rect 13449 8979 13507 8985
rect 15378 8976 15384 8988
rect 15436 8976 15442 9028
rect 15654 8976 15660 9028
rect 15712 9016 15718 9028
rect 16209 9019 16267 9025
rect 16209 9016 16221 9019
rect 15712 8988 16221 9016
rect 15712 8976 15718 8988
rect 16209 8985 16221 8988
rect 16255 8985 16267 9019
rect 20070 9016 20076 9028
rect 20031 8988 20076 9016
rect 16209 8979 16267 8985
rect 20070 8976 20076 8988
rect 20128 8976 20134 9028
rect 20530 9016 20536 9028
rect 20491 8988 20536 9016
rect 20530 8976 20536 8988
rect 20588 8976 20594 9028
rect 11698 8880 11704 8892
rect 11659 8852 11704 8880
rect 11698 8840 11704 8852
rect 11756 8840 11762 8892
rect 13265 8883 13323 8889
rect 13265 8849 13277 8883
rect 13311 8880 13323 8883
rect 13630 8880 13636 8892
rect 13311 8852 13636 8880
rect 13311 8849 13323 8852
rect 13265 8843 13323 8849
rect 13630 8840 13636 8852
rect 13688 8840 13694 8892
rect 16025 8883 16083 8889
rect 16025 8849 16037 8883
rect 16071 8880 16083 8883
rect 16574 8880 16580 8892
rect 16071 8852 16580 8880
rect 16071 8849 16083 8852
rect 16025 8843 16083 8849
rect 16574 8840 16580 8852
rect 16632 8840 16638 8892
rect 19797 8883 19855 8889
rect 19797 8849 19809 8883
rect 19843 8880 19855 8883
rect 20809 8883 20867 8889
rect 20809 8880 20821 8883
rect 19843 8852 20821 8880
rect 19843 8849 19855 8852
rect 19797 8843 19855 8849
rect 20809 8849 20821 8852
rect 20855 8880 20867 8883
rect 22005 8883 22063 8889
rect 22005 8880 22017 8883
rect 20855 8852 22017 8880
rect 20855 8849 20867 8852
rect 20809 8843 20867 8849
rect 22005 8849 22017 8852
rect 22051 8849 22063 8883
rect 22005 8843 22063 8849
rect 16390 8704 16396 8756
rect 16448 8744 16454 8756
rect 20993 8747 21051 8753
rect 20993 8744 21005 8747
rect 16448 8716 21005 8744
rect 16448 8704 16454 8716
rect 20993 8713 21005 8716
rect 21039 8713 21051 8747
rect 20993 8707 21051 8713
rect 1104 8586 21896 8608
rect 1104 8534 4447 8586
rect 4499 8534 4511 8586
rect 4563 8534 4575 8586
rect 4627 8534 4639 8586
rect 4691 8534 11378 8586
rect 11430 8534 11442 8586
rect 11494 8534 11506 8586
rect 11558 8534 11570 8586
rect 11622 8534 18308 8586
rect 18360 8534 18372 8586
rect 18424 8534 18436 8586
rect 18488 8534 18500 8586
rect 18552 8534 21896 8586
rect 1104 8512 21896 8534
rect 16298 8432 16304 8484
rect 16356 8472 16362 8484
rect 21085 8475 21143 8481
rect 21085 8472 21097 8475
rect 16356 8444 21097 8472
rect 16356 8432 16362 8444
rect 21085 8441 21097 8444
rect 21131 8441 21143 8475
rect 21085 8435 21143 8441
rect 11333 8339 11391 8345
rect 11333 8305 11345 8339
rect 11379 8336 11391 8339
rect 11698 8336 11704 8348
rect 11379 8308 11704 8336
rect 11379 8305 11391 8308
rect 11333 8299 11391 8305
rect 11698 8296 11704 8308
rect 11756 8296 11762 8348
rect 13630 8336 13636 8348
rect 13591 8308 13636 8336
rect 13630 8296 13636 8308
rect 13688 8296 13694 8348
rect 16574 8336 16580 8348
rect 16535 8308 16580 8336
rect 16574 8296 16580 8308
rect 16632 8296 16638 8348
rect 11054 8268 11060 8280
rect 11015 8240 11060 8268
rect 11054 8228 11060 8240
rect 11112 8228 11118 8280
rect 13449 8271 13507 8277
rect 13449 8237 13461 8271
rect 13495 8268 13507 8271
rect 14090 8268 14096 8280
rect 13495 8240 14096 8268
rect 13495 8237 13507 8240
rect 13449 8231 13507 8237
rect 14090 8228 14096 8240
rect 14148 8228 14154 8280
rect 16393 8271 16451 8277
rect 16393 8237 16405 8271
rect 16439 8268 16451 8271
rect 16942 8268 16948 8280
rect 16439 8240 16948 8268
rect 16439 8237 16451 8240
rect 16393 8231 16451 8237
rect 16942 8228 16948 8240
rect 17000 8228 17006 8280
rect 20533 8271 20591 8277
rect 20533 8237 20545 8271
rect 20579 8268 20591 8271
rect 20622 8268 20628 8280
rect 20579 8240 20628 8268
rect 20579 8237 20591 8240
rect 20533 8231 20591 8237
rect 20622 8228 20628 8240
rect 20680 8268 20686 8280
rect 20901 8271 20959 8277
rect 20901 8268 20913 8271
rect 20680 8240 20913 8268
rect 20680 8228 20686 8240
rect 20901 8237 20913 8240
rect 20947 8237 20959 8271
rect 22002 8268 22008 8280
rect 21963 8240 22008 8268
rect 20901 8231 20959 8237
rect 22002 8228 22008 8240
rect 22060 8228 22066 8280
rect 14182 8092 14188 8144
rect 14240 8132 14246 8144
rect 21082 8132 21088 8144
rect 14240 8104 21088 8132
rect 14240 8092 14246 8104
rect 21082 8092 21088 8104
rect 21140 8092 21146 8144
rect 1104 8042 21896 8064
rect 1104 7990 7912 8042
rect 7964 7990 7976 8042
rect 8028 7990 8040 8042
rect 8092 7990 8104 8042
rect 8156 7990 14843 8042
rect 14895 7990 14907 8042
rect 14959 7990 14971 8042
rect 15023 7990 15035 8042
rect 15087 7990 21896 8042
rect 1104 7968 21896 7990
rect 11054 7888 11060 7940
rect 11112 7928 11118 7940
rect 11149 7931 11207 7937
rect 11149 7928 11161 7931
rect 11112 7900 11161 7928
rect 11112 7888 11118 7900
rect 11149 7897 11161 7900
rect 11195 7897 11207 7931
rect 16942 7928 16948 7940
rect 16903 7900 16948 7928
rect 11149 7891 11207 7897
rect 16942 7888 16948 7900
rect 17000 7888 17006 7940
rect 19613 7931 19671 7937
rect 17236 7900 18460 7928
rect 15930 7820 15936 7872
rect 15988 7860 15994 7872
rect 17236 7860 17264 7900
rect 15988 7832 17264 7860
rect 17313 7863 17371 7869
rect 15988 7820 15994 7832
rect 17313 7829 17325 7863
rect 17359 7860 17371 7863
rect 18046 7860 18052 7872
rect 17359 7832 18052 7860
rect 17359 7829 17371 7832
rect 17313 7823 17371 7829
rect 18046 7820 18052 7832
rect 18104 7820 18110 7872
rect 18432 7860 18460 7900
rect 19613 7897 19625 7931
rect 19659 7928 19671 7931
rect 19702 7928 19708 7940
rect 19659 7900 19708 7928
rect 19659 7897 19671 7900
rect 19613 7891 19671 7897
rect 19702 7888 19708 7900
rect 19760 7888 19766 7940
rect 20993 7931 21051 7937
rect 20993 7897 21005 7931
rect 21039 7897 21051 7931
rect 20993 7891 21051 7897
rect 21008 7860 21036 7891
rect 18432 7832 21036 7860
rect 10689 7795 10747 7801
rect 10689 7761 10701 7795
rect 10735 7792 10747 7795
rect 11517 7795 11575 7801
rect 11517 7792 11529 7795
rect 10735 7764 11529 7792
rect 10735 7761 10747 7764
rect 10689 7755 10747 7761
rect 11517 7761 11529 7764
rect 11563 7761 11575 7795
rect 11517 7755 11575 7761
rect 12986 7752 12992 7804
rect 13044 7792 13050 7804
rect 13633 7795 13691 7801
rect 13633 7792 13645 7795
rect 13044 7764 13645 7792
rect 13044 7752 13050 7764
rect 13633 7761 13645 7764
rect 13679 7792 13691 7795
rect 13722 7792 13728 7804
rect 13679 7764 13728 7792
rect 13679 7761 13691 7764
rect 13633 7755 13691 7761
rect 13722 7752 13728 7764
rect 13780 7752 13786 7804
rect 13906 7801 13912 7804
rect 13900 7792 13912 7801
rect 13867 7764 13912 7792
rect 13900 7755 13912 7764
rect 13906 7752 13912 7755
rect 13964 7752 13970 7804
rect 18138 7792 18144 7804
rect 17604 7764 18144 7792
rect 11238 7684 11244 7736
rect 11296 7724 11302 7736
rect 11609 7727 11667 7733
rect 11609 7724 11621 7727
rect 11296 7696 11621 7724
rect 11296 7684 11302 7696
rect 11609 7693 11621 7696
rect 11655 7693 11667 7727
rect 11609 7687 11667 7693
rect 11698 7684 11704 7736
rect 11756 7724 11762 7736
rect 15286 7724 15292 7736
rect 11756 7696 11801 7724
rect 15247 7696 15292 7724
rect 11756 7684 11762 7696
rect 15286 7684 15292 7696
rect 15344 7684 15350 7736
rect 17604 7733 17632 7764
rect 18138 7752 18144 7764
rect 18196 7792 18202 7804
rect 18489 7795 18547 7801
rect 18489 7792 18501 7795
rect 18196 7764 18501 7792
rect 18196 7752 18202 7764
rect 18489 7761 18501 7764
rect 18535 7761 18547 7795
rect 18489 7755 18547 7761
rect 20533 7795 20591 7801
rect 20533 7761 20545 7795
rect 20579 7792 20591 7795
rect 20806 7792 20812 7804
rect 20579 7764 20812 7792
rect 20579 7761 20591 7764
rect 20533 7755 20591 7761
rect 20806 7752 20812 7764
rect 20864 7752 20870 7804
rect 17405 7727 17463 7733
rect 17405 7693 17417 7727
rect 17451 7693 17463 7727
rect 17405 7687 17463 7693
rect 17589 7727 17647 7733
rect 17589 7693 17601 7727
rect 17635 7693 17647 7727
rect 17589 7687 17647 7693
rect 15010 7588 15016 7600
rect 14971 7560 15016 7588
rect 15010 7548 15016 7560
rect 15068 7548 15074 7600
rect 17420 7588 17448 7687
rect 17954 7684 17960 7736
rect 18012 7724 18018 7736
rect 18233 7727 18291 7733
rect 18233 7724 18245 7727
rect 18012 7696 18245 7724
rect 18012 7684 18018 7696
rect 18233 7693 18245 7696
rect 18279 7693 18291 7727
rect 18233 7687 18291 7693
rect 18598 7588 18604 7600
rect 17420 7560 18604 7588
rect 18598 7548 18604 7560
rect 18656 7548 18662 7600
rect 1104 7498 21896 7520
rect 1104 7446 4447 7498
rect 4499 7446 4511 7498
rect 4563 7446 4575 7498
rect 4627 7446 4639 7498
rect 4691 7446 11378 7498
rect 11430 7446 11442 7498
rect 11494 7446 11506 7498
rect 11558 7446 11570 7498
rect 11622 7446 18308 7498
rect 18360 7446 18372 7498
rect 18424 7446 18436 7498
rect 18488 7446 18500 7498
rect 18552 7446 21896 7498
rect 1104 7424 21896 7446
rect 11241 7387 11299 7393
rect 11241 7353 11253 7387
rect 11287 7384 11299 7387
rect 11698 7384 11704 7396
rect 11287 7356 11704 7384
rect 11287 7353 11299 7356
rect 11241 7347 11299 7353
rect 11698 7344 11704 7356
rect 11756 7344 11762 7396
rect 11882 7344 11888 7396
rect 11940 7384 11946 7396
rect 17954 7384 17960 7396
rect 11940 7356 13216 7384
rect 11940 7344 11946 7356
rect 8294 7208 8300 7260
rect 8352 7248 8358 7260
rect 9861 7251 9919 7257
rect 9861 7248 9873 7251
rect 8352 7220 9873 7248
rect 8352 7208 8358 7220
rect 9861 7217 9873 7220
rect 9907 7217 9919 7251
rect 11716 7248 11744 7344
rect 11716 7220 12020 7248
rect 9861 7211 9919 7217
rect 11885 7183 11943 7189
rect 11885 7149 11897 7183
rect 11931 7149 11943 7183
rect 11992 7180 12020 7220
rect 12141 7183 12199 7189
rect 12141 7180 12153 7183
rect 11992 7152 12153 7180
rect 11885 7143 11943 7149
rect 12141 7149 12153 7152
rect 12187 7149 12199 7183
rect 13188 7180 13216 7356
rect 17052 7356 17960 7384
rect 13265 7319 13323 7325
rect 13265 7285 13277 7319
rect 13311 7285 13323 7319
rect 13265 7279 13323 7285
rect 13280 7248 13308 7279
rect 13722 7276 13728 7328
rect 13780 7316 13786 7328
rect 13780 7288 15424 7316
rect 13780 7276 13786 7288
rect 13906 7248 13912 7260
rect 13280 7220 13912 7248
rect 13906 7208 13912 7220
rect 13964 7248 13970 7260
rect 15396 7257 15424 7288
rect 14737 7251 14795 7257
rect 14737 7248 14749 7251
rect 13964 7220 14749 7248
rect 13964 7208 13970 7220
rect 14737 7217 14749 7220
rect 14783 7217 14795 7251
rect 14737 7211 14795 7217
rect 15381 7251 15439 7257
rect 15381 7217 15393 7251
rect 15427 7217 15439 7251
rect 15381 7211 15439 7217
rect 14553 7183 14611 7189
rect 13188 7152 13952 7180
rect 12141 7143 12199 7149
rect 10134 7121 10140 7124
rect 10128 7112 10140 7121
rect 10095 7084 10140 7112
rect 10128 7075 10140 7084
rect 10134 7072 10140 7075
rect 10192 7072 10198 7124
rect 11900 7044 11928 7143
rect 12986 7112 12992 7124
rect 12360 7084 12992 7112
rect 12360 7044 12388 7084
rect 12986 7072 12992 7084
rect 13044 7072 13050 7124
rect 13924 7121 13952 7152
rect 14553 7149 14565 7183
rect 14599 7180 14611 7183
rect 15194 7180 15200 7192
rect 14599 7152 15200 7180
rect 14599 7149 14611 7152
rect 14553 7143 14611 7149
rect 15194 7140 15200 7152
rect 15252 7140 15258 7192
rect 15396 7180 15424 7211
rect 17052 7189 17080 7356
rect 17954 7344 17960 7356
rect 18012 7344 18018 7396
rect 18138 7344 18144 7396
rect 18196 7384 18202 7396
rect 18417 7387 18475 7393
rect 18417 7384 18429 7387
rect 18196 7356 18429 7384
rect 18196 7344 18202 7356
rect 18417 7353 18429 7356
rect 18463 7353 18475 7387
rect 18417 7347 18475 7353
rect 18598 7344 18604 7396
rect 18656 7384 18662 7396
rect 18693 7387 18751 7393
rect 18693 7384 18705 7387
rect 18656 7356 18705 7384
rect 18656 7344 18662 7356
rect 18693 7353 18705 7356
rect 18739 7353 18751 7387
rect 21082 7384 21088 7396
rect 21043 7356 21088 7384
rect 18693 7347 18751 7353
rect 21082 7344 21088 7356
rect 21140 7344 21146 7396
rect 18966 7208 18972 7260
rect 19024 7248 19030 7260
rect 19153 7251 19211 7257
rect 19153 7248 19165 7251
rect 19024 7220 19165 7248
rect 19024 7208 19030 7220
rect 19153 7217 19165 7220
rect 19199 7217 19211 7251
rect 19153 7211 19211 7217
rect 19245 7251 19303 7257
rect 19245 7217 19257 7251
rect 19291 7217 19303 7251
rect 19245 7211 19303 7217
rect 17037 7183 17095 7189
rect 17037 7180 17049 7183
rect 15396 7152 17049 7180
rect 17037 7149 17049 7152
rect 17083 7149 17095 7183
rect 17304 7183 17362 7189
rect 17304 7180 17316 7183
rect 17037 7143 17095 7149
rect 17236 7152 17316 7180
rect 13909 7115 13967 7121
rect 13909 7081 13921 7115
rect 13955 7112 13967 7115
rect 13955 7084 14688 7112
rect 13955 7081 13967 7084
rect 13909 7075 13967 7081
rect 14182 7044 14188 7056
rect 11900 7016 12388 7044
rect 14143 7016 14188 7044
rect 14182 7004 14188 7016
rect 14240 7004 14246 7056
rect 14660 7053 14688 7084
rect 14734 7072 14740 7124
rect 14792 7112 14798 7124
rect 15010 7112 15016 7124
rect 14792 7084 15016 7112
rect 14792 7072 14798 7084
rect 15010 7072 15016 7084
rect 15068 7112 15074 7124
rect 15626 7115 15684 7121
rect 15626 7112 15638 7115
rect 15068 7084 15638 7112
rect 15068 7072 15074 7084
rect 15626 7081 15638 7084
rect 15672 7081 15684 7115
rect 15626 7075 15684 7081
rect 14645 7047 14703 7053
rect 14645 7013 14657 7047
rect 14691 7044 14703 7047
rect 15378 7044 15384 7056
rect 14691 7016 15384 7044
rect 14691 7013 14703 7016
rect 14645 7007 14703 7013
rect 15378 7004 15384 7016
rect 15436 7004 15442 7056
rect 16761 7047 16819 7053
rect 16761 7013 16773 7047
rect 16807 7044 16819 7047
rect 17236 7044 17264 7152
rect 17304 7149 17316 7152
rect 17350 7180 17362 7183
rect 19260 7180 19288 7211
rect 17350 7152 19288 7180
rect 20533 7183 20591 7189
rect 17350 7149 17362 7152
rect 17304 7143 17362 7149
rect 20533 7149 20545 7183
rect 20579 7180 20591 7183
rect 20898 7180 20904 7192
rect 20579 7152 20904 7180
rect 20579 7149 20591 7152
rect 20533 7143 20591 7149
rect 20898 7140 20904 7152
rect 20956 7140 20962 7192
rect 19061 7115 19119 7121
rect 19061 7081 19073 7115
rect 19107 7112 19119 7115
rect 19107 7084 19288 7112
rect 19107 7081 19119 7084
rect 19061 7075 19119 7081
rect 19260 7056 19288 7084
rect 16807 7016 17264 7044
rect 16807 7013 16819 7016
rect 16761 7007 16819 7013
rect 19242 7004 19248 7056
rect 19300 7044 19306 7056
rect 19705 7047 19763 7053
rect 19705 7044 19717 7047
rect 19300 7016 19717 7044
rect 19300 7004 19306 7016
rect 19705 7013 19717 7016
rect 19751 7013 19763 7047
rect 19705 7007 19763 7013
rect 1104 6954 21896 6976
rect 1104 6902 7912 6954
rect 7964 6902 7976 6954
rect 8028 6902 8040 6954
rect 8092 6902 8104 6954
rect 8156 6902 14843 6954
rect 14895 6902 14907 6954
rect 14959 6902 14971 6954
rect 15023 6902 15035 6954
rect 15087 6902 21896 6954
rect 1104 6880 21896 6902
rect 11238 6800 11244 6852
rect 11296 6840 11302 6852
rect 11333 6843 11391 6849
rect 11333 6840 11345 6843
rect 11296 6812 11345 6840
rect 11296 6800 11302 6812
rect 11333 6809 11345 6812
rect 11379 6809 11391 6843
rect 11793 6843 11851 6849
rect 11793 6840 11805 6843
rect 11333 6803 11391 6809
rect 11624 6812 11805 6840
rect 8645 6707 8703 6713
rect 8645 6704 8657 6707
rect 8036 6676 8657 6704
rect 4062 6460 4068 6512
rect 4120 6500 4126 6512
rect 8036 6509 8064 6676
rect 8645 6673 8657 6676
rect 8691 6673 8703 6707
rect 8645 6667 8703 6673
rect 11057 6707 11115 6713
rect 11057 6673 11069 6707
rect 11103 6704 11115 6707
rect 11624 6704 11652 6812
rect 11793 6809 11805 6812
rect 11839 6840 11851 6843
rect 11882 6840 11888 6852
rect 11839 6812 11888 6840
rect 11839 6809 11851 6812
rect 11793 6803 11851 6809
rect 11882 6800 11888 6812
rect 11940 6800 11946 6852
rect 14182 6800 14188 6852
rect 14240 6840 14246 6852
rect 14645 6843 14703 6849
rect 14645 6840 14657 6843
rect 14240 6812 14657 6840
rect 14240 6800 14246 6812
rect 14645 6809 14657 6812
rect 14691 6809 14703 6843
rect 14645 6803 14703 6809
rect 15378 6800 15384 6852
rect 15436 6840 15442 6852
rect 18601 6843 18659 6849
rect 18601 6840 18613 6843
rect 15436 6812 18613 6840
rect 15436 6800 15442 6812
rect 18601 6809 18613 6812
rect 18647 6840 18659 6843
rect 18966 6840 18972 6852
rect 18647 6812 18972 6840
rect 18647 6809 18659 6812
rect 18601 6803 18659 6809
rect 18966 6800 18972 6812
rect 19024 6800 19030 6852
rect 11701 6775 11759 6781
rect 11701 6741 11713 6775
rect 11747 6772 11759 6775
rect 12526 6772 12532 6784
rect 11747 6744 12532 6772
rect 11747 6741 11759 6744
rect 11701 6735 11759 6741
rect 12526 6732 12532 6744
rect 12584 6732 12590 6784
rect 14553 6775 14611 6781
rect 14553 6741 14565 6775
rect 14599 6772 14611 6775
rect 15286 6772 15292 6784
rect 14599 6744 15292 6772
rect 14599 6741 14611 6744
rect 14553 6735 14611 6741
rect 15286 6732 15292 6744
rect 15344 6732 15350 6784
rect 18046 6704 18052 6716
rect 11103 6676 11652 6704
rect 18007 6676 18052 6704
rect 11103 6673 11115 6676
rect 11057 6667 11115 6673
rect 18046 6664 18052 6676
rect 18104 6664 18110 6716
rect 8294 6596 8300 6648
rect 8352 6636 8358 6648
rect 8389 6639 8447 6645
rect 8389 6636 8401 6639
rect 8352 6608 8401 6636
rect 8352 6596 8358 6608
rect 8389 6605 8401 6608
rect 8435 6605 8447 6639
rect 8389 6599 8447 6605
rect 11885 6639 11943 6645
rect 11885 6605 11897 6639
rect 11931 6605 11943 6639
rect 14734 6636 14740 6648
rect 14695 6608 14740 6636
rect 11885 6599 11943 6605
rect 9769 6571 9827 6577
rect 9769 6537 9781 6571
rect 9815 6568 9827 6571
rect 10134 6568 10140 6580
rect 9815 6540 10140 6568
rect 9815 6537 9827 6540
rect 9769 6531 9827 6537
rect 10134 6528 10140 6540
rect 10192 6568 10198 6580
rect 11900 6568 11928 6599
rect 14734 6596 14740 6608
rect 14792 6596 14798 6648
rect 10192 6540 11928 6568
rect 10192 6528 10198 6540
rect 14090 6528 14096 6580
rect 14148 6568 14154 6580
rect 14185 6571 14243 6577
rect 14185 6568 14197 6571
rect 14148 6540 14197 6568
rect 14148 6528 14154 6540
rect 14185 6537 14197 6540
rect 14231 6537 14243 6571
rect 14185 6531 14243 6537
rect 8021 6503 8079 6509
rect 8021 6500 8033 6503
rect 4120 6472 8033 6500
rect 4120 6460 4126 6472
rect 8021 6469 8033 6472
rect 8067 6469 8079 6503
rect 12526 6500 12532 6512
rect 12487 6472 12532 6500
rect 8021 6463 8079 6469
rect 12526 6460 12532 6472
rect 12584 6460 12590 6512
rect 15194 6460 15200 6512
rect 15252 6500 15258 6512
rect 15289 6503 15347 6509
rect 15289 6500 15301 6503
rect 15252 6472 15301 6500
rect 15252 6460 15258 6472
rect 15289 6469 15301 6472
rect 15335 6500 15347 6503
rect 17954 6500 17960 6512
rect 15335 6472 17960 6500
rect 15335 6469 15347 6472
rect 15289 6463 15347 6469
rect 17954 6460 17960 6472
rect 18012 6460 18018 6512
rect 21358 6500 21364 6512
rect 21319 6472 21364 6500
rect 21358 6460 21364 6472
rect 21416 6460 21422 6512
rect 1104 6410 21896 6432
rect 1104 6358 4447 6410
rect 4499 6358 4511 6410
rect 4563 6358 4575 6410
rect 4627 6358 4639 6410
rect 4691 6358 11378 6410
rect 11430 6358 11442 6410
rect 11494 6358 11506 6410
rect 11558 6358 11570 6410
rect 11622 6358 18308 6410
rect 18360 6358 18372 6410
rect 18424 6358 18436 6410
rect 18488 6358 18500 6410
rect 18552 6358 21896 6410
rect 1104 6336 21896 6358
rect 12894 6256 12900 6308
rect 12952 6296 12958 6308
rect 21085 6299 21143 6305
rect 21085 6296 21097 6299
rect 12952 6268 21097 6296
rect 12952 6256 12958 6268
rect 21085 6265 21097 6268
rect 21131 6265 21143 6299
rect 21085 6259 21143 6265
rect 20901 6095 20959 6101
rect 20901 6061 20913 6095
rect 20947 6092 20959 6095
rect 21358 6092 21364 6104
rect 20947 6064 21364 6092
rect 20947 6061 20959 6064
rect 20901 6055 20959 6061
rect 21358 6052 21364 6064
rect 21416 6052 21422 6104
rect 1104 5866 21896 5888
rect 1104 5814 7912 5866
rect 7964 5814 7976 5866
rect 8028 5814 8040 5866
rect 8092 5814 8104 5866
rect 8156 5814 14843 5866
rect 14895 5814 14907 5866
rect 14959 5814 14971 5866
rect 15023 5814 15035 5866
rect 15087 5814 21896 5866
rect 1104 5792 21896 5814
rect 12618 5712 12624 5764
rect 12676 5752 12682 5764
rect 20993 5755 21051 5761
rect 20993 5752 21005 5755
rect 12676 5724 21005 5752
rect 12676 5712 12682 5724
rect 20993 5721 21005 5724
rect 21039 5721 21051 5755
rect 20993 5715 21051 5721
rect 20809 5619 20867 5625
rect 20809 5585 20821 5619
rect 20855 5616 20867 5619
rect 21266 5616 21272 5628
rect 20855 5588 21272 5616
rect 20855 5585 20867 5588
rect 20809 5579 20867 5585
rect 21266 5576 21272 5588
rect 21324 5576 21330 5628
rect 1104 5322 21896 5344
rect 1104 5270 4447 5322
rect 4499 5270 4511 5322
rect 4563 5270 4575 5322
rect 4627 5270 4639 5322
rect 4691 5270 11378 5322
rect 11430 5270 11442 5322
rect 11494 5270 11506 5322
rect 11558 5270 11570 5322
rect 11622 5270 18308 5322
rect 18360 5270 18372 5322
rect 18424 5270 18436 5322
rect 18488 5270 18500 5322
rect 18552 5270 21896 5322
rect 1104 5248 21896 5270
rect 12526 5168 12532 5220
rect 12584 5208 12590 5220
rect 17954 5208 17960 5220
rect 12584 5180 17960 5208
rect 12584 5168 12590 5180
rect 17954 5168 17960 5180
rect 18012 5168 18018 5220
rect 21266 5140 21272 5152
rect 21227 5112 21272 5140
rect 21266 5100 21272 5112
rect 21324 5100 21330 5152
rect 1104 4778 21896 4800
rect 1104 4726 7912 4778
rect 7964 4726 7976 4778
rect 8028 4726 8040 4778
rect 8092 4726 8104 4778
rect 8156 4726 14843 4778
rect 14895 4726 14907 4778
rect 14959 4726 14971 4778
rect 15023 4726 15035 4778
rect 15087 4726 21896 4778
rect 1104 4704 21896 4726
rect 20990 4664 20996 4676
rect 20951 4636 20996 4664
rect 20990 4624 20996 4636
rect 21048 4624 21054 4676
rect 20809 4531 20867 4537
rect 20809 4497 20821 4531
rect 20855 4528 20867 4531
rect 21266 4528 21272 4540
rect 20855 4500 21272 4528
rect 20855 4497 20867 4500
rect 20809 4491 20867 4497
rect 21266 4488 21272 4500
rect 21324 4488 21330 4540
rect 1104 4234 21896 4256
rect 1104 4182 4447 4234
rect 4499 4182 4511 4234
rect 4563 4182 4575 4234
rect 4627 4182 4639 4234
rect 4691 4182 11378 4234
rect 11430 4182 11442 4234
rect 11494 4182 11506 4234
rect 11558 4182 11570 4234
rect 11622 4182 18308 4234
rect 18360 4182 18372 4234
rect 18424 4182 18436 4234
rect 18488 4182 18500 4234
rect 18552 4182 21896 4234
rect 1104 4160 21896 4182
rect 21266 4120 21272 4132
rect 21227 4092 21272 4120
rect 21266 4080 21272 4092
rect 21324 4080 21330 4132
rect 16482 3944 16488 3996
rect 16540 3984 16546 3996
rect 18782 3984 18788 3996
rect 16540 3956 18788 3984
rect 16540 3944 16546 3956
rect 18782 3944 18788 3956
rect 18840 3944 18846 3996
rect 1104 3690 21896 3712
rect 1104 3638 7912 3690
rect 7964 3638 7976 3690
rect 8028 3638 8040 3690
rect 8092 3638 8104 3690
rect 8156 3638 14843 3690
rect 14895 3638 14907 3690
rect 14959 3638 14971 3690
rect 15023 3638 15035 3690
rect 15087 3638 21896 3690
rect 1104 3616 21896 3638
rect 1104 3146 21896 3168
rect 1104 3094 4447 3146
rect 4499 3094 4511 3146
rect 4563 3094 4575 3146
rect 4627 3094 4639 3146
rect 4691 3094 11378 3146
rect 11430 3094 11442 3146
rect 11494 3094 11506 3146
rect 11558 3094 11570 3146
rect 11622 3094 18308 3146
rect 18360 3094 18372 3146
rect 18424 3094 18436 3146
rect 18488 3094 18500 3146
rect 18552 3094 21896 3146
rect 1104 3072 21896 3094
rect 18690 2924 18696 2976
rect 18748 2964 18754 2976
rect 18874 2964 18880 2976
rect 18748 2936 18880 2964
rect 18748 2924 18754 2936
rect 18874 2924 18880 2936
rect 18932 2924 18938 2976
rect 1104 2602 21896 2624
rect 1104 2550 7912 2602
rect 7964 2550 7976 2602
rect 8028 2550 8040 2602
rect 8092 2550 8104 2602
rect 8156 2550 14843 2602
rect 14895 2550 14907 2602
rect 14959 2550 14971 2602
rect 15023 2550 15035 2602
rect 15087 2550 21896 2602
rect 1104 2528 21896 2550
rect 14274 2380 14280 2432
rect 14332 2420 14338 2432
rect 18138 2420 18144 2432
rect 14332 2392 18144 2420
rect 14332 2380 14338 2392
rect 18138 2380 18144 2392
rect 18196 2380 18202 2432
rect 1104 2058 21896 2080
rect 1104 2006 4447 2058
rect 4499 2006 4511 2058
rect 4563 2006 4575 2058
rect 4627 2006 4639 2058
rect 4691 2006 11378 2058
rect 11430 2006 11442 2058
rect 11494 2006 11506 2058
rect 11558 2006 11570 2058
rect 11622 2006 18308 2058
rect 18360 2006 18372 2058
rect 18424 2006 18436 2058
rect 18488 2006 18500 2058
rect 18552 2006 21896 2058
rect 1104 1984 21896 2006
rect 13998 1904 14004 1956
rect 14056 1944 14062 1956
rect 18138 1944 18144 1956
rect 14056 1916 18144 1944
rect 14056 1904 14062 1916
rect 18138 1904 18144 1916
rect 18196 1904 18202 1956
rect 14550 1156 14556 1208
rect 14608 1196 14614 1208
rect 17954 1196 17960 1208
rect 14608 1168 17960 1196
rect 14608 1156 14614 1168
rect 17954 1156 17960 1168
rect 18012 1156 18018 1208
<< via1 >>
rect 4447 20502 4499 20554
rect 4511 20502 4563 20554
rect 4575 20502 4627 20554
rect 4639 20502 4691 20554
rect 11378 20502 11430 20554
rect 11442 20502 11494 20554
rect 11506 20502 11558 20554
rect 11570 20502 11622 20554
rect 18308 20502 18360 20554
rect 18372 20502 18424 20554
rect 18436 20502 18488 20554
rect 18500 20502 18552 20554
rect 20168 20443 20220 20452
rect 20168 20409 20177 20443
rect 20177 20409 20211 20443
rect 20211 20409 20220 20443
rect 20168 20400 20220 20409
rect 20536 20400 20588 20452
rect 19984 20239 20036 20248
rect 19984 20205 19993 20239
rect 19993 20205 20027 20239
rect 20027 20205 20036 20239
rect 19984 20196 20036 20205
rect 20076 20196 20128 20248
rect 7912 19958 7964 20010
rect 7976 19958 8028 20010
rect 8040 19958 8092 20010
rect 8104 19958 8156 20010
rect 14843 19958 14895 20010
rect 14907 19958 14959 20010
rect 14971 19958 15023 20010
rect 15035 19958 15087 20010
rect 18604 19856 18656 19908
rect 19248 19856 19300 19908
rect 20628 19856 20680 19908
rect 20076 19831 20128 19840
rect 4896 19720 4948 19772
rect 6552 19720 6604 19772
rect 6828 19763 6880 19772
rect 6828 19729 6837 19763
rect 6837 19729 6871 19763
rect 6871 19729 6880 19763
rect 6828 19720 6880 19729
rect 20076 19797 20085 19831
rect 20085 19797 20119 19831
rect 20119 19797 20128 19831
rect 20076 19788 20128 19797
rect 8300 19763 8352 19772
rect 8300 19729 8334 19763
rect 8334 19729 8352 19763
rect 8300 19720 8352 19729
rect 14188 19720 14240 19772
rect 18052 19763 18104 19772
rect 18052 19729 18061 19763
rect 18061 19729 18095 19763
rect 18095 19729 18104 19763
rect 18052 19720 18104 19729
rect 18144 19720 18196 19772
rect 20168 19720 20220 19772
rect 7748 19652 7800 19704
rect 9680 19695 9732 19704
rect 9680 19661 9689 19695
rect 9689 19661 9723 19695
rect 9723 19661 9732 19695
rect 9680 19652 9732 19661
rect 14740 19584 14792 19636
rect 16396 19584 16448 19636
rect 6276 19516 6328 19568
rect 10232 19516 10284 19568
rect 14004 19559 14056 19568
rect 14004 19525 14013 19559
rect 14013 19525 14047 19559
rect 14047 19525 14056 19559
rect 14004 19516 14056 19525
rect 17040 19516 17092 19568
rect 4447 19414 4499 19466
rect 4511 19414 4563 19466
rect 4575 19414 4627 19466
rect 4639 19414 4691 19466
rect 11378 19414 11430 19466
rect 11442 19414 11494 19466
rect 11506 19414 11558 19466
rect 11570 19414 11622 19466
rect 18308 19414 18360 19466
rect 18372 19414 18424 19466
rect 18436 19414 18488 19466
rect 18500 19414 18552 19466
rect 20444 19355 20496 19364
rect 20444 19321 20453 19355
rect 20453 19321 20487 19355
rect 20487 19321 20496 19355
rect 20444 19312 20496 19321
rect 21088 19355 21140 19364
rect 21088 19321 21097 19355
rect 21097 19321 21131 19355
rect 21131 19321 21140 19355
rect 21088 19312 21140 19321
rect 8300 19176 8352 19228
rect 1952 19108 2004 19160
rect 3884 19108 3936 19160
rect 2504 19040 2556 19092
rect 3976 19040 4028 19092
rect 2412 18972 2464 19024
rect 4896 19108 4948 19160
rect 6276 19108 6328 19160
rect 8668 19108 8720 19160
rect 4252 19040 4304 19092
rect 9956 19176 10008 19228
rect 10232 19219 10284 19228
rect 10232 19185 10241 19219
rect 10241 19185 10275 19219
rect 10275 19185 10284 19219
rect 10232 19176 10284 19185
rect 9680 19108 9732 19160
rect 10140 19108 10192 19160
rect 11060 19151 11112 19160
rect 11060 19117 11069 19151
rect 11069 19117 11103 19151
rect 11103 19117 11112 19151
rect 11060 19108 11112 19117
rect 12532 19108 12584 19160
rect 12992 19151 13044 19160
rect 12992 19117 13015 19151
rect 13015 19117 13044 19151
rect 5448 19015 5500 19024
rect 5448 18981 5457 19015
rect 5457 18981 5491 19015
rect 5491 18981 5500 19015
rect 5448 18972 5500 18981
rect 8300 18972 8352 19024
rect 8760 19015 8812 19024
rect 8760 18981 8769 19015
rect 8769 18981 8803 19015
rect 8803 18981 8812 19015
rect 8760 18972 8812 18981
rect 11152 19040 11204 19092
rect 11612 19040 11664 19092
rect 12992 19108 13044 19117
rect 17040 19151 17092 19160
rect 17040 19117 17049 19151
rect 17049 19117 17083 19151
rect 17083 19117 17092 19151
rect 17040 19108 17092 19117
rect 18052 19108 18104 19160
rect 19248 19176 19300 19228
rect 18328 19108 18380 19160
rect 13544 19040 13596 19092
rect 14740 19040 14792 19092
rect 19064 19083 19116 19092
rect 19064 19049 19073 19083
rect 19073 19049 19107 19083
rect 19107 19049 19116 19083
rect 19064 19040 19116 19049
rect 10416 18972 10468 19024
rect 10968 18972 11020 19024
rect 12532 18972 12584 19024
rect 12900 18972 12952 19024
rect 14096 19015 14148 19024
rect 14096 18981 14105 19015
rect 14105 18981 14139 19015
rect 14139 18981 14148 19015
rect 14096 18972 14148 18981
rect 16396 18972 16448 19024
rect 16764 18972 16816 19024
rect 7912 18870 7964 18922
rect 7976 18870 8028 18922
rect 8040 18870 8092 18922
rect 8104 18870 8156 18922
rect 14843 18870 14895 18922
rect 14907 18870 14959 18922
rect 14971 18870 15023 18922
rect 15035 18870 15087 18922
rect 4160 18768 4212 18820
rect 6828 18811 6880 18820
rect 6828 18777 6837 18811
rect 6837 18777 6871 18811
rect 6871 18777 6880 18811
rect 6828 18768 6880 18777
rect 5816 18700 5868 18752
rect 8576 18768 8628 18820
rect 8668 18768 8720 18820
rect 10140 18768 10192 18820
rect 7012 18700 7064 18752
rect 11428 18768 11480 18820
rect 11612 18811 11664 18820
rect 11612 18777 11621 18811
rect 11621 18777 11655 18811
rect 11655 18777 11664 18811
rect 11612 18768 11664 18777
rect 14740 18768 14792 18820
rect 20996 18811 21048 18820
rect 3148 18632 3200 18684
rect 1768 18564 1820 18616
rect 2412 18607 2464 18616
rect 2412 18573 2421 18607
rect 2421 18573 2455 18607
rect 2455 18573 2464 18607
rect 2412 18564 2464 18573
rect 4252 18496 4304 18548
rect 4344 18428 4396 18480
rect 8760 18632 8812 18684
rect 10968 18632 11020 18684
rect 12440 18632 12492 18684
rect 12716 18632 12768 18684
rect 14096 18700 14148 18752
rect 16764 18700 16816 18752
rect 17132 18700 17184 18752
rect 18420 18743 18472 18752
rect 14280 18632 14332 18684
rect 15660 18632 15712 18684
rect 16856 18675 16908 18684
rect 16856 18641 16865 18675
rect 16865 18641 16899 18675
rect 16899 18641 16908 18675
rect 16856 18632 16908 18641
rect 18420 18709 18429 18743
rect 18429 18709 18463 18743
rect 18463 18709 18472 18743
rect 18420 18700 18472 18709
rect 19984 18700 20036 18752
rect 20168 18743 20220 18752
rect 20168 18709 20177 18743
rect 20177 18709 20211 18743
rect 20211 18709 20220 18743
rect 20168 18700 20220 18709
rect 20996 18777 21005 18811
rect 21005 18777 21039 18811
rect 21039 18777 21048 18811
rect 20996 18768 21048 18777
rect 21732 18700 21784 18752
rect 6644 18564 6696 18616
rect 6276 18496 6328 18548
rect 9680 18564 9732 18616
rect 10140 18564 10192 18616
rect 9772 18428 9824 18480
rect 12992 18607 13044 18616
rect 12992 18573 13001 18607
rect 13001 18573 13035 18607
rect 13035 18573 13044 18607
rect 13544 18607 13596 18616
rect 12992 18564 13044 18573
rect 13544 18573 13553 18607
rect 13553 18573 13587 18607
rect 13587 18573 13596 18607
rect 13544 18564 13596 18573
rect 13912 18428 13964 18480
rect 15476 18428 15528 18480
rect 17040 18607 17092 18616
rect 17040 18573 17049 18607
rect 17049 18573 17083 18607
rect 17083 18573 17092 18607
rect 18604 18607 18656 18616
rect 17040 18564 17092 18573
rect 18604 18573 18613 18607
rect 18613 18573 18647 18607
rect 18647 18573 18656 18607
rect 18604 18564 18656 18573
rect 16212 18496 16264 18548
rect 20812 18675 20864 18684
rect 20812 18641 20821 18675
rect 20821 18641 20855 18675
rect 20855 18641 20864 18675
rect 20812 18632 20864 18641
rect 4447 18326 4499 18378
rect 4511 18326 4563 18378
rect 4575 18326 4627 18378
rect 4639 18326 4691 18378
rect 11378 18326 11430 18378
rect 11442 18326 11494 18378
rect 11506 18326 11558 18378
rect 11570 18326 11622 18378
rect 18308 18326 18360 18378
rect 18372 18326 18424 18378
rect 18436 18326 18488 18378
rect 18500 18326 18552 18378
rect 296 18156 348 18208
rect 6368 18224 6420 18276
rect 6644 18267 6696 18276
rect 6644 18233 6653 18267
rect 6653 18233 6687 18267
rect 6687 18233 6696 18267
rect 6644 18224 6696 18233
rect 5264 18156 5316 18208
rect 8208 18224 8260 18276
rect 1400 18088 1452 18140
rect 6644 18088 6696 18140
rect 7932 18156 7984 18208
rect 10968 18224 11020 18276
rect 12440 18224 12492 18276
rect 12532 18224 12584 18276
rect 15292 18224 15344 18276
rect 16212 18224 16264 18276
rect 17040 18224 17092 18276
rect 17868 18224 17920 18276
rect 21640 18224 21692 18276
rect 6552 18020 6604 18072
rect 11704 18088 11756 18140
rect 13912 18131 13964 18140
rect 13912 18097 13921 18131
rect 13921 18097 13955 18131
rect 13955 18097 13964 18131
rect 13912 18088 13964 18097
rect 14096 18131 14148 18140
rect 14096 18097 14105 18131
rect 14105 18097 14139 18131
rect 14139 18097 14148 18131
rect 14096 18088 14148 18097
rect 18696 18156 18748 18208
rect 21456 18156 21508 18208
rect 18880 18131 18932 18140
rect 9680 18063 9732 18072
rect 9680 18029 9689 18063
rect 9689 18029 9723 18063
rect 9723 18029 9732 18063
rect 9680 18020 9732 18029
rect 9772 18020 9824 18072
rect 9956 18063 10008 18072
rect 9956 18029 9990 18063
rect 9990 18029 10008 18063
rect 9956 18020 10008 18029
rect 10876 18020 10928 18072
rect 15476 18020 15528 18072
rect 6460 17952 6512 18004
rect 11244 17952 11296 18004
rect 12900 17952 12952 18004
rect 13728 17952 13780 18004
rect 14740 17952 14792 18004
rect 16396 18020 16448 18072
rect 17224 18063 17276 18072
rect 17224 18029 17233 18063
rect 17233 18029 17267 18063
rect 17267 18029 17276 18063
rect 17224 18020 17276 18029
rect 18880 18097 18889 18131
rect 18889 18097 18923 18131
rect 18923 18097 18932 18131
rect 18880 18088 18932 18097
rect 20168 18088 20220 18140
rect 21548 18088 21600 18140
rect 20076 18020 20128 18072
rect 18144 17952 18196 18004
rect 18788 17952 18840 18004
rect 19616 17952 19668 18004
rect 20536 17952 20588 18004
rect 22100 17952 22152 18004
rect 3056 17884 3108 17936
rect 4160 17884 4212 17936
rect 4804 17884 4856 17936
rect 6736 17884 6788 17936
rect 7472 17884 7524 17936
rect 8576 17884 8628 17936
rect 11152 17884 11204 17936
rect 11796 17927 11848 17936
rect 11796 17893 11805 17927
rect 11805 17893 11839 17927
rect 11839 17893 11848 17927
rect 11796 17884 11848 17893
rect 11888 17884 11940 17936
rect 12532 17884 12584 17936
rect 12716 17884 12768 17936
rect 15384 17884 15436 17936
rect 15844 17884 15896 17936
rect 18604 17927 18656 17936
rect 18604 17893 18613 17927
rect 18613 17893 18647 17927
rect 18647 17893 18656 17927
rect 18604 17884 18656 17893
rect 19800 17884 19852 17936
rect 20352 17884 20404 17936
rect 21088 17927 21140 17936
rect 21088 17893 21097 17927
rect 21097 17893 21131 17927
rect 21131 17893 21140 17927
rect 21088 17884 21140 17893
rect 21180 17884 21232 17936
rect 22652 17884 22704 17936
rect 7912 17782 7964 17834
rect 7976 17782 8028 17834
rect 8040 17782 8092 17834
rect 8104 17782 8156 17834
rect 14843 17782 14895 17834
rect 14907 17782 14959 17834
rect 14971 17782 15023 17834
rect 15035 17782 15087 17834
rect 4344 17680 4396 17732
rect 9220 17680 9272 17732
rect 11796 17680 11848 17732
rect 12532 17680 12584 17732
rect 15200 17680 15252 17732
rect 19524 17723 19576 17732
rect 19524 17689 19533 17723
rect 19533 17689 19567 17723
rect 19567 17689 19576 17723
rect 19524 17680 19576 17689
rect 4344 17544 4396 17596
rect 9864 17544 9916 17596
rect 5448 17476 5500 17528
rect 10968 17476 11020 17528
rect 18604 17544 18656 17596
rect 18880 17544 18932 17596
rect 20720 17544 20772 17596
rect 4804 17408 4856 17460
rect 4252 17383 4304 17392
rect 4252 17349 4261 17383
rect 4261 17349 4295 17383
rect 4295 17349 4304 17383
rect 4252 17340 4304 17349
rect 8944 17340 8996 17392
rect 20444 17451 20496 17460
rect 20444 17417 20453 17451
rect 20453 17417 20487 17451
rect 20487 17417 20496 17451
rect 20444 17408 20496 17417
rect 20996 17383 21048 17392
rect 20996 17349 21005 17383
rect 21005 17349 21039 17383
rect 21039 17349 21048 17383
rect 20996 17340 21048 17349
rect 4447 17238 4499 17290
rect 4511 17238 4563 17290
rect 4575 17238 4627 17290
rect 4639 17238 4691 17290
rect 11378 17238 11430 17290
rect 11442 17238 11494 17290
rect 11506 17238 11558 17290
rect 11570 17238 11622 17290
rect 18308 17238 18360 17290
rect 18372 17238 18424 17290
rect 18436 17238 18488 17290
rect 18500 17238 18552 17290
rect 3148 17179 3200 17188
rect 3148 17145 3157 17179
rect 3157 17145 3191 17179
rect 3191 17145 3200 17179
rect 3148 17136 3200 17145
rect 3332 17136 3384 17188
rect 3516 17136 3568 17188
rect 6736 17179 6788 17188
rect 6736 17145 6745 17179
rect 6745 17145 6779 17179
rect 6779 17145 6788 17179
rect 6736 17136 6788 17145
rect 19708 17136 19760 17188
rect 4344 17043 4396 17052
rect 4344 17009 4353 17043
rect 4353 17009 4387 17043
rect 4387 17009 4396 17043
rect 4344 17000 4396 17009
rect 9772 17068 9824 17120
rect 10968 17068 11020 17120
rect 20444 17068 20496 17120
rect 7012 17000 7064 17052
rect 8668 17043 8720 17052
rect 8668 17009 8677 17043
rect 8677 17009 8711 17043
rect 8711 17009 8720 17043
rect 8668 17000 8720 17009
rect 12164 17000 12216 17052
rect 14372 17000 14424 17052
rect 18880 17043 18932 17052
rect 1768 16975 1820 16984
rect 1768 16941 1777 16975
rect 1777 16941 1811 16975
rect 1811 16941 1820 16975
rect 1768 16932 1820 16941
rect 4896 16932 4948 16984
rect 5448 16932 5500 16984
rect 6736 16932 6788 16984
rect 3700 16864 3752 16916
rect 9864 16932 9916 16984
rect 10876 16932 10928 16984
rect 12716 16932 12768 16984
rect 15292 16932 15344 16984
rect 15752 16975 15804 16984
rect 15752 16941 15761 16975
rect 15761 16941 15795 16975
rect 15795 16941 15804 16975
rect 15752 16932 15804 16941
rect 18052 16932 18104 16984
rect 18880 17009 18889 17043
rect 18889 17009 18923 17043
rect 18923 17009 18932 17043
rect 18880 17000 18932 17009
rect 20076 17043 20128 17052
rect 20076 17009 20085 17043
rect 20085 17009 20119 17043
rect 20119 17009 20128 17043
rect 20076 17000 20128 17009
rect 10508 16864 10560 16916
rect 12532 16864 12584 16916
rect 3424 16839 3476 16848
rect 3424 16805 3433 16839
rect 3433 16805 3467 16839
rect 3467 16805 3476 16839
rect 3424 16796 3476 16805
rect 8392 16796 8444 16848
rect 11796 16839 11848 16848
rect 11796 16805 11805 16839
rect 11805 16805 11839 16839
rect 11839 16805 11848 16839
rect 11796 16796 11848 16805
rect 19340 16796 19392 16848
rect 19984 16796 20036 16848
rect 21088 16839 21140 16848
rect 21088 16805 21097 16839
rect 21097 16805 21131 16839
rect 21131 16805 21140 16839
rect 21088 16796 21140 16805
rect 7912 16694 7964 16746
rect 7976 16694 8028 16746
rect 8040 16694 8092 16746
rect 8104 16694 8156 16746
rect 14843 16694 14895 16746
rect 14907 16694 14959 16746
rect 14971 16694 15023 16746
rect 15035 16694 15087 16746
rect 3608 16635 3660 16644
rect 3608 16601 3617 16635
rect 3617 16601 3651 16635
rect 3651 16601 3660 16635
rect 3608 16592 3660 16601
rect 10508 16635 10560 16644
rect 7012 16524 7064 16576
rect 10508 16601 10517 16635
rect 10517 16601 10551 16635
rect 10551 16601 10560 16635
rect 10508 16592 10560 16601
rect 10876 16635 10928 16644
rect 10876 16601 10885 16635
rect 10885 16601 10919 16635
rect 10919 16601 10928 16635
rect 10876 16592 10928 16601
rect 10968 16635 11020 16644
rect 10968 16601 10977 16635
rect 10977 16601 11011 16635
rect 11011 16601 11020 16635
rect 11796 16635 11848 16644
rect 10968 16592 11020 16601
rect 11796 16601 11805 16635
rect 11805 16601 11839 16635
rect 11839 16601 11848 16635
rect 11796 16592 11848 16601
rect 18052 16635 18104 16644
rect 8668 16524 8720 16576
rect 4068 16456 4120 16508
rect 4252 16456 4304 16508
rect 12532 16524 12584 16576
rect 11152 16456 11204 16508
rect 15752 16524 15804 16576
rect 16856 16524 16908 16576
rect 14004 16499 14056 16508
rect 14004 16465 14013 16499
rect 14013 16465 14047 16499
rect 14047 16465 14056 16499
rect 14004 16456 14056 16465
rect 14372 16456 14424 16508
rect 16488 16456 16540 16508
rect 18052 16601 18061 16635
rect 18061 16601 18095 16635
rect 18095 16601 18104 16635
rect 18052 16592 18104 16601
rect 18604 16524 18656 16576
rect 20904 16524 20956 16576
rect 19708 16499 19760 16508
rect 19708 16465 19717 16499
rect 19717 16465 19751 16499
rect 19751 16465 19760 16499
rect 19708 16456 19760 16465
rect 20444 16499 20496 16508
rect 20444 16465 20453 16499
rect 20453 16465 20487 16499
rect 20487 16465 20496 16499
rect 20444 16456 20496 16465
rect 20720 16499 20772 16508
rect 20720 16465 20729 16499
rect 20729 16465 20763 16499
rect 20763 16465 20772 16499
rect 20720 16456 20772 16465
rect 3700 16431 3752 16440
rect 3700 16397 3709 16431
rect 3709 16397 3743 16431
rect 3743 16397 3752 16431
rect 3700 16388 3752 16397
rect 4896 16388 4948 16440
rect 6828 16431 6880 16440
rect 6828 16397 6837 16431
rect 6837 16397 6871 16431
rect 6871 16397 6880 16431
rect 6828 16388 6880 16397
rect 3148 16295 3200 16304
rect 3148 16261 3157 16295
rect 3157 16261 3191 16295
rect 3191 16261 3200 16295
rect 3148 16252 3200 16261
rect 6828 16252 6880 16304
rect 13268 16388 13320 16440
rect 14924 16431 14976 16440
rect 14924 16397 14933 16431
rect 14933 16397 14967 16431
rect 14967 16397 14976 16431
rect 14924 16388 14976 16397
rect 16672 16388 16724 16440
rect 18696 16431 18748 16440
rect 18696 16397 18705 16431
rect 18705 16397 18739 16431
rect 18739 16397 18748 16431
rect 18696 16388 18748 16397
rect 9680 16252 9732 16304
rect 10324 16252 10376 16304
rect 4447 16150 4499 16202
rect 4511 16150 4563 16202
rect 4575 16150 4627 16202
rect 4639 16150 4691 16202
rect 11378 16150 11430 16202
rect 11442 16150 11494 16202
rect 11506 16150 11558 16202
rect 11570 16150 11622 16202
rect 18308 16150 18360 16202
rect 18372 16150 18424 16202
rect 18436 16150 18488 16202
rect 18500 16150 18552 16202
rect 3516 16048 3568 16100
rect 6552 16091 6604 16100
rect 6552 16057 6561 16091
rect 6561 16057 6595 16091
rect 6595 16057 6604 16091
rect 6552 16048 6604 16057
rect 6828 16048 6880 16100
rect 13268 16091 13320 16100
rect 13268 16057 13277 16091
rect 13277 16057 13311 16091
rect 13311 16057 13320 16091
rect 13268 16048 13320 16057
rect 14924 16091 14976 16100
rect 14924 16057 14933 16091
rect 14933 16057 14967 16091
rect 14967 16057 14976 16091
rect 14924 16048 14976 16057
rect 16672 16091 16724 16100
rect 16672 16057 16681 16091
rect 16681 16057 16715 16091
rect 16715 16057 16724 16091
rect 16672 16048 16724 16057
rect 18696 16048 18748 16100
rect 21088 16091 21140 16100
rect 21088 16057 21097 16091
rect 21097 16057 21131 16091
rect 21131 16057 21140 16091
rect 21088 16048 21140 16057
rect 3148 15912 3200 15964
rect 3332 15955 3384 15964
rect 3332 15921 3341 15955
rect 3341 15921 3375 15955
rect 3375 15921 3384 15955
rect 3332 15912 3384 15921
rect 4896 15912 4948 15964
rect 7472 15912 7524 15964
rect 8944 15955 8996 15964
rect 8944 15921 8953 15955
rect 8953 15921 8987 15955
rect 8987 15921 8996 15955
rect 8944 15912 8996 15921
rect 9680 15912 9732 15964
rect 18604 15955 18656 15964
rect 4068 15844 4120 15896
rect 8208 15844 8260 15896
rect 8392 15844 8444 15896
rect 10324 15844 10376 15896
rect 13544 15887 13596 15896
rect 13544 15853 13553 15887
rect 13553 15853 13587 15887
rect 13587 15853 13596 15887
rect 13544 15844 13596 15853
rect 18604 15921 18613 15955
rect 18613 15921 18647 15955
rect 18647 15921 18656 15955
rect 18604 15912 18656 15921
rect 20904 15887 20956 15896
rect 3424 15776 3476 15828
rect 7748 15776 7800 15828
rect 12164 15819 12216 15828
rect 12164 15785 12198 15819
rect 12198 15785 12216 15819
rect 12164 15776 12216 15785
rect 14740 15776 14792 15828
rect 20904 15853 20913 15887
rect 20913 15853 20947 15887
rect 20947 15853 20956 15887
rect 20904 15844 20956 15853
rect 17316 15776 17368 15828
rect 7912 15606 7964 15658
rect 7976 15606 8028 15658
rect 8040 15606 8092 15658
rect 8104 15606 8156 15658
rect 14843 15606 14895 15658
rect 14907 15606 14959 15658
rect 14971 15606 15023 15658
rect 15035 15606 15087 15658
rect 3700 15504 3752 15556
rect 7656 15436 7708 15488
rect 18696 15436 18748 15488
rect 1768 15411 1820 15420
rect 1768 15377 1777 15411
rect 1777 15377 1811 15411
rect 1811 15377 1820 15411
rect 1768 15368 1820 15377
rect 4344 15368 4396 15420
rect 8116 15368 8168 15420
rect 17316 15368 17368 15420
rect 20812 15504 20864 15556
rect 20812 15411 20864 15420
rect 20812 15377 20821 15411
rect 20821 15377 20855 15411
rect 20855 15377 20864 15411
rect 20812 15368 20864 15377
rect 7656 15343 7708 15352
rect 7656 15309 7665 15343
rect 7665 15309 7699 15343
rect 7699 15309 7708 15343
rect 7656 15300 7708 15309
rect 7748 15343 7800 15352
rect 7748 15309 7757 15343
rect 7757 15309 7791 15343
rect 7791 15309 7800 15343
rect 7748 15300 7800 15309
rect 19432 15207 19484 15216
rect 19432 15173 19441 15207
rect 19441 15173 19475 15207
rect 19475 15173 19484 15207
rect 19432 15164 19484 15173
rect 20996 15207 21048 15216
rect 20996 15173 21005 15207
rect 21005 15173 21039 15207
rect 21039 15173 21048 15207
rect 20996 15164 21048 15173
rect 4447 15062 4499 15114
rect 4511 15062 4563 15114
rect 4575 15062 4627 15114
rect 4639 15062 4691 15114
rect 11378 15062 11430 15114
rect 11442 15062 11494 15114
rect 11506 15062 11558 15114
rect 11570 15062 11622 15114
rect 18308 15062 18360 15114
rect 18372 15062 18424 15114
rect 18436 15062 18488 15114
rect 18500 15062 18552 15114
rect 7656 14960 7708 15012
rect 4344 14824 4396 14876
rect 7656 14867 7708 14876
rect 7656 14833 7665 14867
rect 7665 14833 7699 14867
rect 7699 14833 7708 14867
rect 7656 14824 7708 14833
rect 8116 14867 8168 14876
rect 8116 14833 8125 14867
rect 8125 14833 8159 14867
rect 8159 14833 8168 14867
rect 8116 14824 8168 14833
rect 3884 14756 3936 14808
rect 7380 14756 7432 14808
rect 7564 14799 7616 14808
rect 7564 14765 7573 14799
rect 7573 14765 7607 14799
rect 7607 14765 7616 14799
rect 7564 14756 7616 14765
rect 10140 14824 10192 14876
rect 20812 14824 20864 14876
rect 8392 14688 8444 14740
rect 10968 14688 11020 14740
rect 16580 14688 16632 14740
rect 20812 14688 20864 14740
rect 4712 14620 4764 14672
rect 8208 14620 8260 14672
rect 12808 14620 12860 14672
rect 14556 14620 14608 14672
rect 21088 14663 21140 14672
rect 21088 14629 21097 14663
rect 21097 14629 21131 14663
rect 21131 14629 21140 14663
rect 21088 14620 21140 14629
rect 7912 14518 7964 14570
rect 7976 14518 8028 14570
rect 8040 14518 8092 14570
rect 8104 14518 8156 14570
rect 14843 14518 14895 14570
rect 14907 14518 14959 14570
rect 14971 14518 15023 14570
rect 15035 14518 15087 14570
rect 4344 14416 4396 14468
rect 4712 14459 4764 14468
rect 4712 14425 4721 14459
rect 4721 14425 4755 14459
rect 4755 14425 4764 14459
rect 4712 14416 4764 14425
rect 7380 14416 7432 14468
rect 7196 14348 7248 14400
rect 7656 14348 7708 14400
rect 15568 14416 15620 14468
rect 21180 14416 21232 14468
rect 8392 14348 8444 14400
rect 10140 14391 10192 14400
rect 9680 14280 9732 14332
rect 3056 14255 3108 14264
rect 3056 14221 3065 14255
rect 3065 14221 3099 14255
rect 3099 14221 3108 14255
rect 3056 14212 3108 14221
rect 4160 14212 4212 14264
rect 5264 14255 5316 14264
rect 5264 14221 5273 14255
rect 5273 14221 5307 14255
rect 5307 14221 5316 14255
rect 6828 14255 6880 14264
rect 5264 14212 5316 14221
rect 6828 14221 6837 14255
rect 6837 14221 6871 14255
rect 6871 14221 6880 14255
rect 6828 14212 6880 14221
rect 8392 14212 8444 14264
rect 9496 14255 9548 14264
rect 9496 14221 9505 14255
rect 9505 14221 9539 14255
rect 9539 14221 9548 14255
rect 9496 14212 9548 14221
rect 7840 14144 7892 14196
rect 10140 14357 10149 14391
rect 10149 14357 10183 14391
rect 10183 14357 10192 14391
rect 10140 14348 10192 14357
rect 12808 14391 12860 14400
rect 12808 14357 12817 14391
rect 12817 14357 12851 14391
rect 12851 14357 12860 14391
rect 12808 14348 12860 14357
rect 18052 14348 18104 14400
rect 13728 14323 13780 14332
rect 13728 14289 13737 14323
rect 13737 14289 13771 14323
rect 13771 14289 13780 14323
rect 13728 14280 13780 14289
rect 14280 14323 14332 14332
rect 14280 14289 14314 14323
rect 14314 14289 14332 14323
rect 14280 14280 14332 14289
rect 15292 14280 15344 14332
rect 18144 14280 18196 14332
rect 18972 14280 19024 14332
rect 20812 14323 20864 14332
rect 20812 14289 20821 14323
rect 20821 14289 20855 14323
rect 20855 14289 20864 14323
rect 20812 14280 20864 14289
rect 13084 14255 13136 14264
rect 3976 14076 4028 14128
rect 8024 14076 8076 14128
rect 9220 14076 9272 14128
rect 13084 14221 13093 14255
rect 13093 14221 13127 14255
rect 13127 14221 13136 14255
rect 13084 14212 13136 14221
rect 16120 14255 16172 14264
rect 13820 14144 13872 14196
rect 12256 14076 12308 14128
rect 13544 14119 13596 14128
rect 13544 14085 13553 14119
rect 13553 14085 13587 14119
rect 13587 14085 13596 14119
rect 16120 14221 16129 14255
rect 16129 14221 16163 14255
rect 16163 14221 16172 14255
rect 16120 14212 16172 14221
rect 19432 14212 19484 14264
rect 20904 14212 20956 14264
rect 13544 14076 13596 14085
rect 15108 14076 15160 14128
rect 16304 14076 16356 14128
rect 18696 14076 18748 14128
rect 20260 14076 20312 14128
rect 4447 13974 4499 14026
rect 4511 13974 4563 14026
rect 4575 13974 4627 14026
rect 4639 13974 4691 14026
rect 11378 13974 11430 14026
rect 11442 13974 11494 14026
rect 11506 13974 11558 14026
rect 11570 13974 11622 14026
rect 18308 13974 18360 14026
rect 18372 13974 18424 14026
rect 18436 13974 18488 14026
rect 18500 13974 18552 14026
rect 4160 13872 4212 13924
rect 3056 13668 3108 13720
rect 6920 13872 6972 13924
rect 7196 13915 7248 13924
rect 7196 13881 7205 13915
rect 7205 13881 7239 13915
rect 7239 13881 7248 13915
rect 7196 13872 7248 13881
rect 8024 13915 8076 13924
rect 8024 13881 8033 13915
rect 8033 13881 8067 13915
rect 8067 13881 8076 13915
rect 8024 13872 8076 13881
rect 8392 13915 8444 13924
rect 8392 13881 8401 13915
rect 8401 13881 8435 13915
rect 8435 13881 8444 13915
rect 8392 13872 8444 13881
rect 8024 13736 8076 13788
rect 9036 13779 9088 13788
rect 9036 13745 9045 13779
rect 9045 13745 9079 13779
rect 9079 13745 9088 13779
rect 9036 13736 9088 13745
rect 9220 13668 9272 13720
rect 15108 13872 15160 13924
rect 15292 13915 15344 13924
rect 15292 13881 15301 13915
rect 15301 13881 15335 13915
rect 15335 13881 15344 13915
rect 15292 13872 15344 13881
rect 18052 13872 18104 13924
rect 18972 13915 19024 13924
rect 12256 13779 12308 13788
rect 12256 13745 12265 13779
rect 12265 13745 12299 13779
rect 12299 13745 12308 13779
rect 12256 13736 12308 13745
rect 16120 13804 16172 13856
rect 18972 13881 18981 13915
rect 18981 13881 19015 13915
rect 19015 13881 19024 13915
rect 18972 13872 19024 13881
rect 20444 13915 20496 13924
rect 20444 13881 20453 13915
rect 20453 13881 20487 13915
rect 20487 13881 20496 13915
rect 20444 13872 20496 13881
rect 20628 13872 20680 13924
rect 13820 13736 13872 13788
rect 16580 13779 16632 13788
rect 14280 13668 14332 13720
rect 16580 13745 16589 13779
rect 16589 13745 16623 13779
rect 16623 13745 16632 13779
rect 16580 13736 16632 13745
rect 17316 13779 17368 13788
rect 17316 13745 17325 13779
rect 17325 13745 17359 13779
rect 17359 13745 17368 13779
rect 17316 13736 17368 13745
rect 18696 13736 18748 13788
rect 15476 13668 15528 13720
rect 16304 13711 16356 13720
rect 16304 13677 16313 13711
rect 16313 13677 16347 13711
rect 16347 13677 16356 13711
rect 16304 13668 16356 13677
rect 19340 13668 19392 13720
rect 20260 13711 20312 13720
rect 20260 13677 20269 13711
rect 20269 13677 20303 13711
rect 20303 13677 20312 13711
rect 20260 13668 20312 13677
rect 20904 13711 20956 13720
rect 20904 13677 20913 13711
rect 20913 13677 20947 13711
rect 20947 13677 20956 13711
rect 20904 13668 20956 13677
rect 12440 13600 12492 13652
rect 12808 13600 12860 13652
rect 8760 13575 8812 13584
rect 8760 13541 8769 13575
rect 8769 13541 8803 13575
rect 8803 13541 8812 13575
rect 8760 13532 8812 13541
rect 10600 13532 10652 13584
rect 14280 13575 14332 13584
rect 14280 13541 14289 13575
rect 14289 13541 14323 13575
rect 14323 13541 14332 13575
rect 14280 13532 14332 13541
rect 16488 13600 16540 13652
rect 19064 13532 19116 13584
rect 19340 13575 19392 13584
rect 19340 13541 19349 13575
rect 19349 13541 19383 13575
rect 19383 13541 19392 13575
rect 19340 13532 19392 13541
rect 7912 13430 7964 13482
rect 7976 13430 8028 13482
rect 8040 13430 8092 13482
rect 8104 13430 8156 13482
rect 14843 13430 14895 13482
rect 14907 13430 14959 13482
rect 14971 13430 15023 13482
rect 15035 13430 15087 13482
rect 5264 13328 5316 13380
rect 8760 13328 8812 13380
rect 9496 13328 9548 13380
rect 10968 13328 11020 13380
rect 14280 13328 14332 13380
rect 15476 13371 15528 13380
rect 15476 13337 15485 13371
rect 15485 13337 15519 13371
rect 15519 13337 15528 13371
rect 15476 13328 15528 13337
rect 16488 13328 16540 13380
rect 19340 13328 19392 13380
rect 20536 13371 20588 13380
rect 20536 13337 20545 13371
rect 20545 13337 20579 13371
rect 20579 13337 20588 13371
rect 20536 13328 20588 13337
rect 21272 13328 21324 13380
rect 9036 13260 9088 13312
rect 12808 13260 12860 13312
rect 12992 13303 13044 13312
rect 12992 13269 13001 13303
rect 13001 13269 13035 13303
rect 13035 13269 13044 13303
rect 13912 13303 13964 13312
rect 12992 13260 13044 13269
rect 13912 13269 13921 13303
rect 13921 13269 13955 13303
rect 13955 13269 13964 13303
rect 13912 13260 13964 13269
rect 15292 13260 15344 13312
rect 3056 13192 3108 13244
rect 6920 13124 6972 13176
rect 7748 13167 7800 13176
rect 7748 13133 7757 13167
rect 7757 13133 7791 13167
rect 7791 13133 7800 13167
rect 7748 13124 7800 13133
rect 9404 13192 9456 13244
rect 12716 13192 12768 13244
rect 12440 13124 12492 13176
rect 13084 13167 13136 13176
rect 13084 13133 13093 13167
rect 13093 13133 13127 13167
rect 13127 13133 13136 13167
rect 13084 13124 13136 13133
rect 18880 13167 18932 13176
rect 18880 13133 18889 13167
rect 18889 13133 18923 13167
rect 18923 13133 18932 13167
rect 18880 13124 18932 13133
rect 19340 13124 19392 13176
rect 20628 13124 20680 13176
rect 13820 12988 13872 13040
rect 4447 12886 4499 12938
rect 4511 12886 4563 12938
rect 4575 12886 4627 12938
rect 4639 12886 4691 12938
rect 11378 12886 11430 12938
rect 11442 12886 11494 12938
rect 11506 12886 11558 12938
rect 11570 12886 11622 12938
rect 18308 12886 18360 12938
rect 18372 12886 18424 12938
rect 18436 12886 18488 12938
rect 18500 12886 18552 12938
rect 7748 12827 7800 12836
rect 7748 12793 7757 12827
rect 7757 12793 7791 12827
rect 7791 12793 7800 12827
rect 7748 12784 7800 12793
rect 9680 12784 9732 12836
rect 10968 12784 11020 12836
rect 10600 12691 10652 12700
rect 10600 12657 10609 12691
rect 10609 12657 10643 12691
rect 10643 12657 10652 12691
rect 10600 12648 10652 12657
rect 8208 12580 8260 12632
rect 10968 12623 11020 12632
rect 10968 12589 10977 12623
rect 10977 12589 11011 12623
rect 11011 12589 11020 12623
rect 10968 12580 11020 12589
rect 12440 12784 12492 12836
rect 13728 12784 13780 12836
rect 18880 12784 18932 12836
rect 19064 12784 19116 12836
rect 20168 12784 20220 12836
rect 20444 12827 20496 12836
rect 20444 12793 20453 12827
rect 20453 12793 20487 12827
rect 20487 12793 20496 12827
rect 20444 12784 20496 12793
rect 21088 12827 21140 12836
rect 21088 12793 21097 12827
rect 21097 12793 21131 12827
rect 21131 12793 21140 12827
rect 21088 12784 21140 12793
rect 11060 12512 11112 12564
rect 19248 12716 19300 12768
rect 16212 12691 16264 12700
rect 16212 12657 16221 12691
rect 16221 12657 16255 12691
rect 16255 12657 16264 12691
rect 16212 12648 16264 12657
rect 17592 12691 17644 12700
rect 17592 12657 17601 12691
rect 17601 12657 17635 12691
rect 17635 12657 17644 12691
rect 17592 12648 17644 12657
rect 17776 12648 17828 12700
rect 19708 12623 19760 12632
rect 19708 12589 19717 12623
rect 19717 12589 19751 12623
rect 19751 12589 19760 12623
rect 19708 12580 19760 12589
rect 20352 12580 20404 12632
rect 16580 12512 16632 12564
rect 17132 12512 17184 12564
rect 7748 12444 7800 12496
rect 8208 12444 8260 12496
rect 11336 12444 11388 12496
rect 14556 12444 14608 12496
rect 16120 12487 16172 12496
rect 16120 12453 16129 12487
rect 16129 12453 16163 12487
rect 16163 12453 16172 12487
rect 16764 12487 16816 12496
rect 16120 12444 16172 12453
rect 16764 12453 16773 12487
rect 16773 12453 16807 12487
rect 16807 12453 16816 12487
rect 16764 12444 16816 12453
rect 17408 12487 17460 12496
rect 17408 12453 17417 12487
rect 17417 12453 17451 12487
rect 17451 12453 17460 12487
rect 17408 12444 17460 12453
rect 18052 12444 18104 12496
rect 18972 12444 19024 12496
rect 7912 12342 7964 12394
rect 7976 12342 8028 12394
rect 8040 12342 8092 12394
rect 8104 12342 8156 12394
rect 14843 12342 14895 12394
rect 14907 12342 14959 12394
rect 14971 12342 15023 12394
rect 15035 12342 15087 12394
rect 10968 12240 11020 12292
rect 13084 12240 13136 12292
rect 14556 12240 14608 12292
rect 16120 12240 16172 12292
rect 16580 12240 16632 12292
rect 16764 12240 16816 12292
rect 18236 12240 18288 12292
rect 18880 12240 18932 12292
rect 19800 12240 19852 12292
rect 10508 12104 10560 12156
rect 15292 12172 15344 12224
rect 17132 12215 17184 12224
rect 8484 12036 8536 12088
rect 11060 12036 11112 12088
rect 848 11968 900 12020
rect 13636 11968 13688 12020
rect 17132 12181 17141 12215
rect 17141 12181 17175 12215
rect 17175 12181 17184 12215
rect 17132 12172 17184 12181
rect 17684 12172 17736 12224
rect 20352 12172 20404 12224
rect 14372 12036 14424 12088
rect 14280 11968 14332 12020
rect 18052 12104 18104 12156
rect 18144 12104 18196 12156
rect 19248 12104 19300 12156
rect 15200 12036 15252 12088
rect 17868 12036 17920 12088
rect 18604 12079 18656 12088
rect 18604 12045 18613 12079
rect 18613 12045 18647 12079
rect 18647 12045 18656 12079
rect 18604 12036 18656 12045
rect 17776 11968 17828 12020
rect 13544 11900 13596 11952
rect 17408 11900 17460 11952
rect 19064 11900 19116 11952
rect 4447 11798 4499 11850
rect 4511 11798 4563 11850
rect 4575 11798 4627 11850
rect 4639 11798 4691 11850
rect 11378 11798 11430 11850
rect 11442 11798 11494 11850
rect 11506 11798 11558 11850
rect 11570 11798 11622 11850
rect 18308 11798 18360 11850
rect 18372 11798 18424 11850
rect 18436 11798 18488 11850
rect 18500 11798 18552 11850
rect 6644 11696 6696 11748
rect 8300 11560 8352 11612
rect 9496 11696 9548 11748
rect 11060 11739 11112 11748
rect 11060 11705 11069 11739
rect 11069 11705 11103 11739
rect 11103 11705 11112 11739
rect 11060 11696 11112 11705
rect 11244 11696 11296 11748
rect 14280 11696 14332 11748
rect 14372 11696 14424 11748
rect 16212 11696 16264 11748
rect 18144 11739 18196 11748
rect 18144 11705 18153 11739
rect 18153 11705 18187 11739
rect 18187 11705 18196 11739
rect 18144 11696 18196 11705
rect 19616 11696 19668 11748
rect 20076 11696 20128 11748
rect 8760 11560 8812 11612
rect 13084 11603 13136 11612
rect 13084 11569 13093 11603
rect 13093 11569 13127 11603
rect 13127 11569 13136 11603
rect 13084 11560 13136 11569
rect 15200 11492 15252 11544
rect 17776 11628 17828 11680
rect 18604 11628 18656 11680
rect 17684 11603 17736 11612
rect 17684 11569 17693 11603
rect 17693 11569 17727 11603
rect 17727 11569 17736 11603
rect 17684 11560 17736 11569
rect 17868 11560 17920 11612
rect 18788 11603 18840 11612
rect 18788 11569 18797 11603
rect 18797 11569 18831 11603
rect 18831 11569 18840 11603
rect 18788 11560 18840 11569
rect 19432 11492 19484 11544
rect 20904 11535 20956 11544
rect 20904 11501 20913 11535
rect 20913 11501 20947 11535
rect 20947 11501 20956 11535
rect 20904 11492 20956 11501
rect 22008 11535 22060 11544
rect 22008 11501 22017 11535
rect 22017 11501 22051 11535
rect 22051 11501 22060 11535
rect 22008 11492 22060 11501
rect 9956 11467 10008 11476
rect 9956 11433 9990 11467
rect 9990 11433 10008 11467
rect 9956 11424 10008 11433
rect 18512 11467 18564 11476
rect 8300 11356 8352 11408
rect 11244 11356 11296 11408
rect 12348 11356 12400 11408
rect 15476 11356 15528 11408
rect 18512 11433 18521 11467
rect 18521 11433 18555 11467
rect 18555 11433 18564 11467
rect 18512 11424 18564 11433
rect 19248 11424 19300 11476
rect 17592 11356 17644 11408
rect 18604 11399 18656 11408
rect 18604 11365 18613 11399
rect 18613 11365 18647 11399
rect 18647 11365 18656 11399
rect 18604 11356 18656 11365
rect 19340 11356 19392 11408
rect 7912 11254 7964 11306
rect 7976 11254 8028 11306
rect 8040 11254 8092 11306
rect 8104 11254 8156 11306
rect 14843 11254 14895 11306
rect 14907 11254 14959 11306
rect 14971 11254 15023 11306
rect 15035 11254 15087 11306
rect 7472 11152 7524 11204
rect 10508 11195 10560 11204
rect 10508 11161 10517 11195
rect 10517 11161 10551 11195
rect 10551 11161 10560 11195
rect 10508 11152 10560 11161
rect 13084 11152 13136 11204
rect 15476 11152 15528 11204
rect 18512 11152 18564 11204
rect 19984 11152 20036 11204
rect 17132 11084 17184 11136
rect 19064 11084 19116 11136
rect 19432 11127 19484 11136
rect 19432 11093 19441 11127
rect 19441 11093 19475 11127
rect 19475 11093 19484 11127
rect 19432 11084 19484 11093
rect 9864 11016 9916 11068
rect 10876 11059 10928 11068
rect 10876 11025 10885 11059
rect 10885 11025 10919 11059
rect 10919 11025 10928 11059
rect 10876 11016 10928 11025
rect 11152 11016 11204 11068
rect 13728 11059 13780 11068
rect 13728 11025 13737 11059
rect 13737 11025 13771 11059
rect 13771 11025 13780 11059
rect 13728 11016 13780 11025
rect 19156 11059 19208 11068
rect 19156 11025 19165 11059
rect 19165 11025 19199 11059
rect 19199 11025 19208 11059
rect 19156 11016 19208 11025
rect 20628 11016 20680 11068
rect 8760 10991 8812 11000
rect 8760 10957 8769 10991
rect 8769 10957 8803 10991
rect 8803 10957 8812 10991
rect 8760 10948 8812 10957
rect 8392 10880 8444 10932
rect 9956 10948 10008 11000
rect 18696 10880 18748 10932
rect 18972 10880 19024 10932
rect 20536 10923 20588 10932
rect 20536 10889 20545 10923
rect 20545 10889 20579 10923
rect 20579 10889 20588 10923
rect 20536 10880 20588 10889
rect 11704 10812 11756 10864
rect 14004 10812 14056 10864
rect 18604 10812 18656 10864
rect 4447 10710 4499 10762
rect 4511 10710 4563 10762
rect 4575 10710 4627 10762
rect 4639 10710 4691 10762
rect 11378 10710 11430 10762
rect 11442 10710 11494 10762
rect 11506 10710 11558 10762
rect 11570 10710 11622 10762
rect 18308 10710 18360 10762
rect 18372 10710 18424 10762
rect 18436 10710 18488 10762
rect 18500 10710 18552 10762
rect 8484 10608 8536 10660
rect 11152 10651 11204 10660
rect 11152 10617 11161 10651
rect 11161 10617 11195 10651
rect 11195 10617 11204 10651
rect 11152 10608 11204 10617
rect 12348 10608 12400 10660
rect 19156 10608 19208 10660
rect 21456 10608 21508 10660
rect 8300 10472 8352 10524
rect 9956 10472 10008 10524
rect 10876 10472 10928 10524
rect 14004 10540 14056 10592
rect 11704 10515 11756 10524
rect 11704 10481 11713 10515
rect 11713 10481 11747 10515
rect 11747 10481 11756 10515
rect 11704 10472 11756 10481
rect 14372 10472 14424 10524
rect 19892 10515 19944 10524
rect 19892 10481 19901 10515
rect 19901 10481 19935 10515
rect 19935 10481 19944 10515
rect 19892 10472 19944 10481
rect 8392 10447 8444 10456
rect 8392 10413 8401 10447
rect 8401 10413 8435 10447
rect 8435 10413 8444 10447
rect 8392 10404 8444 10413
rect 12348 10404 12400 10456
rect 14004 10404 14056 10456
rect 20628 10404 20680 10456
rect 13820 10336 13872 10388
rect 13452 10268 13504 10320
rect 14004 10311 14056 10320
rect 14004 10277 14013 10311
rect 14013 10277 14047 10311
rect 14047 10277 14056 10311
rect 14004 10268 14056 10277
rect 14280 10268 14332 10320
rect 18972 10311 19024 10320
rect 18972 10277 18981 10311
rect 18981 10277 19015 10311
rect 19015 10277 19024 10311
rect 18972 10268 19024 10277
rect 19708 10311 19760 10320
rect 19708 10277 19717 10311
rect 19717 10277 19751 10311
rect 19751 10277 19760 10311
rect 19708 10268 19760 10277
rect 7912 10166 7964 10218
rect 7976 10166 8028 10218
rect 8040 10166 8092 10218
rect 8104 10166 8156 10218
rect 14843 10166 14895 10218
rect 14907 10166 14959 10218
rect 14971 10166 15023 10218
rect 15035 10166 15087 10218
rect 8208 10064 8260 10116
rect 9956 10064 10008 10116
rect 13452 10107 13504 10116
rect 13452 10073 13461 10107
rect 13461 10073 13495 10107
rect 13495 10073 13504 10107
rect 13452 10064 13504 10073
rect 13544 10107 13596 10116
rect 13544 10073 13553 10107
rect 13553 10073 13587 10107
rect 13587 10073 13596 10107
rect 13544 10064 13596 10073
rect 17776 10064 17828 10116
rect 18788 10064 18840 10116
rect 19708 10107 19760 10116
rect 19708 10073 19717 10107
rect 19717 10073 19751 10107
rect 19751 10073 19760 10107
rect 19708 10064 19760 10073
rect 20076 10107 20128 10116
rect 20076 10073 20085 10107
rect 20085 10073 20119 10107
rect 20119 10073 20128 10107
rect 20076 10064 20128 10073
rect 21640 10064 21692 10116
rect 14372 9996 14424 10048
rect 18972 9996 19024 10048
rect 8760 9928 8812 9980
rect 15200 9928 15252 9980
rect 18052 9971 18104 9980
rect 18052 9937 18061 9971
rect 18061 9937 18095 9971
rect 18095 9937 18104 9971
rect 18052 9928 18104 9937
rect 19892 9928 19944 9980
rect 20536 9928 20588 9980
rect 13084 9860 13136 9912
rect 20260 9903 20312 9912
rect 20260 9869 20269 9903
rect 20269 9869 20303 9903
rect 20303 9869 20312 9903
rect 20260 9860 20312 9869
rect 13912 9724 13964 9776
rect 15844 9724 15896 9776
rect 4447 9622 4499 9674
rect 4511 9622 4563 9674
rect 4575 9622 4627 9674
rect 4639 9622 4691 9674
rect 11378 9622 11430 9674
rect 11442 9622 11494 9674
rect 11506 9622 11558 9674
rect 11570 9622 11622 9674
rect 18308 9622 18360 9674
rect 18372 9622 18424 9674
rect 18436 9622 18488 9674
rect 18500 9622 18552 9674
rect 11704 9520 11756 9572
rect 19892 9520 19944 9572
rect 13084 9316 13136 9368
rect 13912 9427 13964 9436
rect 13912 9393 13921 9427
rect 13921 9393 13955 9427
rect 13955 9393 13964 9427
rect 13912 9384 13964 9393
rect 21732 9452 21784 9504
rect 15844 9427 15896 9436
rect 15844 9393 15853 9427
rect 15853 9393 15887 9427
rect 15887 9393 15896 9427
rect 15844 9384 15896 9393
rect 18052 9384 18104 9436
rect 19708 9316 19760 9368
rect 20260 9316 20312 9368
rect 20904 9359 20956 9368
rect 20904 9325 20913 9359
rect 20913 9325 20947 9359
rect 20947 9325 20956 9359
rect 20904 9316 20956 9325
rect 12992 9180 13044 9232
rect 13636 9180 13688 9232
rect 15384 9180 15436 9232
rect 16488 9180 16540 9232
rect 7912 9078 7964 9130
rect 7976 9078 8028 9130
rect 8040 9078 8092 9130
rect 8104 9078 8156 9130
rect 14843 9078 14895 9130
rect 14907 9078 14959 9130
rect 14971 9078 15023 9130
rect 15035 9078 15087 9130
rect 12072 8976 12124 9028
rect 13176 8976 13228 9028
rect 15384 9019 15436 9028
rect 15384 8985 15393 9019
rect 15393 8985 15427 9019
rect 15427 8985 15436 9019
rect 15384 8976 15436 8985
rect 15660 8976 15712 9028
rect 20076 9019 20128 9028
rect 20076 8985 20085 9019
rect 20085 8985 20119 9019
rect 20119 8985 20128 9019
rect 20076 8976 20128 8985
rect 20536 9019 20588 9028
rect 20536 8985 20545 9019
rect 20545 8985 20579 9019
rect 20579 8985 20588 9019
rect 20536 8976 20588 8985
rect 11704 8883 11756 8892
rect 11704 8849 11713 8883
rect 11713 8849 11747 8883
rect 11747 8849 11756 8883
rect 11704 8840 11756 8849
rect 13636 8840 13688 8892
rect 16580 8840 16632 8892
rect 16396 8704 16448 8756
rect 4447 8534 4499 8586
rect 4511 8534 4563 8586
rect 4575 8534 4627 8586
rect 4639 8534 4691 8586
rect 11378 8534 11430 8586
rect 11442 8534 11494 8586
rect 11506 8534 11558 8586
rect 11570 8534 11622 8586
rect 18308 8534 18360 8586
rect 18372 8534 18424 8586
rect 18436 8534 18488 8586
rect 18500 8534 18552 8586
rect 16304 8432 16356 8484
rect 11704 8296 11756 8348
rect 13636 8339 13688 8348
rect 13636 8305 13645 8339
rect 13645 8305 13679 8339
rect 13679 8305 13688 8339
rect 13636 8296 13688 8305
rect 16580 8339 16632 8348
rect 16580 8305 16589 8339
rect 16589 8305 16623 8339
rect 16623 8305 16632 8339
rect 16580 8296 16632 8305
rect 11060 8271 11112 8280
rect 11060 8237 11069 8271
rect 11069 8237 11103 8271
rect 11103 8237 11112 8271
rect 11060 8228 11112 8237
rect 14096 8228 14148 8280
rect 16948 8228 17000 8280
rect 20628 8228 20680 8280
rect 22008 8271 22060 8280
rect 22008 8237 22017 8271
rect 22017 8237 22051 8271
rect 22051 8237 22060 8271
rect 22008 8228 22060 8237
rect 14188 8092 14240 8144
rect 21088 8092 21140 8144
rect 7912 7990 7964 8042
rect 7976 7990 8028 8042
rect 8040 7990 8092 8042
rect 8104 7990 8156 8042
rect 14843 7990 14895 8042
rect 14907 7990 14959 8042
rect 14971 7990 15023 8042
rect 15035 7990 15087 8042
rect 11060 7888 11112 7940
rect 16948 7931 17000 7940
rect 16948 7897 16957 7931
rect 16957 7897 16991 7931
rect 16991 7897 17000 7931
rect 16948 7888 17000 7897
rect 15936 7820 15988 7872
rect 18052 7820 18104 7872
rect 19708 7888 19760 7940
rect 12992 7752 13044 7804
rect 13728 7752 13780 7804
rect 13912 7795 13964 7804
rect 13912 7761 13946 7795
rect 13946 7761 13964 7795
rect 13912 7752 13964 7761
rect 11244 7684 11296 7736
rect 11704 7727 11756 7736
rect 11704 7693 11713 7727
rect 11713 7693 11747 7727
rect 11747 7693 11756 7727
rect 15292 7727 15344 7736
rect 11704 7684 11756 7693
rect 15292 7693 15301 7727
rect 15301 7693 15335 7727
rect 15335 7693 15344 7727
rect 15292 7684 15344 7693
rect 18144 7752 18196 7804
rect 20812 7795 20864 7804
rect 20812 7761 20821 7795
rect 20821 7761 20855 7795
rect 20855 7761 20864 7795
rect 20812 7752 20864 7761
rect 15016 7591 15068 7600
rect 15016 7557 15025 7591
rect 15025 7557 15059 7591
rect 15059 7557 15068 7591
rect 15016 7548 15068 7557
rect 17960 7684 18012 7736
rect 18604 7548 18656 7600
rect 4447 7446 4499 7498
rect 4511 7446 4563 7498
rect 4575 7446 4627 7498
rect 4639 7446 4691 7498
rect 11378 7446 11430 7498
rect 11442 7446 11494 7498
rect 11506 7446 11558 7498
rect 11570 7446 11622 7498
rect 18308 7446 18360 7498
rect 18372 7446 18424 7498
rect 18436 7446 18488 7498
rect 18500 7446 18552 7498
rect 11704 7344 11756 7396
rect 11888 7344 11940 7396
rect 8300 7208 8352 7260
rect 13728 7276 13780 7328
rect 13912 7208 13964 7260
rect 10140 7115 10192 7124
rect 10140 7081 10174 7115
rect 10174 7081 10192 7115
rect 10140 7072 10192 7081
rect 12992 7072 13044 7124
rect 15200 7140 15252 7192
rect 17960 7344 18012 7396
rect 18144 7344 18196 7396
rect 18604 7344 18656 7396
rect 21088 7387 21140 7396
rect 21088 7353 21097 7387
rect 21097 7353 21131 7387
rect 21131 7353 21140 7387
rect 21088 7344 21140 7353
rect 18972 7208 19024 7260
rect 14188 7047 14240 7056
rect 14188 7013 14197 7047
rect 14197 7013 14231 7047
rect 14231 7013 14240 7047
rect 14188 7004 14240 7013
rect 14740 7072 14792 7124
rect 15016 7072 15068 7124
rect 15384 7004 15436 7056
rect 20904 7183 20956 7192
rect 20904 7149 20913 7183
rect 20913 7149 20947 7183
rect 20947 7149 20956 7183
rect 20904 7140 20956 7149
rect 19248 7004 19300 7056
rect 7912 6902 7964 6954
rect 7976 6902 8028 6954
rect 8040 6902 8092 6954
rect 8104 6902 8156 6954
rect 14843 6902 14895 6954
rect 14907 6902 14959 6954
rect 14971 6902 15023 6954
rect 15035 6902 15087 6954
rect 11244 6800 11296 6852
rect 4068 6460 4120 6512
rect 11888 6800 11940 6852
rect 14188 6800 14240 6852
rect 15384 6800 15436 6852
rect 18972 6800 19024 6852
rect 12532 6732 12584 6784
rect 15292 6732 15344 6784
rect 18052 6707 18104 6716
rect 18052 6673 18061 6707
rect 18061 6673 18095 6707
rect 18095 6673 18104 6707
rect 18052 6664 18104 6673
rect 8300 6596 8352 6648
rect 14740 6639 14792 6648
rect 10140 6528 10192 6580
rect 14740 6605 14749 6639
rect 14749 6605 14783 6639
rect 14783 6605 14792 6639
rect 14740 6596 14792 6605
rect 14096 6528 14148 6580
rect 12532 6503 12584 6512
rect 12532 6469 12541 6503
rect 12541 6469 12575 6503
rect 12575 6469 12584 6503
rect 12532 6460 12584 6469
rect 15200 6460 15252 6512
rect 17960 6460 18012 6512
rect 21364 6503 21416 6512
rect 21364 6469 21373 6503
rect 21373 6469 21407 6503
rect 21407 6469 21416 6503
rect 21364 6460 21416 6469
rect 4447 6358 4499 6410
rect 4511 6358 4563 6410
rect 4575 6358 4627 6410
rect 4639 6358 4691 6410
rect 11378 6358 11430 6410
rect 11442 6358 11494 6410
rect 11506 6358 11558 6410
rect 11570 6358 11622 6410
rect 18308 6358 18360 6410
rect 18372 6358 18424 6410
rect 18436 6358 18488 6410
rect 18500 6358 18552 6410
rect 12900 6256 12952 6308
rect 21364 6052 21416 6104
rect 7912 5814 7964 5866
rect 7976 5814 8028 5866
rect 8040 5814 8092 5866
rect 8104 5814 8156 5866
rect 14843 5814 14895 5866
rect 14907 5814 14959 5866
rect 14971 5814 15023 5866
rect 15035 5814 15087 5866
rect 12624 5712 12676 5764
rect 21272 5576 21324 5628
rect 4447 5270 4499 5322
rect 4511 5270 4563 5322
rect 4575 5270 4627 5322
rect 4639 5270 4691 5322
rect 11378 5270 11430 5322
rect 11442 5270 11494 5322
rect 11506 5270 11558 5322
rect 11570 5270 11622 5322
rect 18308 5270 18360 5322
rect 18372 5270 18424 5322
rect 18436 5270 18488 5322
rect 18500 5270 18552 5322
rect 12532 5168 12584 5220
rect 17960 5168 18012 5220
rect 21272 5143 21324 5152
rect 21272 5109 21281 5143
rect 21281 5109 21315 5143
rect 21315 5109 21324 5143
rect 21272 5100 21324 5109
rect 7912 4726 7964 4778
rect 7976 4726 8028 4778
rect 8040 4726 8092 4778
rect 8104 4726 8156 4778
rect 14843 4726 14895 4778
rect 14907 4726 14959 4778
rect 14971 4726 15023 4778
rect 15035 4726 15087 4778
rect 20996 4667 21048 4676
rect 20996 4633 21005 4667
rect 21005 4633 21039 4667
rect 21039 4633 21048 4667
rect 20996 4624 21048 4633
rect 21272 4488 21324 4540
rect 4447 4182 4499 4234
rect 4511 4182 4563 4234
rect 4575 4182 4627 4234
rect 4639 4182 4691 4234
rect 11378 4182 11430 4234
rect 11442 4182 11494 4234
rect 11506 4182 11558 4234
rect 11570 4182 11622 4234
rect 18308 4182 18360 4234
rect 18372 4182 18424 4234
rect 18436 4182 18488 4234
rect 18500 4182 18552 4234
rect 21272 4123 21324 4132
rect 21272 4089 21281 4123
rect 21281 4089 21315 4123
rect 21315 4089 21324 4123
rect 21272 4080 21324 4089
rect 16488 3944 16540 3996
rect 18788 3944 18840 3996
rect 7912 3638 7964 3690
rect 7976 3638 8028 3690
rect 8040 3638 8092 3690
rect 8104 3638 8156 3690
rect 14843 3638 14895 3690
rect 14907 3638 14959 3690
rect 14971 3638 15023 3690
rect 15035 3638 15087 3690
rect 4447 3094 4499 3146
rect 4511 3094 4563 3146
rect 4575 3094 4627 3146
rect 4639 3094 4691 3146
rect 11378 3094 11430 3146
rect 11442 3094 11494 3146
rect 11506 3094 11558 3146
rect 11570 3094 11622 3146
rect 18308 3094 18360 3146
rect 18372 3094 18424 3146
rect 18436 3094 18488 3146
rect 18500 3094 18552 3146
rect 18696 2924 18748 2976
rect 18880 2924 18932 2976
rect 7912 2550 7964 2602
rect 7976 2550 8028 2602
rect 8040 2550 8092 2602
rect 8104 2550 8156 2602
rect 14843 2550 14895 2602
rect 14907 2550 14959 2602
rect 14971 2550 15023 2602
rect 15035 2550 15087 2602
rect 14280 2380 14332 2432
rect 18144 2380 18196 2432
rect 4447 2006 4499 2058
rect 4511 2006 4563 2058
rect 4575 2006 4627 2058
rect 4639 2006 4691 2058
rect 11378 2006 11430 2058
rect 11442 2006 11494 2058
rect 11506 2006 11558 2058
rect 11570 2006 11622 2058
rect 18308 2006 18360 2058
rect 18372 2006 18424 2058
rect 18436 2006 18488 2058
rect 18500 2006 18552 2058
rect 14004 1904 14056 1956
rect 18144 1904 18196 1956
rect 14556 1156 14608 1208
rect 17960 1156 18012 1208
<< metal2 >>
rect 294 22056 350 22856
rect 846 22056 902 22856
rect 1398 22056 1454 22856
rect 1950 22056 2006 22856
rect 2502 22056 2558 22856
rect 3054 22056 3110 22856
rect 3606 22056 3662 22856
rect 4158 22056 4214 22856
rect 4710 22056 4766 22856
rect 5262 22056 5318 22856
rect 5814 22056 5870 22856
rect 6458 22056 6514 22856
rect 7010 22056 7066 22856
rect 7562 22056 7618 22856
rect 8114 22056 8170 22856
rect 8666 22056 8722 22856
rect 9218 22056 9274 22856
rect 9770 22056 9826 22856
rect 10322 22056 10378 22856
rect 10874 22056 10930 22856
rect 11426 22056 11482 22856
rect 12070 22056 12126 22856
rect 12622 22056 12678 22856
rect 13174 22056 13230 22856
rect 13726 22056 13782 22856
rect 14278 22056 14334 22856
rect 14830 22056 14886 22856
rect 15382 22056 15438 22856
rect 15934 22056 15990 22856
rect 16486 22056 16542 22856
rect 17038 22056 17094 22856
rect 17682 22056 17738 22856
rect 18234 22056 18290 22856
rect 18786 22056 18842 22856
rect 19246 22528 19302 22537
rect 19246 22463 19302 22472
rect 308 18214 336 22056
rect 296 18208 348 18214
rect 296 18150 348 18156
rect 860 12026 888 22056
rect 1412 18146 1440 22056
rect 1964 19166 1992 22056
rect 1952 19160 2004 19166
rect 1952 19102 2004 19108
rect 2516 19098 2544 22056
rect 2504 19092 2556 19098
rect 2504 19034 2556 19040
rect 2412 19024 2464 19030
rect 2412 18966 2464 18972
rect 2424 18622 2452 18966
rect 1768 18616 1820 18622
rect 1768 18558 1820 18564
rect 2412 18616 2464 18622
rect 2412 18558 2464 18564
rect 1400 18140 1452 18146
rect 1400 18082 1452 18088
rect 1780 16990 1808 18558
rect 3068 17942 3096 22056
rect 3148 18684 3200 18690
rect 3148 18626 3200 18632
rect 3056 17936 3108 17942
rect 3056 17878 3108 17884
rect 3160 17194 3188 18626
rect 3148 17188 3200 17194
rect 3148 17130 3200 17136
rect 3332 17188 3384 17194
rect 3332 17130 3384 17136
rect 3516 17188 3568 17194
rect 3516 17130 3568 17136
rect 1768 16984 1820 16990
rect 1768 16926 1820 16932
rect 1780 15426 1808 16926
rect 3148 16304 3200 16310
rect 3148 16246 3200 16252
rect 3160 15970 3188 16246
rect 3344 15970 3372 17130
rect 3424 16848 3476 16854
rect 3424 16790 3476 16796
rect 3148 15964 3200 15970
rect 3148 15906 3200 15912
rect 3332 15964 3384 15970
rect 3332 15906 3384 15912
rect 3436 15834 3464 16790
rect 3528 16106 3556 17130
rect 3620 16650 3648 22056
rect 3884 19160 3936 19166
rect 3884 19102 3936 19108
rect 3700 16916 3752 16922
rect 3700 16858 3752 16864
rect 3608 16644 3660 16650
rect 3608 16586 3660 16592
rect 3712 16446 3740 16858
rect 3700 16440 3752 16446
rect 3700 16382 3752 16388
rect 3516 16100 3568 16106
rect 3516 16042 3568 16048
rect 3424 15828 3476 15834
rect 3424 15770 3476 15776
rect 3712 15562 3740 16382
rect 3700 15556 3752 15562
rect 3700 15498 3752 15504
rect 1768 15420 1820 15426
rect 1768 15362 1820 15368
rect 3896 14814 3924 19102
rect 3976 19092 4028 19098
rect 3976 19034 4028 19040
rect 3884 14808 3936 14814
rect 3884 14750 3936 14756
rect 3056 14264 3108 14270
rect 3056 14206 3108 14212
rect 3068 13726 3096 14206
rect 3988 14134 4016 19034
rect 4172 18826 4200 22056
rect 4724 20746 4752 22056
rect 4724 20718 4844 20746
rect 4421 20556 4717 20576
rect 4477 20554 4501 20556
rect 4557 20554 4581 20556
rect 4637 20554 4661 20556
rect 4499 20502 4501 20554
rect 4563 20502 4575 20554
rect 4637 20502 4639 20554
rect 4477 20500 4501 20502
rect 4557 20500 4581 20502
rect 4637 20500 4661 20502
rect 4421 20480 4717 20500
rect 4421 19468 4717 19488
rect 4477 19466 4501 19468
rect 4557 19466 4581 19468
rect 4637 19466 4661 19468
rect 4499 19414 4501 19466
rect 4563 19414 4575 19466
rect 4637 19414 4639 19466
rect 4477 19412 4501 19414
rect 4557 19412 4581 19414
rect 4637 19412 4661 19414
rect 4421 19392 4717 19412
rect 4252 19092 4304 19098
rect 4252 19034 4304 19040
rect 4160 18820 4212 18826
rect 4160 18762 4212 18768
rect 4264 18554 4292 19034
rect 4252 18548 4304 18554
rect 4252 18490 4304 18496
rect 4344 18480 4396 18486
rect 4344 18422 4396 18428
rect 4160 17936 4212 17942
rect 4160 17878 4212 17884
rect 4068 16508 4120 16514
rect 4068 16450 4120 16456
rect 4080 15902 4108 16450
rect 4068 15896 4120 15902
rect 4068 15838 4120 15844
rect 4172 14270 4200 17878
rect 4356 17738 4384 18422
rect 4421 18380 4717 18400
rect 4477 18378 4501 18380
rect 4557 18378 4581 18380
rect 4637 18378 4661 18380
rect 4499 18326 4501 18378
rect 4563 18326 4575 18378
rect 4637 18326 4639 18378
rect 4477 18324 4501 18326
rect 4557 18324 4581 18326
rect 4637 18324 4661 18326
rect 4421 18304 4717 18324
rect 4816 17942 4844 20718
rect 4896 19772 4948 19778
rect 4896 19714 4948 19720
rect 4908 19166 4936 19714
rect 4896 19160 4948 19166
rect 4896 19102 4948 19108
rect 4804 17936 4856 17942
rect 4804 17878 4856 17884
rect 4344 17732 4396 17738
rect 4344 17674 4396 17680
rect 4344 17596 4396 17602
rect 4344 17538 4396 17544
rect 4252 17392 4304 17398
rect 4252 17334 4304 17340
rect 4264 16514 4292 17334
rect 4356 17058 4384 17538
rect 4804 17460 4856 17466
rect 4804 17402 4856 17408
rect 4421 17292 4717 17312
rect 4477 17290 4501 17292
rect 4557 17290 4581 17292
rect 4637 17290 4661 17292
rect 4499 17238 4501 17290
rect 4563 17238 4575 17290
rect 4637 17238 4639 17290
rect 4477 17236 4501 17238
rect 4557 17236 4581 17238
rect 4637 17236 4661 17238
rect 4421 17216 4717 17236
rect 4816 17097 4844 17402
rect 4802 17088 4858 17097
rect 4344 17052 4396 17058
rect 4802 17023 4858 17032
rect 4344 16994 4396 17000
rect 4908 16990 4936 19102
rect 5276 18214 5304 22056
rect 5448 19024 5500 19030
rect 5448 18966 5500 18972
rect 5264 18208 5316 18214
rect 5264 18150 5316 18156
rect 5460 17534 5488 18966
rect 5828 18758 5856 22056
rect 6276 19568 6328 19574
rect 6276 19510 6328 19516
rect 6288 19166 6316 19510
rect 6276 19160 6328 19166
rect 6276 19102 6328 19108
rect 5816 18752 5868 18758
rect 5816 18694 5868 18700
rect 6288 18554 6316 19102
rect 6276 18548 6328 18554
rect 6276 18490 6328 18496
rect 6368 18276 6420 18282
rect 6368 18218 6420 18224
rect 6380 18185 6408 18218
rect 6366 18176 6422 18185
rect 6366 18111 6422 18120
rect 6472 18010 6500 22056
rect 6552 19772 6604 19778
rect 6552 19714 6604 19720
rect 6828 19772 6880 19778
rect 6828 19714 6880 19720
rect 6564 18078 6592 19714
rect 6840 18826 6868 19714
rect 6828 18820 6880 18826
rect 6828 18762 6880 18768
rect 7024 18758 7052 22056
rect 7012 18752 7064 18758
rect 7012 18694 7064 18700
rect 6644 18616 6696 18622
rect 6644 18558 6696 18564
rect 6656 18282 6684 18558
rect 6644 18276 6696 18282
rect 6644 18218 6696 18224
rect 6644 18140 6696 18146
rect 6644 18082 6696 18088
rect 6552 18072 6604 18078
rect 6552 18014 6604 18020
rect 6460 18004 6512 18010
rect 6460 17946 6512 17952
rect 5448 17528 5500 17534
rect 5448 17470 5500 17476
rect 5460 16990 5488 17470
rect 4896 16984 4948 16990
rect 4896 16926 4948 16932
rect 5448 16984 5500 16990
rect 5448 16926 5500 16932
rect 4252 16508 4304 16514
rect 4252 16450 4304 16456
rect 4908 16446 4936 16926
rect 4896 16440 4948 16446
rect 4896 16382 4948 16388
rect 4421 16204 4717 16224
rect 4477 16202 4501 16204
rect 4557 16202 4581 16204
rect 4637 16202 4661 16204
rect 4499 16150 4501 16202
rect 4563 16150 4575 16202
rect 4637 16150 4639 16202
rect 4477 16148 4501 16150
rect 4557 16148 4581 16150
rect 4637 16148 4661 16150
rect 4421 16128 4717 16148
rect 4908 15970 4936 16382
rect 6564 16106 6592 18014
rect 6552 16100 6604 16106
rect 6552 16042 6604 16048
rect 4896 15964 4948 15970
rect 4896 15906 4948 15912
rect 4344 15420 4396 15426
rect 4344 15362 4396 15368
rect 4356 14882 4384 15362
rect 4421 15116 4717 15136
rect 4477 15114 4501 15116
rect 4557 15114 4581 15116
rect 4637 15114 4661 15116
rect 4499 15062 4501 15114
rect 4563 15062 4575 15114
rect 4637 15062 4639 15114
rect 4477 15060 4501 15062
rect 4557 15060 4581 15062
rect 4637 15060 4661 15062
rect 4421 15040 4717 15060
rect 4344 14876 4396 14882
rect 4344 14818 4396 14824
rect 4356 14474 4384 14818
rect 4712 14672 4764 14678
rect 4712 14614 4764 14620
rect 4724 14474 4752 14614
rect 4344 14468 4396 14474
rect 4344 14410 4396 14416
rect 4712 14468 4764 14474
rect 4712 14410 4764 14416
rect 4160 14264 4212 14270
rect 4160 14206 4212 14212
rect 5264 14264 5316 14270
rect 5264 14206 5316 14212
rect 3976 14128 4028 14134
rect 3976 14070 4028 14076
rect 4172 13930 4200 14206
rect 4421 14028 4717 14048
rect 4477 14026 4501 14028
rect 4557 14026 4581 14028
rect 4637 14026 4661 14028
rect 4499 13974 4501 14026
rect 4563 13974 4575 14026
rect 4637 13974 4639 14026
rect 4477 13972 4501 13974
rect 4557 13972 4581 13974
rect 4637 13972 4661 13974
rect 4421 13952 4717 13972
rect 4160 13924 4212 13930
rect 4160 13866 4212 13872
rect 3056 13720 3108 13726
rect 3056 13662 3108 13668
rect 3068 13250 3096 13662
rect 5276 13386 5304 14206
rect 5264 13380 5316 13386
rect 5264 13322 5316 13328
rect 3056 13244 3108 13250
rect 3056 13186 3108 13192
rect 4421 12940 4717 12960
rect 4477 12938 4501 12940
rect 4557 12938 4581 12940
rect 4637 12938 4661 12940
rect 4499 12886 4501 12938
rect 4563 12886 4575 12938
rect 4637 12886 4639 12938
rect 4477 12884 4501 12886
rect 4557 12884 4581 12886
rect 4637 12884 4661 12886
rect 4421 12864 4717 12884
rect 848 12020 900 12026
rect 848 11962 900 11968
rect 4421 11852 4717 11872
rect 4477 11850 4501 11852
rect 4557 11850 4581 11852
rect 4637 11850 4661 11852
rect 4499 11798 4501 11850
rect 4563 11798 4575 11850
rect 4637 11798 4639 11850
rect 4477 11796 4501 11798
rect 4557 11796 4581 11798
rect 4637 11796 4661 11798
rect 4421 11776 4717 11796
rect 6656 11754 6684 18082
rect 6736 17936 6788 17942
rect 6736 17878 6788 17884
rect 7472 17936 7524 17942
rect 7472 17878 7524 17884
rect 6748 17194 6776 17878
rect 6736 17188 6788 17194
rect 6736 17130 6788 17136
rect 6748 16990 6776 17130
rect 7012 17052 7064 17058
rect 7012 16994 7064 17000
rect 6736 16984 6788 16990
rect 6736 16926 6788 16932
rect 7024 16582 7052 16994
rect 7012 16576 7064 16582
rect 7012 16518 7064 16524
rect 6828 16440 6880 16446
rect 6828 16382 6880 16388
rect 6840 16310 6868 16382
rect 6828 16304 6880 16310
rect 6828 16246 6880 16252
rect 6840 16106 6868 16246
rect 6828 16100 6880 16106
rect 6828 16042 6880 16048
rect 7484 15970 7512 17878
rect 7576 15986 7604 22056
rect 8128 20202 8156 22056
rect 8128 20174 8248 20202
rect 7886 20012 8182 20032
rect 7942 20010 7966 20012
rect 8022 20010 8046 20012
rect 8102 20010 8126 20012
rect 7964 19958 7966 20010
rect 8028 19958 8040 20010
rect 8102 19958 8104 20010
rect 7942 19956 7966 19958
rect 8022 19956 8046 19958
rect 8102 19956 8126 19958
rect 7886 19936 8182 19956
rect 7748 19704 7800 19710
rect 7748 19646 7800 19652
rect 7760 18706 7788 19646
rect 7886 18924 8182 18944
rect 7942 18922 7966 18924
rect 8022 18922 8046 18924
rect 8102 18922 8126 18924
rect 7964 18870 7966 18922
rect 8028 18870 8040 18922
rect 8102 18870 8104 18922
rect 7942 18868 7966 18870
rect 8022 18868 8046 18870
rect 8102 18868 8126 18870
rect 7886 18848 8182 18868
rect 7760 18678 7972 18706
rect 7944 18214 7972 18678
rect 8220 18282 8248 20174
rect 8300 19772 8352 19778
rect 8300 19714 8352 19720
rect 8312 19234 8340 19714
rect 8300 19228 8352 19234
rect 8300 19170 8352 19176
rect 8312 19030 8340 19170
rect 8680 19166 8708 22056
rect 8668 19160 8720 19166
rect 8668 19102 8720 19108
rect 8300 19024 8352 19030
rect 8300 18966 8352 18972
rect 8680 18826 8708 19102
rect 8760 19024 8812 19030
rect 8760 18966 8812 18972
rect 8576 18820 8628 18826
rect 8576 18762 8628 18768
rect 8668 18820 8720 18826
rect 8668 18762 8720 18768
rect 8208 18276 8260 18282
rect 8208 18218 8260 18224
rect 7932 18208 7984 18214
rect 7932 18150 7984 18156
rect 8588 17942 8616 18762
rect 8772 18690 8800 18966
rect 8760 18684 8812 18690
rect 8760 18626 8812 18632
rect 8576 17936 8628 17942
rect 8576 17878 8628 17884
rect 7886 17836 8182 17856
rect 7942 17834 7966 17836
rect 8022 17834 8046 17836
rect 8102 17834 8126 17836
rect 7964 17782 7966 17834
rect 8028 17782 8040 17834
rect 8102 17782 8104 17834
rect 7942 17780 7966 17782
rect 8022 17780 8046 17782
rect 8102 17780 8126 17782
rect 7886 17760 8182 17780
rect 9232 17738 9260 22056
rect 9680 19704 9732 19710
rect 9680 19646 9732 19652
rect 9692 19166 9720 19646
rect 9680 19160 9732 19166
rect 9680 19102 9732 19108
rect 9680 18616 9732 18622
rect 9680 18558 9732 18564
rect 9692 18078 9720 18558
rect 9784 18486 9812 22056
rect 10232 19568 10284 19574
rect 10232 19510 10284 19516
rect 10244 19234 10272 19510
rect 9956 19228 10008 19234
rect 9956 19170 10008 19176
rect 10232 19228 10284 19234
rect 10232 19170 10284 19176
rect 9772 18480 9824 18486
rect 9772 18422 9824 18428
rect 9968 18078 9996 19170
rect 10140 19160 10192 19166
rect 10140 19102 10192 19108
rect 10152 18826 10180 19102
rect 10336 19001 10364 22056
rect 10416 19024 10468 19030
rect 10322 18992 10378 19001
rect 10416 18966 10468 18972
rect 10322 18927 10378 18936
rect 10140 18820 10192 18826
rect 10140 18762 10192 18768
rect 10140 18616 10192 18622
rect 10428 18604 10456 18966
rect 10192 18576 10456 18604
rect 10140 18558 10192 18564
rect 10888 18078 10916 22056
rect 11440 20746 11468 22056
rect 11440 20718 11928 20746
rect 11352 20556 11648 20576
rect 11408 20554 11432 20556
rect 11488 20554 11512 20556
rect 11568 20554 11592 20556
rect 11430 20502 11432 20554
rect 11494 20502 11506 20554
rect 11568 20502 11570 20554
rect 11408 20500 11432 20502
rect 11488 20500 11512 20502
rect 11568 20500 11592 20502
rect 11352 20480 11648 20500
rect 11352 19468 11648 19488
rect 11408 19466 11432 19468
rect 11488 19466 11512 19468
rect 11568 19466 11592 19468
rect 11430 19414 11432 19466
rect 11494 19414 11506 19466
rect 11568 19414 11570 19466
rect 11408 19412 11432 19414
rect 11488 19412 11512 19414
rect 11568 19412 11592 19414
rect 11352 19392 11648 19412
rect 11060 19160 11112 19166
rect 10980 19120 11060 19148
rect 10980 19030 11008 19120
rect 11060 19102 11112 19108
rect 11150 19128 11206 19137
rect 11150 19063 11152 19072
rect 11204 19063 11206 19072
rect 11612 19092 11664 19098
rect 11152 19034 11204 19040
rect 11612 19034 11664 19040
rect 10968 19024 11020 19030
rect 10968 18966 11020 18972
rect 11624 18826 11652 19034
rect 11428 18820 11480 18826
rect 11428 18762 11480 18768
rect 11612 18820 11664 18826
rect 11612 18762 11664 18768
rect 11440 18729 11468 18762
rect 11426 18720 11482 18729
rect 10968 18684 11020 18690
rect 11426 18655 11482 18664
rect 10968 18626 11020 18632
rect 10980 18282 11008 18626
rect 11242 18584 11298 18593
rect 11624 18570 11652 18762
rect 11624 18542 11744 18570
rect 11242 18519 11298 18528
rect 10968 18276 11020 18282
rect 10968 18218 11020 18224
rect 9680 18072 9732 18078
rect 9680 18014 9732 18020
rect 9772 18072 9824 18078
rect 9772 18014 9824 18020
rect 9956 18072 10008 18078
rect 9956 18014 10008 18020
rect 10876 18072 10928 18078
rect 10876 18014 10928 18020
rect 9220 17732 9272 17738
rect 9220 17674 9272 17680
rect 8944 17392 8996 17398
rect 8944 17334 8996 17340
rect 8668 17052 8720 17058
rect 8668 16994 8720 17000
rect 8392 16848 8444 16854
rect 8392 16790 8444 16796
rect 7886 16748 8182 16768
rect 7942 16746 7966 16748
rect 8022 16746 8046 16748
rect 8102 16746 8126 16748
rect 7964 16694 7966 16746
rect 8028 16694 8040 16746
rect 8102 16694 8104 16746
rect 7942 16692 7966 16694
rect 8022 16692 8046 16694
rect 8102 16692 8126 16694
rect 7886 16672 8182 16692
rect 7472 15964 7524 15970
rect 7576 15958 7696 15986
rect 7472 15906 7524 15912
rect 7380 14808 7432 14814
rect 7380 14750 7432 14756
rect 7392 14474 7420 14750
rect 7380 14468 7432 14474
rect 7380 14410 7432 14416
rect 7196 14400 7248 14406
rect 7196 14342 7248 14348
rect 6828 14264 6880 14270
rect 6880 14212 6960 14218
rect 6828 14206 6960 14212
rect 6840 14190 6960 14206
rect 6932 13930 6960 14190
rect 7208 13930 7236 14342
rect 6920 13924 6972 13930
rect 6920 13866 6972 13872
rect 7196 13924 7248 13930
rect 7196 13866 7248 13872
rect 6932 13182 6960 13866
rect 6920 13176 6972 13182
rect 6920 13118 6972 13124
rect 6644 11748 6696 11754
rect 6644 11690 6696 11696
rect 7484 11210 7512 15906
rect 7668 15494 7696 15958
rect 8404 15902 8432 16790
rect 8680 16582 8708 16994
rect 8668 16576 8720 16582
rect 8668 16518 8720 16524
rect 8956 15970 8984 17334
rect 9692 16310 9720 18014
rect 9784 17126 9812 18014
rect 9864 17596 9916 17602
rect 9864 17538 9916 17544
rect 9772 17120 9824 17126
rect 9772 17062 9824 17068
rect 9876 16990 9904 17538
rect 10980 17534 11008 18218
rect 11256 18010 11284 18519
rect 11352 18380 11648 18400
rect 11408 18378 11432 18380
rect 11488 18378 11512 18380
rect 11568 18378 11592 18380
rect 11430 18326 11432 18378
rect 11494 18326 11506 18378
rect 11568 18326 11570 18378
rect 11408 18324 11432 18326
rect 11488 18324 11512 18326
rect 11568 18324 11592 18326
rect 11352 18304 11648 18324
rect 11610 18176 11666 18185
rect 11716 18146 11744 18542
rect 11610 18111 11666 18120
rect 11704 18140 11756 18146
rect 11624 18026 11652 18111
rect 11704 18082 11756 18088
rect 11244 18004 11296 18010
rect 11624 17998 11744 18026
rect 11244 17946 11296 17952
rect 11152 17936 11204 17942
rect 11152 17878 11204 17884
rect 10968 17528 11020 17534
rect 10968 17470 11020 17476
rect 10968 17120 11020 17126
rect 10968 17062 11020 17068
rect 9864 16984 9916 16990
rect 9864 16926 9916 16932
rect 10876 16984 10928 16990
rect 10876 16926 10928 16932
rect 9680 16304 9732 16310
rect 9680 16246 9732 16252
rect 9692 15970 9720 16246
rect 8944 15964 8996 15970
rect 8944 15906 8996 15912
rect 9680 15964 9732 15970
rect 9680 15906 9732 15912
rect 8208 15896 8260 15902
rect 8208 15838 8260 15844
rect 8392 15896 8444 15902
rect 8392 15838 8444 15844
rect 7748 15828 7800 15834
rect 7748 15770 7800 15776
rect 7656 15488 7708 15494
rect 7576 15436 7656 15442
rect 7576 15430 7708 15436
rect 7576 15414 7696 15430
rect 7576 14814 7604 15414
rect 7760 15358 7788 15770
rect 7886 15660 8182 15680
rect 7942 15658 7966 15660
rect 8022 15658 8046 15660
rect 8102 15658 8126 15660
rect 7964 15606 7966 15658
rect 8028 15606 8040 15658
rect 8102 15606 8104 15658
rect 7942 15604 7966 15606
rect 8022 15604 8046 15606
rect 8102 15604 8126 15606
rect 7886 15584 8182 15604
rect 8116 15420 8168 15426
rect 8116 15362 8168 15368
rect 7656 15352 7708 15358
rect 7656 15294 7708 15300
rect 7748 15352 7800 15358
rect 7748 15294 7800 15300
rect 7668 15018 7696 15294
rect 7656 15012 7708 15018
rect 7656 14954 7708 14960
rect 7656 14876 7708 14882
rect 7656 14818 7708 14824
rect 7564 14808 7616 14814
rect 7564 14750 7616 14756
rect 7668 14406 7696 14818
rect 7656 14400 7708 14406
rect 7656 14342 7708 14348
rect 7760 14218 7788 15294
rect 8128 14882 8156 15362
rect 8116 14876 8168 14882
rect 8116 14818 8168 14824
rect 8220 14678 8248 15838
rect 8392 14740 8444 14746
rect 8392 14682 8444 14688
rect 8208 14672 8260 14678
rect 8208 14614 8260 14620
rect 7886 14572 8182 14592
rect 7942 14570 7966 14572
rect 8022 14570 8046 14572
rect 8102 14570 8126 14572
rect 7964 14518 7966 14570
rect 8028 14518 8040 14570
rect 8102 14518 8104 14570
rect 7942 14516 7966 14518
rect 8022 14516 8046 14518
rect 8102 14516 8126 14518
rect 7886 14496 8182 14516
rect 7760 14202 7880 14218
rect 7760 14196 7892 14202
rect 7760 14190 7840 14196
rect 7840 14138 7892 14144
rect 8024 14128 8076 14134
rect 8024 14070 8076 14076
rect 8036 13930 8064 14070
rect 8024 13924 8076 13930
rect 8024 13866 8076 13872
rect 8036 13794 8064 13866
rect 8024 13788 8076 13794
rect 8024 13730 8076 13736
rect 7886 13484 8182 13504
rect 7942 13482 7966 13484
rect 8022 13482 8046 13484
rect 8102 13482 8126 13484
rect 7964 13430 7966 13482
rect 8028 13430 8040 13482
rect 8102 13430 8104 13482
rect 7942 13428 7966 13430
rect 8022 13428 8046 13430
rect 8102 13428 8126 13430
rect 7886 13408 8182 13428
rect 7748 13176 7800 13182
rect 7748 13118 7800 13124
rect 7760 12842 7788 13118
rect 7748 12836 7800 12842
rect 7748 12778 7800 12784
rect 7760 12502 7788 12778
rect 8220 12638 8248 14614
rect 8404 14406 8432 14682
rect 8392 14400 8444 14406
rect 8392 14342 8444 14348
rect 9680 14332 9732 14338
rect 9680 14274 9732 14280
rect 8392 14264 8444 14270
rect 8392 14206 8444 14212
rect 9496 14264 9548 14270
rect 9496 14206 9548 14212
rect 8404 13930 8432 14206
rect 9220 14128 9272 14134
rect 9220 14070 9272 14076
rect 8392 13924 8444 13930
rect 8392 13866 8444 13872
rect 9036 13788 9088 13794
rect 9036 13730 9088 13736
rect 8760 13584 8812 13590
rect 8760 13526 8812 13532
rect 8772 13386 8800 13526
rect 8760 13380 8812 13386
rect 8760 13322 8812 13328
rect 9048 13318 9076 13730
rect 9232 13726 9260 14070
rect 9220 13720 9272 13726
rect 9220 13662 9272 13668
rect 9508 13538 9536 14206
rect 9416 13510 9536 13538
rect 9036 13312 9088 13318
rect 9036 13254 9088 13260
rect 9416 13250 9444 13510
rect 9496 13380 9548 13386
rect 9496 13322 9548 13328
rect 9404 13244 9456 13250
rect 9404 13186 9456 13192
rect 8208 12632 8260 12638
rect 8208 12574 8260 12580
rect 7748 12496 7800 12502
rect 7748 12438 7800 12444
rect 8208 12496 8260 12502
rect 8208 12438 8260 12444
rect 7886 12396 8182 12416
rect 7942 12394 7966 12396
rect 8022 12394 8046 12396
rect 8102 12394 8126 12396
rect 7964 12342 7966 12394
rect 8028 12342 8040 12394
rect 8102 12342 8104 12394
rect 7942 12340 7966 12342
rect 8022 12340 8046 12342
rect 8102 12340 8126 12342
rect 7886 12320 8182 12340
rect 8220 11634 8248 12438
rect 8484 12088 8536 12094
rect 8484 12030 8536 12036
rect 8220 11618 8340 11634
rect 8220 11612 8352 11618
rect 8220 11606 8300 11612
rect 7886 11308 8182 11328
rect 7942 11306 7966 11308
rect 8022 11306 8046 11308
rect 8102 11306 8126 11308
rect 7964 11254 7966 11306
rect 8028 11254 8040 11306
rect 8102 11254 8104 11306
rect 7942 11252 7966 11254
rect 8022 11252 8046 11254
rect 8102 11252 8126 11254
rect 7886 11232 8182 11252
rect 7472 11204 7524 11210
rect 7472 11146 7524 11152
rect 4421 10764 4717 10784
rect 4477 10762 4501 10764
rect 4557 10762 4581 10764
rect 4637 10762 4661 10764
rect 4499 10710 4501 10762
rect 4563 10710 4575 10762
rect 4637 10710 4639 10762
rect 4477 10708 4501 10710
rect 4557 10708 4581 10710
rect 4637 10708 4661 10710
rect 4421 10688 4717 10708
rect 7886 10220 8182 10240
rect 7942 10218 7966 10220
rect 8022 10218 8046 10220
rect 8102 10218 8126 10220
rect 7964 10166 7966 10218
rect 8028 10166 8040 10218
rect 8102 10166 8104 10218
rect 7942 10164 7966 10166
rect 8022 10164 8046 10166
rect 8102 10164 8126 10166
rect 7886 10144 8182 10164
rect 8220 10122 8248 11606
rect 8300 11554 8352 11560
rect 8300 11408 8352 11414
rect 8300 11350 8352 11356
rect 8312 10530 8340 11350
rect 8392 10932 8444 10938
rect 8392 10874 8444 10880
rect 8300 10524 8352 10530
rect 8300 10466 8352 10472
rect 8404 10462 8432 10874
rect 8496 10666 8524 12030
rect 9508 11754 9536 13322
rect 9692 12842 9720 14274
rect 9680 12836 9732 12842
rect 9680 12778 9732 12784
rect 9496 11748 9548 11754
rect 9496 11690 9548 11696
rect 8760 11612 8812 11618
rect 8760 11554 8812 11560
rect 8772 11006 8800 11554
rect 9876 11074 9904 16926
rect 10508 16916 10560 16922
rect 10508 16858 10560 16864
rect 10520 16650 10548 16858
rect 10888 16650 10916 16926
rect 10980 16650 11008 17062
rect 10508 16644 10560 16650
rect 10508 16586 10560 16592
rect 10876 16644 10928 16650
rect 10876 16586 10928 16592
rect 10968 16644 11020 16650
rect 10968 16586 11020 16592
rect 11164 16514 11192 17878
rect 11352 17292 11648 17312
rect 11408 17290 11432 17292
rect 11488 17290 11512 17292
rect 11568 17290 11592 17292
rect 11430 17238 11432 17290
rect 11494 17238 11506 17290
rect 11568 17238 11570 17290
rect 11408 17236 11432 17238
rect 11488 17236 11512 17238
rect 11568 17236 11592 17238
rect 11352 17216 11648 17236
rect 11152 16508 11204 16514
rect 11152 16450 11204 16456
rect 10324 16304 10376 16310
rect 10324 16246 10376 16252
rect 10336 15902 10364 16246
rect 11352 16204 11648 16224
rect 11408 16202 11432 16204
rect 11488 16202 11512 16204
rect 11568 16202 11592 16204
rect 11430 16150 11432 16202
rect 11494 16150 11506 16202
rect 11568 16150 11570 16202
rect 11408 16148 11432 16150
rect 11488 16148 11512 16150
rect 11568 16148 11592 16150
rect 11352 16128 11648 16148
rect 10324 15896 10376 15902
rect 10324 15838 10376 15844
rect 11352 15116 11648 15136
rect 11408 15114 11432 15116
rect 11488 15114 11512 15116
rect 11568 15114 11592 15116
rect 11430 15062 11432 15114
rect 11494 15062 11506 15114
rect 11568 15062 11570 15114
rect 11408 15060 11432 15062
rect 11488 15060 11512 15062
rect 11568 15060 11592 15062
rect 11352 15040 11648 15060
rect 10140 14876 10192 14882
rect 10140 14818 10192 14824
rect 10152 14406 10180 14818
rect 10968 14740 11020 14746
rect 10968 14682 11020 14688
rect 10140 14400 10192 14406
rect 10140 14342 10192 14348
rect 10600 13584 10652 13590
rect 10600 13526 10652 13532
rect 10612 12706 10640 13526
rect 10980 13386 11008 14682
rect 11352 14028 11648 14048
rect 11408 14026 11432 14028
rect 11488 14026 11512 14028
rect 11568 14026 11592 14028
rect 11430 13974 11432 14026
rect 11494 13974 11506 14026
rect 11568 13974 11570 14026
rect 11408 13972 11432 13974
rect 11488 13972 11512 13974
rect 11568 13972 11592 13974
rect 11352 13952 11648 13972
rect 10968 13380 11020 13386
rect 10968 13322 11020 13328
rect 10980 12842 11008 13322
rect 11352 12940 11648 12960
rect 11408 12938 11432 12940
rect 11488 12938 11512 12940
rect 11568 12938 11592 12940
rect 11430 12886 11432 12938
rect 11494 12886 11506 12938
rect 11568 12886 11570 12938
rect 11408 12884 11432 12886
rect 11488 12884 11512 12886
rect 11568 12884 11592 12886
rect 11352 12864 11648 12884
rect 10968 12836 11020 12842
rect 10968 12778 11020 12784
rect 10600 12700 10652 12706
rect 10600 12642 10652 12648
rect 10968 12632 11020 12638
rect 10968 12574 11020 12580
rect 10980 12298 11008 12574
rect 11060 12564 11112 12570
rect 11060 12506 11112 12512
rect 10968 12292 11020 12298
rect 10968 12234 11020 12240
rect 10508 12156 10560 12162
rect 10508 12098 10560 12104
rect 9956 11476 10008 11482
rect 9956 11418 10008 11424
rect 9864 11068 9916 11074
rect 9864 11010 9916 11016
rect 9968 11006 9996 11418
rect 10520 11210 10548 12098
rect 11072 12094 11100 12506
rect 11336 12496 11388 12502
rect 11336 12438 11388 12444
rect 11060 12088 11112 12094
rect 11348 12042 11376 12438
rect 11060 12030 11112 12036
rect 11072 11754 11100 12030
rect 11256 12014 11376 12042
rect 11256 11754 11284 12014
rect 11352 11852 11648 11872
rect 11408 11850 11432 11852
rect 11488 11850 11512 11852
rect 11568 11850 11592 11852
rect 11430 11798 11432 11850
rect 11494 11798 11506 11850
rect 11568 11798 11570 11850
rect 11408 11796 11432 11798
rect 11488 11796 11512 11798
rect 11568 11796 11592 11798
rect 11352 11776 11648 11796
rect 11060 11748 11112 11754
rect 11060 11690 11112 11696
rect 11244 11748 11296 11754
rect 11244 11690 11296 11696
rect 11256 11414 11284 11690
rect 11244 11408 11296 11414
rect 11244 11350 11296 11356
rect 10508 11204 10560 11210
rect 10508 11146 10560 11152
rect 10876 11068 10928 11074
rect 10876 11010 10928 11016
rect 11152 11068 11204 11074
rect 11152 11010 11204 11016
rect 8760 11000 8812 11006
rect 8760 10942 8812 10948
rect 9956 11000 10008 11006
rect 9956 10942 10008 10948
rect 8484 10660 8536 10666
rect 8484 10602 8536 10608
rect 8392 10456 8444 10462
rect 8392 10398 8444 10404
rect 8208 10116 8260 10122
rect 8208 10058 8260 10064
rect 4421 9676 4717 9696
rect 4477 9674 4501 9676
rect 4557 9674 4581 9676
rect 4637 9674 4661 9676
rect 4499 9622 4501 9674
rect 4563 9622 4575 9674
rect 4637 9622 4639 9674
rect 4477 9620 4501 9622
rect 4557 9620 4581 9622
rect 4637 9620 4661 9622
rect 4421 9600 4717 9620
rect 8220 9594 8248 10058
rect 8772 9986 8800 10942
rect 9968 10530 9996 10942
rect 10888 10530 10916 11010
rect 11164 10666 11192 11010
rect 11716 10954 11744 17998
rect 11900 17942 11928 20718
rect 11796 17936 11848 17942
rect 11796 17878 11848 17884
rect 11888 17936 11940 17942
rect 11888 17878 11940 17884
rect 11808 17738 11836 17878
rect 11796 17732 11848 17738
rect 11796 17674 11848 17680
rect 11796 16848 11848 16854
rect 11796 16790 11848 16796
rect 11808 16650 11836 16790
rect 11796 16644 11848 16650
rect 11796 16586 11848 16592
rect 11716 10926 11928 10954
rect 11704 10864 11756 10870
rect 11704 10806 11756 10812
rect 11352 10764 11648 10784
rect 11408 10762 11432 10764
rect 11488 10762 11512 10764
rect 11568 10762 11592 10764
rect 11430 10710 11432 10762
rect 11494 10710 11506 10762
rect 11568 10710 11570 10762
rect 11408 10708 11432 10710
rect 11488 10708 11512 10710
rect 11568 10708 11592 10710
rect 11352 10688 11648 10708
rect 11152 10660 11204 10666
rect 11152 10602 11204 10608
rect 11716 10530 11744 10806
rect 9956 10524 10008 10530
rect 9956 10466 10008 10472
rect 10876 10524 10928 10530
rect 10876 10466 10928 10472
rect 11704 10524 11756 10530
rect 11704 10466 11756 10472
rect 9968 10122 9996 10466
rect 9956 10116 10008 10122
rect 9956 10058 10008 10064
rect 8760 9980 8812 9986
rect 8760 9922 8812 9928
rect 11352 9676 11648 9696
rect 11408 9674 11432 9676
rect 11488 9674 11512 9676
rect 11568 9674 11592 9676
rect 11430 9622 11432 9674
rect 11494 9622 11506 9674
rect 11568 9622 11570 9674
rect 11408 9620 11432 9622
rect 11488 9620 11512 9622
rect 11568 9620 11592 9622
rect 11352 9600 11648 9620
rect 8220 9566 8340 9594
rect 11716 9578 11744 10466
rect 7886 9132 8182 9152
rect 7942 9130 7966 9132
rect 8022 9130 8046 9132
rect 8102 9130 8126 9132
rect 7964 9078 7966 9130
rect 8028 9078 8040 9130
rect 8102 9078 8104 9130
rect 7942 9076 7966 9078
rect 8022 9076 8046 9078
rect 8102 9076 8126 9078
rect 7886 9056 8182 9076
rect 4421 8588 4717 8608
rect 4477 8586 4501 8588
rect 4557 8586 4581 8588
rect 4637 8586 4661 8588
rect 4499 8534 4501 8586
rect 4563 8534 4575 8586
rect 4637 8534 4639 8586
rect 4477 8532 4501 8534
rect 4557 8532 4581 8534
rect 4637 8532 4661 8534
rect 4421 8512 4717 8532
rect 7886 8044 8182 8064
rect 7942 8042 7966 8044
rect 8022 8042 8046 8044
rect 8102 8042 8126 8044
rect 7964 7990 7966 8042
rect 8028 7990 8040 8042
rect 8102 7990 8104 8042
rect 7942 7988 7966 7990
rect 8022 7988 8046 7990
rect 8102 7988 8126 7990
rect 7886 7968 8182 7988
rect 4421 7500 4717 7520
rect 4477 7498 4501 7500
rect 4557 7498 4581 7500
rect 4637 7498 4661 7500
rect 4499 7446 4501 7498
rect 4563 7446 4575 7498
rect 4637 7446 4639 7498
rect 4477 7444 4501 7446
rect 4557 7444 4581 7446
rect 4637 7444 4661 7446
rect 4421 7424 4717 7444
rect 8312 7266 8340 9566
rect 11704 9572 11756 9578
rect 11704 9514 11756 9520
rect 11704 8892 11756 8898
rect 11704 8834 11756 8840
rect 11352 8588 11648 8608
rect 11408 8586 11432 8588
rect 11488 8586 11512 8588
rect 11568 8586 11592 8588
rect 11430 8534 11432 8586
rect 11494 8534 11506 8586
rect 11568 8534 11570 8586
rect 11408 8532 11432 8534
rect 11488 8532 11512 8534
rect 11568 8532 11592 8534
rect 11352 8512 11648 8532
rect 11716 8354 11744 8834
rect 11704 8348 11756 8354
rect 11704 8290 11756 8296
rect 11060 8280 11112 8286
rect 11060 8222 11112 8228
rect 11072 7946 11100 8222
rect 11060 7940 11112 7946
rect 11060 7882 11112 7888
rect 11244 7736 11296 7742
rect 11244 7678 11296 7684
rect 11704 7736 11756 7742
rect 11704 7678 11756 7684
rect 8300 7260 8352 7266
rect 8300 7202 8352 7208
rect 7886 6956 8182 6976
rect 7942 6954 7966 6956
rect 8022 6954 8046 6956
rect 8102 6954 8126 6956
rect 7964 6902 7966 6954
rect 8028 6902 8040 6954
rect 8102 6902 8104 6954
rect 7942 6900 7966 6902
rect 8022 6900 8046 6902
rect 8102 6900 8126 6902
rect 7886 6880 8182 6900
rect 8312 6654 8340 7202
rect 10140 7124 10192 7130
rect 10140 7066 10192 7072
rect 8300 6648 8352 6654
rect 8300 6590 8352 6596
rect 10152 6586 10180 7066
rect 11256 6858 11284 7678
rect 11352 7500 11648 7520
rect 11408 7498 11432 7500
rect 11488 7498 11512 7500
rect 11568 7498 11592 7500
rect 11430 7446 11432 7498
rect 11494 7446 11506 7498
rect 11568 7446 11570 7498
rect 11408 7444 11432 7446
rect 11488 7444 11512 7446
rect 11568 7444 11592 7446
rect 11352 7424 11648 7444
rect 11716 7402 11744 7678
rect 11900 7402 11928 10926
rect 12084 9034 12112 22056
rect 12532 19160 12584 19166
rect 12532 19102 12584 19108
rect 12544 19030 12572 19102
rect 12532 19024 12584 19030
rect 12532 18966 12584 18972
rect 12440 18684 12492 18690
rect 12440 18626 12492 18632
rect 12452 18282 12480 18626
rect 12530 18584 12586 18593
rect 12530 18519 12586 18528
rect 12544 18282 12572 18519
rect 12440 18276 12492 18282
rect 12440 18218 12492 18224
rect 12532 18276 12584 18282
rect 12532 18218 12584 18224
rect 12532 17936 12584 17942
rect 12532 17878 12584 17884
rect 12544 17738 12572 17878
rect 12532 17732 12584 17738
rect 12532 17674 12584 17680
rect 12164 17052 12216 17058
rect 12164 16994 12216 17000
rect 12176 15834 12204 16994
rect 12532 16916 12584 16922
rect 12532 16858 12584 16864
rect 12544 16582 12572 16858
rect 12532 16576 12584 16582
rect 12532 16518 12584 16524
rect 12164 15828 12216 15834
rect 12164 15770 12216 15776
rect 12256 14128 12308 14134
rect 12256 14070 12308 14076
rect 12268 13794 12296 14070
rect 12256 13788 12308 13794
rect 12256 13730 12308 13736
rect 12440 13652 12492 13658
rect 12440 13594 12492 13600
rect 12452 13182 12480 13594
rect 12440 13176 12492 13182
rect 12440 13118 12492 13124
rect 12452 12842 12480 13118
rect 12440 12836 12492 12842
rect 12440 12778 12492 12784
rect 12348 11408 12400 11414
rect 12348 11350 12400 11356
rect 12360 10666 12388 11350
rect 12348 10660 12400 10666
rect 12348 10602 12400 10608
rect 12360 10462 12388 10602
rect 12348 10456 12400 10462
rect 12348 10398 12400 10404
rect 12072 9028 12124 9034
rect 12072 8970 12124 8976
rect 11704 7396 11756 7402
rect 11704 7338 11756 7344
rect 11888 7396 11940 7402
rect 11888 7338 11940 7344
rect 11900 6858 11928 7338
rect 11244 6852 11296 6858
rect 11244 6794 11296 6800
rect 11888 6852 11940 6858
rect 11888 6794 11940 6800
rect 12532 6784 12584 6790
rect 12532 6726 12584 6732
rect 10140 6580 10192 6586
rect 10140 6522 10192 6528
rect 12544 6518 12572 6726
rect 4068 6512 4120 6518
rect 4068 6454 4120 6460
rect 12532 6512 12584 6518
rect 12532 6454 12584 6460
rect 4080 5673 4108 6454
rect 4421 6412 4717 6432
rect 4477 6410 4501 6412
rect 4557 6410 4581 6412
rect 4637 6410 4661 6412
rect 4499 6358 4501 6410
rect 4563 6358 4575 6410
rect 4637 6358 4639 6410
rect 4477 6356 4501 6358
rect 4557 6356 4581 6358
rect 4637 6356 4661 6358
rect 4421 6336 4717 6356
rect 11352 6412 11648 6432
rect 11408 6410 11432 6412
rect 11488 6410 11512 6412
rect 11568 6410 11592 6412
rect 11430 6358 11432 6410
rect 11494 6358 11506 6410
rect 11568 6358 11570 6410
rect 11408 6356 11432 6358
rect 11488 6356 11512 6358
rect 11568 6356 11592 6358
rect 11352 6336 11648 6356
rect 7886 5868 8182 5888
rect 7942 5866 7966 5868
rect 8022 5866 8046 5868
rect 8102 5866 8126 5868
rect 7964 5814 7966 5866
rect 8028 5814 8040 5866
rect 8102 5814 8104 5866
rect 7942 5812 7966 5814
rect 8022 5812 8046 5814
rect 8102 5812 8126 5814
rect 7886 5792 8182 5812
rect 4066 5664 4122 5673
rect 4066 5599 4122 5608
rect 4421 5324 4717 5344
rect 4477 5322 4501 5324
rect 4557 5322 4581 5324
rect 4637 5322 4661 5324
rect 4499 5270 4501 5322
rect 4563 5270 4575 5322
rect 4637 5270 4639 5322
rect 4477 5268 4501 5270
rect 4557 5268 4581 5270
rect 4637 5268 4661 5270
rect 4421 5248 4717 5268
rect 11352 5324 11648 5344
rect 11408 5322 11432 5324
rect 11488 5322 11512 5324
rect 11568 5322 11592 5324
rect 11430 5270 11432 5322
rect 11494 5270 11506 5322
rect 11568 5270 11570 5322
rect 11408 5268 11432 5270
rect 11488 5268 11512 5270
rect 11568 5268 11592 5270
rect 11352 5248 11648 5268
rect 12544 5226 12572 6454
rect 12636 5770 12664 22056
rect 12992 19160 13044 19166
rect 12992 19102 13044 19108
rect 12900 19024 12952 19030
rect 12900 18966 12952 18972
rect 12716 18684 12768 18690
rect 12716 18626 12768 18632
rect 12728 17942 12756 18626
rect 12912 18162 12940 18966
rect 13004 18622 13032 19102
rect 12992 18616 13044 18622
rect 12992 18558 13044 18564
rect 12912 18134 13032 18162
rect 12900 18004 12952 18010
rect 12900 17946 12952 17952
rect 12716 17936 12768 17942
rect 12716 17878 12768 17884
rect 12728 16990 12756 17878
rect 12716 16984 12768 16990
rect 12716 16926 12768 16932
rect 12728 13250 12756 16926
rect 12808 14672 12860 14678
rect 12808 14614 12860 14620
rect 12820 14406 12848 14614
rect 12808 14400 12860 14406
rect 12808 14342 12860 14348
rect 12808 13652 12860 13658
rect 12808 13594 12860 13600
rect 12820 13318 12848 13594
rect 12808 13312 12860 13318
rect 12808 13254 12860 13260
rect 12716 13244 12768 13250
rect 12716 13186 12768 13192
rect 12912 6314 12940 17946
rect 13004 13318 13032 18134
rect 13084 14264 13136 14270
rect 13084 14206 13136 14212
rect 12992 13312 13044 13318
rect 12992 13254 13044 13260
rect 13096 13182 13124 14206
rect 13084 13176 13136 13182
rect 13084 13118 13136 13124
rect 13084 12292 13136 12298
rect 13084 12234 13136 12240
rect 13096 11618 13124 12234
rect 13084 11612 13136 11618
rect 13084 11554 13136 11560
rect 13096 11210 13124 11554
rect 13084 11204 13136 11210
rect 13084 11146 13136 11152
rect 13096 10002 13124 11146
rect 13004 9974 13124 10002
rect 13004 9238 13032 9974
rect 13084 9912 13136 9918
rect 13084 9854 13136 9860
rect 13096 9374 13124 9854
rect 13084 9368 13136 9374
rect 13084 9310 13136 9316
rect 12992 9232 13044 9238
rect 12992 9174 13044 9180
rect 13004 7810 13032 9174
rect 13188 9034 13216 22056
rect 13544 19092 13596 19098
rect 13544 19034 13596 19040
rect 13556 18622 13584 19034
rect 13544 18616 13596 18622
rect 13544 18558 13596 18564
rect 13268 16440 13320 16446
rect 13268 16382 13320 16388
rect 13280 16106 13308 16382
rect 13268 16100 13320 16106
rect 13268 16042 13320 16048
rect 13556 15902 13584 18558
rect 13740 18010 13768 22056
rect 14188 19772 14240 19778
rect 14188 19714 14240 19720
rect 14004 19568 14056 19574
rect 14004 19510 14056 19516
rect 14016 19001 14044 19510
rect 14096 19024 14148 19030
rect 14002 18992 14058 19001
rect 14096 18966 14148 18972
rect 14002 18927 14058 18936
rect 14108 18758 14136 18966
rect 14096 18752 14148 18758
rect 14096 18694 14148 18700
rect 13912 18480 13964 18486
rect 13912 18422 13964 18428
rect 13924 18146 13952 18422
rect 14108 18146 14136 18694
rect 13912 18140 13964 18146
rect 13912 18082 13964 18088
rect 14096 18140 14148 18146
rect 14096 18082 14148 18088
rect 14200 18026 14228 19714
rect 14292 18690 14320 22056
rect 14844 20202 14872 22056
rect 14384 20174 14872 20202
rect 14280 18684 14332 18690
rect 14280 18626 14332 18632
rect 13728 18004 13780 18010
rect 13728 17946 13780 17952
rect 14016 17998 14228 18026
rect 14016 16514 14044 17998
rect 14384 17210 14412 20174
rect 14817 20012 15113 20032
rect 14873 20010 14897 20012
rect 14953 20010 14977 20012
rect 15033 20010 15057 20012
rect 14895 19958 14897 20010
rect 14959 19958 14971 20010
rect 15033 19958 15035 20010
rect 14873 19956 14897 19958
rect 14953 19956 14977 19958
rect 15033 19956 15057 19958
rect 14817 19936 15113 19956
rect 14740 19636 14792 19642
rect 14740 19578 14792 19584
rect 14752 19098 14780 19578
rect 14740 19092 14792 19098
rect 14740 19034 14792 19040
rect 14752 18826 14780 19034
rect 14817 18924 15113 18944
rect 14873 18922 14897 18924
rect 14953 18922 14977 18924
rect 15033 18922 15057 18924
rect 14895 18870 14897 18922
rect 14959 18870 14971 18922
rect 15033 18870 15035 18922
rect 14873 18868 14897 18870
rect 14953 18868 14977 18870
rect 15033 18868 15057 18870
rect 14817 18848 15113 18868
rect 14740 18820 14792 18826
rect 14740 18762 14792 18768
rect 15292 18276 15344 18282
rect 15292 18218 15344 18224
rect 14740 18004 14792 18010
rect 14740 17946 14792 17952
rect 14200 17182 14412 17210
rect 14004 16508 14056 16514
rect 14004 16450 14056 16456
rect 13544 15896 13596 15902
rect 13544 15838 13596 15844
rect 13556 14134 13584 15838
rect 13728 14332 13780 14338
rect 13728 14274 13780 14280
rect 13544 14128 13596 14134
rect 13544 14070 13596 14076
rect 13740 12842 13768 14274
rect 13820 14196 13872 14202
rect 13820 14138 13872 14144
rect 13832 13794 13860 14138
rect 13820 13788 13872 13794
rect 13820 13730 13872 13736
rect 13912 13312 13964 13318
rect 13912 13254 13964 13260
rect 13820 13040 13872 13046
rect 13820 12982 13872 12988
rect 13728 12836 13780 12842
rect 13728 12778 13780 12784
rect 13636 12020 13688 12026
rect 13636 11962 13688 11968
rect 13544 11952 13596 11958
rect 13544 11894 13596 11900
rect 13452 10320 13504 10326
rect 13452 10262 13504 10268
rect 13464 10122 13492 10262
rect 13556 10122 13584 11894
rect 13452 10116 13504 10122
rect 13452 10058 13504 10064
rect 13544 10116 13596 10122
rect 13544 10058 13596 10064
rect 13648 9238 13676 11962
rect 13740 11074 13768 12778
rect 13728 11068 13780 11074
rect 13728 11010 13780 11016
rect 13832 10394 13860 12982
rect 13924 10444 13952 13254
rect 14016 10870 14044 16450
rect 14004 10864 14056 10870
rect 14004 10806 14056 10812
rect 14016 10598 14044 10806
rect 14004 10592 14056 10598
rect 14004 10534 14056 10540
rect 14004 10456 14056 10462
rect 13924 10416 14004 10444
rect 14004 10398 14056 10404
rect 13820 10388 13872 10394
rect 13820 10330 13872 10336
rect 14016 10326 14044 10398
rect 14004 10320 14056 10326
rect 14004 10262 14056 10268
rect 13912 9776 13964 9782
rect 13912 9718 13964 9724
rect 13924 9442 13952 9718
rect 13912 9436 13964 9442
rect 13912 9378 13964 9384
rect 13636 9232 13688 9238
rect 13636 9174 13688 9180
rect 13176 9028 13228 9034
rect 13176 8970 13228 8976
rect 13636 8892 13688 8898
rect 13636 8834 13688 8840
rect 13648 8354 13676 8834
rect 13636 8348 13688 8354
rect 13636 8290 13688 8296
rect 12992 7804 13044 7810
rect 12992 7746 13044 7752
rect 13728 7804 13780 7810
rect 13728 7746 13780 7752
rect 13912 7804 13964 7810
rect 13912 7746 13964 7752
rect 13004 7130 13032 7746
rect 13740 7334 13768 7746
rect 13728 7328 13780 7334
rect 13728 7270 13780 7276
rect 13924 7266 13952 7746
rect 13912 7260 13964 7266
rect 13912 7202 13964 7208
rect 12992 7124 13044 7130
rect 12992 7066 13044 7072
rect 12900 6308 12952 6314
rect 12900 6250 12952 6256
rect 12624 5764 12676 5770
rect 12624 5706 12676 5712
rect 12532 5220 12584 5226
rect 12532 5162 12584 5168
rect 7886 4780 8182 4800
rect 7942 4778 7966 4780
rect 8022 4778 8046 4780
rect 8102 4778 8126 4780
rect 7964 4726 7966 4778
rect 8028 4726 8040 4778
rect 8102 4726 8104 4778
rect 7942 4724 7966 4726
rect 8022 4724 8046 4726
rect 8102 4724 8126 4726
rect 7886 4704 8182 4724
rect 4421 4236 4717 4256
rect 4477 4234 4501 4236
rect 4557 4234 4581 4236
rect 4637 4234 4661 4236
rect 4499 4182 4501 4234
rect 4563 4182 4575 4234
rect 4637 4182 4639 4234
rect 4477 4180 4501 4182
rect 4557 4180 4581 4182
rect 4637 4180 4661 4182
rect 4421 4160 4717 4180
rect 11352 4236 11648 4256
rect 11408 4234 11432 4236
rect 11488 4234 11512 4236
rect 11568 4234 11592 4236
rect 11430 4182 11432 4234
rect 11494 4182 11506 4234
rect 11568 4182 11570 4234
rect 11408 4180 11432 4182
rect 11488 4180 11512 4182
rect 11568 4180 11592 4182
rect 11352 4160 11648 4180
rect 7886 3692 8182 3712
rect 7942 3690 7966 3692
rect 8022 3690 8046 3692
rect 8102 3690 8126 3692
rect 7964 3638 7966 3690
rect 8028 3638 8040 3690
rect 8102 3638 8104 3690
rect 7942 3636 7966 3638
rect 8022 3636 8046 3638
rect 8102 3636 8126 3638
rect 7886 3616 8182 3636
rect 4421 3148 4717 3168
rect 4477 3146 4501 3148
rect 4557 3146 4581 3148
rect 4637 3146 4661 3148
rect 4499 3094 4501 3146
rect 4563 3094 4575 3146
rect 4637 3094 4639 3146
rect 4477 3092 4501 3094
rect 4557 3092 4581 3094
rect 4637 3092 4661 3094
rect 4421 3072 4717 3092
rect 11352 3148 11648 3168
rect 11408 3146 11432 3148
rect 11488 3146 11512 3148
rect 11568 3146 11592 3148
rect 11430 3094 11432 3146
rect 11494 3094 11506 3146
rect 11568 3094 11570 3146
rect 11408 3092 11432 3094
rect 11488 3092 11512 3094
rect 11568 3092 11592 3094
rect 11352 3072 11648 3092
rect 7886 2604 8182 2624
rect 7942 2602 7966 2604
rect 8022 2602 8046 2604
rect 8102 2602 8126 2604
rect 7964 2550 7966 2602
rect 8028 2550 8040 2602
rect 8102 2550 8104 2602
rect 7942 2548 7966 2550
rect 8022 2548 8046 2550
rect 8102 2548 8126 2550
rect 7886 2528 8182 2548
rect 4421 2060 4717 2080
rect 4477 2058 4501 2060
rect 4557 2058 4581 2060
rect 4637 2058 4661 2060
rect 4499 2006 4501 2058
rect 4563 2006 4575 2058
rect 4637 2006 4639 2058
rect 4477 2004 4501 2006
rect 4557 2004 4581 2006
rect 4637 2004 4661 2006
rect 4421 1984 4717 2004
rect 11352 2060 11648 2080
rect 11408 2058 11432 2060
rect 11488 2058 11512 2060
rect 11568 2058 11592 2060
rect 11430 2006 11432 2058
rect 11494 2006 11506 2058
rect 11568 2006 11570 2058
rect 11408 2004 11432 2006
rect 11488 2004 11512 2006
rect 11568 2004 11592 2006
rect 11352 1984 11648 2004
rect 14016 1962 14044 10262
rect 14096 8280 14148 8286
rect 14096 8222 14148 8228
rect 14108 6586 14136 8222
rect 14200 8150 14228 17182
rect 14372 17052 14424 17058
rect 14372 16994 14424 17000
rect 14384 16514 14412 16994
rect 14372 16508 14424 16514
rect 14372 16450 14424 16456
rect 14752 15834 14780 17946
rect 14817 17836 15113 17856
rect 14873 17834 14897 17836
rect 14953 17834 14977 17836
rect 15033 17834 15057 17836
rect 14895 17782 14897 17834
rect 14959 17782 14971 17834
rect 15033 17782 15035 17834
rect 14873 17780 14897 17782
rect 14953 17780 14977 17782
rect 15033 17780 15057 17782
rect 14817 17760 15113 17780
rect 15200 17732 15252 17738
rect 15200 17674 15252 17680
rect 14817 16748 15113 16768
rect 14873 16746 14897 16748
rect 14953 16746 14977 16748
rect 15033 16746 15057 16748
rect 14895 16694 14897 16746
rect 14959 16694 14971 16746
rect 15033 16694 15035 16746
rect 14873 16692 14897 16694
rect 14953 16692 14977 16694
rect 15033 16692 15057 16694
rect 14817 16672 15113 16692
rect 14924 16440 14976 16446
rect 14924 16382 14976 16388
rect 14936 16106 14964 16382
rect 14924 16100 14976 16106
rect 14924 16042 14976 16048
rect 14740 15828 14792 15834
rect 14740 15770 14792 15776
rect 14817 15660 15113 15680
rect 14873 15658 14897 15660
rect 14953 15658 14977 15660
rect 15033 15658 15057 15660
rect 14895 15606 14897 15658
rect 14959 15606 14971 15658
rect 15033 15606 15035 15658
rect 14873 15604 14897 15606
rect 14953 15604 14977 15606
rect 15033 15604 15057 15606
rect 14817 15584 15113 15604
rect 14556 14672 14608 14678
rect 14556 14614 14608 14620
rect 14280 14332 14332 14338
rect 14280 14274 14332 14280
rect 14292 13726 14320 14274
rect 14280 13720 14332 13726
rect 14280 13662 14332 13668
rect 14280 13584 14332 13590
rect 14280 13526 14332 13532
rect 14292 13386 14320 13526
rect 14280 13380 14332 13386
rect 14280 13322 14332 13328
rect 14568 12502 14596 14614
rect 14817 14572 15113 14592
rect 14873 14570 14897 14572
rect 14953 14570 14977 14572
rect 15033 14570 15057 14572
rect 14895 14518 14897 14570
rect 14959 14518 14971 14570
rect 15033 14518 15035 14570
rect 14873 14516 14897 14518
rect 14953 14516 14977 14518
rect 15033 14516 15057 14518
rect 14817 14496 15113 14516
rect 15108 14128 15160 14134
rect 15108 14070 15160 14076
rect 15120 13930 15148 14070
rect 15108 13924 15160 13930
rect 15108 13866 15160 13872
rect 14817 13484 15113 13504
rect 14873 13482 14897 13484
rect 14953 13482 14977 13484
rect 15033 13482 15057 13484
rect 14895 13430 14897 13482
rect 14959 13430 14971 13482
rect 15033 13430 15035 13482
rect 14873 13428 14897 13430
rect 14953 13428 14977 13430
rect 15033 13428 15057 13430
rect 14817 13408 15113 13428
rect 14556 12496 14608 12502
rect 14556 12438 14608 12444
rect 14568 12298 14596 12438
rect 14817 12396 15113 12416
rect 14873 12394 14897 12396
rect 14953 12394 14977 12396
rect 15033 12394 15057 12396
rect 14895 12342 14897 12394
rect 14959 12342 14971 12394
rect 15033 12342 15035 12394
rect 14873 12340 14897 12342
rect 14953 12340 14977 12342
rect 15033 12340 15057 12342
rect 14817 12320 15113 12340
rect 14556 12292 14608 12298
rect 14556 12234 14608 12240
rect 14372 12088 14424 12094
rect 14372 12030 14424 12036
rect 14280 12020 14332 12026
rect 14280 11962 14332 11968
rect 14292 11754 14320 11962
rect 14384 11754 14412 12030
rect 14280 11748 14332 11754
rect 14280 11690 14332 11696
rect 14372 11748 14424 11754
rect 14372 11690 14424 11696
rect 14384 10530 14412 11690
rect 14372 10524 14424 10530
rect 14372 10466 14424 10472
rect 14280 10320 14332 10326
rect 14280 10262 14332 10268
rect 14188 8144 14240 8150
rect 14188 8086 14240 8092
rect 14188 7056 14240 7062
rect 14188 6998 14240 7004
rect 14200 6858 14228 6998
rect 14188 6852 14240 6858
rect 14188 6794 14240 6800
rect 14096 6580 14148 6586
rect 14096 6522 14148 6528
rect 14292 2438 14320 10262
rect 14384 10054 14412 10466
rect 14372 10048 14424 10054
rect 14372 9990 14424 9996
rect 14280 2432 14332 2438
rect 14280 2374 14332 2380
rect 14004 1956 14056 1962
rect 14004 1898 14056 1904
rect 14568 1214 14596 12234
rect 15212 12094 15240 17674
rect 15304 16990 15332 18218
rect 15396 17942 15424 22056
rect 15566 18720 15622 18729
rect 15566 18655 15622 18664
rect 15660 18684 15712 18690
rect 15476 18480 15528 18486
rect 15476 18422 15528 18428
rect 15488 18078 15516 18422
rect 15476 18072 15528 18078
rect 15476 18014 15528 18020
rect 15384 17936 15436 17942
rect 15384 17878 15436 17884
rect 15292 16984 15344 16990
rect 15292 16926 15344 16932
rect 15580 14474 15608 18655
rect 15660 18626 15712 18632
rect 15568 14468 15620 14474
rect 15568 14410 15620 14416
rect 15292 14332 15344 14338
rect 15292 14274 15344 14280
rect 15304 13930 15332 14274
rect 15292 13924 15344 13930
rect 15292 13866 15344 13872
rect 15476 13720 15528 13726
rect 15476 13662 15528 13668
rect 15488 13386 15516 13662
rect 15476 13380 15528 13386
rect 15476 13322 15528 13328
rect 15292 13312 15344 13318
rect 15292 13254 15344 13260
rect 15304 12230 15332 13254
rect 15292 12224 15344 12230
rect 15292 12166 15344 12172
rect 15200 12088 15252 12094
rect 15200 12030 15252 12036
rect 15200 11544 15252 11550
rect 15200 11486 15252 11492
rect 14817 11308 15113 11328
rect 14873 11306 14897 11308
rect 14953 11306 14977 11308
rect 15033 11306 15057 11308
rect 14895 11254 14897 11306
rect 14959 11254 14971 11306
rect 15033 11254 15035 11306
rect 14873 11252 14897 11254
rect 14953 11252 14977 11254
rect 15033 11252 15057 11254
rect 14817 11232 15113 11252
rect 14817 10220 15113 10240
rect 14873 10218 14897 10220
rect 14953 10218 14977 10220
rect 15033 10218 15057 10220
rect 14895 10166 14897 10218
rect 14959 10166 14971 10218
rect 15033 10166 15035 10218
rect 14873 10164 14897 10166
rect 14953 10164 14977 10166
rect 15033 10164 15057 10166
rect 14817 10144 15113 10164
rect 15212 9986 15240 11486
rect 15476 11408 15528 11414
rect 15476 11350 15528 11356
rect 15488 11210 15516 11350
rect 15476 11204 15528 11210
rect 15476 11146 15528 11152
rect 15200 9980 15252 9986
rect 15200 9922 15252 9928
rect 15384 9232 15436 9238
rect 15384 9174 15436 9180
rect 14817 9132 15113 9152
rect 14873 9130 14897 9132
rect 14953 9130 14977 9132
rect 15033 9130 15057 9132
rect 14895 9078 14897 9130
rect 14959 9078 14971 9130
rect 15033 9078 15035 9130
rect 14873 9076 14897 9078
rect 14953 9076 14977 9078
rect 15033 9076 15057 9078
rect 14817 9056 15113 9076
rect 15396 9034 15424 9174
rect 15672 9034 15700 18626
rect 15844 17936 15896 17942
rect 15844 17878 15896 17884
rect 15752 16984 15804 16990
rect 15752 16926 15804 16932
rect 15764 16582 15792 16926
rect 15752 16576 15804 16582
rect 15752 16518 15804 16524
rect 15856 9866 15884 17878
rect 15948 13538 15976 22056
rect 16396 19636 16448 19642
rect 16396 19578 16448 19584
rect 16408 19030 16436 19578
rect 16396 19024 16448 19030
rect 16396 18966 16448 18972
rect 16212 18548 16264 18554
rect 16212 18490 16264 18496
rect 16224 18282 16252 18490
rect 16212 18276 16264 18282
rect 16212 18218 16264 18224
rect 16408 18078 16436 18966
rect 16396 18072 16448 18078
rect 16396 18014 16448 18020
rect 16500 17210 16528 22056
rect 17052 19658 17080 22056
rect 17052 19630 17172 19658
rect 17040 19568 17092 19574
rect 17040 19510 17092 19516
rect 17052 19166 17080 19510
rect 17040 19160 17092 19166
rect 17040 19102 17092 19108
rect 16764 19024 16816 19030
rect 16764 18966 16816 18972
rect 16776 18758 16804 18966
rect 17144 18758 17172 19630
rect 16764 18752 16816 18758
rect 16764 18694 16816 18700
rect 17132 18752 17184 18758
rect 17132 18694 17184 18700
rect 16856 18684 16908 18690
rect 16856 18626 16908 18632
rect 16408 17182 16528 17210
rect 16120 14264 16172 14270
rect 16120 14206 16172 14212
rect 16132 13862 16160 14206
rect 16304 14128 16356 14134
rect 16304 14070 16356 14076
rect 16120 13856 16172 13862
rect 16120 13798 16172 13804
rect 16316 13726 16344 14070
rect 16304 13720 16356 13726
rect 16304 13662 16356 13668
rect 15948 13510 16344 13538
rect 16212 12700 16264 12706
rect 16212 12642 16264 12648
rect 16120 12496 16172 12502
rect 16120 12438 16172 12444
rect 16132 12298 16160 12438
rect 16120 12292 16172 12298
rect 16120 12234 16172 12240
rect 16224 11754 16252 12642
rect 16212 11748 16264 11754
rect 16212 11690 16264 11696
rect 15856 9838 15976 9866
rect 15844 9776 15896 9782
rect 15844 9718 15896 9724
rect 15856 9442 15884 9718
rect 15844 9436 15896 9442
rect 15844 9378 15896 9384
rect 15384 9028 15436 9034
rect 15384 8970 15436 8976
rect 15660 9028 15712 9034
rect 15660 8970 15712 8976
rect 14817 8044 15113 8064
rect 14873 8042 14897 8044
rect 14953 8042 14977 8044
rect 15033 8042 15057 8044
rect 14895 7990 14897 8042
rect 14959 7990 14971 8042
rect 15033 7990 15035 8042
rect 14873 7988 14897 7990
rect 14953 7988 14977 7990
rect 15033 7988 15057 7990
rect 14817 7968 15113 7988
rect 15948 7878 15976 9838
rect 16316 8490 16344 13510
rect 16408 8762 16436 17182
rect 16868 16582 16896 18626
rect 17040 18616 17092 18622
rect 17040 18558 17092 18564
rect 17052 18282 17080 18558
rect 17696 18298 17724 22056
rect 18248 21698 18276 22056
rect 18248 21670 18736 21698
rect 18602 21576 18658 21585
rect 18602 21511 18658 21520
rect 18282 20556 18578 20576
rect 18338 20554 18362 20556
rect 18418 20554 18442 20556
rect 18498 20554 18522 20556
rect 18360 20502 18362 20554
rect 18424 20502 18436 20554
rect 18498 20502 18500 20554
rect 18338 20500 18362 20502
rect 18418 20500 18442 20502
rect 18498 20500 18522 20502
rect 18282 20480 18578 20500
rect 18616 19914 18644 21511
rect 18604 19908 18656 19914
rect 18604 19850 18656 19856
rect 18052 19772 18104 19778
rect 18052 19714 18104 19720
rect 18144 19772 18196 19778
rect 18144 19714 18196 19720
rect 18064 19166 18092 19714
rect 18052 19160 18104 19166
rect 18052 19102 18104 19108
rect 17696 18282 17908 18298
rect 17040 18276 17092 18282
rect 17696 18276 17920 18282
rect 17696 18270 17868 18276
rect 17040 18218 17092 18224
rect 17868 18218 17920 18224
rect 17224 18072 17276 18078
rect 17276 18032 17356 18060
rect 17224 18014 17276 18020
rect 16856 16576 16908 16582
rect 16856 16518 16908 16524
rect 16488 16508 16540 16514
rect 16488 16450 16540 16456
rect 16500 13658 16528 16450
rect 16672 16440 16724 16446
rect 16672 16382 16724 16388
rect 16684 16106 16712 16382
rect 16672 16100 16724 16106
rect 16672 16042 16724 16048
rect 17328 15834 17356 18032
rect 18156 18010 18184 19714
rect 18282 19468 18578 19488
rect 18338 19466 18362 19468
rect 18418 19466 18442 19468
rect 18498 19466 18522 19468
rect 18360 19414 18362 19466
rect 18424 19414 18436 19466
rect 18498 19414 18500 19466
rect 18338 19412 18362 19414
rect 18418 19412 18442 19414
rect 18498 19412 18522 19414
rect 18282 19392 18578 19412
rect 18328 19160 18380 19166
rect 18326 19128 18328 19137
rect 18380 19128 18382 19137
rect 18326 19063 18382 19072
rect 18420 18752 18472 18758
rect 18420 18694 18472 18700
rect 18432 18593 18460 18694
rect 18604 18616 18656 18622
rect 18418 18584 18474 18593
rect 18604 18558 18656 18564
rect 18418 18519 18474 18528
rect 18282 18380 18578 18400
rect 18338 18378 18362 18380
rect 18418 18378 18442 18380
rect 18498 18378 18522 18380
rect 18360 18326 18362 18378
rect 18424 18326 18436 18378
rect 18498 18326 18500 18378
rect 18338 18324 18362 18326
rect 18418 18324 18442 18326
rect 18498 18324 18522 18326
rect 18282 18304 18578 18324
rect 18144 18004 18196 18010
rect 18144 17946 18196 17952
rect 18616 17942 18644 18558
rect 18708 18214 18736 21670
rect 18696 18208 18748 18214
rect 18696 18150 18748 18156
rect 18800 18010 18828 22056
rect 19260 19914 19288 22463
rect 19338 22056 19394 22856
rect 19890 22056 19946 22856
rect 20166 22120 20222 22129
rect 19248 19908 19300 19914
rect 19248 19850 19300 19856
rect 19260 19234 19288 19850
rect 19248 19228 19300 19234
rect 19248 19170 19300 19176
rect 19064 19092 19116 19098
rect 19064 19034 19116 19040
rect 18878 18584 18934 18593
rect 18878 18519 18934 18528
rect 18892 18146 18920 18519
rect 18880 18140 18932 18146
rect 18880 18082 18932 18088
rect 18788 18004 18840 18010
rect 18788 17946 18840 17952
rect 18604 17936 18656 17942
rect 18604 17878 18656 17884
rect 18616 17602 18644 17878
rect 18604 17596 18656 17602
rect 18604 17538 18656 17544
rect 18880 17596 18932 17602
rect 18880 17538 18932 17544
rect 18282 17292 18578 17312
rect 18338 17290 18362 17292
rect 18418 17290 18442 17292
rect 18498 17290 18522 17292
rect 18360 17238 18362 17290
rect 18424 17238 18436 17290
rect 18498 17238 18500 17290
rect 18338 17236 18362 17238
rect 18418 17236 18442 17238
rect 18498 17236 18522 17238
rect 18282 17216 18578 17236
rect 18892 17058 18920 17538
rect 18880 17052 18932 17058
rect 18880 16994 18932 17000
rect 18052 16984 18104 16990
rect 18052 16926 18104 16932
rect 18064 16650 18092 16926
rect 18052 16644 18104 16650
rect 18052 16586 18104 16592
rect 18604 16576 18656 16582
rect 18604 16518 18656 16524
rect 18282 16204 18578 16224
rect 18338 16202 18362 16204
rect 18418 16202 18442 16204
rect 18498 16202 18522 16204
rect 18360 16150 18362 16202
rect 18424 16150 18436 16202
rect 18498 16150 18500 16202
rect 18338 16148 18362 16150
rect 18418 16148 18442 16150
rect 18498 16148 18522 16150
rect 18282 16128 18578 16148
rect 18616 15970 18644 16518
rect 18696 16440 18748 16446
rect 18696 16382 18748 16388
rect 18708 16106 18736 16382
rect 18696 16100 18748 16106
rect 18696 16042 18748 16048
rect 18604 15964 18656 15970
rect 18604 15906 18656 15912
rect 17316 15828 17368 15834
rect 17316 15770 17368 15776
rect 17328 15426 17356 15770
rect 18708 15494 18736 16042
rect 18696 15488 18748 15494
rect 18696 15430 18748 15436
rect 17316 15420 17368 15426
rect 17316 15362 17368 15368
rect 16580 14740 16632 14746
rect 16580 14682 16632 14688
rect 16592 13794 16620 14682
rect 17328 13794 17356 15362
rect 18282 15116 18578 15136
rect 18338 15114 18362 15116
rect 18418 15114 18442 15116
rect 18498 15114 18522 15116
rect 18360 15062 18362 15114
rect 18424 15062 18436 15114
rect 18498 15062 18500 15114
rect 18338 15060 18362 15062
rect 18418 15060 18442 15062
rect 18498 15060 18522 15062
rect 18282 15040 18578 15060
rect 18052 14400 18104 14406
rect 18052 14342 18104 14348
rect 18064 13930 18092 14342
rect 18144 14332 18196 14338
rect 18144 14274 18196 14280
rect 18972 14332 19024 14338
rect 18972 14274 19024 14280
rect 18052 13924 18104 13930
rect 18052 13866 18104 13872
rect 16580 13788 16632 13794
rect 16580 13730 16632 13736
rect 17316 13788 17368 13794
rect 17316 13730 17368 13736
rect 16488 13652 16540 13658
rect 16488 13594 16540 13600
rect 16500 13386 16528 13594
rect 16488 13380 16540 13386
rect 16488 13322 16540 13328
rect 16500 9238 16528 13322
rect 18156 12722 18184 14274
rect 18696 14128 18748 14134
rect 18696 14070 18748 14076
rect 18282 14028 18578 14048
rect 18338 14026 18362 14028
rect 18418 14026 18442 14028
rect 18498 14026 18522 14028
rect 18360 13974 18362 14026
rect 18424 13974 18436 14026
rect 18498 13974 18500 14026
rect 18338 13972 18362 13974
rect 18418 13972 18442 13974
rect 18498 13972 18522 13974
rect 18282 13952 18578 13972
rect 18708 13794 18736 14070
rect 18984 13930 19012 14274
rect 18972 13924 19024 13930
rect 18972 13866 19024 13872
rect 18696 13788 18748 13794
rect 18696 13730 18748 13736
rect 19076 13590 19104 19034
rect 19352 16854 19380 22056
rect 19522 18448 19578 18457
rect 19522 18383 19578 18392
rect 19536 17738 19564 18383
rect 19616 18004 19668 18010
rect 19616 17946 19668 17952
rect 19524 17732 19576 17738
rect 19524 17674 19576 17680
rect 19340 16848 19392 16854
rect 19340 16790 19392 16796
rect 19432 15216 19484 15222
rect 19432 15158 19484 15164
rect 19444 14270 19472 15158
rect 19432 14264 19484 14270
rect 19432 14206 19484 14212
rect 19340 13720 19392 13726
rect 19444 13708 19472 14206
rect 19392 13680 19472 13708
rect 19340 13662 19392 13668
rect 19064 13584 19116 13590
rect 19064 13526 19116 13532
rect 19340 13584 19392 13590
rect 19340 13526 19392 13532
rect 19352 13386 19380 13526
rect 19340 13380 19392 13386
rect 19340 13322 19392 13328
rect 19444 13266 19472 13680
rect 19352 13238 19472 13266
rect 19352 13182 19380 13238
rect 18880 13176 18932 13182
rect 18880 13118 18932 13124
rect 19340 13176 19392 13182
rect 19340 13118 19392 13124
rect 18282 12940 18578 12960
rect 18338 12938 18362 12940
rect 18418 12938 18442 12940
rect 18498 12938 18522 12940
rect 18360 12886 18362 12938
rect 18424 12886 18436 12938
rect 18498 12886 18500 12938
rect 18338 12884 18362 12886
rect 18418 12884 18442 12886
rect 18498 12884 18522 12886
rect 18282 12864 18578 12884
rect 18892 12842 18920 13118
rect 18880 12836 18932 12842
rect 18880 12778 18932 12784
rect 19064 12836 19116 12842
rect 19064 12778 19116 12784
rect 17592 12700 17644 12706
rect 17592 12642 17644 12648
rect 17776 12700 17828 12706
rect 18156 12694 18276 12722
rect 17776 12642 17828 12648
rect 16580 12564 16632 12570
rect 16580 12506 16632 12512
rect 17132 12564 17184 12570
rect 17132 12506 17184 12512
rect 16592 12298 16620 12506
rect 16764 12496 16816 12502
rect 16764 12438 16816 12444
rect 16776 12298 16804 12438
rect 16580 12292 16632 12298
rect 16580 12234 16632 12240
rect 16764 12292 16816 12298
rect 16764 12234 16816 12240
rect 17144 12230 17172 12506
rect 17408 12496 17460 12502
rect 17408 12438 17460 12444
rect 17132 12224 17184 12230
rect 17132 12166 17184 12172
rect 17144 11142 17172 12166
rect 17420 11958 17448 12438
rect 17408 11952 17460 11958
rect 17408 11894 17460 11900
rect 17604 11414 17632 12642
rect 17684 12224 17736 12230
rect 17684 12166 17736 12172
rect 17696 11618 17724 12166
rect 17788 12026 17816 12642
rect 18052 12496 18104 12502
rect 18052 12438 18104 12444
rect 18064 12162 18092 12438
rect 18248 12298 18276 12694
rect 18972 12496 19024 12502
rect 18972 12438 19024 12444
rect 18236 12292 18288 12298
rect 18236 12234 18288 12240
rect 18880 12292 18932 12298
rect 18880 12234 18932 12240
rect 18052 12156 18104 12162
rect 18052 12098 18104 12104
rect 18144 12156 18196 12162
rect 18144 12098 18196 12104
rect 17868 12088 17920 12094
rect 17868 12030 17920 12036
rect 17776 12020 17828 12026
rect 17776 11962 17828 11968
rect 17776 11680 17828 11686
rect 17776 11622 17828 11628
rect 17684 11612 17736 11618
rect 17684 11554 17736 11560
rect 17592 11408 17644 11414
rect 17592 11350 17644 11356
rect 17132 11136 17184 11142
rect 17132 11078 17184 11084
rect 17788 10122 17816 11622
rect 17880 11618 17908 12030
rect 18156 11754 18184 12098
rect 18604 12088 18656 12094
rect 18604 12030 18656 12036
rect 18282 11852 18578 11872
rect 18338 11850 18362 11852
rect 18418 11850 18442 11852
rect 18498 11850 18522 11852
rect 18360 11798 18362 11850
rect 18424 11798 18436 11850
rect 18498 11798 18500 11850
rect 18338 11796 18362 11798
rect 18418 11796 18442 11798
rect 18498 11796 18522 11798
rect 18282 11776 18578 11796
rect 18144 11748 18196 11754
rect 18144 11690 18196 11696
rect 18616 11686 18644 12030
rect 18604 11680 18656 11686
rect 18604 11622 18656 11628
rect 17868 11612 17920 11618
rect 17868 11554 17920 11560
rect 18788 11612 18840 11618
rect 18788 11554 18840 11560
rect 18512 11476 18564 11482
rect 18512 11418 18564 11424
rect 18524 11210 18552 11418
rect 18604 11408 18656 11414
rect 18604 11350 18656 11356
rect 18512 11204 18564 11210
rect 18512 11146 18564 11152
rect 18616 10870 18644 11350
rect 18696 10932 18748 10938
rect 18696 10874 18748 10880
rect 18604 10864 18656 10870
rect 18604 10806 18656 10812
rect 18282 10764 18578 10784
rect 18338 10762 18362 10764
rect 18418 10762 18442 10764
rect 18498 10762 18522 10764
rect 18360 10710 18362 10762
rect 18424 10710 18436 10762
rect 18498 10710 18500 10762
rect 18338 10708 18362 10710
rect 18418 10708 18442 10710
rect 18498 10708 18522 10710
rect 18282 10688 18578 10708
rect 17776 10116 17828 10122
rect 17776 10058 17828 10064
rect 18052 9980 18104 9986
rect 18052 9922 18104 9928
rect 18064 9442 18092 9922
rect 18282 9676 18578 9696
rect 18338 9674 18362 9676
rect 18418 9674 18442 9676
rect 18498 9674 18522 9676
rect 18360 9622 18362 9674
rect 18424 9622 18436 9674
rect 18498 9622 18500 9674
rect 18338 9620 18362 9622
rect 18418 9620 18442 9622
rect 18498 9620 18522 9622
rect 18282 9600 18578 9620
rect 18052 9436 18104 9442
rect 18052 9378 18104 9384
rect 16488 9232 16540 9238
rect 16488 9174 16540 9180
rect 16396 8756 16448 8762
rect 16396 8698 16448 8704
rect 16304 8484 16356 8490
rect 16304 8426 16356 8432
rect 15936 7872 15988 7878
rect 15936 7814 15988 7820
rect 15292 7736 15344 7742
rect 15292 7678 15344 7684
rect 15016 7600 15068 7606
rect 15016 7542 15068 7548
rect 15028 7130 15056 7542
rect 15200 7192 15252 7198
rect 15200 7134 15252 7140
rect 14740 7124 14792 7130
rect 14740 7066 14792 7072
rect 15016 7124 15068 7130
rect 15016 7066 15068 7072
rect 14752 6654 14780 7066
rect 14817 6956 15113 6976
rect 14873 6954 14897 6956
rect 14953 6954 14977 6956
rect 15033 6954 15057 6956
rect 14895 6902 14897 6954
rect 14959 6902 14971 6954
rect 15033 6902 15035 6954
rect 14873 6900 14897 6902
rect 14953 6900 14977 6902
rect 15033 6900 15057 6902
rect 14817 6880 15113 6900
rect 14740 6648 14792 6654
rect 14740 6590 14792 6596
rect 15212 6518 15240 7134
rect 15304 6790 15332 7678
rect 15384 7056 15436 7062
rect 15384 6998 15436 7004
rect 15396 6858 15424 6998
rect 15384 6852 15436 6858
rect 15384 6794 15436 6800
rect 15292 6784 15344 6790
rect 15292 6726 15344 6732
rect 15200 6512 15252 6518
rect 15200 6454 15252 6460
rect 14817 5868 15113 5888
rect 14873 5866 14897 5868
rect 14953 5866 14977 5868
rect 15033 5866 15057 5868
rect 14895 5814 14897 5866
rect 14959 5814 14971 5866
rect 15033 5814 15035 5866
rect 14873 5812 14897 5814
rect 14953 5812 14977 5814
rect 15033 5812 15057 5814
rect 14817 5792 15113 5812
rect 14817 4780 15113 4800
rect 14873 4778 14897 4780
rect 14953 4778 14977 4780
rect 15033 4778 15057 4780
rect 14895 4726 14897 4778
rect 14959 4726 14971 4778
rect 15033 4726 15035 4778
rect 14873 4724 14897 4726
rect 14953 4724 14977 4726
rect 15033 4724 15057 4726
rect 14817 4704 15113 4724
rect 16500 4002 16528 9174
rect 16580 8892 16632 8898
rect 16580 8834 16632 8840
rect 16592 8354 16620 8834
rect 18282 8588 18578 8608
rect 18338 8586 18362 8588
rect 18418 8586 18442 8588
rect 18498 8586 18522 8588
rect 18360 8534 18362 8586
rect 18424 8534 18436 8586
rect 18498 8534 18500 8586
rect 18338 8532 18362 8534
rect 18418 8532 18442 8534
rect 18498 8532 18522 8534
rect 18282 8512 18578 8532
rect 16580 8348 16632 8354
rect 16580 8290 16632 8296
rect 16948 8280 17000 8286
rect 16948 8222 17000 8228
rect 16960 7946 16988 8222
rect 16948 7940 17000 7946
rect 16948 7882 17000 7888
rect 18052 7872 18104 7878
rect 18052 7814 18104 7820
rect 17960 7736 18012 7742
rect 17960 7678 18012 7684
rect 17972 7402 18000 7678
rect 17960 7396 18012 7402
rect 17960 7338 18012 7344
rect 18064 6722 18092 7814
rect 18144 7804 18196 7810
rect 18144 7746 18196 7752
rect 18156 7402 18184 7746
rect 18604 7600 18656 7606
rect 18604 7542 18656 7548
rect 18282 7500 18578 7520
rect 18338 7498 18362 7500
rect 18418 7498 18442 7500
rect 18498 7498 18522 7500
rect 18360 7446 18362 7498
rect 18424 7446 18436 7498
rect 18498 7446 18500 7498
rect 18338 7444 18362 7446
rect 18418 7444 18442 7446
rect 18498 7444 18522 7446
rect 18282 7424 18578 7444
rect 18616 7402 18644 7542
rect 18144 7396 18196 7402
rect 18144 7338 18196 7344
rect 18604 7396 18656 7402
rect 18604 7338 18656 7344
rect 18052 6716 18104 6722
rect 18052 6658 18104 6664
rect 17960 6512 18012 6518
rect 17960 6454 18012 6460
rect 17972 5537 18000 6454
rect 18282 6412 18578 6432
rect 18338 6410 18362 6412
rect 18418 6410 18442 6412
rect 18498 6410 18522 6412
rect 18360 6358 18362 6410
rect 18424 6358 18436 6410
rect 18498 6358 18500 6410
rect 18338 6356 18362 6358
rect 18418 6356 18442 6358
rect 18498 6356 18522 6358
rect 18282 6336 18578 6356
rect 17958 5528 18014 5537
rect 17958 5463 18014 5472
rect 18282 5324 18578 5344
rect 18338 5322 18362 5324
rect 18418 5322 18442 5324
rect 18498 5322 18522 5324
rect 18360 5270 18362 5322
rect 18424 5270 18436 5322
rect 18498 5270 18500 5322
rect 18338 5268 18362 5270
rect 18418 5268 18442 5270
rect 18498 5268 18522 5270
rect 18282 5248 18578 5268
rect 17960 5220 18012 5226
rect 17960 5162 18012 5168
rect 17972 4585 18000 5162
rect 17958 4576 18014 4585
rect 17958 4511 18014 4520
rect 18282 4236 18578 4256
rect 18338 4234 18362 4236
rect 18418 4234 18442 4236
rect 18498 4234 18522 4236
rect 18360 4182 18362 4234
rect 18424 4182 18436 4234
rect 18498 4182 18500 4234
rect 18338 4180 18362 4182
rect 18418 4180 18442 4182
rect 18498 4180 18522 4182
rect 18282 4160 18578 4180
rect 16488 3996 16540 4002
rect 16488 3938 16540 3944
rect 14817 3692 15113 3712
rect 14873 3690 14897 3692
rect 14953 3690 14977 3692
rect 15033 3690 15057 3692
rect 14895 3638 14897 3690
rect 14959 3638 14971 3690
rect 15033 3638 15035 3690
rect 14873 3636 14897 3638
rect 14953 3636 14977 3638
rect 15033 3636 15057 3638
rect 14817 3616 15113 3636
rect 18282 3148 18578 3168
rect 18338 3146 18362 3148
rect 18418 3146 18442 3148
rect 18498 3146 18522 3148
rect 18360 3094 18362 3146
rect 18424 3094 18436 3146
rect 18498 3094 18500 3146
rect 18338 3092 18362 3094
rect 18418 3092 18442 3094
rect 18498 3092 18522 3094
rect 18282 3072 18578 3092
rect 18708 2982 18736 10874
rect 18800 10122 18828 11554
rect 18788 10116 18840 10122
rect 18788 10058 18840 10064
rect 18788 3996 18840 4002
rect 18788 3938 18840 3944
rect 18800 3225 18828 3938
rect 18786 3216 18842 3225
rect 18786 3151 18842 3160
rect 18892 3066 18920 12234
rect 18984 10938 19012 12438
rect 19076 11958 19104 12778
rect 19248 12768 19300 12774
rect 19248 12710 19300 12716
rect 19260 12162 19288 12710
rect 19248 12156 19300 12162
rect 19248 12098 19300 12104
rect 19064 11952 19116 11958
rect 19064 11894 19116 11900
rect 19076 11226 19104 11894
rect 19628 11754 19656 17946
rect 19800 17936 19852 17942
rect 19800 17878 19852 17884
rect 19708 17188 19760 17194
rect 19708 17130 19760 17136
rect 19720 16514 19748 17130
rect 19708 16508 19760 16514
rect 19708 16450 19760 16456
rect 19708 12632 19760 12638
rect 19708 12574 19760 12580
rect 19720 12473 19748 12574
rect 19706 12464 19762 12473
rect 19706 12399 19762 12408
rect 19812 12298 19840 17878
rect 19904 16938 19932 22056
rect 20166 22055 20222 22064
rect 20442 22056 20498 22856
rect 20994 22056 21050 22856
rect 21546 22056 21602 22856
rect 22098 22056 22154 22856
rect 22650 22056 22706 22856
rect 20180 20458 20208 22055
rect 20168 20452 20220 20458
rect 20168 20394 20220 20400
rect 20456 20338 20484 22056
rect 20534 21168 20590 21177
rect 20534 21103 20590 21112
rect 20548 20458 20576 21103
rect 20626 20760 20682 20769
rect 20626 20695 20682 20704
rect 20536 20452 20588 20458
rect 20536 20394 20588 20400
rect 20364 20310 20484 20338
rect 19984 20248 20036 20254
rect 19984 20190 20036 20196
rect 20076 20248 20128 20254
rect 20076 20190 20128 20196
rect 19996 18758 20024 20190
rect 20088 19846 20116 20190
rect 20076 19840 20128 19846
rect 20076 19782 20128 19788
rect 20168 19772 20220 19778
rect 20168 19714 20220 19720
rect 20180 18758 20208 19714
rect 19984 18752 20036 18758
rect 19984 18694 20036 18700
rect 20168 18752 20220 18758
rect 20168 18694 20220 18700
rect 20168 18140 20220 18146
rect 20168 18082 20220 18088
rect 20076 18072 20128 18078
rect 20076 18014 20128 18020
rect 20088 17058 20116 18014
rect 20076 17052 20128 17058
rect 20076 16994 20128 17000
rect 19904 16910 20116 16938
rect 19984 16848 20036 16854
rect 19984 16790 20036 16796
rect 19800 12292 19852 12298
rect 19800 12234 19852 12240
rect 19616 11748 19668 11754
rect 19616 11690 19668 11696
rect 19432 11544 19484 11550
rect 19432 11486 19484 11492
rect 19248 11476 19300 11482
rect 19248 11418 19300 11424
rect 19260 11226 19288 11418
rect 19340 11408 19392 11414
rect 19340 11350 19392 11356
rect 19076 11198 19288 11226
rect 19064 11136 19116 11142
rect 19064 11078 19116 11084
rect 18972 10932 19024 10938
rect 18972 10874 19024 10880
rect 18972 10320 19024 10326
rect 18972 10262 19024 10268
rect 18984 10054 19012 10262
rect 18972 10048 19024 10054
rect 18972 9990 19024 9996
rect 18984 7266 19012 9990
rect 18972 7260 19024 7266
rect 18972 7202 19024 7208
rect 18984 6858 19012 7202
rect 18972 6852 19024 6858
rect 18972 6794 19024 6800
rect 19076 3610 19104 11078
rect 19156 11068 19208 11074
rect 19156 11010 19208 11016
rect 19168 10666 19196 11010
rect 19156 10660 19208 10666
rect 19156 10602 19208 10608
rect 19260 10546 19288 11198
rect 19168 10518 19288 10546
rect 19168 3769 19196 10518
rect 19352 10444 19380 11350
rect 19444 11142 19472 11486
rect 19996 11210 20024 16790
rect 20088 11754 20116 16910
rect 20180 12842 20208 18082
rect 20364 17942 20392 20310
rect 20442 20216 20498 20225
rect 20442 20151 20498 20160
rect 20456 19370 20484 20151
rect 20640 19914 20668 20695
rect 21008 19930 21036 22056
rect 20628 19908 20680 19914
rect 21008 19902 21312 19930
rect 20628 19850 20680 19856
rect 21086 19808 21142 19817
rect 21086 19743 21142 19752
rect 21100 19370 21128 19743
rect 20444 19364 20496 19370
rect 20444 19306 20496 19312
rect 21088 19364 21140 19370
rect 21088 19306 21140 19312
rect 20994 19264 21050 19273
rect 20994 19199 21050 19208
rect 20626 18856 20682 18865
rect 21008 18826 21036 19199
rect 20626 18791 20682 18800
rect 20996 18820 21048 18826
rect 20536 18004 20588 18010
rect 20536 17946 20588 17952
rect 20352 17936 20404 17942
rect 20352 17878 20404 17884
rect 20442 17496 20498 17505
rect 20442 17431 20444 17440
rect 20496 17431 20498 17440
rect 20444 17402 20496 17408
rect 20444 17120 20496 17126
rect 20444 17062 20496 17068
rect 20456 16514 20484 17062
rect 20444 16508 20496 16514
rect 20444 16450 20496 16456
rect 20548 16394 20576 17946
rect 20456 16366 20576 16394
rect 20260 14128 20312 14134
rect 20260 14070 20312 14076
rect 20272 13726 20300 14070
rect 20456 13930 20484 16366
rect 20534 14232 20590 14241
rect 20534 14167 20590 14176
rect 20444 13924 20496 13930
rect 20444 13866 20496 13872
rect 20442 13824 20498 13833
rect 20442 13759 20498 13768
rect 20260 13720 20312 13726
rect 20260 13662 20312 13668
rect 20272 12881 20300 13662
rect 20258 12872 20314 12881
rect 20168 12836 20220 12842
rect 20456 12842 20484 13759
rect 20548 13386 20576 14167
rect 20640 13930 20668 18791
rect 20996 18762 21048 18768
rect 20812 18684 20864 18690
rect 20812 18626 20864 18632
rect 20720 17596 20772 17602
rect 20720 17538 20772 17544
rect 20732 16514 20760 17538
rect 20720 16508 20772 16514
rect 20720 16450 20772 16456
rect 20824 15562 20852 18626
rect 21088 17936 21140 17942
rect 21086 17904 21088 17913
rect 21180 17936 21232 17942
rect 21140 17904 21142 17913
rect 21180 17878 21232 17884
rect 21086 17839 21142 17848
rect 20996 17392 21048 17398
rect 20996 17334 21048 17340
rect 21008 17097 21036 17334
rect 20994 17088 21050 17097
rect 20994 17023 21050 17032
rect 21088 16848 21140 16854
rect 21088 16790 21140 16796
rect 20904 16576 20956 16582
rect 21100 16553 21128 16790
rect 20904 16518 20956 16524
rect 21086 16544 21142 16553
rect 20916 15902 20944 16518
rect 21086 16479 21142 16488
rect 21086 16136 21142 16145
rect 21086 16071 21088 16080
rect 21140 16071 21142 16080
rect 21088 16042 21140 16048
rect 20904 15896 20956 15902
rect 20904 15838 20956 15844
rect 21192 15714 21220 17878
rect 21100 15686 21220 15714
rect 20812 15556 20864 15562
rect 20812 15498 20864 15504
rect 20812 15420 20864 15426
rect 20812 15362 20864 15368
rect 20824 14882 20852 15362
rect 20996 15216 21048 15222
rect 20994 15184 20996 15193
rect 21048 15184 21050 15193
rect 20994 15119 21050 15128
rect 21100 15034 21128 15686
rect 21178 15592 21234 15601
rect 21178 15527 21234 15536
rect 21008 15006 21128 15034
rect 20812 14876 20864 14882
rect 20812 14818 20864 14824
rect 20812 14740 20864 14746
rect 20812 14682 20864 14688
rect 20824 14338 20852 14682
rect 20812 14332 20864 14338
rect 20812 14274 20864 14280
rect 20904 14264 20956 14270
rect 20904 14206 20956 14212
rect 20628 13924 20680 13930
rect 20628 13866 20680 13872
rect 20916 13726 20944 14206
rect 20904 13720 20956 13726
rect 20904 13662 20956 13668
rect 20536 13380 20588 13386
rect 20536 13322 20588 13328
rect 20628 13176 20680 13182
rect 20628 13118 20680 13124
rect 20258 12807 20314 12816
rect 20444 12836 20496 12842
rect 20168 12778 20220 12784
rect 20444 12778 20496 12784
rect 20352 12632 20404 12638
rect 20352 12574 20404 12580
rect 20364 12230 20392 12574
rect 20352 12224 20404 12230
rect 20352 12166 20404 12172
rect 20640 11929 20668 13118
rect 20626 11920 20682 11929
rect 20626 11855 20682 11864
rect 20076 11748 20128 11754
rect 20076 11690 20128 11696
rect 20904 11544 20956 11550
rect 20904 11486 20956 11492
rect 19984 11204 20036 11210
rect 19984 11146 20036 11152
rect 19432 11136 19484 11142
rect 20916 11113 20944 11486
rect 19432 11078 19484 11084
rect 20902 11104 20958 11113
rect 20628 11068 20680 11074
rect 20902 11039 20958 11048
rect 20628 11010 20680 11016
rect 20536 10932 20588 10938
rect 20536 10874 20588 10880
rect 19892 10524 19944 10530
rect 19892 10466 19944 10472
rect 19260 10416 19380 10444
rect 19260 7146 19288 10416
rect 19708 10320 19760 10326
rect 19708 10262 19760 10268
rect 19720 10122 19748 10262
rect 19708 10116 19760 10122
rect 19708 10058 19760 10064
rect 19904 9986 19932 10466
rect 20548 10444 20576 10874
rect 20640 10569 20668 11010
rect 20626 10560 20682 10569
rect 20626 10495 20682 10504
rect 20628 10456 20680 10462
rect 20548 10416 20628 10444
rect 20628 10398 20680 10404
rect 20074 10152 20130 10161
rect 20074 10087 20076 10096
rect 20128 10087 20130 10096
rect 20076 10058 20128 10064
rect 19892 9980 19944 9986
rect 19892 9922 19944 9928
rect 19904 9578 19932 9922
rect 19892 9572 19944 9578
rect 19892 9514 19944 9520
rect 19708 9368 19760 9374
rect 19708 9310 19760 9316
rect 19720 7946 19748 9310
rect 20088 9034 20116 10058
rect 20536 9980 20588 9986
rect 20536 9922 20588 9928
rect 20260 9912 20312 9918
rect 20260 9854 20312 9860
rect 20272 9374 20300 9854
rect 20260 9368 20312 9374
rect 20260 9310 20312 9316
rect 20548 9209 20576 9922
rect 20640 9617 20668 10398
rect 20626 9608 20682 9617
rect 20626 9543 20682 9552
rect 20904 9368 20956 9374
rect 20904 9310 20956 9316
rect 20534 9200 20590 9209
rect 20534 9135 20590 9144
rect 20548 9034 20576 9135
rect 20076 9028 20128 9034
rect 20076 8970 20128 8976
rect 20536 9028 20588 9034
rect 20536 8970 20588 8976
rect 20916 8801 20944 9310
rect 20902 8792 20958 8801
rect 20902 8727 20958 8736
rect 20628 8280 20680 8286
rect 20628 8222 20680 8228
rect 19708 7940 19760 7946
rect 19708 7882 19760 7888
rect 20640 7849 20668 8222
rect 20626 7840 20682 7849
rect 20626 7775 20682 7784
rect 20812 7804 20864 7810
rect 20812 7746 20864 7752
rect 20824 7441 20852 7746
rect 20810 7432 20866 7441
rect 20810 7367 20866 7376
rect 20904 7192 20956 7198
rect 19260 7118 19380 7146
rect 20904 7134 20956 7140
rect 19248 7056 19300 7062
rect 19248 6998 19300 7004
rect 19260 6489 19288 6998
rect 19246 6480 19302 6489
rect 19246 6415 19302 6424
rect 19352 6330 19380 7118
rect 20916 6897 20944 7134
rect 20902 6888 20958 6897
rect 20902 6823 20958 6832
rect 19260 6302 19380 6330
rect 19154 3760 19210 3769
rect 19154 3695 19210 3704
rect 19076 3582 19196 3610
rect 18800 3038 18920 3066
rect 18696 2976 18748 2982
rect 18696 2918 18748 2924
rect 14817 2604 15113 2624
rect 14873 2602 14897 2604
rect 14953 2602 14977 2604
rect 15033 2602 15057 2604
rect 14895 2550 14897 2602
rect 14959 2550 14971 2602
rect 15033 2550 15035 2602
rect 14873 2548 14897 2550
rect 14953 2548 14977 2550
rect 15033 2548 15057 2550
rect 14817 2528 15113 2548
rect 18144 2432 18196 2438
rect 18144 2374 18196 2380
rect 18156 2273 18184 2374
rect 18142 2264 18198 2273
rect 18142 2199 18198 2208
rect 18282 2060 18578 2080
rect 18338 2058 18362 2060
rect 18418 2058 18442 2060
rect 18498 2058 18522 2060
rect 18360 2006 18362 2058
rect 18424 2006 18436 2058
rect 18498 2006 18500 2058
rect 18338 2004 18362 2006
rect 18418 2004 18442 2006
rect 18498 2004 18522 2006
rect 18282 1984 18578 2004
rect 18144 1956 18196 1962
rect 18144 1898 18196 1904
rect 18156 1457 18184 1898
rect 18142 1448 18198 1457
rect 18142 1383 18198 1392
rect 14556 1208 14608 1214
rect 14556 1150 14608 1156
rect 17960 1208 18012 1214
rect 17960 1150 18012 1156
rect 17972 505 18000 1150
rect 17958 496 18014 505
rect 17958 431 18014 440
rect 18800 97 18828 3038
rect 18880 2976 18932 2982
rect 18880 2918 18932 2924
rect 18892 1865 18920 2918
rect 18878 1856 18934 1865
rect 18878 1791 18934 1800
rect 19168 913 19196 3582
rect 19260 2817 19288 6302
rect 21008 4682 21036 15006
rect 21086 14776 21142 14785
rect 21086 14711 21142 14720
rect 21100 14678 21128 14711
rect 21088 14672 21140 14678
rect 21088 14614 21140 14620
rect 21192 14474 21220 15527
rect 21180 14468 21232 14474
rect 21180 14410 21232 14416
rect 21086 13416 21142 13425
rect 21284 13386 21312 19902
rect 21456 18208 21508 18214
rect 21456 18150 21508 18156
rect 21086 13351 21142 13360
rect 21272 13380 21324 13386
rect 21100 12842 21128 13351
rect 21272 13322 21324 13328
rect 21088 12836 21140 12842
rect 21088 12778 21140 12784
rect 21468 10666 21496 18150
rect 21560 18146 21588 22056
rect 21732 18752 21784 18758
rect 21732 18694 21784 18700
rect 21640 18276 21692 18282
rect 21640 18218 21692 18224
rect 21548 18140 21600 18146
rect 21548 18082 21600 18088
rect 21456 10660 21508 10666
rect 21456 10602 21508 10608
rect 21652 10122 21680 18218
rect 21640 10116 21692 10122
rect 21640 10058 21692 10064
rect 21744 9510 21772 18694
rect 22112 18010 22140 22056
rect 22100 18004 22152 18010
rect 22100 17946 22152 17952
rect 22664 17942 22692 22056
rect 22652 17936 22704 17942
rect 22652 17878 22704 17884
rect 22008 11544 22060 11550
rect 22006 11512 22008 11521
rect 22060 11512 22062 11521
rect 22006 11447 22062 11456
rect 21732 9504 21784 9510
rect 21732 9446 21784 9452
rect 22008 8280 22060 8286
rect 22006 8248 22008 8257
rect 22060 8248 22062 8257
rect 22006 8183 22062 8192
rect 21088 8144 21140 8150
rect 21088 8086 21140 8092
rect 21100 7402 21128 8086
rect 21088 7396 21140 7402
rect 21088 7338 21140 7344
rect 21364 6512 21416 6518
rect 21364 6454 21416 6460
rect 21376 6110 21404 6454
rect 21364 6104 21416 6110
rect 21364 6046 21416 6052
rect 21376 5945 21404 6046
rect 21362 5936 21418 5945
rect 21362 5871 21418 5880
rect 21272 5628 21324 5634
rect 21272 5570 21324 5576
rect 21284 5158 21312 5570
rect 21272 5152 21324 5158
rect 21270 5120 21272 5129
rect 21324 5120 21326 5129
rect 21270 5055 21326 5064
rect 20996 4676 21048 4682
rect 20996 4618 21048 4624
rect 21272 4540 21324 4546
rect 21272 4482 21324 4488
rect 21284 4177 21312 4482
rect 21270 4168 21326 4177
rect 21270 4103 21272 4112
rect 21324 4103 21326 4112
rect 21272 4074 21324 4080
rect 19246 2808 19302 2817
rect 19246 2743 19302 2752
rect 19154 904 19210 913
rect 19154 839 19210 848
rect 18786 88 18842 97
rect 18786 23 18842 32
<< via2 >>
rect 19246 22472 19302 22528
rect 4421 20554 4477 20556
rect 4501 20554 4557 20556
rect 4581 20554 4637 20556
rect 4661 20554 4717 20556
rect 4421 20502 4447 20554
rect 4447 20502 4477 20554
rect 4501 20502 4511 20554
rect 4511 20502 4557 20554
rect 4581 20502 4627 20554
rect 4627 20502 4637 20554
rect 4661 20502 4691 20554
rect 4691 20502 4717 20554
rect 4421 20500 4477 20502
rect 4501 20500 4557 20502
rect 4581 20500 4637 20502
rect 4661 20500 4717 20502
rect 4421 19466 4477 19468
rect 4501 19466 4557 19468
rect 4581 19466 4637 19468
rect 4661 19466 4717 19468
rect 4421 19414 4447 19466
rect 4447 19414 4477 19466
rect 4501 19414 4511 19466
rect 4511 19414 4557 19466
rect 4581 19414 4627 19466
rect 4627 19414 4637 19466
rect 4661 19414 4691 19466
rect 4691 19414 4717 19466
rect 4421 19412 4477 19414
rect 4501 19412 4557 19414
rect 4581 19412 4637 19414
rect 4661 19412 4717 19414
rect 4421 18378 4477 18380
rect 4501 18378 4557 18380
rect 4581 18378 4637 18380
rect 4661 18378 4717 18380
rect 4421 18326 4447 18378
rect 4447 18326 4477 18378
rect 4501 18326 4511 18378
rect 4511 18326 4557 18378
rect 4581 18326 4627 18378
rect 4627 18326 4637 18378
rect 4661 18326 4691 18378
rect 4691 18326 4717 18378
rect 4421 18324 4477 18326
rect 4501 18324 4557 18326
rect 4581 18324 4637 18326
rect 4661 18324 4717 18326
rect 4421 17290 4477 17292
rect 4501 17290 4557 17292
rect 4581 17290 4637 17292
rect 4661 17290 4717 17292
rect 4421 17238 4447 17290
rect 4447 17238 4477 17290
rect 4501 17238 4511 17290
rect 4511 17238 4557 17290
rect 4581 17238 4627 17290
rect 4627 17238 4637 17290
rect 4661 17238 4691 17290
rect 4691 17238 4717 17290
rect 4421 17236 4477 17238
rect 4501 17236 4557 17238
rect 4581 17236 4637 17238
rect 4661 17236 4717 17238
rect 4802 17032 4858 17088
rect 6366 18120 6422 18176
rect 4421 16202 4477 16204
rect 4501 16202 4557 16204
rect 4581 16202 4637 16204
rect 4661 16202 4717 16204
rect 4421 16150 4447 16202
rect 4447 16150 4477 16202
rect 4501 16150 4511 16202
rect 4511 16150 4557 16202
rect 4581 16150 4627 16202
rect 4627 16150 4637 16202
rect 4661 16150 4691 16202
rect 4691 16150 4717 16202
rect 4421 16148 4477 16150
rect 4501 16148 4557 16150
rect 4581 16148 4637 16150
rect 4661 16148 4717 16150
rect 4421 15114 4477 15116
rect 4501 15114 4557 15116
rect 4581 15114 4637 15116
rect 4661 15114 4717 15116
rect 4421 15062 4447 15114
rect 4447 15062 4477 15114
rect 4501 15062 4511 15114
rect 4511 15062 4557 15114
rect 4581 15062 4627 15114
rect 4627 15062 4637 15114
rect 4661 15062 4691 15114
rect 4691 15062 4717 15114
rect 4421 15060 4477 15062
rect 4501 15060 4557 15062
rect 4581 15060 4637 15062
rect 4661 15060 4717 15062
rect 4421 14026 4477 14028
rect 4501 14026 4557 14028
rect 4581 14026 4637 14028
rect 4661 14026 4717 14028
rect 4421 13974 4447 14026
rect 4447 13974 4477 14026
rect 4501 13974 4511 14026
rect 4511 13974 4557 14026
rect 4581 13974 4627 14026
rect 4627 13974 4637 14026
rect 4661 13974 4691 14026
rect 4691 13974 4717 14026
rect 4421 13972 4477 13974
rect 4501 13972 4557 13974
rect 4581 13972 4637 13974
rect 4661 13972 4717 13974
rect 4421 12938 4477 12940
rect 4501 12938 4557 12940
rect 4581 12938 4637 12940
rect 4661 12938 4717 12940
rect 4421 12886 4447 12938
rect 4447 12886 4477 12938
rect 4501 12886 4511 12938
rect 4511 12886 4557 12938
rect 4581 12886 4627 12938
rect 4627 12886 4637 12938
rect 4661 12886 4691 12938
rect 4691 12886 4717 12938
rect 4421 12884 4477 12886
rect 4501 12884 4557 12886
rect 4581 12884 4637 12886
rect 4661 12884 4717 12886
rect 4421 11850 4477 11852
rect 4501 11850 4557 11852
rect 4581 11850 4637 11852
rect 4661 11850 4717 11852
rect 4421 11798 4447 11850
rect 4447 11798 4477 11850
rect 4501 11798 4511 11850
rect 4511 11798 4557 11850
rect 4581 11798 4627 11850
rect 4627 11798 4637 11850
rect 4661 11798 4691 11850
rect 4691 11798 4717 11850
rect 4421 11796 4477 11798
rect 4501 11796 4557 11798
rect 4581 11796 4637 11798
rect 4661 11796 4717 11798
rect 7886 20010 7942 20012
rect 7966 20010 8022 20012
rect 8046 20010 8102 20012
rect 8126 20010 8182 20012
rect 7886 19958 7912 20010
rect 7912 19958 7942 20010
rect 7966 19958 7976 20010
rect 7976 19958 8022 20010
rect 8046 19958 8092 20010
rect 8092 19958 8102 20010
rect 8126 19958 8156 20010
rect 8156 19958 8182 20010
rect 7886 19956 7942 19958
rect 7966 19956 8022 19958
rect 8046 19956 8102 19958
rect 8126 19956 8182 19958
rect 7886 18922 7942 18924
rect 7966 18922 8022 18924
rect 8046 18922 8102 18924
rect 8126 18922 8182 18924
rect 7886 18870 7912 18922
rect 7912 18870 7942 18922
rect 7966 18870 7976 18922
rect 7976 18870 8022 18922
rect 8046 18870 8092 18922
rect 8092 18870 8102 18922
rect 8126 18870 8156 18922
rect 8156 18870 8182 18922
rect 7886 18868 7942 18870
rect 7966 18868 8022 18870
rect 8046 18868 8102 18870
rect 8126 18868 8182 18870
rect 7886 17834 7942 17836
rect 7966 17834 8022 17836
rect 8046 17834 8102 17836
rect 8126 17834 8182 17836
rect 7886 17782 7912 17834
rect 7912 17782 7942 17834
rect 7966 17782 7976 17834
rect 7976 17782 8022 17834
rect 8046 17782 8092 17834
rect 8092 17782 8102 17834
rect 8126 17782 8156 17834
rect 8156 17782 8182 17834
rect 7886 17780 7942 17782
rect 7966 17780 8022 17782
rect 8046 17780 8102 17782
rect 8126 17780 8182 17782
rect 10322 18936 10378 18992
rect 11352 20554 11408 20556
rect 11432 20554 11488 20556
rect 11512 20554 11568 20556
rect 11592 20554 11648 20556
rect 11352 20502 11378 20554
rect 11378 20502 11408 20554
rect 11432 20502 11442 20554
rect 11442 20502 11488 20554
rect 11512 20502 11558 20554
rect 11558 20502 11568 20554
rect 11592 20502 11622 20554
rect 11622 20502 11648 20554
rect 11352 20500 11408 20502
rect 11432 20500 11488 20502
rect 11512 20500 11568 20502
rect 11592 20500 11648 20502
rect 11352 19466 11408 19468
rect 11432 19466 11488 19468
rect 11512 19466 11568 19468
rect 11592 19466 11648 19468
rect 11352 19414 11378 19466
rect 11378 19414 11408 19466
rect 11432 19414 11442 19466
rect 11442 19414 11488 19466
rect 11512 19414 11558 19466
rect 11558 19414 11568 19466
rect 11592 19414 11622 19466
rect 11622 19414 11648 19466
rect 11352 19412 11408 19414
rect 11432 19412 11488 19414
rect 11512 19412 11568 19414
rect 11592 19412 11648 19414
rect 11150 19092 11206 19128
rect 11150 19072 11152 19092
rect 11152 19072 11204 19092
rect 11204 19072 11206 19092
rect 11426 18664 11482 18720
rect 11242 18528 11298 18584
rect 7886 16746 7942 16748
rect 7966 16746 8022 16748
rect 8046 16746 8102 16748
rect 8126 16746 8182 16748
rect 7886 16694 7912 16746
rect 7912 16694 7942 16746
rect 7966 16694 7976 16746
rect 7976 16694 8022 16746
rect 8046 16694 8092 16746
rect 8092 16694 8102 16746
rect 8126 16694 8156 16746
rect 8156 16694 8182 16746
rect 7886 16692 7942 16694
rect 7966 16692 8022 16694
rect 8046 16692 8102 16694
rect 8126 16692 8182 16694
rect 11352 18378 11408 18380
rect 11432 18378 11488 18380
rect 11512 18378 11568 18380
rect 11592 18378 11648 18380
rect 11352 18326 11378 18378
rect 11378 18326 11408 18378
rect 11432 18326 11442 18378
rect 11442 18326 11488 18378
rect 11512 18326 11558 18378
rect 11558 18326 11568 18378
rect 11592 18326 11622 18378
rect 11622 18326 11648 18378
rect 11352 18324 11408 18326
rect 11432 18324 11488 18326
rect 11512 18324 11568 18326
rect 11592 18324 11648 18326
rect 11610 18120 11666 18176
rect 7886 15658 7942 15660
rect 7966 15658 8022 15660
rect 8046 15658 8102 15660
rect 8126 15658 8182 15660
rect 7886 15606 7912 15658
rect 7912 15606 7942 15658
rect 7966 15606 7976 15658
rect 7976 15606 8022 15658
rect 8046 15606 8092 15658
rect 8092 15606 8102 15658
rect 8126 15606 8156 15658
rect 8156 15606 8182 15658
rect 7886 15604 7942 15606
rect 7966 15604 8022 15606
rect 8046 15604 8102 15606
rect 8126 15604 8182 15606
rect 7886 14570 7942 14572
rect 7966 14570 8022 14572
rect 8046 14570 8102 14572
rect 8126 14570 8182 14572
rect 7886 14518 7912 14570
rect 7912 14518 7942 14570
rect 7966 14518 7976 14570
rect 7976 14518 8022 14570
rect 8046 14518 8092 14570
rect 8092 14518 8102 14570
rect 8126 14518 8156 14570
rect 8156 14518 8182 14570
rect 7886 14516 7942 14518
rect 7966 14516 8022 14518
rect 8046 14516 8102 14518
rect 8126 14516 8182 14518
rect 7886 13482 7942 13484
rect 7966 13482 8022 13484
rect 8046 13482 8102 13484
rect 8126 13482 8182 13484
rect 7886 13430 7912 13482
rect 7912 13430 7942 13482
rect 7966 13430 7976 13482
rect 7976 13430 8022 13482
rect 8046 13430 8092 13482
rect 8092 13430 8102 13482
rect 8126 13430 8156 13482
rect 8156 13430 8182 13482
rect 7886 13428 7942 13430
rect 7966 13428 8022 13430
rect 8046 13428 8102 13430
rect 8126 13428 8182 13430
rect 7886 12394 7942 12396
rect 7966 12394 8022 12396
rect 8046 12394 8102 12396
rect 8126 12394 8182 12396
rect 7886 12342 7912 12394
rect 7912 12342 7942 12394
rect 7966 12342 7976 12394
rect 7976 12342 8022 12394
rect 8046 12342 8092 12394
rect 8092 12342 8102 12394
rect 8126 12342 8156 12394
rect 8156 12342 8182 12394
rect 7886 12340 7942 12342
rect 7966 12340 8022 12342
rect 8046 12340 8102 12342
rect 8126 12340 8182 12342
rect 7886 11306 7942 11308
rect 7966 11306 8022 11308
rect 8046 11306 8102 11308
rect 8126 11306 8182 11308
rect 7886 11254 7912 11306
rect 7912 11254 7942 11306
rect 7966 11254 7976 11306
rect 7976 11254 8022 11306
rect 8046 11254 8092 11306
rect 8092 11254 8102 11306
rect 8126 11254 8156 11306
rect 8156 11254 8182 11306
rect 7886 11252 7942 11254
rect 7966 11252 8022 11254
rect 8046 11252 8102 11254
rect 8126 11252 8182 11254
rect 4421 10762 4477 10764
rect 4501 10762 4557 10764
rect 4581 10762 4637 10764
rect 4661 10762 4717 10764
rect 4421 10710 4447 10762
rect 4447 10710 4477 10762
rect 4501 10710 4511 10762
rect 4511 10710 4557 10762
rect 4581 10710 4627 10762
rect 4627 10710 4637 10762
rect 4661 10710 4691 10762
rect 4691 10710 4717 10762
rect 4421 10708 4477 10710
rect 4501 10708 4557 10710
rect 4581 10708 4637 10710
rect 4661 10708 4717 10710
rect 7886 10218 7942 10220
rect 7966 10218 8022 10220
rect 8046 10218 8102 10220
rect 8126 10218 8182 10220
rect 7886 10166 7912 10218
rect 7912 10166 7942 10218
rect 7966 10166 7976 10218
rect 7976 10166 8022 10218
rect 8046 10166 8092 10218
rect 8092 10166 8102 10218
rect 8126 10166 8156 10218
rect 8156 10166 8182 10218
rect 7886 10164 7942 10166
rect 7966 10164 8022 10166
rect 8046 10164 8102 10166
rect 8126 10164 8182 10166
rect 11352 17290 11408 17292
rect 11432 17290 11488 17292
rect 11512 17290 11568 17292
rect 11592 17290 11648 17292
rect 11352 17238 11378 17290
rect 11378 17238 11408 17290
rect 11432 17238 11442 17290
rect 11442 17238 11488 17290
rect 11512 17238 11558 17290
rect 11558 17238 11568 17290
rect 11592 17238 11622 17290
rect 11622 17238 11648 17290
rect 11352 17236 11408 17238
rect 11432 17236 11488 17238
rect 11512 17236 11568 17238
rect 11592 17236 11648 17238
rect 11352 16202 11408 16204
rect 11432 16202 11488 16204
rect 11512 16202 11568 16204
rect 11592 16202 11648 16204
rect 11352 16150 11378 16202
rect 11378 16150 11408 16202
rect 11432 16150 11442 16202
rect 11442 16150 11488 16202
rect 11512 16150 11558 16202
rect 11558 16150 11568 16202
rect 11592 16150 11622 16202
rect 11622 16150 11648 16202
rect 11352 16148 11408 16150
rect 11432 16148 11488 16150
rect 11512 16148 11568 16150
rect 11592 16148 11648 16150
rect 11352 15114 11408 15116
rect 11432 15114 11488 15116
rect 11512 15114 11568 15116
rect 11592 15114 11648 15116
rect 11352 15062 11378 15114
rect 11378 15062 11408 15114
rect 11432 15062 11442 15114
rect 11442 15062 11488 15114
rect 11512 15062 11558 15114
rect 11558 15062 11568 15114
rect 11592 15062 11622 15114
rect 11622 15062 11648 15114
rect 11352 15060 11408 15062
rect 11432 15060 11488 15062
rect 11512 15060 11568 15062
rect 11592 15060 11648 15062
rect 11352 14026 11408 14028
rect 11432 14026 11488 14028
rect 11512 14026 11568 14028
rect 11592 14026 11648 14028
rect 11352 13974 11378 14026
rect 11378 13974 11408 14026
rect 11432 13974 11442 14026
rect 11442 13974 11488 14026
rect 11512 13974 11558 14026
rect 11558 13974 11568 14026
rect 11592 13974 11622 14026
rect 11622 13974 11648 14026
rect 11352 13972 11408 13974
rect 11432 13972 11488 13974
rect 11512 13972 11568 13974
rect 11592 13972 11648 13974
rect 11352 12938 11408 12940
rect 11432 12938 11488 12940
rect 11512 12938 11568 12940
rect 11592 12938 11648 12940
rect 11352 12886 11378 12938
rect 11378 12886 11408 12938
rect 11432 12886 11442 12938
rect 11442 12886 11488 12938
rect 11512 12886 11558 12938
rect 11558 12886 11568 12938
rect 11592 12886 11622 12938
rect 11622 12886 11648 12938
rect 11352 12884 11408 12886
rect 11432 12884 11488 12886
rect 11512 12884 11568 12886
rect 11592 12884 11648 12886
rect 11352 11850 11408 11852
rect 11432 11850 11488 11852
rect 11512 11850 11568 11852
rect 11592 11850 11648 11852
rect 11352 11798 11378 11850
rect 11378 11798 11408 11850
rect 11432 11798 11442 11850
rect 11442 11798 11488 11850
rect 11512 11798 11558 11850
rect 11558 11798 11568 11850
rect 11592 11798 11622 11850
rect 11622 11798 11648 11850
rect 11352 11796 11408 11798
rect 11432 11796 11488 11798
rect 11512 11796 11568 11798
rect 11592 11796 11648 11798
rect 4421 9674 4477 9676
rect 4501 9674 4557 9676
rect 4581 9674 4637 9676
rect 4661 9674 4717 9676
rect 4421 9622 4447 9674
rect 4447 9622 4477 9674
rect 4501 9622 4511 9674
rect 4511 9622 4557 9674
rect 4581 9622 4627 9674
rect 4627 9622 4637 9674
rect 4661 9622 4691 9674
rect 4691 9622 4717 9674
rect 4421 9620 4477 9622
rect 4501 9620 4557 9622
rect 4581 9620 4637 9622
rect 4661 9620 4717 9622
rect 11352 10762 11408 10764
rect 11432 10762 11488 10764
rect 11512 10762 11568 10764
rect 11592 10762 11648 10764
rect 11352 10710 11378 10762
rect 11378 10710 11408 10762
rect 11432 10710 11442 10762
rect 11442 10710 11488 10762
rect 11512 10710 11558 10762
rect 11558 10710 11568 10762
rect 11592 10710 11622 10762
rect 11622 10710 11648 10762
rect 11352 10708 11408 10710
rect 11432 10708 11488 10710
rect 11512 10708 11568 10710
rect 11592 10708 11648 10710
rect 11352 9674 11408 9676
rect 11432 9674 11488 9676
rect 11512 9674 11568 9676
rect 11592 9674 11648 9676
rect 11352 9622 11378 9674
rect 11378 9622 11408 9674
rect 11432 9622 11442 9674
rect 11442 9622 11488 9674
rect 11512 9622 11558 9674
rect 11558 9622 11568 9674
rect 11592 9622 11622 9674
rect 11622 9622 11648 9674
rect 11352 9620 11408 9622
rect 11432 9620 11488 9622
rect 11512 9620 11568 9622
rect 11592 9620 11648 9622
rect 7886 9130 7942 9132
rect 7966 9130 8022 9132
rect 8046 9130 8102 9132
rect 8126 9130 8182 9132
rect 7886 9078 7912 9130
rect 7912 9078 7942 9130
rect 7966 9078 7976 9130
rect 7976 9078 8022 9130
rect 8046 9078 8092 9130
rect 8092 9078 8102 9130
rect 8126 9078 8156 9130
rect 8156 9078 8182 9130
rect 7886 9076 7942 9078
rect 7966 9076 8022 9078
rect 8046 9076 8102 9078
rect 8126 9076 8182 9078
rect 4421 8586 4477 8588
rect 4501 8586 4557 8588
rect 4581 8586 4637 8588
rect 4661 8586 4717 8588
rect 4421 8534 4447 8586
rect 4447 8534 4477 8586
rect 4501 8534 4511 8586
rect 4511 8534 4557 8586
rect 4581 8534 4627 8586
rect 4627 8534 4637 8586
rect 4661 8534 4691 8586
rect 4691 8534 4717 8586
rect 4421 8532 4477 8534
rect 4501 8532 4557 8534
rect 4581 8532 4637 8534
rect 4661 8532 4717 8534
rect 7886 8042 7942 8044
rect 7966 8042 8022 8044
rect 8046 8042 8102 8044
rect 8126 8042 8182 8044
rect 7886 7990 7912 8042
rect 7912 7990 7942 8042
rect 7966 7990 7976 8042
rect 7976 7990 8022 8042
rect 8046 7990 8092 8042
rect 8092 7990 8102 8042
rect 8126 7990 8156 8042
rect 8156 7990 8182 8042
rect 7886 7988 7942 7990
rect 7966 7988 8022 7990
rect 8046 7988 8102 7990
rect 8126 7988 8182 7990
rect 4421 7498 4477 7500
rect 4501 7498 4557 7500
rect 4581 7498 4637 7500
rect 4661 7498 4717 7500
rect 4421 7446 4447 7498
rect 4447 7446 4477 7498
rect 4501 7446 4511 7498
rect 4511 7446 4557 7498
rect 4581 7446 4627 7498
rect 4627 7446 4637 7498
rect 4661 7446 4691 7498
rect 4691 7446 4717 7498
rect 4421 7444 4477 7446
rect 4501 7444 4557 7446
rect 4581 7444 4637 7446
rect 4661 7444 4717 7446
rect 11352 8586 11408 8588
rect 11432 8586 11488 8588
rect 11512 8586 11568 8588
rect 11592 8586 11648 8588
rect 11352 8534 11378 8586
rect 11378 8534 11408 8586
rect 11432 8534 11442 8586
rect 11442 8534 11488 8586
rect 11512 8534 11558 8586
rect 11558 8534 11568 8586
rect 11592 8534 11622 8586
rect 11622 8534 11648 8586
rect 11352 8532 11408 8534
rect 11432 8532 11488 8534
rect 11512 8532 11568 8534
rect 11592 8532 11648 8534
rect 7886 6954 7942 6956
rect 7966 6954 8022 6956
rect 8046 6954 8102 6956
rect 8126 6954 8182 6956
rect 7886 6902 7912 6954
rect 7912 6902 7942 6954
rect 7966 6902 7976 6954
rect 7976 6902 8022 6954
rect 8046 6902 8092 6954
rect 8092 6902 8102 6954
rect 8126 6902 8156 6954
rect 8156 6902 8182 6954
rect 7886 6900 7942 6902
rect 7966 6900 8022 6902
rect 8046 6900 8102 6902
rect 8126 6900 8182 6902
rect 11352 7498 11408 7500
rect 11432 7498 11488 7500
rect 11512 7498 11568 7500
rect 11592 7498 11648 7500
rect 11352 7446 11378 7498
rect 11378 7446 11408 7498
rect 11432 7446 11442 7498
rect 11442 7446 11488 7498
rect 11512 7446 11558 7498
rect 11558 7446 11568 7498
rect 11592 7446 11622 7498
rect 11622 7446 11648 7498
rect 11352 7444 11408 7446
rect 11432 7444 11488 7446
rect 11512 7444 11568 7446
rect 11592 7444 11648 7446
rect 12530 18528 12586 18584
rect 4421 6410 4477 6412
rect 4501 6410 4557 6412
rect 4581 6410 4637 6412
rect 4661 6410 4717 6412
rect 4421 6358 4447 6410
rect 4447 6358 4477 6410
rect 4501 6358 4511 6410
rect 4511 6358 4557 6410
rect 4581 6358 4627 6410
rect 4627 6358 4637 6410
rect 4661 6358 4691 6410
rect 4691 6358 4717 6410
rect 4421 6356 4477 6358
rect 4501 6356 4557 6358
rect 4581 6356 4637 6358
rect 4661 6356 4717 6358
rect 11352 6410 11408 6412
rect 11432 6410 11488 6412
rect 11512 6410 11568 6412
rect 11592 6410 11648 6412
rect 11352 6358 11378 6410
rect 11378 6358 11408 6410
rect 11432 6358 11442 6410
rect 11442 6358 11488 6410
rect 11512 6358 11558 6410
rect 11558 6358 11568 6410
rect 11592 6358 11622 6410
rect 11622 6358 11648 6410
rect 11352 6356 11408 6358
rect 11432 6356 11488 6358
rect 11512 6356 11568 6358
rect 11592 6356 11648 6358
rect 7886 5866 7942 5868
rect 7966 5866 8022 5868
rect 8046 5866 8102 5868
rect 8126 5866 8182 5868
rect 7886 5814 7912 5866
rect 7912 5814 7942 5866
rect 7966 5814 7976 5866
rect 7976 5814 8022 5866
rect 8046 5814 8092 5866
rect 8092 5814 8102 5866
rect 8126 5814 8156 5866
rect 8156 5814 8182 5866
rect 7886 5812 7942 5814
rect 7966 5812 8022 5814
rect 8046 5812 8102 5814
rect 8126 5812 8182 5814
rect 4066 5608 4122 5664
rect 4421 5322 4477 5324
rect 4501 5322 4557 5324
rect 4581 5322 4637 5324
rect 4661 5322 4717 5324
rect 4421 5270 4447 5322
rect 4447 5270 4477 5322
rect 4501 5270 4511 5322
rect 4511 5270 4557 5322
rect 4581 5270 4627 5322
rect 4627 5270 4637 5322
rect 4661 5270 4691 5322
rect 4691 5270 4717 5322
rect 4421 5268 4477 5270
rect 4501 5268 4557 5270
rect 4581 5268 4637 5270
rect 4661 5268 4717 5270
rect 11352 5322 11408 5324
rect 11432 5322 11488 5324
rect 11512 5322 11568 5324
rect 11592 5322 11648 5324
rect 11352 5270 11378 5322
rect 11378 5270 11408 5322
rect 11432 5270 11442 5322
rect 11442 5270 11488 5322
rect 11512 5270 11558 5322
rect 11558 5270 11568 5322
rect 11592 5270 11622 5322
rect 11622 5270 11648 5322
rect 11352 5268 11408 5270
rect 11432 5268 11488 5270
rect 11512 5268 11568 5270
rect 11592 5268 11648 5270
rect 14002 18936 14058 18992
rect 14817 20010 14873 20012
rect 14897 20010 14953 20012
rect 14977 20010 15033 20012
rect 15057 20010 15113 20012
rect 14817 19958 14843 20010
rect 14843 19958 14873 20010
rect 14897 19958 14907 20010
rect 14907 19958 14953 20010
rect 14977 19958 15023 20010
rect 15023 19958 15033 20010
rect 15057 19958 15087 20010
rect 15087 19958 15113 20010
rect 14817 19956 14873 19958
rect 14897 19956 14953 19958
rect 14977 19956 15033 19958
rect 15057 19956 15113 19958
rect 14817 18922 14873 18924
rect 14897 18922 14953 18924
rect 14977 18922 15033 18924
rect 15057 18922 15113 18924
rect 14817 18870 14843 18922
rect 14843 18870 14873 18922
rect 14897 18870 14907 18922
rect 14907 18870 14953 18922
rect 14977 18870 15023 18922
rect 15023 18870 15033 18922
rect 15057 18870 15087 18922
rect 15087 18870 15113 18922
rect 14817 18868 14873 18870
rect 14897 18868 14953 18870
rect 14977 18868 15033 18870
rect 15057 18868 15113 18870
rect 7886 4778 7942 4780
rect 7966 4778 8022 4780
rect 8046 4778 8102 4780
rect 8126 4778 8182 4780
rect 7886 4726 7912 4778
rect 7912 4726 7942 4778
rect 7966 4726 7976 4778
rect 7976 4726 8022 4778
rect 8046 4726 8092 4778
rect 8092 4726 8102 4778
rect 8126 4726 8156 4778
rect 8156 4726 8182 4778
rect 7886 4724 7942 4726
rect 7966 4724 8022 4726
rect 8046 4724 8102 4726
rect 8126 4724 8182 4726
rect 4421 4234 4477 4236
rect 4501 4234 4557 4236
rect 4581 4234 4637 4236
rect 4661 4234 4717 4236
rect 4421 4182 4447 4234
rect 4447 4182 4477 4234
rect 4501 4182 4511 4234
rect 4511 4182 4557 4234
rect 4581 4182 4627 4234
rect 4627 4182 4637 4234
rect 4661 4182 4691 4234
rect 4691 4182 4717 4234
rect 4421 4180 4477 4182
rect 4501 4180 4557 4182
rect 4581 4180 4637 4182
rect 4661 4180 4717 4182
rect 11352 4234 11408 4236
rect 11432 4234 11488 4236
rect 11512 4234 11568 4236
rect 11592 4234 11648 4236
rect 11352 4182 11378 4234
rect 11378 4182 11408 4234
rect 11432 4182 11442 4234
rect 11442 4182 11488 4234
rect 11512 4182 11558 4234
rect 11558 4182 11568 4234
rect 11592 4182 11622 4234
rect 11622 4182 11648 4234
rect 11352 4180 11408 4182
rect 11432 4180 11488 4182
rect 11512 4180 11568 4182
rect 11592 4180 11648 4182
rect 7886 3690 7942 3692
rect 7966 3690 8022 3692
rect 8046 3690 8102 3692
rect 8126 3690 8182 3692
rect 7886 3638 7912 3690
rect 7912 3638 7942 3690
rect 7966 3638 7976 3690
rect 7976 3638 8022 3690
rect 8046 3638 8092 3690
rect 8092 3638 8102 3690
rect 8126 3638 8156 3690
rect 8156 3638 8182 3690
rect 7886 3636 7942 3638
rect 7966 3636 8022 3638
rect 8046 3636 8102 3638
rect 8126 3636 8182 3638
rect 4421 3146 4477 3148
rect 4501 3146 4557 3148
rect 4581 3146 4637 3148
rect 4661 3146 4717 3148
rect 4421 3094 4447 3146
rect 4447 3094 4477 3146
rect 4501 3094 4511 3146
rect 4511 3094 4557 3146
rect 4581 3094 4627 3146
rect 4627 3094 4637 3146
rect 4661 3094 4691 3146
rect 4691 3094 4717 3146
rect 4421 3092 4477 3094
rect 4501 3092 4557 3094
rect 4581 3092 4637 3094
rect 4661 3092 4717 3094
rect 11352 3146 11408 3148
rect 11432 3146 11488 3148
rect 11512 3146 11568 3148
rect 11592 3146 11648 3148
rect 11352 3094 11378 3146
rect 11378 3094 11408 3146
rect 11432 3094 11442 3146
rect 11442 3094 11488 3146
rect 11512 3094 11558 3146
rect 11558 3094 11568 3146
rect 11592 3094 11622 3146
rect 11622 3094 11648 3146
rect 11352 3092 11408 3094
rect 11432 3092 11488 3094
rect 11512 3092 11568 3094
rect 11592 3092 11648 3094
rect 7886 2602 7942 2604
rect 7966 2602 8022 2604
rect 8046 2602 8102 2604
rect 8126 2602 8182 2604
rect 7886 2550 7912 2602
rect 7912 2550 7942 2602
rect 7966 2550 7976 2602
rect 7976 2550 8022 2602
rect 8046 2550 8092 2602
rect 8092 2550 8102 2602
rect 8126 2550 8156 2602
rect 8156 2550 8182 2602
rect 7886 2548 7942 2550
rect 7966 2548 8022 2550
rect 8046 2548 8102 2550
rect 8126 2548 8182 2550
rect 4421 2058 4477 2060
rect 4501 2058 4557 2060
rect 4581 2058 4637 2060
rect 4661 2058 4717 2060
rect 4421 2006 4447 2058
rect 4447 2006 4477 2058
rect 4501 2006 4511 2058
rect 4511 2006 4557 2058
rect 4581 2006 4627 2058
rect 4627 2006 4637 2058
rect 4661 2006 4691 2058
rect 4691 2006 4717 2058
rect 4421 2004 4477 2006
rect 4501 2004 4557 2006
rect 4581 2004 4637 2006
rect 4661 2004 4717 2006
rect 11352 2058 11408 2060
rect 11432 2058 11488 2060
rect 11512 2058 11568 2060
rect 11592 2058 11648 2060
rect 11352 2006 11378 2058
rect 11378 2006 11408 2058
rect 11432 2006 11442 2058
rect 11442 2006 11488 2058
rect 11512 2006 11558 2058
rect 11558 2006 11568 2058
rect 11592 2006 11622 2058
rect 11622 2006 11648 2058
rect 11352 2004 11408 2006
rect 11432 2004 11488 2006
rect 11512 2004 11568 2006
rect 11592 2004 11648 2006
rect 14817 17834 14873 17836
rect 14897 17834 14953 17836
rect 14977 17834 15033 17836
rect 15057 17834 15113 17836
rect 14817 17782 14843 17834
rect 14843 17782 14873 17834
rect 14897 17782 14907 17834
rect 14907 17782 14953 17834
rect 14977 17782 15023 17834
rect 15023 17782 15033 17834
rect 15057 17782 15087 17834
rect 15087 17782 15113 17834
rect 14817 17780 14873 17782
rect 14897 17780 14953 17782
rect 14977 17780 15033 17782
rect 15057 17780 15113 17782
rect 14817 16746 14873 16748
rect 14897 16746 14953 16748
rect 14977 16746 15033 16748
rect 15057 16746 15113 16748
rect 14817 16694 14843 16746
rect 14843 16694 14873 16746
rect 14897 16694 14907 16746
rect 14907 16694 14953 16746
rect 14977 16694 15023 16746
rect 15023 16694 15033 16746
rect 15057 16694 15087 16746
rect 15087 16694 15113 16746
rect 14817 16692 14873 16694
rect 14897 16692 14953 16694
rect 14977 16692 15033 16694
rect 15057 16692 15113 16694
rect 14817 15658 14873 15660
rect 14897 15658 14953 15660
rect 14977 15658 15033 15660
rect 15057 15658 15113 15660
rect 14817 15606 14843 15658
rect 14843 15606 14873 15658
rect 14897 15606 14907 15658
rect 14907 15606 14953 15658
rect 14977 15606 15023 15658
rect 15023 15606 15033 15658
rect 15057 15606 15087 15658
rect 15087 15606 15113 15658
rect 14817 15604 14873 15606
rect 14897 15604 14953 15606
rect 14977 15604 15033 15606
rect 15057 15604 15113 15606
rect 14817 14570 14873 14572
rect 14897 14570 14953 14572
rect 14977 14570 15033 14572
rect 15057 14570 15113 14572
rect 14817 14518 14843 14570
rect 14843 14518 14873 14570
rect 14897 14518 14907 14570
rect 14907 14518 14953 14570
rect 14977 14518 15023 14570
rect 15023 14518 15033 14570
rect 15057 14518 15087 14570
rect 15087 14518 15113 14570
rect 14817 14516 14873 14518
rect 14897 14516 14953 14518
rect 14977 14516 15033 14518
rect 15057 14516 15113 14518
rect 14817 13482 14873 13484
rect 14897 13482 14953 13484
rect 14977 13482 15033 13484
rect 15057 13482 15113 13484
rect 14817 13430 14843 13482
rect 14843 13430 14873 13482
rect 14897 13430 14907 13482
rect 14907 13430 14953 13482
rect 14977 13430 15023 13482
rect 15023 13430 15033 13482
rect 15057 13430 15087 13482
rect 15087 13430 15113 13482
rect 14817 13428 14873 13430
rect 14897 13428 14953 13430
rect 14977 13428 15033 13430
rect 15057 13428 15113 13430
rect 14817 12394 14873 12396
rect 14897 12394 14953 12396
rect 14977 12394 15033 12396
rect 15057 12394 15113 12396
rect 14817 12342 14843 12394
rect 14843 12342 14873 12394
rect 14897 12342 14907 12394
rect 14907 12342 14953 12394
rect 14977 12342 15023 12394
rect 15023 12342 15033 12394
rect 15057 12342 15087 12394
rect 15087 12342 15113 12394
rect 14817 12340 14873 12342
rect 14897 12340 14953 12342
rect 14977 12340 15033 12342
rect 15057 12340 15113 12342
rect 15566 18664 15622 18720
rect 14817 11306 14873 11308
rect 14897 11306 14953 11308
rect 14977 11306 15033 11308
rect 15057 11306 15113 11308
rect 14817 11254 14843 11306
rect 14843 11254 14873 11306
rect 14897 11254 14907 11306
rect 14907 11254 14953 11306
rect 14977 11254 15023 11306
rect 15023 11254 15033 11306
rect 15057 11254 15087 11306
rect 15087 11254 15113 11306
rect 14817 11252 14873 11254
rect 14897 11252 14953 11254
rect 14977 11252 15033 11254
rect 15057 11252 15113 11254
rect 14817 10218 14873 10220
rect 14897 10218 14953 10220
rect 14977 10218 15033 10220
rect 15057 10218 15113 10220
rect 14817 10166 14843 10218
rect 14843 10166 14873 10218
rect 14897 10166 14907 10218
rect 14907 10166 14953 10218
rect 14977 10166 15023 10218
rect 15023 10166 15033 10218
rect 15057 10166 15087 10218
rect 15087 10166 15113 10218
rect 14817 10164 14873 10166
rect 14897 10164 14953 10166
rect 14977 10164 15033 10166
rect 15057 10164 15113 10166
rect 14817 9130 14873 9132
rect 14897 9130 14953 9132
rect 14977 9130 15033 9132
rect 15057 9130 15113 9132
rect 14817 9078 14843 9130
rect 14843 9078 14873 9130
rect 14897 9078 14907 9130
rect 14907 9078 14953 9130
rect 14977 9078 15023 9130
rect 15023 9078 15033 9130
rect 15057 9078 15087 9130
rect 15087 9078 15113 9130
rect 14817 9076 14873 9078
rect 14897 9076 14953 9078
rect 14977 9076 15033 9078
rect 15057 9076 15113 9078
rect 14817 8042 14873 8044
rect 14897 8042 14953 8044
rect 14977 8042 15033 8044
rect 15057 8042 15113 8044
rect 14817 7990 14843 8042
rect 14843 7990 14873 8042
rect 14897 7990 14907 8042
rect 14907 7990 14953 8042
rect 14977 7990 15023 8042
rect 15023 7990 15033 8042
rect 15057 7990 15087 8042
rect 15087 7990 15113 8042
rect 14817 7988 14873 7990
rect 14897 7988 14953 7990
rect 14977 7988 15033 7990
rect 15057 7988 15113 7990
rect 18602 21520 18658 21576
rect 18282 20554 18338 20556
rect 18362 20554 18418 20556
rect 18442 20554 18498 20556
rect 18522 20554 18578 20556
rect 18282 20502 18308 20554
rect 18308 20502 18338 20554
rect 18362 20502 18372 20554
rect 18372 20502 18418 20554
rect 18442 20502 18488 20554
rect 18488 20502 18498 20554
rect 18522 20502 18552 20554
rect 18552 20502 18578 20554
rect 18282 20500 18338 20502
rect 18362 20500 18418 20502
rect 18442 20500 18498 20502
rect 18522 20500 18578 20502
rect 18282 19466 18338 19468
rect 18362 19466 18418 19468
rect 18442 19466 18498 19468
rect 18522 19466 18578 19468
rect 18282 19414 18308 19466
rect 18308 19414 18338 19466
rect 18362 19414 18372 19466
rect 18372 19414 18418 19466
rect 18442 19414 18488 19466
rect 18488 19414 18498 19466
rect 18522 19414 18552 19466
rect 18552 19414 18578 19466
rect 18282 19412 18338 19414
rect 18362 19412 18418 19414
rect 18442 19412 18498 19414
rect 18522 19412 18578 19414
rect 18326 19108 18328 19128
rect 18328 19108 18380 19128
rect 18380 19108 18382 19128
rect 18326 19072 18382 19108
rect 18418 18528 18474 18584
rect 18282 18378 18338 18380
rect 18362 18378 18418 18380
rect 18442 18378 18498 18380
rect 18522 18378 18578 18380
rect 18282 18326 18308 18378
rect 18308 18326 18338 18378
rect 18362 18326 18372 18378
rect 18372 18326 18418 18378
rect 18442 18326 18488 18378
rect 18488 18326 18498 18378
rect 18522 18326 18552 18378
rect 18552 18326 18578 18378
rect 18282 18324 18338 18326
rect 18362 18324 18418 18326
rect 18442 18324 18498 18326
rect 18522 18324 18578 18326
rect 20166 22064 20222 22120
rect 18878 18528 18934 18584
rect 18282 17290 18338 17292
rect 18362 17290 18418 17292
rect 18442 17290 18498 17292
rect 18522 17290 18578 17292
rect 18282 17238 18308 17290
rect 18308 17238 18338 17290
rect 18362 17238 18372 17290
rect 18372 17238 18418 17290
rect 18442 17238 18488 17290
rect 18488 17238 18498 17290
rect 18522 17238 18552 17290
rect 18552 17238 18578 17290
rect 18282 17236 18338 17238
rect 18362 17236 18418 17238
rect 18442 17236 18498 17238
rect 18522 17236 18578 17238
rect 18282 16202 18338 16204
rect 18362 16202 18418 16204
rect 18442 16202 18498 16204
rect 18522 16202 18578 16204
rect 18282 16150 18308 16202
rect 18308 16150 18338 16202
rect 18362 16150 18372 16202
rect 18372 16150 18418 16202
rect 18442 16150 18488 16202
rect 18488 16150 18498 16202
rect 18522 16150 18552 16202
rect 18552 16150 18578 16202
rect 18282 16148 18338 16150
rect 18362 16148 18418 16150
rect 18442 16148 18498 16150
rect 18522 16148 18578 16150
rect 18282 15114 18338 15116
rect 18362 15114 18418 15116
rect 18442 15114 18498 15116
rect 18522 15114 18578 15116
rect 18282 15062 18308 15114
rect 18308 15062 18338 15114
rect 18362 15062 18372 15114
rect 18372 15062 18418 15114
rect 18442 15062 18488 15114
rect 18488 15062 18498 15114
rect 18522 15062 18552 15114
rect 18552 15062 18578 15114
rect 18282 15060 18338 15062
rect 18362 15060 18418 15062
rect 18442 15060 18498 15062
rect 18522 15060 18578 15062
rect 18282 14026 18338 14028
rect 18362 14026 18418 14028
rect 18442 14026 18498 14028
rect 18522 14026 18578 14028
rect 18282 13974 18308 14026
rect 18308 13974 18338 14026
rect 18362 13974 18372 14026
rect 18372 13974 18418 14026
rect 18442 13974 18488 14026
rect 18488 13974 18498 14026
rect 18522 13974 18552 14026
rect 18552 13974 18578 14026
rect 18282 13972 18338 13974
rect 18362 13972 18418 13974
rect 18442 13972 18498 13974
rect 18522 13972 18578 13974
rect 19522 18392 19578 18448
rect 18282 12938 18338 12940
rect 18362 12938 18418 12940
rect 18442 12938 18498 12940
rect 18522 12938 18578 12940
rect 18282 12886 18308 12938
rect 18308 12886 18338 12938
rect 18362 12886 18372 12938
rect 18372 12886 18418 12938
rect 18442 12886 18488 12938
rect 18488 12886 18498 12938
rect 18522 12886 18552 12938
rect 18552 12886 18578 12938
rect 18282 12884 18338 12886
rect 18362 12884 18418 12886
rect 18442 12884 18498 12886
rect 18522 12884 18578 12886
rect 18282 11850 18338 11852
rect 18362 11850 18418 11852
rect 18442 11850 18498 11852
rect 18522 11850 18578 11852
rect 18282 11798 18308 11850
rect 18308 11798 18338 11850
rect 18362 11798 18372 11850
rect 18372 11798 18418 11850
rect 18442 11798 18488 11850
rect 18488 11798 18498 11850
rect 18522 11798 18552 11850
rect 18552 11798 18578 11850
rect 18282 11796 18338 11798
rect 18362 11796 18418 11798
rect 18442 11796 18498 11798
rect 18522 11796 18578 11798
rect 18282 10762 18338 10764
rect 18362 10762 18418 10764
rect 18442 10762 18498 10764
rect 18522 10762 18578 10764
rect 18282 10710 18308 10762
rect 18308 10710 18338 10762
rect 18362 10710 18372 10762
rect 18372 10710 18418 10762
rect 18442 10710 18488 10762
rect 18488 10710 18498 10762
rect 18522 10710 18552 10762
rect 18552 10710 18578 10762
rect 18282 10708 18338 10710
rect 18362 10708 18418 10710
rect 18442 10708 18498 10710
rect 18522 10708 18578 10710
rect 18282 9674 18338 9676
rect 18362 9674 18418 9676
rect 18442 9674 18498 9676
rect 18522 9674 18578 9676
rect 18282 9622 18308 9674
rect 18308 9622 18338 9674
rect 18362 9622 18372 9674
rect 18372 9622 18418 9674
rect 18442 9622 18488 9674
rect 18488 9622 18498 9674
rect 18522 9622 18552 9674
rect 18552 9622 18578 9674
rect 18282 9620 18338 9622
rect 18362 9620 18418 9622
rect 18442 9620 18498 9622
rect 18522 9620 18578 9622
rect 14817 6954 14873 6956
rect 14897 6954 14953 6956
rect 14977 6954 15033 6956
rect 15057 6954 15113 6956
rect 14817 6902 14843 6954
rect 14843 6902 14873 6954
rect 14897 6902 14907 6954
rect 14907 6902 14953 6954
rect 14977 6902 15023 6954
rect 15023 6902 15033 6954
rect 15057 6902 15087 6954
rect 15087 6902 15113 6954
rect 14817 6900 14873 6902
rect 14897 6900 14953 6902
rect 14977 6900 15033 6902
rect 15057 6900 15113 6902
rect 14817 5866 14873 5868
rect 14897 5866 14953 5868
rect 14977 5866 15033 5868
rect 15057 5866 15113 5868
rect 14817 5814 14843 5866
rect 14843 5814 14873 5866
rect 14897 5814 14907 5866
rect 14907 5814 14953 5866
rect 14977 5814 15023 5866
rect 15023 5814 15033 5866
rect 15057 5814 15087 5866
rect 15087 5814 15113 5866
rect 14817 5812 14873 5814
rect 14897 5812 14953 5814
rect 14977 5812 15033 5814
rect 15057 5812 15113 5814
rect 14817 4778 14873 4780
rect 14897 4778 14953 4780
rect 14977 4778 15033 4780
rect 15057 4778 15113 4780
rect 14817 4726 14843 4778
rect 14843 4726 14873 4778
rect 14897 4726 14907 4778
rect 14907 4726 14953 4778
rect 14977 4726 15023 4778
rect 15023 4726 15033 4778
rect 15057 4726 15087 4778
rect 15087 4726 15113 4778
rect 14817 4724 14873 4726
rect 14897 4724 14953 4726
rect 14977 4724 15033 4726
rect 15057 4724 15113 4726
rect 18282 8586 18338 8588
rect 18362 8586 18418 8588
rect 18442 8586 18498 8588
rect 18522 8586 18578 8588
rect 18282 8534 18308 8586
rect 18308 8534 18338 8586
rect 18362 8534 18372 8586
rect 18372 8534 18418 8586
rect 18442 8534 18488 8586
rect 18488 8534 18498 8586
rect 18522 8534 18552 8586
rect 18552 8534 18578 8586
rect 18282 8532 18338 8534
rect 18362 8532 18418 8534
rect 18442 8532 18498 8534
rect 18522 8532 18578 8534
rect 18282 7498 18338 7500
rect 18362 7498 18418 7500
rect 18442 7498 18498 7500
rect 18522 7498 18578 7500
rect 18282 7446 18308 7498
rect 18308 7446 18338 7498
rect 18362 7446 18372 7498
rect 18372 7446 18418 7498
rect 18442 7446 18488 7498
rect 18488 7446 18498 7498
rect 18522 7446 18552 7498
rect 18552 7446 18578 7498
rect 18282 7444 18338 7446
rect 18362 7444 18418 7446
rect 18442 7444 18498 7446
rect 18522 7444 18578 7446
rect 18282 6410 18338 6412
rect 18362 6410 18418 6412
rect 18442 6410 18498 6412
rect 18522 6410 18578 6412
rect 18282 6358 18308 6410
rect 18308 6358 18338 6410
rect 18362 6358 18372 6410
rect 18372 6358 18418 6410
rect 18442 6358 18488 6410
rect 18488 6358 18498 6410
rect 18522 6358 18552 6410
rect 18552 6358 18578 6410
rect 18282 6356 18338 6358
rect 18362 6356 18418 6358
rect 18442 6356 18498 6358
rect 18522 6356 18578 6358
rect 17958 5472 18014 5528
rect 18282 5322 18338 5324
rect 18362 5322 18418 5324
rect 18442 5322 18498 5324
rect 18522 5322 18578 5324
rect 18282 5270 18308 5322
rect 18308 5270 18338 5322
rect 18362 5270 18372 5322
rect 18372 5270 18418 5322
rect 18442 5270 18488 5322
rect 18488 5270 18498 5322
rect 18522 5270 18552 5322
rect 18552 5270 18578 5322
rect 18282 5268 18338 5270
rect 18362 5268 18418 5270
rect 18442 5268 18498 5270
rect 18522 5268 18578 5270
rect 17958 4520 18014 4576
rect 18282 4234 18338 4236
rect 18362 4234 18418 4236
rect 18442 4234 18498 4236
rect 18522 4234 18578 4236
rect 18282 4182 18308 4234
rect 18308 4182 18338 4234
rect 18362 4182 18372 4234
rect 18372 4182 18418 4234
rect 18442 4182 18488 4234
rect 18488 4182 18498 4234
rect 18522 4182 18552 4234
rect 18552 4182 18578 4234
rect 18282 4180 18338 4182
rect 18362 4180 18418 4182
rect 18442 4180 18498 4182
rect 18522 4180 18578 4182
rect 14817 3690 14873 3692
rect 14897 3690 14953 3692
rect 14977 3690 15033 3692
rect 15057 3690 15113 3692
rect 14817 3638 14843 3690
rect 14843 3638 14873 3690
rect 14897 3638 14907 3690
rect 14907 3638 14953 3690
rect 14977 3638 15023 3690
rect 15023 3638 15033 3690
rect 15057 3638 15087 3690
rect 15087 3638 15113 3690
rect 14817 3636 14873 3638
rect 14897 3636 14953 3638
rect 14977 3636 15033 3638
rect 15057 3636 15113 3638
rect 18282 3146 18338 3148
rect 18362 3146 18418 3148
rect 18442 3146 18498 3148
rect 18522 3146 18578 3148
rect 18282 3094 18308 3146
rect 18308 3094 18338 3146
rect 18362 3094 18372 3146
rect 18372 3094 18418 3146
rect 18442 3094 18488 3146
rect 18488 3094 18498 3146
rect 18522 3094 18552 3146
rect 18552 3094 18578 3146
rect 18282 3092 18338 3094
rect 18362 3092 18418 3094
rect 18442 3092 18498 3094
rect 18522 3092 18578 3094
rect 18786 3160 18842 3216
rect 19706 12408 19762 12464
rect 20534 21112 20590 21168
rect 20626 20704 20682 20760
rect 20442 20160 20498 20216
rect 21086 19752 21142 19808
rect 20994 19208 21050 19264
rect 20626 18800 20682 18856
rect 20442 17460 20498 17496
rect 20442 17440 20444 17460
rect 20444 17440 20496 17460
rect 20496 17440 20498 17460
rect 20534 14176 20590 14232
rect 20442 13768 20498 13824
rect 20258 12816 20314 12872
rect 21086 17884 21088 17904
rect 21088 17884 21140 17904
rect 21140 17884 21142 17904
rect 21086 17848 21142 17884
rect 20994 17032 21050 17088
rect 21086 16488 21142 16544
rect 21086 16100 21142 16136
rect 21086 16080 21088 16100
rect 21088 16080 21140 16100
rect 21140 16080 21142 16100
rect 20994 15164 20996 15184
rect 20996 15164 21048 15184
rect 21048 15164 21050 15184
rect 20994 15128 21050 15164
rect 21178 15536 21234 15592
rect 20626 11864 20682 11920
rect 20902 11048 20958 11104
rect 20626 10504 20682 10560
rect 20074 10116 20130 10152
rect 20074 10096 20076 10116
rect 20076 10096 20128 10116
rect 20128 10096 20130 10116
rect 20626 9552 20682 9608
rect 20534 9144 20590 9200
rect 20902 8736 20958 8792
rect 20626 7784 20682 7840
rect 20810 7376 20866 7432
rect 19246 6424 19302 6480
rect 20902 6832 20958 6888
rect 19154 3704 19210 3760
rect 14817 2602 14873 2604
rect 14897 2602 14953 2604
rect 14977 2602 15033 2604
rect 15057 2602 15113 2604
rect 14817 2550 14843 2602
rect 14843 2550 14873 2602
rect 14897 2550 14907 2602
rect 14907 2550 14953 2602
rect 14977 2550 15023 2602
rect 15023 2550 15033 2602
rect 15057 2550 15087 2602
rect 15087 2550 15113 2602
rect 14817 2548 14873 2550
rect 14897 2548 14953 2550
rect 14977 2548 15033 2550
rect 15057 2548 15113 2550
rect 18142 2208 18198 2264
rect 18282 2058 18338 2060
rect 18362 2058 18418 2060
rect 18442 2058 18498 2060
rect 18522 2058 18578 2060
rect 18282 2006 18308 2058
rect 18308 2006 18338 2058
rect 18362 2006 18372 2058
rect 18372 2006 18418 2058
rect 18442 2006 18488 2058
rect 18488 2006 18498 2058
rect 18522 2006 18552 2058
rect 18552 2006 18578 2058
rect 18282 2004 18338 2006
rect 18362 2004 18418 2006
rect 18442 2004 18498 2006
rect 18522 2004 18578 2006
rect 18142 1392 18198 1448
rect 17958 440 18014 496
rect 18878 1800 18934 1856
rect 21086 14720 21142 14776
rect 21086 13360 21142 13416
rect 22006 11492 22008 11512
rect 22008 11492 22060 11512
rect 22060 11492 22062 11512
rect 22006 11456 22062 11492
rect 22006 8228 22008 8248
rect 22008 8228 22060 8248
rect 22060 8228 22062 8248
rect 22006 8192 22062 8228
rect 21362 5880 21418 5936
rect 21270 5100 21272 5120
rect 21272 5100 21324 5120
rect 21324 5100 21326 5120
rect 21270 5064 21326 5100
rect 21270 4132 21326 4168
rect 21270 4112 21272 4132
rect 21272 4112 21324 4132
rect 21324 4112 21326 4132
rect 19246 2752 19302 2808
rect 19154 848 19210 904
rect 18786 32 18842 88
<< metal3 >>
rect 19241 22530 19307 22533
rect 22200 22530 23000 22560
rect 19241 22528 23000 22530
rect 19241 22472 19246 22528
rect 19302 22472 23000 22528
rect 19241 22470 23000 22472
rect 19241 22467 19307 22470
rect 22200 22440 23000 22470
rect 20161 22122 20227 22125
rect 22200 22122 23000 22152
rect 20161 22120 23000 22122
rect 20161 22064 20166 22120
rect 20222 22064 23000 22120
rect 20161 22062 23000 22064
rect 20161 22059 20227 22062
rect 22200 22032 23000 22062
rect 18597 21578 18663 21581
rect 22200 21578 23000 21608
rect 18597 21576 23000 21578
rect 18597 21520 18602 21576
rect 18658 21520 23000 21576
rect 18597 21518 23000 21520
rect 18597 21515 18663 21518
rect 22200 21488 23000 21518
rect 20529 21170 20595 21173
rect 22200 21170 23000 21200
rect 20529 21168 23000 21170
rect 20529 21112 20534 21168
rect 20590 21112 23000 21168
rect 20529 21110 23000 21112
rect 20529 21107 20595 21110
rect 22200 21080 23000 21110
rect 20621 20762 20687 20765
rect 22200 20762 23000 20792
rect 20621 20760 23000 20762
rect 20621 20704 20626 20760
rect 20682 20704 23000 20760
rect 20621 20702 23000 20704
rect 20621 20699 20687 20702
rect 22200 20672 23000 20702
rect 4409 20560 4729 20561
rect 4409 20496 4417 20560
rect 4481 20496 4497 20560
rect 4561 20496 4577 20560
rect 4641 20496 4657 20560
rect 4721 20496 4729 20560
rect 4409 20495 4729 20496
rect 11340 20560 11660 20561
rect 11340 20496 11348 20560
rect 11412 20496 11428 20560
rect 11492 20496 11508 20560
rect 11572 20496 11588 20560
rect 11652 20496 11660 20560
rect 11340 20495 11660 20496
rect 18270 20560 18590 20561
rect 18270 20496 18278 20560
rect 18342 20496 18358 20560
rect 18422 20496 18438 20560
rect 18502 20496 18518 20560
rect 18582 20496 18590 20560
rect 18270 20495 18590 20496
rect 20437 20218 20503 20221
rect 22200 20218 23000 20248
rect 20437 20216 23000 20218
rect 20437 20160 20442 20216
rect 20498 20160 23000 20216
rect 20437 20158 23000 20160
rect 20437 20155 20503 20158
rect 22200 20128 23000 20158
rect 7874 20016 8194 20017
rect 7874 19952 7882 20016
rect 7946 19952 7962 20016
rect 8026 19952 8042 20016
rect 8106 19952 8122 20016
rect 8186 19952 8194 20016
rect 7874 19951 8194 19952
rect 14805 20016 15125 20017
rect 14805 19952 14813 20016
rect 14877 19952 14893 20016
rect 14957 19952 14973 20016
rect 15037 19952 15053 20016
rect 15117 19952 15125 20016
rect 14805 19951 15125 19952
rect 21081 19810 21147 19813
rect 22200 19810 23000 19840
rect 21081 19808 23000 19810
rect 21081 19752 21086 19808
rect 21142 19752 23000 19808
rect 21081 19750 23000 19752
rect 21081 19747 21147 19750
rect 22200 19720 23000 19750
rect 4409 19472 4729 19473
rect 4409 19408 4417 19472
rect 4481 19408 4497 19472
rect 4561 19408 4577 19472
rect 4641 19408 4657 19472
rect 4721 19408 4729 19472
rect 4409 19407 4729 19408
rect 11340 19472 11660 19473
rect 11340 19408 11348 19472
rect 11412 19408 11428 19472
rect 11492 19408 11508 19472
rect 11572 19408 11588 19472
rect 11652 19408 11660 19472
rect 11340 19407 11660 19408
rect 18270 19472 18590 19473
rect 18270 19408 18278 19472
rect 18342 19408 18358 19472
rect 18422 19408 18438 19472
rect 18502 19408 18518 19472
rect 18582 19408 18590 19472
rect 18270 19407 18590 19408
rect 20989 19266 21055 19269
rect 22200 19266 23000 19296
rect 20989 19264 23000 19266
rect 20989 19208 20994 19264
rect 21050 19208 23000 19264
rect 20989 19206 23000 19208
rect 20989 19203 21055 19206
rect 22200 19176 23000 19206
rect 11145 19130 11211 19133
rect 18321 19130 18387 19133
rect 11145 19128 18387 19130
rect 11145 19072 11150 19128
rect 11206 19072 18326 19128
rect 18382 19072 18387 19128
rect 11145 19070 18387 19072
rect 11145 19067 11211 19070
rect 18321 19067 18387 19070
rect 10317 18994 10383 18997
rect 13997 18994 14063 18997
rect 10317 18992 14063 18994
rect 10317 18936 10322 18992
rect 10378 18936 14002 18992
rect 14058 18936 14063 18992
rect 10317 18934 14063 18936
rect 10317 18931 10383 18934
rect 13997 18931 14063 18934
rect 7874 18928 8194 18929
rect 7874 18864 7882 18928
rect 7946 18864 7962 18928
rect 8026 18864 8042 18928
rect 8106 18864 8122 18928
rect 8186 18864 8194 18928
rect 7874 18863 8194 18864
rect 14805 18928 15125 18929
rect 14805 18864 14813 18928
rect 14877 18864 14893 18928
rect 14957 18864 14973 18928
rect 15037 18864 15053 18928
rect 15117 18864 15125 18928
rect 14805 18863 15125 18864
rect 20621 18858 20687 18861
rect 22200 18858 23000 18888
rect 20621 18856 23000 18858
rect 20621 18800 20626 18856
rect 20682 18800 23000 18856
rect 20621 18798 23000 18800
rect 20621 18795 20687 18798
rect 22200 18768 23000 18798
rect 11421 18722 11487 18725
rect 15561 18722 15627 18725
rect 11421 18720 15627 18722
rect 11421 18664 11426 18720
rect 11482 18664 15566 18720
rect 15622 18664 15627 18720
rect 11421 18662 15627 18664
rect 11421 18659 11487 18662
rect 15561 18659 15627 18662
rect 11237 18586 11303 18589
rect 12525 18586 12591 18589
rect 11237 18584 12591 18586
rect 11237 18528 11242 18584
rect 11298 18528 12530 18584
rect 12586 18528 12591 18584
rect 11237 18526 12591 18528
rect 11237 18523 11303 18526
rect 12525 18523 12591 18526
rect 18413 18586 18479 18589
rect 18873 18586 18939 18589
rect 18413 18584 18939 18586
rect 18413 18528 18418 18584
rect 18474 18528 18878 18584
rect 18934 18528 18939 18584
rect 18413 18526 18939 18528
rect 18413 18523 18479 18526
rect 18873 18523 18939 18526
rect 19517 18450 19583 18453
rect 22200 18450 23000 18480
rect 19517 18448 23000 18450
rect 19517 18392 19522 18448
rect 19578 18392 23000 18448
rect 19517 18390 23000 18392
rect 19517 18387 19583 18390
rect 4409 18384 4729 18385
rect 4409 18320 4417 18384
rect 4481 18320 4497 18384
rect 4561 18320 4577 18384
rect 4641 18320 4657 18384
rect 4721 18320 4729 18384
rect 4409 18319 4729 18320
rect 11340 18384 11660 18385
rect 11340 18320 11348 18384
rect 11412 18320 11428 18384
rect 11492 18320 11508 18384
rect 11572 18320 11588 18384
rect 11652 18320 11660 18384
rect 11340 18319 11660 18320
rect 18270 18384 18590 18385
rect 18270 18320 18278 18384
rect 18342 18320 18358 18384
rect 18422 18320 18438 18384
rect 18502 18320 18518 18384
rect 18582 18320 18590 18384
rect 22200 18360 23000 18390
rect 18270 18319 18590 18320
rect 6361 18178 6427 18181
rect 11605 18178 11671 18181
rect 6361 18176 11671 18178
rect 6361 18120 6366 18176
rect 6422 18120 11610 18176
rect 11666 18120 11671 18176
rect 6361 18118 11671 18120
rect 6361 18115 6427 18118
rect 11605 18115 11671 18118
rect 21081 17906 21147 17909
rect 22200 17906 23000 17936
rect 21081 17904 23000 17906
rect 21081 17848 21086 17904
rect 21142 17848 23000 17904
rect 21081 17846 23000 17848
rect 21081 17843 21147 17846
rect 7874 17840 8194 17841
rect 7874 17776 7882 17840
rect 7946 17776 7962 17840
rect 8026 17776 8042 17840
rect 8106 17776 8122 17840
rect 8186 17776 8194 17840
rect 7874 17775 8194 17776
rect 14805 17840 15125 17841
rect 14805 17776 14813 17840
rect 14877 17776 14893 17840
rect 14957 17776 14973 17840
rect 15037 17776 15053 17840
rect 15117 17776 15125 17840
rect 22200 17816 23000 17846
rect 14805 17775 15125 17776
rect 20437 17498 20503 17501
rect 22200 17498 23000 17528
rect 20437 17496 23000 17498
rect 20437 17440 20442 17496
rect 20498 17440 23000 17496
rect 20437 17438 23000 17440
rect 20437 17435 20503 17438
rect 22200 17408 23000 17438
rect 4409 17296 4729 17297
rect 4409 17232 4417 17296
rect 4481 17232 4497 17296
rect 4561 17232 4577 17296
rect 4641 17232 4657 17296
rect 4721 17232 4729 17296
rect 4409 17231 4729 17232
rect 11340 17296 11660 17297
rect 11340 17232 11348 17296
rect 11412 17232 11428 17296
rect 11492 17232 11508 17296
rect 11572 17232 11588 17296
rect 11652 17232 11660 17296
rect 11340 17231 11660 17232
rect 18270 17296 18590 17297
rect 18270 17232 18278 17296
rect 18342 17232 18358 17296
rect 18422 17232 18438 17296
rect 18502 17232 18518 17296
rect 18582 17232 18590 17296
rect 18270 17231 18590 17232
rect 0 17090 800 17120
rect 4797 17090 4863 17093
rect 0 17088 4863 17090
rect 0 17032 4802 17088
rect 4858 17032 4863 17088
rect 0 17030 4863 17032
rect 0 17000 800 17030
rect 4797 17027 4863 17030
rect 20989 17090 21055 17093
rect 22200 17090 23000 17120
rect 20989 17088 23000 17090
rect 20989 17032 20994 17088
rect 21050 17032 23000 17088
rect 20989 17030 23000 17032
rect 20989 17027 21055 17030
rect 22200 17000 23000 17030
rect 7874 16752 8194 16753
rect 7874 16688 7882 16752
rect 7946 16688 7962 16752
rect 8026 16688 8042 16752
rect 8106 16688 8122 16752
rect 8186 16688 8194 16752
rect 7874 16687 8194 16688
rect 14805 16752 15125 16753
rect 14805 16688 14813 16752
rect 14877 16688 14893 16752
rect 14957 16688 14973 16752
rect 15037 16688 15053 16752
rect 15117 16688 15125 16752
rect 14805 16687 15125 16688
rect 21081 16546 21147 16549
rect 22200 16546 23000 16576
rect 21081 16544 23000 16546
rect 21081 16488 21086 16544
rect 21142 16488 23000 16544
rect 21081 16486 23000 16488
rect 21081 16483 21147 16486
rect 22200 16456 23000 16486
rect 4409 16208 4729 16209
rect 4409 16144 4417 16208
rect 4481 16144 4497 16208
rect 4561 16144 4577 16208
rect 4641 16144 4657 16208
rect 4721 16144 4729 16208
rect 4409 16143 4729 16144
rect 11340 16208 11660 16209
rect 11340 16144 11348 16208
rect 11412 16144 11428 16208
rect 11492 16144 11508 16208
rect 11572 16144 11588 16208
rect 11652 16144 11660 16208
rect 11340 16143 11660 16144
rect 18270 16208 18590 16209
rect 18270 16144 18278 16208
rect 18342 16144 18358 16208
rect 18422 16144 18438 16208
rect 18502 16144 18518 16208
rect 18582 16144 18590 16208
rect 18270 16143 18590 16144
rect 21081 16138 21147 16141
rect 22200 16138 23000 16168
rect 21081 16136 23000 16138
rect 21081 16080 21086 16136
rect 21142 16080 23000 16136
rect 21081 16078 23000 16080
rect 21081 16075 21147 16078
rect 22200 16048 23000 16078
rect 7874 15664 8194 15665
rect 7874 15600 7882 15664
rect 7946 15600 7962 15664
rect 8026 15600 8042 15664
rect 8106 15600 8122 15664
rect 8186 15600 8194 15664
rect 7874 15599 8194 15600
rect 14805 15664 15125 15665
rect 14805 15600 14813 15664
rect 14877 15600 14893 15664
rect 14957 15600 14973 15664
rect 15037 15600 15053 15664
rect 15117 15600 15125 15664
rect 14805 15599 15125 15600
rect 21173 15594 21239 15597
rect 22200 15594 23000 15624
rect 21173 15592 23000 15594
rect 21173 15536 21178 15592
rect 21234 15536 23000 15592
rect 21173 15534 23000 15536
rect 21173 15531 21239 15534
rect 22200 15504 23000 15534
rect 20989 15186 21055 15189
rect 22200 15186 23000 15216
rect 20989 15184 23000 15186
rect 20989 15128 20994 15184
rect 21050 15128 23000 15184
rect 20989 15126 23000 15128
rect 20989 15123 21055 15126
rect 4409 15120 4729 15121
rect 4409 15056 4417 15120
rect 4481 15056 4497 15120
rect 4561 15056 4577 15120
rect 4641 15056 4657 15120
rect 4721 15056 4729 15120
rect 4409 15055 4729 15056
rect 11340 15120 11660 15121
rect 11340 15056 11348 15120
rect 11412 15056 11428 15120
rect 11492 15056 11508 15120
rect 11572 15056 11588 15120
rect 11652 15056 11660 15120
rect 11340 15055 11660 15056
rect 18270 15120 18590 15121
rect 18270 15056 18278 15120
rect 18342 15056 18358 15120
rect 18422 15056 18438 15120
rect 18502 15056 18518 15120
rect 18582 15056 18590 15120
rect 22200 15096 23000 15126
rect 18270 15055 18590 15056
rect 21081 14778 21147 14781
rect 22200 14778 23000 14808
rect 21081 14776 23000 14778
rect 21081 14720 21086 14776
rect 21142 14720 23000 14776
rect 21081 14718 23000 14720
rect 21081 14715 21147 14718
rect 22200 14688 23000 14718
rect 7874 14576 8194 14577
rect 7874 14512 7882 14576
rect 7946 14512 7962 14576
rect 8026 14512 8042 14576
rect 8106 14512 8122 14576
rect 8186 14512 8194 14576
rect 7874 14511 8194 14512
rect 14805 14576 15125 14577
rect 14805 14512 14813 14576
rect 14877 14512 14893 14576
rect 14957 14512 14973 14576
rect 15037 14512 15053 14576
rect 15117 14512 15125 14576
rect 14805 14511 15125 14512
rect 20529 14234 20595 14237
rect 22200 14234 23000 14264
rect 20529 14232 23000 14234
rect 20529 14176 20534 14232
rect 20590 14176 23000 14232
rect 20529 14174 23000 14176
rect 20529 14171 20595 14174
rect 22200 14144 23000 14174
rect 4409 14032 4729 14033
rect 4409 13968 4417 14032
rect 4481 13968 4497 14032
rect 4561 13968 4577 14032
rect 4641 13968 4657 14032
rect 4721 13968 4729 14032
rect 4409 13967 4729 13968
rect 11340 14032 11660 14033
rect 11340 13968 11348 14032
rect 11412 13968 11428 14032
rect 11492 13968 11508 14032
rect 11572 13968 11588 14032
rect 11652 13968 11660 14032
rect 11340 13967 11660 13968
rect 18270 14032 18590 14033
rect 18270 13968 18278 14032
rect 18342 13968 18358 14032
rect 18422 13968 18438 14032
rect 18502 13968 18518 14032
rect 18582 13968 18590 14032
rect 18270 13967 18590 13968
rect 20437 13826 20503 13829
rect 22200 13826 23000 13856
rect 20437 13824 23000 13826
rect 20437 13768 20442 13824
rect 20498 13768 23000 13824
rect 20437 13766 23000 13768
rect 20437 13763 20503 13766
rect 22200 13736 23000 13766
rect 7874 13488 8194 13489
rect 7874 13424 7882 13488
rect 7946 13424 7962 13488
rect 8026 13424 8042 13488
rect 8106 13424 8122 13488
rect 8186 13424 8194 13488
rect 7874 13423 8194 13424
rect 14805 13488 15125 13489
rect 14805 13424 14813 13488
rect 14877 13424 14893 13488
rect 14957 13424 14973 13488
rect 15037 13424 15053 13488
rect 15117 13424 15125 13488
rect 14805 13423 15125 13424
rect 21081 13418 21147 13421
rect 22200 13418 23000 13448
rect 21081 13416 23000 13418
rect 21081 13360 21086 13416
rect 21142 13360 23000 13416
rect 21081 13358 23000 13360
rect 21081 13355 21147 13358
rect 22200 13328 23000 13358
rect 4409 12944 4729 12945
rect 4409 12880 4417 12944
rect 4481 12880 4497 12944
rect 4561 12880 4577 12944
rect 4641 12880 4657 12944
rect 4721 12880 4729 12944
rect 4409 12879 4729 12880
rect 11340 12944 11660 12945
rect 11340 12880 11348 12944
rect 11412 12880 11428 12944
rect 11492 12880 11508 12944
rect 11572 12880 11588 12944
rect 11652 12880 11660 12944
rect 11340 12879 11660 12880
rect 18270 12944 18590 12945
rect 18270 12880 18278 12944
rect 18342 12880 18358 12944
rect 18422 12880 18438 12944
rect 18502 12880 18518 12944
rect 18582 12880 18590 12944
rect 18270 12879 18590 12880
rect 20253 12874 20319 12877
rect 22200 12874 23000 12904
rect 20253 12872 23000 12874
rect 20253 12816 20258 12872
rect 20314 12816 23000 12872
rect 20253 12814 23000 12816
rect 20253 12811 20319 12814
rect 22200 12784 23000 12814
rect 19701 12466 19767 12469
rect 22200 12466 23000 12496
rect 19701 12464 23000 12466
rect 19701 12408 19706 12464
rect 19762 12408 23000 12464
rect 19701 12406 23000 12408
rect 19701 12403 19767 12406
rect 7874 12400 8194 12401
rect 7874 12336 7882 12400
rect 7946 12336 7962 12400
rect 8026 12336 8042 12400
rect 8106 12336 8122 12400
rect 8186 12336 8194 12400
rect 7874 12335 8194 12336
rect 14805 12400 15125 12401
rect 14805 12336 14813 12400
rect 14877 12336 14893 12400
rect 14957 12336 14973 12400
rect 15037 12336 15053 12400
rect 15117 12336 15125 12400
rect 22200 12376 23000 12406
rect 14805 12335 15125 12336
rect 20621 11922 20687 11925
rect 22200 11922 23000 11952
rect 20621 11920 23000 11922
rect 20621 11864 20626 11920
rect 20682 11864 23000 11920
rect 20621 11862 23000 11864
rect 20621 11859 20687 11862
rect 4409 11856 4729 11857
rect 4409 11792 4417 11856
rect 4481 11792 4497 11856
rect 4561 11792 4577 11856
rect 4641 11792 4657 11856
rect 4721 11792 4729 11856
rect 4409 11791 4729 11792
rect 11340 11856 11660 11857
rect 11340 11792 11348 11856
rect 11412 11792 11428 11856
rect 11492 11792 11508 11856
rect 11572 11792 11588 11856
rect 11652 11792 11660 11856
rect 11340 11791 11660 11792
rect 18270 11856 18590 11857
rect 18270 11792 18278 11856
rect 18342 11792 18358 11856
rect 18422 11792 18438 11856
rect 18502 11792 18518 11856
rect 18582 11792 18590 11856
rect 22200 11832 23000 11862
rect 18270 11791 18590 11792
rect 22001 11514 22067 11517
rect 22200 11514 23000 11544
rect 22001 11512 23000 11514
rect 22001 11456 22006 11512
rect 22062 11456 23000 11512
rect 22001 11454 23000 11456
rect 22001 11451 22067 11454
rect 22200 11424 23000 11454
rect 7874 11312 8194 11313
rect 7874 11248 7882 11312
rect 7946 11248 7962 11312
rect 8026 11248 8042 11312
rect 8106 11248 8122 11312
rect 8186 11248 8194 11312
rect 7874 11247 8194 11248
rect 14805 11312 15125 11313
rect 14805 11248 14813 11312
rect 14877 11248 14893 11312
rect 14957 11248 14973 11312
rect 15037 11248 15053 11312
rect 15117 11248 15125 11312
rect 14805 11247 15125 11248
rect 20897 11106 20963 11109
rect 22200 11106 23000 11136
rect 20897 11104 23000 11106
rect 20897 11048 20902 11104
rect 20958 11048 23000 11104
rect 20897 11046 23000 11048
rect 20897 11043 20963 11046
rect 22200 11016 23000 11046
rect 4409 10768 4729 10769
rect 4409 10704 4417 10768
rect 4481 10704 4497 10768
rect 4561 10704 4577 10768
rect 4641 10704 4657 10768
rect 4721 10704 4729 10768
rect 4409 10703 4729 10704
rect 11340 10768 11660 10769
rect 11340 10704 11348 10768
rect 11412 10704 11428 10768
rect 11492 10704 11508 10768
rect 11572 10704 11588 10768
rect 11652 10704 11660 10768
rect 11340 10703 11660 10704
rect 18270 10768 18590 10769
rect 18270 10704 18278 10768
rect 18342 10704 18358 10768
rect 18422 10704 18438 10768
rect 18502 10704 18518 10768
rect 18582 10704 18590 10768
rect 18270 10703 18590 10704
rect 20621 10562 20687 10565
rect 22200 10562 23000 10592
rect 20621 10560 23000 10562
rect 20621 10504 20626 10560
rect 20682 10504 23000 10560
rect 20621 10502 23000 10504
rect 20621 10499 20687 10502
rect 22200 10472 23000 10502
rect 7874 10224 8194 10225
rect 7874 10160 7882 10224
rect 7946 10160 7962 10224
rect 8026 10160 8042 10224
rect 8106 10160 8122 10224
rect 8186 10160 8194 10224
rect 7874 10159 8194 10160
rect 14805 10224 15125 10225
rect 14805 10160 14813 10224
rect 14877 10160 14893 10224
rect 14957 10160 14973 10224
rect 15037 10160 15053 10224
rect 15117 10160 15125 10224
rect 14805 10159 15125 10160
rect 20069 10154 20135 10157
rect 22200 10154 23000 10184
rect 20069 10152 23000 10154
rect 20069 10096 20074 10152
rect 20130 10096 23000 10152
rect 20069 10094 23000 10096
rect 20069 10091 20135 10094
rect 22200 10064 23000 10094
rect 4409 9680 4729 9681
rect 4409 9616 4417 9680
rect 4481 9616 4497 9680
rect 4561 9616 4577 9680
rect 4641 9616 4657 9680
rect 4721 9616 4729 9680
rect 4409 9615 4729 9616
rect 11340 9680 11660 9681
rect 11340 9616 11348 9680
rect 11412 9616 11428 9680
rect 11492 9616 11508 9680
rect 11572 9616 11588 9680
rect 11652 9616 11660 9680
rect 11340 9615 11660 9616
rect 18270 9680 18590 9681
rect 18270 9616 18278 9680
rect 18342 9616 18358 9680
rect 18422 9616 18438 9680
rect 18502 9616 18518 9680
rect 18582 9616 18590 9680
rect 18270 9615 18590 9616
rect 20621 9610 20687 9613
rect 22200 9610 23000 9640
rect 20621 9608 23000 9610
rect 20621 9552 20626 9608
rect 20682 9552 23000 9608
rect 20621 9550 23000 9552
rect 20621 9547 20687 9550
rect 22200 9520 23000 9550
rect 20529 9202 20595 9205
rect 22200 9202 23000 9232
rect 20529 9200 23000 9202
rect 20529 9144 20534 9200
rect 20590 9144 23000 9200
rect 20529 9142 23000 9144
rect 20529 9139 20595 9142
rect 7874 9136 8194 9137
rect 7874 9072 7882 9136
rect 7946 9072 7962 9136
rect 8026 9072 8042 9136
rect 8106 9072 8122 9136
rect 8186 9072 8194 9136
rect 7874 9071 8194 9072
rect 14805 9136 15125 9137
rect 14805 9072 14813 9136
rect 14877 9072 14893 9136
rect 14957 9072 14973 9136
rect 15037 9072 15053 9136
rect 15117 9072 15125 9136
rect 22200 9112 23000 9142
rect 14805 9071 15125 9072
rect 20897 8794 20963 8797
rect 22200 8794 23000 8824
rect 20897 8792 23000 8794
rect 20897 8736 20902 8792
rect 20958 8736 23000 8792
rect 20897 8734 23000 8736
rect 20897 8731 20963 8734
rect 22200 8704 23000 8734
rect 4409 8592 4729 8593
rect 4409 8528 4417 8592
rect 4481 8528 4497 8592
rect 4561 8528 4577 8592
rect 4641 8528 4657 8592
rect 4721 8528 4729 8592
rect 4409 8527 4729 8528
rect 11340 8592 11660 8593
rect 11340 8528 11348 8592
rect 11412 8528 11428 8592
rect 11492 8528 11508 8592
rect 11572 8528 11588 8592
rect 11652 8528 11660 8592
rect 11340 8527 11660 8528
rect 18270 8592 18590 8593
rect 18270 8528 18278 8592
rect 18342 8528 18358 8592
rect 18422 8528 18438 8592
rect 18502 8528 18518 8592
rect 18582 8528 18590 8592
rect 18270 8527 18590 8528
rect 22001 8250 22067 8253
rect 22200 8250 23000 8280
rect 22001 8248 23000 8250
rect 22001 8192 22006 8248
rect 22062 8192 23000 8248
rect 22001 8190 23000 8192
rect 22001 8187 22067 8190
rect 22200 8160 23000 8190
rect 7874 8048 8194 8049
rect 7874 7984 7882 8048
rect 7946 7984 7962 8048
rect 8026 7984 8042 8048
rect 8106 7984 8122 8048
rect 8186 7984 8194 8048
rect 7874 7983 8194 7984
rect 14805 8048 15125 8049
rect 14805 7984 14813 8048
rect 14877 7984 14893 8048
rect 14957 7984 14973 8048
rect 15037 7984 15053 8048
rect 15117 7984 15125 8048
rect 14805 7983 15125 7984
rect 20621 7842 20687 7845
rect 22200 7842 23000 7872
rect 20621 7840 23000 7842
rect 20621 7784 20626 7840
rect 20682 7784 23000 7840
rect 20621 7782 23000 7784
rect 20621 7779 20687 7782
rect 22200 7752 23000 7782
rect 4409 7504 4729 7505
rect 4409 7440 4417 7504
rect 4481 7440 4497 7504
rect 4561 7440 4577 7504
rect 4641 7440 4657 7504
rect 4721 7440 4729 7504
rect 4409 7439 4729 7440
rect 11340 7504 11660 7505
rect 11340 7440 11348 7504
rect 11412 7440 11428 7504
rect 11492 7440 11508 7504
rect 11572 7440 11588 7504
rect 11652 7440 11660 7504
rect 11340 7439 11660 7440
rect 18270 7504 18590 7505
rect 18270 7440 18278 7504
rect 18342 7440 18358 7504
rect 18422 7440 18438 7504
rect 18502 7440 18518 7504
rect 18582 7440 18590 7504
rect 18270 7439 18590 7440
rect 20805 7434 20871 7437
rect 22200 7434 23000 7464
rect 20805 7432 23000 7434
rect 20805 7376 20810 7432
rect 20866 7376 23000 7432
rect 20805 7374 23000 7376
rect 20805 7371 20871 7374
rect 22200 7344 23000 7374
rect 7874 6960 8194 6961
rect 7874 6896 7882 6960
rect 7946 6896 7962 6960
rect 8026 6896 8042 6960
rect 8106 6896 8122 6960
rect 8186 6896 8194 6960
rect 7874 6895 8194 6896
rect 14805 6960 15125 6961
rect 14805 6896 14813 6960
rect 14877 6896 14893 6960
rect 14957 6896 14973 6960
rect 15037 6896 15053 6960
rect 15117 6896 15125 6960
rect 14805 6895 15125 6896
rect 20897 6890 20963 6893
rect 22200 6890 23000 6920
rect 20897 6888 23000 6890
rect 20897 6832 20902 6888
rect 20958 6832 23000 6888
rect 20897 6830 23000 6832
rect 20897 6827 20963 6830
rect 22200 6800 23000 6830
rect 19241 6482 19307 6485
rect 22200 6482 23000 6512
rect 19241 6480 23000 6482
rect 19241 6424 19246 6480
rect 19302 6424 23000 6480
rect 19241 6422 23000 6424
rect 19241 6419 19307 6422
rect 4409 6416 4729 6417
rect 4409 6352 4417 6416
rect 4481 6352 4497 6416
rect 4561 6352 4577 6416
rect 4641 6352 4657 6416
rect 4721 6352 4729 6416
rect 4409 6351 4729 6352
rect 11340 6416 11660 6417
rect 11340 6352 11348 6416
rect 11412 6352 11428 6416
rect 11492 6352 11508 6416
rect 11572 6352 11588 6416
rect 11652 6352 11660 6416
rect 11340 6351 11660 6352
rect 18270 6416 18590 6417
rect 18270 6352 18278 6416
rect 18342 6352 18358 6416
rect 18422 6352 18438 6416
rect 18502 6352 18518 6416
rect 18582 6352 18590 6416
rect 22200 6392 23000 6422
rect 18270 6351 18590 6352
rect 21357 5938 21423 5941
rect 22200 5938 23000 5968
rect 21357 5936 23000 5938
rect 21357 5880 21362 5936
rect 21418 5880 23000 5936
rect 21357 5878 23000 5880
rect 21357 5875 21423 5878
rect 7874 5872 8194 5873
rect 7874 5808 7882 5872
rect 7946 5808 7962 5872
rect 8026 5808 8042 5872
rect 8106 5808 8122 5872
rect 8186 5808 8194 5872
rect 7874 5807 8194 5808
rect 14805 5872 15125 5873
rect 14805 5808 14813 5872
rect 14877 5808 14893 5872
rect 14957 5808 14973 5872
rect 15037 5808 15053 5872
rect 15117 5808 15125 5872
rect 22200 5848 23000 5878
rect 14805 5807 15125 5808
rect 0 5666 800 5696
rect 4061 5666 4127 5669
rect 0 5664 4127 5666
rect 0 5608 4066 5664
rect 4122 5608 4127 5664
rect 0 5606 4127 5608
rect 0 5576 800 5606
rect 4061 5603 4127 5606
rect 17953 5530 18019 5533
rect 22200 5530 23000 5560
rect 17953 5528 23000 5530
rect 17953 5472 17958 5528
rect 18014 5472 23000 5528
rect 17953 5470 23000 5472
rect 17953 5467 18019 5470
rect 22200 5440 23000 5470
rect 4409 5328 4729 5329
rect 4409 5264 4417 5328
rect 4481 5264 4497 5328
rect 4561 5264 4577 5328
rect 4641 5264 4657 5328
rect 4721 5264 4729 5328
rect 4409 5263 4729 5264
rect 11340 5328 11660 5329
rect 11340 5264 11348 5328
rect 11412 5264 11428 5328
rect 11492 5264 11508 5328
rect 11572 5264 11588 5328
rect 11652 5264 11660 5328
rect 11340 5263 11660 5264
rect 18270 5328 18590 5329
rect 18270 5264 18278 5328
rect 18342 5264 18358 5328
rect 18422 5264 18438 5328
rect 18502 5264 18518 5328
rect 18582 5264 18590 5328
rect 18270 5263 18590 5264
rect 21265 5122 21331 5125
rect 22200 5122 23000 5152
rect 21265 5120 23000 5122
rect 21265 5064 21270 5120
rect 21326 5064 23000 5120
rect 21265 5062 23000 5064
rect 21265 5059 21331 5062
rect 22200 5032 23000 5062
rect 7874 4784 8194 4785
rect 7874 4720 7882 4784
rect 7946 4720 7962 4784
rect 8026 4720 8042 4784
rect 8106 4720 8122 4784
rect 8186 4720 8194 4784
rect 7874 4719 8194 4720
rect 14805 4784 15125 4785
rect 14805 4720 14813 4784
rect 14877 4720 14893 4784
rect 14957 4720 14973 4784
rect 15037 4720 15053 4784
rect 15117 4720 15125 4784
rect 14805 4719 15125 4720
rect 17953 4578 18019 4581
rect 22200 4578 23000 4608
rect 17953 4576 23000 4578
rect 17953 4520 17958 4576
rect 18014 4520 23000 4576
rect 17953 4518 23000 4520
rect 17953 4515 18019 4518
rect 22200 4488 23000 4518
rect 4409 4240 4729 4241
rect 4409 4176 4417 4240
rect 4481 4176 4497 4240
rect 4561 4176 4577 4240
rect 4641 4176 4657 4240
rect 4721 4176 4729 4240
rect 4409 4175 4729 4176
rect 11340 4240 11660 4241
rect 11340 4176 11348 4240
rect 11412 4176 11428 4240
rect 11492 4176 11508 4240
rect 11572 4176 11588 4240
rect 11652 4176 11660 4240
rect 11340 4175 11660 4176
rect 18270 4240 18590 4241
rect 18270 4176 18278 4240
rect 18342 4176 18358 4240
rect 18422 4176 18438 4240
rect 18502 4176 18518 4240
rect 18582 4176 18590 4240
rect 18270 4175 18590 4176
rect 21265 4170 21331 4173
rect 22200 4170 23000 4200
rect 21265 4168 23000 4170
rect 21265 4112 21270 4168
rect 21326 4112 23000 4168
rect 21265 4110 23000 4112
rect 21265 4107 21331 4110
rect 22200 4080 23000 4110
rect 19149 3762 19215 3765
rect 22200 3762 23000 3792
rect 19149 3760 23000 3762
rect 19149 3704 19154 3760
rect 19210 3704 23000 3760
rect 19149 3702 23000 3704
rect 19149 3699 19215 3702
rect 7874 3696 8194 3697
rect 7874 3632 7882 3696
rect 7946 3632 7962 3696
rect 8026 3632 8042 3696
rect 8106 3632 8122 3696
rect 8186 3632 8194 3696
rect 7874 3631 8194 3632
rect 14805 3696 15125 3697
rect 14805 3632 14813 3696
rect 14877 3632 14893 3696
rect 14957 3632 14973 3696
rect 15037 3632 15053 3696
rect 15117 3632 15125 3696
rect 22200 3672 23000 3702
rect 14805 3631 15125 3632
rect 18781 3218 18847 3221
rect 22200 3218 23000 3248
rect 18781 3216 23000 3218
rect 18781 3160 18786 3216
rect 18842 3160 23000 3216
rect 18781 3158 23000 3160
rect 18781 3155 18847 3158
rect 4409 3152 4729 3153
rect 4409 3088 4417 3152
rect 4481 3088 4497 3152
rect 4561 3088 4577 3152
rect 4641 3088 4657 3152
rect 4721 3088 4729 3152
rect 4409 3087 4729 3088
rect 11340 3152 11660 3153
rect 11340 3088 11348 3152
rect 11412 3088 11428 3152
rect 11492 3088 11508 3152
rect 11572 3088 11588 3152
rect 11652 3088 11660 3152
rect 11340 3087 11660 3088
rect 18270 3152 18590 3153
rect 18270 3088 18278 3152
rect 18342 3088 18358 3152
rect 18422 3088 18438 3152
rect 18502 3088 18518 3152
rect 18582 3088 18590 3152
rect 22200 3128 23000 3158
rect 18270 3087 18590 3088
rect 19241 2810 19307 2813
rect 22200 2810 23000 2840
rect 19241 2808 23000 2810
rect 19241 2752 19246 2808
rect 19302 2752 23000 2808
rect 19241 2750 23000 2752
rect 19241 2747 19307 2750
rect 22200 2720 23000 2750
rect 7874 2608 8194 2609
rect 7874 2544 7882 2608
rect 7946 2544 7962 2608
rect 8026 2544 8042 2608
rect 8106 2544 8122 2608
rect 8186 2544 8194 2608
rect 7874 2543 8194 2544
rect 14805 2608 15125 2609
rect 14805 2544 14813 2608
rect 14877 2544 14893 2608
rect 14957 2544 14973 2608
rect 15037 2544 15053 2608
rect 15117 2544 15125 2608
rect 14805 2543 15125 2544
rect 18137 2266 18203 2269
rect 22200 2266 23000 2296
rect 18137 2264 23000 2266
rect 18137 2208 18142 2264
rect 18198 2208 23000 2264
rect 18137 2206 23000 2208
rect 18137 2203 18203 2206
rect 22200 2176 23000 2206
rect 4409 2064 4729 2065
rect 4409 2000 4417 2064
rect 4481 2000 4497 2064
rect 4561 2000 4577 2064
rect 4641 2000 4657 2064
rect 4721 2000 4729 2064
rect 4409 1999 4729 2000
rect 11340 2064 11660 2065
rect 11340 2000 11348 2064
rect 11412 2000 11428 2064
rect 11492 2000 11508 2064
rect 11572 2000 11588 2064
rect 11652 2000 11660 2064
rect 11340 1999 11660 2000
rect 18270 2064 18590 2065
rect 18270 2000 18278 2064
rect 18342 2000 18358 2064
rect 18422 2000 18438 2064
rect 18502 2000 18518 2064
rect 18582 2000 18590 2064
rect 18270 1999 18590 2000
rect 18873 1858 18939 1861
rect 22200 1858 23000 1888
rect 18873 1856 23000 1858
rect 18873 1800 18878 1856
rect 18934 1800 23000 1856
rect 18873 1798 23000 1800
rect 18873 1795 18939 1798
rect 22200 1768 23000 1798
rect 18137 1450 18203 1453
rect 22200 1450 23000 1480
rect 18137 1448 23000 1450
rect 18137 1392 18142 1448
rect 18198 1392 23000 1448
rect 18137 1390 23000 1392
rect 18137 1387 18203 1390
rect 22200 1360 23000 1390
rect 19149 906 19215 909
rect 22200 906 23000 936
rect 19149 904 23000 906
rect 19149 848 19154 904
rect 19210 848 23000 904
rect 19149 846 23000 848
rect 19149 843 19215 846
rect 22200 816 23000 846
rect 17953 498 18019 501
rect 22200 498 23000 528
rect 17953 496 23000 498
rect 17953 440 17958 496
rect 18014 440 23000 496
rect 17953 438 23000 440
rect 17953 435 18019 438
rect 22200 408 23000 438
rect 18781 90 18847 93
rect 22200 90 23000 120
rect 18781 88 23000 90
rect 18781 32 18786 88
rect 18842 32 23000 88
rect 18781 30 23000 32
rect 18781 27 18847 30
rect 22200 0 23000 30
<< via3 >>
rect 4417 20556 4481 20560
rect 4417 20500 4421 20556
rect 4421 20500 4477 20556
rect 4477 20500 4481 20556
rect 4417 20496 4481 20500
rect 4497 20556 4561 20560
rect 4497 20500 4501 20556
rect 4501 20500 4557 20556
rect 4557 20500 4561 20556
rect 4497 20496 4561 20500
rect 4577 20556 4641 20560
rect 4577 20500 4581 20556
rect 4581 20500 4637 20556
rect 4637 20500 4641 20556
rect 4577 20496 4641 20500
rect 4657 20556 4721 20560
rect 4657 20500 4661 20556
rect 4661 20500 4717 20556
rect 4717 20500 4721 20556
rect 4657 20496 4721 20500
rect 11348 20556 11412 20560
rect 11348 20500 11352 20556
rect 11352 20500 11408 20556
rect 11408 20500 11412 20556
rect 11348 20496 11412 20500
rect 11428 20556 11492 20560
rect 11428 20500 11432 20556
rect 11432 20500 11488 20556
rect 11488 20500 11492 20556
rect 11428 20496 11492 20500
rect 11508 20556 11572 20560
rect 11508 20500 11512 20556
rect 11512 20500 11568 20556
rect 11568 20500 11572 20556
rect 11508 20496 11572 20500
rect 11588 20556 11652 20560
rect 11588 20500 11592 20556
rect 11592 20500 11648 20556
rect 11648 20500 11652 20556
rect 11588 20496 11652 20500
rect 18278 20556 18342 20560
rect 18278 20500 18282 20556
rect 18282 20500 18338 20556
rect 18338 20500 18342 20556
rect 18278 20496 18342 20500
rect 18358 20556 18422 20560
rect 18358 20500 18362 20556
rect 18362 20500 18418 20556
rect 18418 20500 18422 20556
rect 18358 20496 18422 20500
rect 18438 20556 18502 20560
rect 18438 20500 18442 20556
rect 18442 20500 18498 20556
rect 18498 20500 18502 20556
rect 18438 20496 18502 20500
rect 18518 20556 18582 20560
rect 18518 20500 18522 20556
rect 18522 20500 18578 20556
rect 18578 20500 18582 20556
rect 18518 20496 18582 20500
rect 7882 20012 7946 20016
rect 7882 19956 7886 20012
rect 7886 19956 7942 20012
rect 7942 19956 7946 20012
rect 7882 19952 7946 19956
rect 7962 20012 8026 20016
rect 7962 19956 7966 20012
rect 7966 19956 8022 20012
rect 8022 19956 8026 20012
rect 7962 19952 8026 19956
rect 8042 20012 8106 20016
rect 8042 19956 8046 20012
rect 8046 19956 8102 20012
rect 8102 19956 8106 20012
rect 8042 19952 8106 19956
rect 8122 20012 8186 20016
rect 8122 19956 8126 20012
rect 8126 19956 8182 20012
rect 8182 19956 8186 20012
rect 8122 19952 8186 19956
rect 14813 20012 14877 20016
rect 14813 19956 14817 20012
rect 14817 19956 14873 20012
rect 14873 19956 14877 20012
rect 14813 19952 14877 19956
rect 14893 20012 14957 20016
rect 14893 19956 14897 20012
rect 14897 19956 14953 20012
rect 14953 19956 14957 20012
rect 14893 19952 14957 19956
rect 14973 20012 15037 20016
rect 14973 19956 14977 20012
rect 14977 19956 15033 20012
rect 15033 19956 15037 20012
rect 14973 19952 15037 19956
rect 15053 20012 15117 20016
rect 15053 19956 15057 20012
rect 15057 19956 15113 20012
rect 15113 19956 15117 20012
rect 15053 19952 15117 19956
rect 4417 19468 4481 19472
rect 4417 19412 4421 19468
rect 4421 19412 4477 19468
rect 4477 19412 4481 19468
rect 4417 19408 4481 19412
rect 4497 19468 4561 19472
rect 4497 19412 4501 19468
rect 4501 19412 4557 19468
rect 4557 19412 4561 19468
rect 4497 19408 4561 19412
rect 4577 19468 4641 19472
rect 4577 19412 4581 19468
rect 4581 19412 4637 19468
rect 4637 19412 4641 19468
rect 4577 19408 4641 19412
rect 4657 19468 4721 19472
rect 4657 19412 4661 19468
rect 4661 19412 4717 19468
rect 4717 19412 4721 19468
rect 4657 19408 4721 19412
rect 11348 19468 11412 19472
rect 11348 19412 11352 19468
rect 11352 19412 11408 19468
rect 11408 19412 11412 19468
rect 11348 19408 11412 19412
rect 11428 19468 11492 19472
rect 11428 19412 11432 19468
rect 11432 19412 11488 19468
rect 11488 19412 11492 19468
rect 11428 19408 11492 19412
rect 11508 19468 11572 19472
rect 11508 19412 11512 19468
rect 11512 19412 11568 19468
rect 11568 19412 11572 19468
rect 11508 19408 11572 19412
rect 11588 19468 11652 19472
rect 11588 19412 11592 19468
rect 11592 19412 11648 19468
rect 11648 19412 11652 19468
rect 11588 19408 11652 19412
rect 18278 19468 18342 19472
rect 18278 19412 18282 19468
rect 18282 19412 18338 19468
rect 18338 19412 18342 19468
rect 18278 19408 18342 19412
rect 18358 19468 18422 19472
rect 18358 19412 18362 19468
rect 18362 19412 18418 19468
rect 18418 19412 18422 19468
rect 18358 19408 18422 19412
rect 18438 19468 18502 19472
rect 18438 19412 18442 19468
rect 18442 19412 18498 19468
rect 18498 19412 18502 19468
rect 18438 19408 18502 19412
rect 18518 19468 18582 19472
rect 18518 19412 18522 19468
rect 18522 19412 18578 19468
rect 18578 19412 18582 19468
rect 18518 19408 18582 19412
rect 7882 18924 7946 18928
rect 7882 18868 7886 18924
rect 7886 18868 7942 18924
rect 7942 18868 7946 18924
rect 7882 18864 7946 18868
rect 7962 18924 8026 18928
rect 7962 18868 7966 18924
rect 7966 18868 8022 18924
rect 8022 18868 8026 18924
rect 7962 18864 8026 18868
rect 8042 18924 8106 18928
rect 8042 18868 8046 18924
rect 8046 18868 8102 18924
rect 8102 18868 8106 18924
rect 8042 18864 8106 18868
rect 8122 18924 8186 18928
rect 8122 18868 8126 18924
rect 8126 18868 8182 18924
rect 8182 18868 8186 18924
rect 8122 18864 8186 18868
rect 14813 18924 14877 18928
rect 14813 18868 14817 18924
rect 14817 18868 14873 18924
rect 14873 18868 14877 18924
rect 14813 18864 14877 18868
rect 14893 18924 14957 18928
rect 14893 18868 14897 18924
rect 14897 18868 14953 18924
rect 14953 18868 14957 18924
rect 14893 18864 14957 18868
rect 14973 18924 15037 18928
rect 14973 18868 14977 18924
rect 14977 18868 15033 18924
rect 15033 18868 15037 18924
rect 14973 18864 15037 18868
rect 15053 18924 15117 18928
rect 15053 18868 15057 18924
rect 15057 18868 15113 18924
rect 15113 18868 15117 18924
rect 15053 18864 15117 18868
rect 4417 18380 4481 18384
rect 4417 18324 4421 18380
rect 4421 18324 4477 18380
rect 4477 18324 4481 18380
rect 4417 18320 4481 18324
rect 4497 18380 4561 18384
rect 4497 18324 4501 18380
rect 4501 18324 4557 18380
rect 4557 18324 4561 18380
rect 4497 18320 4561 18324
rect 4577 18380 4641 18384
rect 4577 18324 4581 18380
rect 4581 18324 4637 18380
rect 4637 18324 4641 18380
rect 4577 18320 4641 18324
rect 4657 18380 4721 18384
rect 4657 18324 4661 18380
rect 4661 18324 4717 18380
rect 4717 18324 4721 18380
rect 4657 18320 4721 18324
rect 11348 18380 11412 18384
rect 11348 18324 11352 18380
rect 11352 18324 11408 18380
rect 11408 18324 11412 18380
rect 11348 18320 11412 18324
rect 11428 18380 11492 18384
rect 11428 18324 11432 18380
rect 11432 18324 11488 18380
rect 11488 18324 11492 18380
rect 11428 18320 11492 18324
rect 11508 18380 11572 18384
rect 11508 18324 11512 18380
rect 11512 18324 11568 18380
rect 11568 18324 11572 18380
rect 11508 18320 11572 18324
rect 11588 18380 11652 18384
rect 11588 18324 11592 18380
rect 11592 18324 11648 18380
rect 11648 18324 11652 18380
rect 11588 18320 11652 18324
rect 18278 18380 18342 18384
rect 18278 18324 18282 18380
rect 18282 18324 18338 18380
rect 18338 18324 18342 18380
rect 18278 18320 18342 18324
rect 18358 18380 18422 18384
rect 18358 18324 18362 18380
rect 18362 18324 18418 18380
rect 18418 18324 18422 18380
rect 18358 18320 18422 18324
rect 18438 18380 18502 18384
rect 18438 18324 18442 18380
rect 18442 18324 18498 18380
rect 18498 18324 18502 18380
rect 18438 18320 18502 18324
rect 18518 18380 18582 18384
rect 18518 18324 18522 18380
rect 18522 18324 18578 18380
rect 18578 18324 18582 18380
rect 18518 18320 18582 18324
rect 7882 17836 7946 17840
rect 7882 17780 7886 17836
rect 7886 17780 7942 17836
rect 7942 17780 7946 17836
rect 7882 17776 7946 17780
rect 7962 17836 8026 17840
rect 7962 17780 7966 17836
rect 7966 17780 8022 17836
rect 8022 17780 8026 17836
rect 7962 17776 8026 17780
rect 8042 17836 8106 17840
rect 8042 17780 8046 17836
rect 8046 17780 8102 17836
rect 8102 17780 8106 17836
rect 8042 17776 8106 17780
rect 8122 17836 8186 17840
rect 8122 17780 8126 17836
rect 8126 17780 8182 17836
rect 8182 17780 8186 17836
rect 8122 17776 8186 17780
rect 14813 17836 14877 17840
rect 14813 17780 14817 17836
rect 14817 17780 14873 17836
rect 14873 17780 14877 17836
rect 14813 17776 14877 17780
rect 14893 17836 14957 17840
rect 14893 17780 14897 17836
rect 14897 17780 14953 17836
rect 14953 17780 14957 17836
rect 14893 17776 14957 17780
rect 14973 17836 15037 17840
rect 14973 17780 14977 17836
rect 14977 17780 15033 17836
rect 15033 17780 15037 17836
rect 14973 17776 15037 17780
rect 15053 17836 15117 17840
rect 15053 17780 15057 17836
rect 15057 17780 15113 17836
rect 15113 17780 15117 17836
rect 15053 17776 15117 17780
rect 4417 17292 4481 17296
rect 4417 17236 4421 17292
rect 4421 17236 4477 17292
rect 4477 17236 4481 17292
rect 4417 17232 4481 17236
rect 4497 17292 4561 17296
rect 4497 17236 4501 17292
rect 4501 17236 4557 17292
rect 4557 17236 4561 17292
rect 4497 17232 4561 17236
rect 4577 17292 4641 17296
rect 4577 17236 4581 17292
rect 4581 17236 4637 17292
rect 4637 17236 4641 17292
rect 4577 17232 4641 17236
rect 4657 17292 4721 17296
rect 4657 17236 4661 17292
rect 4661 17236 4717 17292
rect 4717 17236 4721 17292
rect 4657 17232 4721 17236
rect 11348 17292 11412 17296
rect 11348 17236 11352 17292
rect 11352 17236 11408 17292
rect 11408 17236 11412 17292
rect 11348 17232 11412 17236
rect 11428 17292 11492 17296
rect 11428 17236 11432 17292
rect 11432 17236 11488 17292
rect 11488 17236 11492 17292
rect 11428 17232 11492 17236
rect 11508 17292 11572 17296
rect 11508 17236 11512 17292
rect 11512 17236 11568 17292
rect 11568 17236 11572 17292
rect 11508 17232 11572 17236
rect 11588 17292 11652 17296
rect 11588 17236 11592 17292
rect 11592 17236 11648 17292
rect 11648 17236 11652 17292
rect 11588 17232 11652 17236
rect 18278 17292 18342 17296
rect 18278 17236 18282 17292
rect 18282 17236 18338 17292
rect 18338 17236 18342 17292
rect 18278 17232 18342 17236
rect 18358 17292 18422 17296
rect 18358 17236 18362 17292
rect 18362 17236 18418 17292
rect 18418 17236 18422 17292
rect 18358 17232 18422 17236
rect 18438 17292 18502 17296
rect 18438 17236 18442 17292
rect 18442 17236 18498 17292
rect 18498 17236 18502 17292
rect 18438 17232 18502 17236
rect 18518 17292 18582 17296
rect 18518 17236 18522 17292
rect 18522 17236 18578 17292
rect 18578 17236 18582 17292
rect 18518 17232 18582 17236
rect 7882 16748 7946 16752
rect 7882 16692 7886 16748
rect 7886 16692 7942 16748
rect 7942 16692 7946 16748
rect 7882 16688 7946 16692
rect 7962 16748 8026 16752
rect 7962 16692 7966 16748
rect 7966 16692 8022 16748
rect 8022 16692 8026 16748
rect 7962 16688 8026 16692
rect 8042 16748 8106 16752
rect 8042 16692 8046 16748
rect 8046 16692 8102 16748
rect 8102 16692 8106 16748
rect 8042 16688 8106 16692
rect 8122 16748 8186 16752
rect 8122 16692 8126 16748
rect 8126 16692 8182 16748
rect 8182 16692 8186 16748
rect 8122 16688 8186 16692
rect 14813 16748 14877 16752
rect 14813 16692 14817 16748
rect 14817 16692 14873 16748
rect 14873 16692 14877 16748
rect 14813 16688 14877 16692
rect 14893 16748 14957 16752
rect 14893 16692 14897 16748
rect 14897 16692 14953 16748
rect 14953 16692 14957 16748
rect 14893 16688 14957 16692
rect 14973 16748 15037 16752
rect 14973 16692 14977 16748
rect 14977 16692 15033 16748
rect 15033 16692 15037 16748
rect 14973 16688 15037 16692
rect 15053 16748 15117 16752
rect 15053 16692 15057 16748
rect 15057 16692 15113 16748
rect 15113 16692 15117 16748
rect 15053 16688 15117 16692
rect 4417 16204 4481 16208
rect 4417 16148 4421 16204
rect 4421 16148 4477 16204
rect 4477 16148 4481 16204
rect 4417 16144 4481 16148
rect 4497 16204 4561 16208
rect 4497 16148 4501 16204
rect 4501 16148 4557 16204
rect 4557 16148 4561 16204
rect 4497 16144 4561 16148
rect 4577 16204 4641 16208
rect 4577 16148 4581 16204
rect 4581 16148 4637 16204
rect 4637 16148 4641 16204
rect 4577 16144 4641 16148
rect 4657 16204 4721 16208
rect 4657 16148 4661 16204
rect 4661 16148 4717 16204
rect 4717 16148 4721 16204
rect 4657 16144 4721 16148
rect 11348 16204 11412 16208
rect 11348 16148 11352 16204
rect 11352 16148 11408 16204
rect 11408 16148 11412 16204
rect 11348 16144 11412 16148
rect 11428 16204 11492 16208
rect 11428 16148 11432 16204
rect 11432 16148 11488 16204
rect 11488 16148 11492 16204
rect 11428 16144 11492 16148
rect 11508 16204 11572 16208
rect 11508 16148 11512 16204
rect 11512 16148 11568 16204
rect 11568 16148 11572 16204
rect 11508 16144 11572 16148
rect 11588 16204 11652 16208
rect 11588 16148 11592 16204
rect 11592 16148 11648 16204
rect 11648 16148 11652 16204
rect 11588 16144 11652 16148
rect 18278 16204 18342 16208
rect 18278 16148 18282 16204
rect 18282 16148 18338 16204
rect 18338 16148 18342 16204
rect 18278 16144 18342 16148
rect 18358 16204 18422 16208
rect 18358 16148 18362 16204
rect 18362 16148 18418 16204
rect 18418 16148 18422 16204
rect 18358 16144 18422 16148
rect 18438 16204 18502 16208
rect 18438 16148 18442 16204
rect 18442 16148 18498 16204
rect 18498 16148 18502 16204
rect 18438 16144 18502 16148
rect 18518 16204 18582 16208
rect 18518 16148 18522 16204
rect 18522 16148 18578 16204
rect 18578 16148 18582 16204
rect 18518 16144 18582 16148
rect 7882 15660 7946 15664
rect 7882 15604 7886 15660
rect 7886 15604 7942 15660
rect 7942 15604 7946 15660
rect 7882 15600 7946 15604
rect 7962 15660 8026 15664
rect 7962 15604 7966 15660
rect 7966 15604 8022 15660
rect 8022 15604 8026 15660
rect 7962 15600 8026 15604
rect 8042 15660 8106 15664
rect 8042 15604 8046 15660
rect 8046 15604 8102 15660
rect 8102 15604 8106 15660
rect 8042 15600 8106 15604
rect 8122 15660 8186 15664
rect 8122 15604 8126 15660
rect 8126 15604 8182 15660
rect 8182 15604 8186 15660
rect 8122 15600 8186 15604
rect 14813 15660 14877 15664
rect 14813 15604 14817 15660
rect 14817 15604 14873 15660
rect 14873 15604 14877 15660
rect 14813 15600 14877 15604
rect 14893 15660 14957 15664
rect 14893 15604 14897 15660
rect 14897 15604 14953 15660
rect 14953 15604 14957 15660
rect 14893 15600 14957 15604
rect 14973 15660 15037 15664
rect 14973 15604 14977 15660
rect 14977 15604 15033 15660
rect 15033 15604 15037 15660
rect 14973 15600 15037 15604
rect 15053 15660 15117 15664
rect 15053 15604 15057 15660
rect 15057 15604 15113 15660
rect 15113 15604 15117 15660
rect 15053 15600 15117 15604
rect 4417 15116 4481 15120
rect 4417 15060 4421 15116
rect 4421 15060 4477 15116
rect 4477 15060 4481 15116
rect 4417 15056 4481 15060
rect 4497 15116 4561 15120
rect 4497 15060 4501 15116
rect 4501 15060 4557 15116
rect 4557 15060 4561 15116
rect 4497 15056 4561 15060
rect 4577 15116 4641 15120
rect 4577 15060 4581 15116
rect 4581 15060 4637 15116
rect 4637 15060 4641 15116
rect 4577 15056 4641 15060
rect 4657 15116 4721 15120
rect 4657 15060 4661 15116
rect 4661 15060 4717 15116
rect 4717 15060 4721 15116
rect 4657 15056 4721 15060
rect 11348 15116 11412 15120
rect 11348 15060 11352 15116
rect 11352 15060 11408 15116
rect 11408 15060 11412 15116
rect 11348 15056 11412 15060
rect 11428 15116 11492 15120
rect 11428 15060 11432 15116
rect 11432 15060 11488 15116
rect 11488 15060 11492 15116
rect 11428 15056 11492 15060
rect 11508 15116 11572 15120
rect 11508 15060 11512 15116
rect 11512 15060 11568 15116
rect 11568 15060 11572 15116
rect 11508 15056 11572 15060
rect 11588 15116 11652 15120
rect 11588 15060 11592 15116
rect 11592 15060 11648 15116
rect 11648 15060 11652 15116
rect 11588 15056 11652 15060
rect 18278 15116 18342 15120
rect 18278 15060 18282 15116
rect 18282 15060 18338 15116
rect 18338 15060 18342 15116
rect 18278 15056 18342 15060
rect 18358 15116 18422 15120
rect 18358 15060 18362 15116
rect 18362 15060 18418 15116
rect 18418 15060 18422 15116
rect 18358 15056 18422 15060
rect 18438 15116 18502 15120
rect 18438 15060 18442 15116
rect 18442 15060 18498 15116
rect 18498 15060 18502 15116
rect 18438 15056 18502 15060
rect 18518 15116 18582 15120
rect 18518 15060 18522 15116
rect 18522 15060 18578 15116
rect 18578 15060 18582 15116
rect 18518 15056 18582 15060
rect 7882 14572 7946 14576
rect 7882 14516 7886 14572
rect 7886 14516 7942 14572
rect 7942 14516 7946 14572
rect 7882 14512 7946 14516
rect 7962 14572 8026 14576
rect 7962 14516 7966 14572
rect 7966 14516 8022 14572
rect 8022 14516 8026 14572
rect 7962 14512 8026 14516
rect 8042 14572 8106 14576
rect 8042 14516 8046 14572
rect 8046 14516 8102 14572
rect 8102 14516 8106 14572
rect 8042 14512 8106 14516
rect 8122 14572 8186 14576
rect 8122 14516 8126 14572
rect 8126 14516 8182 14572
rect 8182 14516 8186 14572
rect 8122 14512 8186 14516
rect 14813 14572 14877 14576
rect 14813 14516 14817 14572
rect 14817 14516 14873 14572
rect 14873 14516 14877 14572
rect 14813 14512 14877 14516
rect 14893 14572 14957 14576
rect 14893 14516 14897 14572
rect 14897 14516 14953 14572
rect 14953 14516 14957 14572
rect 14893 14512 14957 14516
rect 14973 14572 15037 14576
rect 14973 14516 14977 14572
rect 14977 14516 15033 14572
rect 15033 14516 15037 14572
rect 14973 14512 15037 14516
rect 15053 14572 15117 14576
rect 15053 14516 15057 14572
rect 15057 14516 15113 14572
rect 15113 14516 15117 14572
rect 15053 14512 15117 14516
rect 4417 14028 4481 14032
rect 4417 13972 4421 14028
rect 4421 13972 4477 14028
rect 4477 13972 4481 14028
rect 4417 13968 4481 13972
rect 4497 14028 4561 14032
rect 4497 13972 4501 14028
rect 4501 13972 4557 14028
rect 4557 13972 4561 14028
rect 4497 13968 4561 13972
rect 4577 14028 4641 14032
rect 4577 13972 4581 14028
rect 4581 13972 4637 14028
rect 4637 13972 4641 14028
rect 4577 13968 4641 13972
rect 4657 14028 4721 14032
rect 4657 13972 4661 14028
rect 4661 13972 4717 14028
rect 4717 13972 4721 14028
rect 4657 13968 4721 13972
rect 11348 14028 11412 14032
rect 11348 13972 11352 14028
rect 11352 13972 11408 14028
rect 11408 13972 11412 14028
rect 11348 13968 11412 13972
rect 11428 14028 11492 14032
rect 11428 13972 11432 14028
rect 11432 13972 11488 14028
rect 11488 13972 11492 14028
rect 11428 13968 11492 13972
rect 11508 14028 11572 14032
rect 11508 13972 11512 14028
rect 11512 13972 11568 14028
rect 11568 13972 11572 14028
rect 11508 13968 11572 13972
rect 11588 14028 11652 14032
rect 11588 13972 11592 14028
rect 11592 13972 11648 14028
rect 11648 13972 11652 14028
rect 11588 13968 11652 13972
rect 18278 14028 18342 14032
rect 18278 13972 18282 14028
rect 18282 13972 18338 14028
rect 18338 13972 18342 14028
rect 18278 13968 18342 13972
rect 18358 14028 18422 14032
rect 18358 13972 18362 14028
rect 18362 13972 18418 14028
rect 18418 13972 18422 14028
rect 18358 13968 18422 13972
rect 18438 14028 18502 14032
rect 18438 13972 18442 14028
rect 18442 13972 18498 14028
rect 18498 13972 18502 14028
rect 18438 13968 18502 13972
rect 18518 14028 18582 14032
rect 18518 13972 18522 14028
rect 18522 13972 18578 14028
rect 18578 13972 18582 14028
rect 18518 13968 18582 13972
rect 7882 13484 7946 13488
rect 7882 13428 7886 13484
rect 7886 13428 7942 13484
rect 7942 13428 7946 13484
rect 7882 13424 7946 13428
rect 7962 13484 8026 13488
rect 7962 13428 7966 13484
rect 7966 13428 8022 13484
rect 8022 13428 8026 13484
rect 7962 13424 8026 13428
rect 8042 13484 8106 13488
rect 8042 13428 8046 13484
rect 8046 13428 8102 13484
rect 8102 13428 8106 13484
rect 8042 13424 8106 13428
rect 8122 13484 8186 13488
rect 8122 13428 8126 13484
rect 8126 13428 8182 13484
rect 8182 13428 8186 13484
rect 8122 13424 8186 13428
rect 14813 13484 14877 13488
rect 14813 13428 14817 13484
rect 14817 13428 14873 13484
rect 14873 13428 14877 13484
rect 14813 13424 14877 13428
rect 14893 13484 14957 13488
rect 14893 13428 14897 13484
rect 14897 13428 14953 13484
rect 14953 13428 14957 13484
rect 14893 13424 14957 13428
rect 14973 13484 15037 13488
rect 14973 13428 14977 13484
rect 14977 13428 15033 13484
rect 15033 13428 15037 13484
rect 14973 13424 15037 13428
rect 15053 13484 15117 13488
rect 15053 13428 15057 13484
rect 15057 13428 15113 13484
rect 15113 13428 15117 13484
rect 15053 13424 15117 13428
rect 4417 12940 4481 12944
rect 4417 12884 4421 12940
rect 4421 12884 4477 12940
rect 4477 12884 4481 12940
rect 4417 12880 4481 12884
rect 4497 12940 4561 12944
rect 4497 12884 4501 12940
rect 4501 12884 4557 12940
rect 4557 12884 4561 12940
rect 4497 12880 4561 12884
rect 4577 12940 4641 12944
rect 4577 12884 4581 12940
rect 4581 12884 4637 12940
rect 4637 12884 4641 12940
rect 4577 12880 4641 12884
rect 4657 12940 4721 12944
rect 4657 12884 4661 12940
rect 4661 12884 4717 12940
rect 4717 12884 4721 12940
rect 4657 12880 4721 12884
rect 11348 12940 11412 12944
rect 11348 12884 11352 12940
rect 11352 12884 11408 12940
rect 11408 12884 11412 12940
rect 11348 12880 11412 12884
rect 11428 12940 11492 12944
rect 11428 12884 11432 12940
rect 11432 12884 11488 12940
rect 11488 12884 11492 12940
rect 11428 12880 11492 12884
rect 11508 12940 11572 12944
rect 11508 12884 11512 12940
rect 11512 12884 11568 12940
rect 11568 12884 11572 12940
rect 11508 12880 11572 12884
rect 11588 12940 11652 12944
rect 11588 12884 11592 12940
rect 11592 12884 11648 12940
rect 11648 12884 11652 12940
rect 11588 12880 11652 12884
rect 18278 12940 18342 12944
rect 18278 12884 18282 12940
rect 18282 12884 18338 12940
rect 18338 12884 18342 12940
rect 18278 12880 18342 12884
rect 18358 12940 18422 12944
rect 18358 12884 18362 12940
rect 18362 12884 18418 12940
rect 18418 12884 18422 12940
rect 18358 12880 18422 12884
rect 18438 12940 18502 12944
rect 18438 12884 18442 12940
rect 18442 12884 18498 12940
rect 18498 12884 18502 12940
rect 18438 12880 18502 12884
rect 18518 12940 18582 12944
rect 18518 12884 18522 12940
rect 18522 12884 18578 12940
rect 18578 12884 18582 12940
rect 18518 12880 18582 12884
rect 7882 12396 7946 12400
rect 7882 12340 7886 12396
rect 7886 12340 7942 12396
rect 7942 12340 7946 12396
rect 7882 12336 7946 12340
rect 7962 12396 8026 12400
rect 7962 12340 7966 12396
rect 7966 12340 8022 12396
rect 8022 12340 8026 12396
rect 7962 12336 8026 12340
rect 8042 12396 8106 12400
rect 8042 12340 8046 12396
rect 8046 12340 8102 12396
rect 8102 12340 8106 12396
rect 8042 12336 8106 12340
rect 8122 12396 8186 12400
rect 8122 12340 8126 12396
rect 8126 12340 8182 12396
rect 8182 12340 8186 12396
rect 8122 12336 8186 12340
rect 14813 12396 14877 12400
rect 14813 12340 14817 12396
rect 14817 12340 14873 12396
rect 14873 12340 14877 12396
rect 14813 12336 14877 12340
rect 14893 12396 14957 12400
rect 14893 12340 14897 12396
rect 14897 12340 14953 12396
rect 14953 12340 14957 12396
rect 14893 12336 14957 12340
rect 14973 12396 15037 12400
rect 14973 12340 14977 12396
rect 14977 12340 15033 12396
rect 15033 12340 15037 12396
rect 14973 12336 15037 12340
rect 15053 12396 15117 12400
rect 15053 12340 15057 12396
rect 15057 12340 15113 12396
rect 15113 12340 15117 12396
rect 15053 12336 15117 12340
rect 4417 11852 4481 11856
rect 4417 11796 4421 11852
rect 4421 11796 4477 11852
rect 4477 11796 4481 11852
rect 4417 11792 4481 11796
rect 4497 11852 4561 11856
rect 4497 11796 4501 11852
rect 4501 11796 4557 11852
rect 4557 11796 4561 11852
rect 4497 11792 4561 11796
rect 4577 11852 4641 11856
rect 4577 11796 4581 11852
rect 4581 11796 4637 11852
rect 4637 11796 4641 11852
rect 4577 11792 4641 11796
rect 4657 11852 4721 11856
rect 4657 11796 4661 11852
rect 4661 11796 4717 11852
rect 4717 11796 4721 11852
rect 4657 11792 4721 11796
rect 11348 11852 11412 11856
rect 11348 11796 11352 11852
rect 11352 11796 11408 11852
rect 11408 11796 11412 11852
rect 11348 11792 11412 11796
rect 11428 11852 11492 11856
rect 11428 11796 11432 11852
rect 11432 11796 11488 11852
rect 11488 11796 11492 11852
rect 11428 11792 11492 11796
rect 11508 11852 11572 11856
rect 11508 11796 11512 11852
rect 11512 11796 11568 11852
rect 11568 11796 11572 11852
rect 11508 11792 11572 11796
rect 11588 11852 11652 11856
rect 11588 11796 11592 11852
rect 11592 11796 11648 11852
rect 11648 11796 11652 11852
rect 11588 11792 11652 11796
rect 18278 11852 18342 11856
rect 18278 11796 18282 11852
rect 18282 11796 18338 11852
rect 18338 11796 18342 11852
rect 18278 11792 18342 11796
rect 18358 11852 18422 11856
rect 18358 11796 18362 11852
rect 18362 11796 18418 11852
rect 18418 11796 18422 11852
rect 18358 11792 18422 11796
rect 18438 11852 18502 11856
rect 18438 11796 18442 11852
rect 18442 11796 18498 11852
rect 18498 11796 18502 11852
rect 18438 11792 18502 11796
rect 18518 11852 18582 11856
rect 18518 11796 18522 11852
rect 18522 11796 18578 11852
rect 18578 11796 18582 11852
rect 18518 11792 18582 11796
rect 7882 11308 7946 11312
rect 7882 11252 7886 11308
rect 7886 11252 7942 11308
rect 7942 11252 7946 11308
rect 7882 11248 7946 11252
rect 7962 11308 8026 11312
rect 7962 11252 7966 11308
rect 7966 11252 8022 11308
rect 8022 11252 8026 11308
rect 7962 11248 8026 11252
rect 8042 11308 8106 11312
rect 8042 11252 8046 11308
rect 8046 11252 8102 11308
rect 8102 11252 8106 11308
rect 8042 11248 8106 11252
rect 8122 11308 8186 11312
rect 8122 11252 8126 11308
rect 8126 11252 8182 11308
rect 8182 11252 8186 11308
rect 8122 11248 8186 11252
rect 14813 11308 14877 11312
rect 14813 11252 14817 11308
rect 14817 11252 14873 11308
rect 14873 11252 14877 11308
rect 14813 11248 14877 11252
rect 14893 11308 14957 11312
rect 14893 11252 14897 11308
rect 14897 11252 14953 11308
rect 14953 11252 14957 11308
rect 14893 11248 14957 11252
rect 14973 11308 15037 11312
rect 14973 11252 14977 11308
rect 14977 11252 15033 11308
rect 15033 11252 15037 11308
rect 14973 11248 15037 11252
rect 15053 11308 15117 11312
rect 15053 11252 15057 11308
rect 15057 11252 15113 11308
rect 15113 11252 15117 11308
rect 15053 11248 15117 11252
rect 4417 10764 4481 10768
rect 4417 10708 4421 10764
rect 4421 10708 4477 10764
rect 4477 10708 4481 10764
rect 4417 10704 4481 10708
rect 4497 10764 4561 10768
rect 4497 10708 4501 10764
rect 4501 10708 4557 10764
rect 4557 10708 4561 10764
rect 4497 10704 4561 10708
rect 4577 10764 4641 10768
rect 4577 10708 4581 10764
rect 4581 10708 4637 10764
rect 4637 10708 4641 10764
rect 4577 10704 4641 10708
rect 4657 10764 4721 10768
rect 4657 10708 4661 10764
rect 4661 10708 4717 10764
rect 4717 10708 4721 10764
rect 4657 10704 4721 10708
rect 11348 10764 11412 10768
rect 11348 10708 11352 10764
rect 11352 10708 11408 10764
rect 11408 10708 11412 10764
rect 11348 10704 11412 10708
rect 11428 10764 11492 10768
rect 11428 10708 11432 10764
rect 11432 10708 11488 10764
rect 11488 10708 11492 10764
rect 11428 10704 11492 10708
rect 11508 10764 11572 10768
rect 11508 10708 11512 10764
rect 11512 10708 11568 10764
rect 11568 10708 11572 10764
rect 11508 10704 11572 10708
rect 11588 10764 11652 10768
rect 11588 10708 11592 10764
rect 11592 10708 11648 10764
rect 11648 10708 11652 10764
rect 11588 10704 11652 10708
rect 18278 10764 18342 10768
rect 18278 10708 18282 10764
rect 18282 10708 18338 10764
rect 18338 10708 18342 10764
rect 18278 10704 18342 10708
rect 18358 10764 18422 10768
rect 18358 10708 18362 10764
rect 18362 10708 18418 10764
rect 18418 10708 18422 10764
rect 18358 10704 18422 10708
rect 18438 10764 18502 10768
rect 18438 10708 18442 10764
rect 18442 10708 18498 10764
rect 18498 10708 18502 10764
rect 18438 10704 18502 10708
rect 18518 10764 18582 10768
rect 18518 10708 18522 10764
rect 18522 10708 18578 10764
rect 18578 10708 18582 10764
rect 18518 10704 18582 10708
rect 7882 10220 7946 10224
rect 7882 10164 7886 10220
rect 7886 10164 7942 10220
rect 7942 10164 7946 10220
rect 7882 10160 7946 10164
rect 7962 10220 8026 10224
rect 7962 10164 7966 10220
rect 7966 10164 8022 10220
rect 8022 10164 8026 10220
rect 7962 10160 8026 10164
rect 8042 10220 8106 10224
rect 8042 10164 8046 10220
rect 8046 10164 8102 10220
rect 8102 10164 8106 10220
rect 8042 10160 8106 10164
rect 8122 10220 8186 10224
rect 8122 10164 8126 10220
rect 8126 10164 8182 10220
rect 8182 10164 8186 10220
rect 8122 10160 8186 10164
rect 14813 10220 14877 10224
rect 14813 10164 14817 10220
rect 14817 10164 14873 10220
rect 14873 10164 14877 10220
rect 14813 10160 14877 10164
rect 14893 10220 14957 10224
rect 14893 10164 14897 10220
rect 14897 10164 14953 10220
rect 14953 10164 14957 10220
rect 14893 10160 14957 10164
rect 14973 10220 15037 10224
rect 14973 10164 14977 10220
rect 14977 10164 15033 10220
rect 15033 10164 15037 10220
rect 14973 10160 15037 10164
rect 15053 10220 15117 10224
rect 15053 10164 15057 10220
rect 15057 10164 15113 10220
rect 15113 10164 15117 10220
rect 15053 10160 15117 10164
rect 4417 9676 4481 9680
rect 4417 9620 4421 9676
rect 4421 9620 4477 9676
rect 4477 9620 4481 9676
rect 4417 9616 4481 9620
rect 4497 9676 4561 9680
rect 4497 9620 4501 9676
rect 4501 9620 4557 9676
rect 4557 9620 4561 9676
rect 4497 9616 4561 9620
rect 4577 9676 4641 9680
rect 4577 9620 4581 9676
rect 4581 9620 4637 9676
rect 4637 9620 4641 9676
rect 4577 9616 4641 9620
rect 4657 9676 4721 9680
rect 4657 9620 4661 9676
rect 4661 9620 4717 9676
rect 4717 9620 4721 9676
rect 4657 9616 4721 9620
rect 11348 9676 11412 9680
rect 11348 9620 11352 9676
rect 11352 9620 11408 9676
rect 11408 9620 11412 9676
rect 11348 9616 11412 9620
rect 11428 9676 11492 9680
rect 11428 9620 11432 9676
rect 11432 9620 11488 9676
rect 11488 9620 11492 9676
rect 11428 9616 11492 9620
rect 11508 9676 11572 9680
rect 11508 9620 11512 9676
rect 11512 9620 11568 9676
rect 11568 9620 11572 9676
rect 11508 9616 11572 9620
rect 11588 9676 11652 9680
rect 11588 9620 11592 9676
rect 11592 9620 11648 9676
rect 11648 9620 11652 9676
rect 11588 9616 11652 9620
rect 18278 9676 18342 9680
rect 18278 9620 18282 9676
rect 18282 9620 18338 9676
rect 18338 9620 18342 9676
rect 18278 9616 18342 9620
rect 18358 9676 18422 9680
rect 18358 9620 18362 9676
rect 18362 9620 18418 9676
rect 18418 9620 18422 9676
rect 18358 9616 18422 9620
rect 18438 9676 18502 9680
rect 18438 9620 18442 9676
rect 18442 9620 18498 9676
rect 18498 9620 18502 9676
rect 18438 9616 18502 9620
rect 18518 9676 18582 9680
rect 18518 9620 18522 9676
rect 18522 9620 18578 9676
rect 18578 9620 18582 9676
rect 18518 9616 18582 9620
rect 7882 9132 7946 9136
rect 7882 9076 7886 9132
rect 7886 9076 7942 9132
rect 7942 9076 7946 9132
rect 7882 9072 7946 9076
rect 7962 9132 8026 9136
rect 7962 9076 7966 9132
rect 7966 9076 8022 9132
rect 8022 9076 8026 9132
rect 7962 9072 8026 9076
rect 8042 9132 8106 9136
rect 8042 9076 8046 9132
rect 8046 9076 8102 9132
rect 8102 9076 8106 9132
rect 8042 9072 8106 9076
rect 8122 9132 8186 9136
rect 8122 9076 8126 9132
rect 8126 9076 8182 9132
rect 8182 9076 8186 9132
rect 8122 9072 8186 9076
rect 14813 9132 14877 9136
rect 14813 9076 14817 9132
rect 14817 9076 14873 9132
rect 14873 9076 14877 9132
rect 14813 9072 14877 9076
rect 14893 9132 14957 9136
rect 14893 9076 14897 9132
rect 14897 9076 14953 9132
rect 14953 9076 14957 9132
rect 14893 9072 14957 9076
rect 14973 9132 15037 9136
rect 14973 9076 14977 9132
rect 14977 9076 15033 9132
rect 15033 9076 15037 9132
rect 14973 9072 15037 9076
rect 15053 9132 15117 9136
rect 15053 9076 15057 9132
rect 15057 9076 15113 9132
rect 15113 9076 15117 9132
rect 15053 9072 15117 9076
rect 4417 8588 4481 8592
rect 4417 8532 4421 8588
rect 4421 8532 4477 8588
rect 4477 8532 4481 8588
rect 4417 8528 4481 8532
rect 4497 8588 4561 8592
rect 4497 8532 4501 8588
rect 4501 8532 4557 8588
rect 4557 8532 4561 8588
rect 4497 8528 4561 8532
rect 4577 8588 4641 8592
rect 4577 8532 4581 8588
rect 4581 8532 4637 8588
rect 4637 8532 4641 8588
rect 4577 8528 4641 8532
rect 4657 8588 4721 8592
rect 4657 8532 4661 8588
rect 4661 8532 4717 8588
rect 4717 8532 4721 8588
rect 4657 8528 4721 8532
rect 11348 8588 11412 8592
rect 11348 8532 11352 8588
rect 11352 8532 11408 8588
rect 11408 8532 11412 8588
rect 11348 8528 11412 8532
rect 11428 8588 11492 8592
rect 11428 8532 11432 8588
rect 11432 8532 11488 8588
rect 11488 8532 11492 8588
rect 11428 8528 11492 8532
rect 11508 8588 11572 8592
rect 11508 8532 11512 8588
rect 11512 8532 11568 8588
rect 11568 8532 11572 8588
rect 11508 8528 11572 8532
rect 11588 8588 11652 8592
rect 11588 8532 11592 8588
rect 11592 8532 11648 8588
rect 11648 8532 11652 8588
rect 11588 8528 11652 8532
rect 18278 8588 18342 8592
rect 18278 8532 18282 8588
rect 18282 8532 18338 8588
rect 18338 8532 18342 8588
rect 18278 8528 18342 8532
rect 18358 8588 18422 8592
rect 18358 8532 18362 8588
rect 18362 8532 18418 8588
rect 18418 8532 18422 8588
rect 18358 8528 18422 8532
rect 18438 8588 18502 8592
rect 18438 8532 18442 8588
rect 18442 8532 18498 8588
rect 18498 8532 18502 8588
rect 18438 8528 18502 8532
rect 18518 8588 18582 8592
rect 18518 8532 18522 8588
rect 18522 8532 18578 8588
rect 18578 8532 18582 8588
rect 18518 8528 18582 8532
rect 7882 8044 7946 8048
rect 7882 7988 7886 8044
rect 7886 7988 7942 8044
rect 7942 7988 7946 8044
rect 7882 7984 7946 7988
rect 7962 8044 8026 8048
rect 7962 7988 7966 8044
rect 7966 7988 8022 8044
rect 8022 7988 8026 8044
rect 7962 7984 8026 7988
rect 8042 8044 8106 8048
rect 8042 7988 8046 8044
rect 8046 7988 8102 8044
rect 8102 7988 8106 8044
rect 8042 7984 8106 7988
rect 8122 8044 8186 8048
rect 8122 7988 8126 8044
rect 8126 7988 8182 8044
rect 8182 7988 8186 8044
rect 8122 7984 8186 7988
rect 14813 8044 14877 8048
rect 14813 7988 14817 8044
rect 14817 7988 14873 8044
rect 14873 7988 14877 8044
rect 14813 7984 14877 7988
rect 14893 8044 14957 8048
rect 14893 7988 14897 8044
rect 14897 7988 14953 8044
rect 14953 7988 14957 8044
rect 14893 7984 14957 7988
rect 14973 8044 15037 8048
rect 14973 7988 14977 8044
rect 14977 7988 15033 8044
rect 15033 7988 15037 8044
rect 14973 7984 15037 7988
rect 15053 8044 15117 8048
rect 15053 7988 15057 8044
rect 15057 7988 15113 8044
rect 15113 7988 15117 8044
rect 15053 7984 15117 7988
rect 4417 7500 4481 7504
rect 4417 7444 4421 7500
rect 4421 7444 4477 7500
rect 4477 7444 4481 7500
rect 4417 7440 4481 7444
rect 4497 7500 4561 7504
rect 4497 7444 4501 7500
rect 4501 7444 4557 7500
rect 4557 7444 4561 7500
rect 4497 7440 4561 7444
rect 4577 7500 4641 7504
rect 4577 7444 4581 7500
rect 4581 7444 4637 7500
rect 4637 7444 4641 7500
rect 4577 7440 4641 7444
rect 4657 7500 4721 7504
rect 4657 7444 4661 7500
rect 4661 7444 4717 7500
rect 4717 7444 4721 7500
rect 4657 7440 4721 7444
rect 11348 7500 11412 7504
rect 11348 7444 11352 7500
rect 11352 7444 11408 7500
rect 11408 7444 11412 7500
rect 11348 7440 11412 7444
rect 11428 7500 11492 7504
rect 11428 7444 11432 7500
rect 11432 7444 11488 7500
rect 11488 7444 11492 7500
rect 11428 7440 11492 7444
rect 11508 7500 11572 7504
rect 11508 7444 11512 7500
rect 11512 7444 11568 7500
rect 11568 7444 11572 7500
rect 11508 7440 11572 7444
rect 11588 7500 11652 7504
rect 11588 7444 11592 7500
rect 11592 7444 11648 7500
rect 11648 7444 11652 7500
rect 11588 7440 11652 7444
rect 18278 7500 18342 7504
rect 18278 7444 18282 7500
rect 18282 7444 18338 7500
rect 18338 7444 18342 7500
rect 18278 7440 18342 7444
rect 18358 7500 18422 7504
rect 18358 7444 18362 7500
rect 18362 7444 18418 7500
rect 18418 7444 18422 7500
rect 18358 7440 18422 7444
rect 18438 7500 18502 7504
rect 18438 7444 18442 7500
rect 18442 7444 18498 7500
rect 18498 7444 18502 7500
rect 18438 7440 18502 7444
rect 18518 7500 18582 7504
rect 18518 7444 18522 7500
rect 18522 7444 18578 7500
rect 18578 7444 18582 7500
rect 18518 7440 18582 7444
rect 7882 6956 7946 6960
rect 7882 6900 7886 6956
rect 7886 6900 7942 6956
rect 7942 6900 7946 6956
rect 7882 6896 7946 6900
rect 7962 6956 8026 6960
rect 7962 6900 7966 6956
rect 7966 6900 8022 6956
rect 8022 6900 8026 6956
rect 7962 6896 8026 6900
rect 8042 6956 8106 6960
rect 8042 6900 8046 6956
rect 8046 6900 8102 6956
rect 8102 6900 8106 6956
rect 8042 6896 8106 6900
rect 8122 6956 8186 6960
rect 8122 6900 8126 6956
rect 8126 6900 8182 6956
rect 8182 6900 8186 6956
rect 8122 6896 8186 6900
rect 14813 6956 14877 6960
rect 14813 6900 14817 6956
rect 14817 6900 14873 6956
rect 14873 6900 14877 6956
rect 14813 6896 14877 6900
rect 14893 6956 14957 6960
rect 14893 6900 14897 6956
rect 14897 6900 14953 6956
rect 14953 6900 14957 6956
rect 14893 6896 14957 6900
rect 14973 6956 15037 6960
rect 14973 6900 14977 6956
rect 14977 6900 15033 6956
rect 15033 6900 15037 6956
rect 14973 6896 15037 6900
rect 15053 6956 15117 6960
rect 15053 6900 15057 6956
rect 15057 6900 15113 6956
rect 15113 6900 15117 6956
rect 15053 6896 15117 6900
rect 4417 6412 4481 6416
rect 4417 6356 4421 6412
rect 4421 6356 4477 6412
rect 4477 6356 4481 6412
rect 4417 6352 4481 6356
rect 4497 6412 4561 6416
rect 4497 6356 4501 6412
rect 4501 6356 4557 6412
rect 4557 6356 4561 6412
rect 4497 6352 4561 6356
rect 4577 6412 4641 6416
rect 4577 6356 4581 6412
rect 4581 6356 4637 6412
rect 4637 6356 4641 6412
rect 4577 6352 4641 6356
rect 4657 6412 4721 6416
rect 4657 6356 4661 6412
rect 4661 6356 4717 6412
rect 4717 6356 4721 6412
rect 4657 6352 4721 6356
rect 11348 6412 11412 6416
rect 11348 6356 11352 6412
rect 11352 6356 11408 6412
rect 11408 6356 11412 6412
rect 11348 6352 11412 6356
rect 11428 6412 11492 6416
rect 11428 6356 11432 6412
rect 11432 6356 11488 6412
rect 11488 6356 11492 6412
rect 11428 6352 11492 6356
rect 11508 6412 11572 6416
rect 11508 6356 11512 6412
rect 11512 6356 11568 6412
rect 11568 6356 11572 6412
rect 11508 6352 11572 6356
rect 11588 6412 11652 6416
rect 11588 6356 11592 6412
rect 11592 6356 11648 6412
rect 11648 6356 11652 6412
rect 11588 6352 11652 6356
rect 18278 6412 18342 6416
rect 18278 6356 18282 6412
rect 18282 6356 18338 6412
rect 18338 6356 18342 6412
rect 18278 6352 18342 6356
rect 18358 6412 18422 6416
rect 18358 6356 18362 6412
rect 18362 6356 18418 6412
rect 18418 6356 18422 6412
rect 18358 6352 18422 6356
rect 18438 6412 18502 6416
rect 18438 6356 18442 6412
rect 18442 6356 18498 6412
rect 18498 6356 18502 6412
rect 18438 6352 18502 6356
rect 18518 6412 18582 6416
rect 18518 6356 18522 6412
rect 18522 6356 18578 6412
rect 18578 6356 18582 6412
rect 18518 6352 18582 6356
rect 7882 5868 7946 5872
rect 7882 5812 7886 5868
rect 7886 5812 7942 5868
rect 7942 5812 7946 5868
rect 7882 5808 7946 5812
rect 7962 5868 8026 5872
rect 7962 5812 7966 5868
rect 7966 5812 8022 5868
rect 8022 5812 8026 5868
rect 7962 5808 8026 5812
rect 8042 5868 8106 5872
rect 8042 5812 8046 5868
rect 8046 5812 8102 5868
rect 8102 5812 8106 5868
rect 8042 5808 8106 5812
rect 8122 5868 8186 5872
rect 8122 5812 8126 5868
rect 8126 5812 8182 5868
rect 8182 5812 8186 5868
rect 8122 5808 8186 5812
rect 14813 5868 14877 5872
rect 14813 5812 14817 5868
rect 14817 5812 14873 5868
rect 14873 5812 14877 5868
rect 14813 5808 14877 5812
rect 14893 5868 14957 5872
rect 14893 5812 14897 5868
rect 14897 5812 14953 5868
rect 14953 5812 14957 5868
rect 14893 5808 14957 5812
rect 14973 5868 15037 5872
rect 14973 5812 14977 5868
rect 14977 5812 15033 5868
rect 15033 5812 15037 5868
rect 14973 5808 15037 5812
rect 15053 5868 15117 5872
rect 15053 5812 15057 5868
rect 15057 5812 15113 5868
rect 15113 5812 15117 5868
rect 15053 5808 15117 5812
rect 4417 5324 4481 5328
rect 4417 5268 4421 5324
rect 4421 5268 4477 5324
rect 4477 5268 4481 5324
rect 4417 5264 4481 5268
rect 4497 5324 4561 5328
rect 4497 5268 4501 5324
rect 4501 5268 4557 5324
rect 4557 5268 4561 5324
rect 4497 5264 4561 5268
rect 4577 5324 4641 5328
rect 4577 5268 4581 5324
rect 4581 5268 4637 5324
rect 4637 5268 4641 5324
rect 4577 5264 4641 5268
rect 4657 5324 4721 5328
rect 4657 5268 4661 5324
rect 4661 5268 4717 5324
rect 4717 5268 4721 5324
rect 4657 5264 4721 5268
rect 11348 5324 11412 5328
rect 11348 5268 11352 5324
rect 11352 5268 11408 5324
rect 11408 5268 11412 5324
rect 11348 5264 11412 5268
rect 11428 5324 11492 5328
rect 11428 5268 11432 5324
rect 11432 5268 11488 5324
rect 11488 5268 11492 5324
rect 11428 5264 11492 5268
rect 11508 5324 11572 5328
rect 11508 5268 11512 5324
rect 11512 5268 11568 5324
rect 11568 5268 11572 5324
rect 11508 5264 11572 5268
rect 11588 5324 11652 5328
rect 11588 5268 11592 5324
rect 11592 5268 11648 5324
rect 11648 5268 11652 5324
rect 11588 5264 11652 5268
rect 18278 5324 18342 5328
rect 18278 5268 18282 5324
rect 18282 5268 18338 5324
rect 18338 5268 18342 5324
rect 18278 5264 18342 5268
rect 18358 5324 18422 5328
rect 18358 5268 18362 5324
rect 18362 5268 18418 5324
rect 18418 5268 18422 5324
rect 18358 5264 18422 5268
rect 18438 5324 18502 5328
rect 18438 5268 18442 5324
rect 18442 5268 18498 5324
rect 18498 5268 18502 5324
rect 18438 5264 18502 5268
rect 18518 5324 18582 5328
rect 18518 5268 18522 5324
rect 18522 5268 18578 5324
rect 18578 5268 18582 5324
rect 18518 5264 18582 5268
rect 7882 4780 7946 4784
rect 7882 4724 7886 4780
rect 7886 4724 7942 4780
rect 7942 4724 7946 4780
rect 7882 4720 7946 4724
rect 7962 4780 8026 4784
rect 7962 4724 7966 4780
rect 7966 4724 8022 4780
rect 8022 4724 8026 4780
rect 7962 4720 8026 4724
rect 8042 4780 8106 4784
rect 8042 4724 8046 4780
rect 8046 4724 8102 4780
rect 8102 4724 8106 4780
rect 8042 4720 8106 4724
rect 8122 4780 8186 4784
rect 8122 4724 8126 4780
rect 8126 4724 8182 4780
rect 8182 4724 8186 4780
rect 8122 4720 8186 4724
rect 14813 4780 14877 4784
rect 14813 4724 14817 4780
rect 14817 4724 14873 4780
rect 14873 4724 14877 4780
rect 14813 4720 14877 4724
rect 14893 4780 14957 4784
rect 14893 4724 14897 4780
rect 14897 4724 14953 4780
rect 14953 4724 14957 4780
rect 14893 4720 14957 4724
rect 14973 4780 15037 4784
rect 14973 4724 14977 4780
rect 14977 4724 15033 4780
rect 15033 4724 15037 4780
rect 14973 4720 15037 4724
rect 15053 4780 15117 4784
rect 15053 4724 15057 4780
rect 15057 4724 15113 4780
rect 15113 4724 15117 4780
rect 15053 4720 15117 4724
rect 4417 4236 4481 4240
rect 4417 4180 4421 4236
rect 4421 4180 4477 4236
rect 4477 4180 4481 4236
rect 4417 4176 4481 4180
rect 4497 4236 4561 4240
rect 4497 4180 4501 4236
rect 4501 4180 4557 4236
rect 4557 4180 4561 4236
rect 4497 4176 4561 4180
rect 4577 4236 4641 4240
rect 4577 4180 4581 4236
rect 4581 4180 4637 4236
rect 4637 4180 4641 4236
rect 4577 4176 4641 4180
rect 4657 4236 4721 4240
rect 4657 4180 4661 4236
rect 4661 4180 4717 4236
rect 4717 4180 4721 4236
rect 4657 4176 4721 4180
rect 11348 4236 11412 4240
rect 11348 4180 11352 4236
rect 11352 4180 11408 4236
rect 11408 4180 11412 4236
rect 11348 4176 11412 4180
rect 11428 4236 11492 4240
rect 11428 4180 11432 4236
rect 11432 4180 11488 4236
rect 11488 4180 11492 4236
rect 11428 4176 11492 4180
rect 11508 4236 11572 4240
rect 11508 4180 11512 4236
rect 11512 4180 11568 4236
rect 11568 4180 11572 4236
rect 11508 4176 11572 4180
rect 11588 4236 11652 4240
rect 11588 4180 11592 4236
rect 11592 4180 11648 4236
rect 11648 4180 11652 4236
rect 11588 4176 11652 4180
rect 18278 4236 18342 4240
rect 18278 4180 18282 4236
rect 18282 4180 18338 4236
rect 18338 4180 18342 4236
rect 18278 4176 18342 4180
rect 18358 4236 18422 4240
rect 18358 4180 18362 4236
rect 18362 4180 18418 4236
rect 18418 4180 18422 4236
rect 18358 4176 18422 4180
rect 18438 4236 18502 4240
rect 18438 4180 18442 4236
rect 18442 4180 18498 4236
rect 18498 4180 18502 4236
rect 18438 4176 18502 4180
rect 18518 4236 18582 4240
rect 18518 4180 18522 4236
rect 18522 4180 18578 4236
rect 18578 4180 18582 4236
rect 18518 4176 18582 4180
rect 7882 3692 7946 3696
rect 7882 3636 7886 3692
rect 7886 3636 7942 3692
rect 7942 3636 7946 3692
rect 7882 3632 7946 3636
rect 7962 3692 8026 3696
rect 7962 3636 7966 3692
rect 7966 3636 8022 3692
rect 8022 3636 8026 3692
rect 7962 3632 8026 3636
rect 8042 3692 8106 3696
rect 8042 3636 8046 3692
rect 8046 3636 8102 3692
rect 8102 3636 8106 3692
rect 8042 3632 8106 3636
rect 8122 3692 8186 3696
rect 8122 3636 8126 3692
rect 8126 3636 8182 3692
rect 8182 3636 8186 3692
rect 8122 3632 8186 3636
rect 14813 3692 14877 3696
rect 14813 3636 14817 3692
rect 14817 3636 14873 3692
rect 14873 3636 14877 3692
rect 14813 3632 14877 3636
rect 14893 3692 14957 3696
rect 14893 3636 14897 3692
rect 14897 3636 14953 3692
rect 14953 3636 14957 3692
rect 14893 3632 14957 3636
rect 14973 3692 15037 3696
rect 14973 3636 14977 3692
rect 14977 3636 15033 3692
rect 15033 3636 15037 3692
rect 14973 3632 15037 3636
rect 15053 3692 15117 3696
rect 15053 3636 15057 3692
rect 15057 3636 15113 3692
rect 15113 3636 15117 3692
rect 15053 3632 15117 3636
rect 4417 3148 4481 3152
rect 4417 3092 4421 3148
rect 4421 3092 4477 3148
rect 4477 3092 4481 3148
rect 4417 3088 4481 3092
rect 4497 3148 4561 3152
rect 4497 3092 4501 3148
rect 4501 3092 4557 3148
rect 4557 3092 4561 3148
rect 4497 3088 4561 3092
rect 4577 3148 4641 3152
rect 4577 3092 4581 3148
rect 4581 3092 4637 3148
rect 4637 3092 4641 3148
rect 4577 3088 4641 3092
rect 4657 3148 4721 3152
rect 4657 3092 4661 3148
rect 4661 3092 4717 3148
rect 4717 3092 4721 3148
rect 4657 3088 4721 3092
rect 11348 3148 11412 3152
rect 11348 3092 11352 3148
rect 11352 3092 11408 3148
rect 11408 3092 11412 3148
rect 11348 3088 11412 3092
rect 11428 3148 11492 3152
rect 11428 3092 11432 3148
rect 11432 3092 11488 3148
rect 11488 3092 11492 3148
rect 11428 3088 11492 3092
rect 11508 3148 11572 3152
rect 11508 3092 11512 3148
rect 11512 3092 11568 3148
rect 11568 3092 11572 3148
rect 11508 3088 11572 3092
rect 11588 3148 11652 3152
rect 11588 3092 11592 3148
rect 11592 3092 11648 3148
rect 11648 3092 11652 3148
rect 11588 3088 11652 3092
rect 18278 3148 18342 3152
rect 18278 3092 18282 3148
rect 18282 3092 18338 3148
rect 18338 3092 18342 3148
rect 18278 3088 18342 3092
rect 18358 3148 18422 3152
rect 18358 3092 18362 3148
rect 18362 3092 18418 3148
rect 18418 3092 18422 3148
rect 18358 3088 18422 3092
rect 18438 3148 18502 3152
rect 18438 3092 18442 3148
rect 18442 3092 18498 3148
rect 18498 3092 18502 3148
rect 18438 3088 18502 3092
rect 18518 3148 18582 3152
rect 18518 3092 18522 3148
rect 18522 3092 18578 3148
rect 18578 3092 18582 3148
rect 18518 3088 18582 3092
rect 7882 2604 7946 2608
rect 7882 2548 7886 2604
rect 7886 2548 7942 2604
rect 7942 2548 7946 2604
rect 7882 2544 7946 2548
rect 7962 2604 8026 2608
rect 7962 2548 7966 2604
rect 7966 2548 8022 2604
rect 8022 2548 8026 2604
rect 7962 2544 8026 2548
rect 8042 2604 8106 2608
rect 8042 2548 8046 2604
rect 8046 2548 8102 2604
rect 8102 2548 8106 2604
rect 8042 2544 8106 2548
rect 8122 2604 8186 2608
rect 8122 2548 8126 2604
rect 8126 2548 8182 2604
rect 8182 2548 8186 2604
rect 8122 2544 8186 2548
rect 14813 2604 14877 2608
rect 14813 2548 14817 2604
rect 14817 2548 14873 2604
rect 14873 2548 14877 2604
rect 14813 2544 14877 2548
rect 14893 2604 14957 2608
rect 14893 2548 14897 2604
rect 14897 2548 14953 2604
rect 14953 2548 14957 2604
rect 14893 2544 14957 2548
rect 14973 2604 15037 2608
rect 14973 2548 14977 2604
rect 14977 2548 15033 2604
rect 15033 2548 15037 2604
rect 14973 2544 15037 2548
rect 15053 2604 15117 2608
rect 15053 2548 15057 2604
rect 15057 2548 15113 2604
rect 15113 2548 15117 2604
rect 15053 2544 15117 2548
rect 4417 2060 4481 2064
rect 4417 2004 4421 2060
rect 4421 2004 4477 2060
rect 4477 2004 4481 2060
rect 4417 2000 4481 2004
rect 4497 2060 4561 2064
rect 4497 2004 4501 2060
rect 4501 2004 4557 2060
rect 4557 2004 4561 2060
rect 4497 2000 4561 2004
rect 4577 2060 4641 2064
rect 4577 2004 4581 2060
rect 4581 2004 4637 2060
rect 4637 2004 4641 2060
rect 4577 2000 4641 2004
rect 4657 2060 4721 2064
rect 4657 2004 4661 2060
rect 4661 2004 4717 2060
rect 4717 2004 4721 2060
rect 4657 2000 4721 2004
rect 11348 2060 11412 2064
rect 11348 2004 11352 2060
rect 11352 2004 11408 2060
rect 11408 2004 11412 2060
rect 11348 2000 11412 2004
rect 11428 2060 11492 2064
rect 11428 2004 11432 2060
rect 11432 2004 11488 2060
rect 11488 2004 11492 2060
rect 11428 2000 11492 2004
rect 11508 2060 11572 2064
rect 11508 2004 11512 2060
rect 11512 2004 11568 2060
rect 11568 2004 11572 2060
rect 11508 2000 11572 2004
rect 11588 2060 11652 2064
rect 11588 2004 11592 2060
rect 11592 2004 11648 2060
rect 11648 2004 11652 2060
rect 11588 2000 11652 2004
rect 18278 2060 18342 2064
rect 18278 2004 18282 2060
rect 18282 2004 18338 2060
rect 18338 2004 18342 2060
rect 18278 2000 18342 2004
rect 18358 2060 18422 2064
rect 18358 2004 18362 2060
rect 18362 2004 18418 2060
rect 18418 2004 18422 2060
rect 18358 2000 18422 2004
rect 18438 2060 18502 2064
rect 18438 2004 18442 2060
rect 18442 2004 18498 2060
rect 18498 2004 18502 2060
rect 18438 2000 18502 2004
rect 18518 2060 18582 2064
rect 18518 2004 18522 2060
rect 18522 2004 18578 2060
rect 18578 2004 18582 2060
rect 18518 2000 18582 2004
<< metal4 >>
rect 4409 20560 4729 20576
rect 4409 20496 4417 20560
rect 4481 20496 4497 20560
rect 4561 20496 4577 20560
rect 4641 20496 4657 20560
rect 4721 20496 4729 20560
rect 4409 19472 4729 20496
rect 4409 19408 4417 19472
rect 4481 19408 4497 19472
rect 4561 19408 4577 19472
rect 4641 19408 4657 19472
rect 4721 19408 4729 19472
rect 4409 18384 4729 19408
rect 4409 18320 4417 18384
rect 4481 18320 4497 18384
rect 4561 18320 4577 18384
rect 4641 18320 4657 18384
rect 4721 18320 4729 18384
rect 4409 17296 4729 18320
rect 4409 17232 4417 17296
rect 4481 17232 4497 17296
rect 4561 17232 4577 17296
rect 4641 17232 4657 17296
rect 4721 17232 4729 17296
rect 4409 16208 4729 17232
rect 4409 16144 4417 16208
rect 4481 16144 4497 16208
rect 4561 16144 4577 16208
rect 4641 16144 4657 16208
rect 4721 16144 4729 16208
rect 4409 15120 4729 16144
rect 4409 15056 4417 15120
rect 4481 15056 4497 15120
rect 4561 15056 4577 15120
rect 4641 15056 4657 15120
rect 4721 15056 4729 15120
rect 4409 14032 4729 15056
rect 4409 13968 4417 14032
rect 4481 13968 4497 14032
rect 4561 13968 4577 14032
rect 4641 13968 4657 14032
rect 4721 13968 4729 14032
rect 4409 12944 4729 13968
rect 4409 12880 4417 12944
rect 4481 12880 4497 12944
rect 4561 12880 4577 12944
rect 4641 12880 4657 12944
rect 4721 12880 4729 12944
rect 4409 11856 4729 12880
rect 4409 11792 4417 11856
rect 4481 11792 4497 11856
rect 4561 11792 4577 11856
rect 4641 11792 4657 11856
rect 4721 11792 4729 11856
rect 4409 10768 4729 11792
rect 4409 10704 4417 10768
rect 4481 10704 4497 10768
rect 4561 10704 4577 10768
rect 4641 10704 4657 10768
rect 4721 10704 4729 10768
rect 4409 9680 4729 10704
rect 4409 9616 4417 9680
rect 4481 9616 4497 9680
rect 4561 9616 4577 9680
rect 4641 9616 4657 9680
rect 4721 9616 4729 9680
rect 4409 8592 4729 9616
rect 4409 8528 4417 8592
rect 4481 8528 4497 8592
rect 4561 8528 4577 8592
rect 4641 8528 4657 8592
rect 4721 8528 4729 8592
rect 4409 7504 4729 8528
rect 4409 7440 4417 7504
rect 4481 7440 4497 7504
rect 4561 7440 4577 7504
rect 4641 7440 4657 7504
rect 4721 7440 4729 7504
rect 4409 6416 4729 7440
rect 4409 6352 4417 6416
rect 4481 6352 4497 6416
rect 4561 6352 4577 6416
rect 4641 6352 4657 6416
rect 4721 6352 4729 6416
rect 4409 5328 4729 6352
rect 4409 5264 4417 5328
rect 4481 5264 4497 5328
rect 4561 5264 4577 5328
rect 4641 5264 4657 5328
rect 4721 5264 4729 5328
rect 4409 4240 4729 5264
rect 4409 4176 4417 4240
rect 4481 4176 4497 4240
rect 4561 4176 4577 4240
rect 4641 4176 4657 4240
rect 4721 4176 4729 4240
rect 4409 3152 4729 4176
rect 4409 3088 4417 3152
rect 4481 3088 4497 3152
rect 4561 3088 4577 3152
rect 4641 3088 4657 3152
rect 4721 3088 4729 3152
rect 4409 2064 4729 3088
rect 4409 2000 4417 2064
rect 4481 2000 4497 2064
rect 4561 2000 4577 2064
rect 4641 2000 4657 2064
rect 4721 2000 4729 2064
rect 4409 1984 4729 2000
rect 7874 20016 8195 20576
rect 7874 19952 7882 20016
rect 7946 19952 7962 20016
rect 8026 19952 8042 20016
rect 8106 19952 8122 20016
rect 8186 19952 8195 20016
rect 7874 18928 8195 19952
rect 7874 18864 7882 18928
rect 7946 18864 7962 18928
rect 8026 18864 8042 18928
rect 8106 18864 8122 18928
rect 8186 18864 8195 18928
rect 7874 17840 8195 18864
rect 7874 17776 7882 17840
rect 7946 17776 7962 17840
rect 8026 17776 8042 17840
rect 8106 17776 8122 17840
rect 8186 17776 8195 17840
rect 7874 16752 8195 17776
rect 7874 16688 7882 16752
rect 7946 16688 7962 16752
rect 8026 16688 8042 16752
rect 8106 16688 8122 16752
rect 8186 16688 8195 16752
rect 7874 15664 8195 16688
rect 7874 15600 7882 15664
rect 7946 15600 7962 15664
rect 8026 15600 8042 15664
rect 8106 15600 8122 15664
rect 8186 15600 8195 15664
rect 7874 14576 8195 15600
rect 7874 14512 7882 14576
rect 7946 14512 7962 14576
rect 8026 14512 8042 14576
rect 8106 14512 8122 14576
rect 8186 14512 8195 14576
rect 7874 13488 8195 14512
rect 7874 13424 7882 13488
rect 7946 13424 7962 13488
rect 8026 13424 8042 13488
rect 8106 13424 8122 13488
rect 8186 13424 8195 13488
rect 7874 12400 8195 13424
rect 7874 12336 7882 12400
rect 7946 12336 7962 12400
rect 8026 12336 8042 12400
rect 8106 12336 8122 12400
rect 8186 12336 8195 12400
rect 7874 11312 8195 12336
rect 7874 11248 7882 11312
rect 7946 11248 7962 11312
rect 8026 11248 8042 11312
rect 8106 11248 8122 11312
rect 8186 11248 8195 11312
rect 7874 10224 8195 11248
rect 7874 10160 7882 10224
rect 7946 10160 7962 10224
rect 8026 10160 8042 10224
rect 8106 10160 8122 10224
rect 8186 10160 8195 10224
rect 7874 9136 8195 10160
rect 7874 9072 7882 9136
rect 7946 9072 7962 9136
rect 8026 9072 8042 9136
rect 8106 9072 8122 9136
rect 8186 9072 8195 9136
rect 7874 8048 8195 9072
rect 7874 7984 7882 8048
rect 7946 7984 7962 8048
rect 8026 7984 8042 8048
rect 8106 7984 8122 8048
rect 8186 7984 8195 8048
rect 7874 6960 8195 7984
rect 7874 6896 7882 6960
rect 7946 6896 7962 6960
rect 8026 6896 8042 6960
rect 8106 6896 8122 6960
rect 8186 6896 8195 6960
rect 7874 5872 8195 6896
rect 7874 5808 7882 5872
rect 7946 5808 7962 5872
rect 8026 5808 8042 5872
rect 8106 5808 8122 5872
rect 8186 5808 8195 5872
rect 7874 4784 8195 5808
rect 7874 4720 7882 4784
rect 7946 4720 7962 4784
rect 8026 4720 8042 4784
rect 8106 4720 8122 4784
rect 8186 4720 8195 4784
rect 7874 3696 8195 4720
rect 7874 3632 7882 3696
rect 7946 3632 7962 3696
rect 8026 3632 8042 3696
rect 8106 3632 8122 3696
rect 8186 3632 8195 3696
rect 7874 2608 8195 3632
rect 7874 2544 7882 2608
rect 7946 2544 7962 2608
rect 8026 2544 8042 2608
rect 8106 2544 8122 2608
rect 8186 2544 8195 2608
rect 7874 1984 8195 2544
rect 11340 20560 11660 20576
rect 11340 20496 11348 20560
rect 11412 20496 11428 20560
rect 11492 20496 11508 20560
rect 11572 20496 11588 20560
rect 11652 20496 11660 20560
rect 11340 19472 11660 20496
rect 11340 19408 11348 19472
rect 11412 19408 11428 19472
rect 11492 19408 11508 19472
rect 11572 19408 11588 19472
rect 11652 19408 11660 19472
rect 11340 18384 11660 19408
rect 11340 18320 11348 18384
rect 11412 18320 11428 18384
rect 11492 18320 11508 18384
rect 11572 18320 11588 18384
rect 11652 18320 11660 18384
rect 11340 17296 11660 18320
rect 11340 17232 11348 17296
rect 11412 17232 11428 17296
rect 11492 17232 11508 17296
rect 11572 17232 11588 17296
rect 11652 17232 11660 17296
rect 11340 16208 11660 17232
rect 11340 16144 11348 16208
rect 11412 16144 11428 16208
rect 11492 16144 11508 16208
rect 11572 16144 11588 16208
rect 11652 16144 11660 16208
rect 11340 15120 11660 16144
rect 11340 15056 11348 15120
rect 11412 15056 11428 15120
rect 11492 15056 11508 15120
rect 11572 15056 11588 15120
rect 11652 15056 11660 15120
rect 11340 14032 11660 15056
rect 11340 13968 11348 14032
rect 11412 13968 11428 14032
rect 11492 13968 11508 14032
rect 11572 13968 11588 14032
rect 11652 13968 11660 14032
rect 11340 12944 11660 13968
rect 11340 12880 11348 12944
rect 11412 12880 11428 12944
rect 11492 12880 11508 12944
rect 11572 12880 11588 12944
rect 11652 12880 11660 12944
rect 11340 11856 11660 12880
rect 11340 11792 11348 11856
rect 11412 11792 11428 11856
rect 11492 11792 11508 11856
rect 11572 11792 11588 11856
rect 11652 11792 11660 11856
rect 11340 10768 11660 11792
rect 11340 10704 11348 10768
rect 11412 10704 11428 10768
rect 11492 10704 11508 10768
rect 11572 10704 11588 10768
rect 11652 10704 11660 10768
rect 11340 9680 11660 10704
rect 11340 9616 11348 9680
rect 11412 9616 11428 9680
rect 11492 9616 11508 9680
rect 11572 9616 11588 9680
rect 11652 9616 11660 9680
rect 11340 8592 11660 9616
rect 11340 8528 11348 8592
rect 11412 8528 11428 8592
rect 11492 8528 11508 8592
rect 11572 8528 11588 8592
rect 11652 8528 11660 8592
rect 11340 7504 11660 8528
rect 11340 7440 11348 7504
rect 11412 7440 11428 7504
rect 11492 7440 11508 7504
rect 11572 7440 11588 7504
rect 11652 7440 11660 7504
rect 11340 6416 11660 7440
rect 11340 6352 11348 6416
rect 11412 6352 11428 6416
rect 11492 6352 11508 6416
rect 11572 6352 11588 6416
rect 11652 6352 11660 6416
rect 11340 5328 11660 6352
rect 11340 5264 11348 5328
rect 11412 5264 11428 5328
rect 11492 5264 11508 5328
rect 11572 5264 11588 5328
rect 11652 5264 11660 5328
rect 11340 4240 11660 5264
rect 11340 4176 11348 4240
rect 11412 4176 11428 4240
rect 11492 4176 11508 4240
rect 11572 4176 11588 4240
rect 11652 4176 11660 4240
rect 11340 3152 11660 4176
rect 11340 3088 11348 3152
rect 11412 3088 11428 3152
rect 11492 3088 11508 3152
rect 11572 3088 11588 3152
rect 11652 3088 11660 3152
rect 11340 2064 11660 3088
rect 11340 2000 11348 2064
rect 11412 2000 11428 2064
rect 11492 2000 11508 2064
rect 11572 2000 11588 2064
rect 11652 2000 11660 2064
rect 11340 1984 11660 2000
rect 14805 20016 15125 20576
rect 14805 19952 14813 20016
rect 14877 19952 14893 20016
rect 14957 19952 14973 20016
rect 15037 19952 15053 20016
rect 15117 19952 15125 20016
rect 14805 18928 15125 19952
rect 14805 18864 14813 18928
rect 14877 18864 14893 18928
rect 14957 18864 14973 18928
rect 15037 18864 15053 18928
rect 15117 18864 15125 18928
rect 14805 17840 15125 18864
rect 14805 17776 14813 17840
rect 14877 17776 14893 17840
rect 14957 17776 14973 17840
rect 15037 17776 15053 17840
rect 15117 17776 15125 17840
rect 14805 16752 15125 17776
rect 14805 16688 14813 16752
rect 14877 16688 14893 16752
rect 14957 16688 14973 16752
rect 15037 16688 15053 16752
rect 15117 16688 15125 16752
rect 14805 15664 15125 16688
rect 14805 15600 14813 15664
rect 14877 15600 14893 15664
rect 14957 15600 14973 15664
rect 15037 15600 15053 15664
rect 15117 15600 15125 15664
rect 14805 14576 15125 15600
rect 14805 14512 14813 14576
rect 14877 14512 14893 14576
rect 14957 14512 14973 14576
rect 15037 14512 15053 14576
rect 15117 14512 15125 14576
rect 14805 13488 15125 14512
rect 14805 13424 14813 13488
rect 14877 13424 14893 13488
rect 14957 13424 14973 13488
rect 15037 13424 15053 13488
rect 15117 13424 15125 13488
rect 14805 12400 15125 13424
rect 14805 12336 14813 12400
rect 14877 12336 14893 12400
rect 14957 12336 14973 12400
rect 15037 12336 15053 12400
rect 15117 12336 15125 12400
rect 14805 11312 15125 12336
rect 14805 11248 14813 11312
rect 14877 11248 14893 11312
rect 14957 11248 14973 11312
rect 15037 11248 15053 11312
rect 15117 11248 15125 11312
rect 14805 10224 15125 11248
rect 14805 10160 14813 10224
rect 14877 10160 14893 10224
rect 14957 10160 14973 10224
rect 15037 10160 15053 10224
rect 15117 10160 15125 10224
rect 14805 9136 15125 10160
rect 14805 9072 14813 9136
rect 14877 9072 14893 9136
rect 14957 9072 14973 9136
rect 15037 9072 15053 9136
rect 15117 9072 15125 9136
rect 14805 8048 15125 9072
rect 14805 7984 14813 8048
rect 14877 7984 14893 8048
rect 14957 7984 14973 8048
rect 15037 7984 15053 8048
rect 15117 7984 15125 8048
rect 14805 6960 15125 7984
rect 14805 6896 14813 6960
rect 14877 6896 14893 6960
rect 14957 6896 14973 6960
rect 15037 6896 15053 6960
rect 15117 6896 15125 6960
rect 14805 5872 15125 6896
rect 14805 5808 14813 5872
rect 14877 5808 14893 5872
rect 14957 5808 14973 5872
rect 15037 5808 15053 5872
rect 15117 5808 15125 5872
rect 14805 4784 15125 5808
rect 14805 4720 14813 4784
rect 14877 4720 14893 4784
rect 14957 4720 14973 4784
rect 15037 4720 15053 4784
rect 15117 4720 15125 4784
rect 14805 3696 15125 4720
rect 14805 3632 14813 3696
rect 14877 3632 14893 3696
rect 14957 3632 14973 3696
rect 15037 3632 15053 3696
rect 15117 3632 15125 3696
rect 14805 2608 15125 3632
rect 14805 2544 14813 2608
rect 14877 2544 14893 2608
rect 14957 2544 14973 2608
rect 15037 2544 15053 2608
rect 15117 2544 15125 2608
rect 14805 1984 15125 2544
rect 18270 20560 18591 20576
rect 18270 20496 18278 20560
rect 18342 20496 18358 20560
rect 18422 20496 18438 20560
rect 18502 20496 18518 20560
rect 18582 20496 18591 20560
rect 18270 19472 18591 20496
rect 18270 19408 18278 19472
rect 18342 19408 18358 19472
rect 18422 19408 18438 19472
rect 18502 19408 18518 19472
rect 18582 19408 18591 19472
rect 18270 18384 18591 19408
rect 18270 18320 18278 18384
rect 18342 18320 18358 18384
rect 18422 18320 18438 18384
rect 18502 18320 18518 18384
rect 18582 18320 18591 18384
rect 18270 17296 18591 18320
rect 18270 17232 18278 17296
rect 18342 17232 18358 17296
rect 18422 17232 18438 17296
rect 18502 17232 18518 17296
rect 18582 17232 18591 17296
rect 18270 16208 18591 17232
rect 18270 16144 18278 16208
rect 18342 16144 18358 16208
rect 18422 16144 18438 16208
rect 18502 16144 18518 16208
rect 18582 16144 18591 16208
rect 18270 15120 18591 16144
rect 18270 15056 18278 15120
rect 18342 15056 18358 15120
rect 18422 15056 18438 15120
rect 18502 15056 18518 15120
rect 18582 15056 18591 15120
rect 18270 14032 18591 15056
rect 18270 13968 18278 14032
rect 18342 13968 18358 14032
rect 18422 13968 18438 14032
rect 18502 13968 18518 14032
rect 18582 13968 18591 14032
rect 18270 12944 18591 13968
rect 18270 12880 18278 12944
rect 18342 12880 18358 12944
rect 18422 12880 18438 12944
rect 18502 12880 18518 12944
rect 18582 12880 18591 12944
rect 18270 11856 18591 12880
rect 18270 11792 18278 11856
rect 18342 11792 18358 11856
rect 18422 11792 18438 11856
rect 18502 11792 18518 11856
rect 18582 11792 18591 11856
rect 18270 10768 18591 11792
rect 18270 10704 18278 10768
rect 18342 10704 18358 10768
rect 18422 10704 18438 10768
rect 18502 10704 18518 10768
rect 18582 10704 18591 10768
rect 18270 9680 18591 10704
rect 18270 9616 18278 9680
rect 18342 9616 18358 9680
rect 18422 9616 18438 9680
rect 18502 9616 18518 9680
rect 18582 9616 18591 9680
rect 18270 8592 18591 9616
rect 18270 8528 18278 8592
rect 18342 8528 18358 8592
rect 18422 8528 18438 8592
rect 18502 8528 18518 8592
rect 18582 8528 18591 8592
rect 18270 7504 18591 8528
rect 18270 7440 18278 7504
rect 18342 7440 18358 7504
rect 18422 7440 18438 7504
rect 18502 7440 18518 7504
rect 18582 7440 18591 7504
rect 18270 6416 18591 7440
rect 18270 6352 18278 6416
rect 18342 6352 18358 6416
rect 18422 6352 18438 6416
rect 18502 6352 18518 6416
rect 18582 6352 18591 6416
rect 18270 5328 18591 6352
rect 18270 5264 18278 5328
rect 18342 5264 18358 5328
rect 18422 5264 18438 5328
rect 18502 5264 18518 5328
rect 18582 5264 18591 5328
rect 18270 4240 18591 5264
rect 18270 4176 18278 4240
rect 18342 4176 18358 4240
rect 18422 4176 18438 4240
rect 18502 4176 18518 4240
rect 18582 4176 18591 4240
rect 18270 3152 18591 4176
rect 18270 3088 18278 3152
rect 18342 3088 18358 3152
rect 18422 3088 18438 3152
rect 18502 3088 18518 3152
rect 18582 3088 18591 3152
rect 18270 2064 18591 3088
rect 18270 2000 18278 2064
rect 18342 2000 18358 2064
rect 18422 2000 18438 2064
rect 18502 2000 18518 2064
rect 18582 2000 18591 2064
rect 18270 1984 18591 2000
use sky130_fd_sc_hd__decap_12  FILLER_1_15 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 2484 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1608910539
transform 1 0 1380 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1608910539
transform 1 0 2484 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1608910539
transform 1 0 1380 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1104 0 1 2576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608910539
transform 1 0 1104 0 -1 2576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_32
timestamp 1608910539
transform 1 0 4048 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3588 0 1 2576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1608910539
transform 1 0 4048 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1608910539
transform 1 0 3588 0 -1 2576
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3956 0 1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1608910539
transform 1 0 3956 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_56
timestamp 1608910539
transform 1 0 6256 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_44
timestamp 1608910539
transform 1 0 5152 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 6256 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1608910539
transform 1 0 5152 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608910539
transform 1 0 6808 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_80
timestamp 1608910539
transform 1 0 8464 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_68
timestamp 1608910539
transform 1 0 7360 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1608910539
transform 1 0 8004 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1608910539
transform 1 0 6900 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_93
timestamp 1608910539
transform 1 0 9660 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1608910539
transform 1 0 9752 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1608910539
transform 1 0 9108 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608910539
transform 1 0 9568 0 1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608910539
transform 1 0 9660 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_117
timestamp 1608910539
transform 1 0 11868 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_105
timestamp 1608910539
transform 1 0 10764 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1608910539
transform 1 0 12604 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1608910539
transform 1 0 11960 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1608910539
transform 1 0 10856 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608910539
transform 1 0 12512 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_141
timestamp 1608910539
transform 1 0 14076 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_129
timestamp 1608910539
transform 1 0 12972 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1608910539
transform 1 0 13708 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_166
timestamp 1608910539
transform 1 0 16376 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_154
timestamp 1608910539
transform 1 0 15272 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1608910539
transform 1 0 15456 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1608910539
transform 1 0 14812 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608910539
transform 1 0 15180 0 1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608910539
transform 1 0 15364 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_178
timestamp 1608910539
transform 1 0 17480 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1608910539
transform 1 0 18308 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1608910539
transform 1 0 17664 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1608910539
transform 1 0 16560 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608910539
transform 1 0 18216 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_202
timestamp 1608910539
transform 1 0 19688 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_190
timestamp 1608910539
transform 1 0 18584 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1608910539
transform 1 0 19412 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_215 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 20884 0 1 2576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_222 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 21528 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_218
timestamp 1608910539
transform 1 0 21160 0 -1 2576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1608910539
transform 1 0 20516 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608910539
transform 1 0 20792 0 1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608910539
transform 1 0 21068 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608910539
transform -1 0 21896 0 1 2576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608910539
transform -1 0 21896 0 -1 2576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1608910539
transform 1 0 2484 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1608910539
transform 1 0 1380 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608910539
transform 1 0 1104 0 -1 3664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_39
timestamp 1608910539
transform 1 0 4692 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_27
timestamp 1608910539
transform 1 0 3588 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_62
timestamp 1608910539
transform 1 0 6808 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 6532 0 -1 3664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_51
timestamp 1608910539
transform 1 0 5796 0 -1 3664
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608910539
transform 1 0 6716 0 -1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_74
timestamp 1608910539
transform 1 0 7912 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_98
timestamp 1608910539
transform 1 0 10120 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_86
timestamp 1608910539
transform 1 0 9016 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_123
timestamp 1608910539
transform 1 0 12420 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_110
timestamp 1608910539
transform 1 0 11224 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608910539
transform 1 0 12328 0 -1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_135
timestamp 1608910539
transform 1 0 13524 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_159
timestamp 1608910539
transform 1 0 15732 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_147
timestamp 1608910539
transform 1 0 14628 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_184
timestamp 1608910539
transform 1 0 18032 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_171
timestamp 1608910539
transform 1 0 16836 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608910539
transform 1 0 17940 0 -1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_208
timestamp 1608910539
transform 1 0 20240 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_196
timestamp 1608910539
transform 1 0 19136 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_220
timestamp 1608910539
transform 1 0 21344 0 -1 3664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608910539
transform -1 0 21896 0 -1 3664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1608910539
transform 1 0 2484 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1608910539
transform 1 0 1380 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608910539
transform 1 0 1104 0 1 3664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_32
timestamp 1608910539
transform 1 0 4048 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 1608910539
transform 1 0 3588 0 1 3664
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608910539
transform 1 0 3956 0 1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_56
timestamp 1608910539
transform 1 0 6256 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_44
timestamp 1608910539
transform 1 0 5152 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_80
timestamp 1608910539
transform 1 0 8464 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_68
timestamp 1608910539
transform 1 0 7360 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_93
timestamp 1608910539
transform 1 0 9660 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608910539
transform 1 0 9568 0 1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_117
timestamp 1608910539
transform 1 0 11868 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_105
timestamp 1608910539
transform 1 0 10764 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_141
timestamp 1608910539
transform 1 0 14076 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_129
timestamp 1608910539
transform 1 0 12972 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_166
timestamp 1608910539
transform 1 0 16376 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_154
timestamp 1608910539
transform 1 0 15272 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608910539
transform 1 0 15180 0 1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_178
timestamp 1608910539
transform 1 0 17480 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_202
timestamp 1608910539
transform 1 0 19688 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_190
timestamp 1608910539
transform 1 0 18584 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_220
timestamp 1608910539
transform 1 0 21344 0 1 3664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_215
timestamp 1608910539
transform 1 0 20884 0 1 3664
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__87__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 21160 0 1 3664
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608910539
transform 1 0 20792 0 1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608910539
transform -1 0 21896 0 1 3664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1608910539
transform 1 0 2484 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1608910539
transform 1 0 1380 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608910539
transform 1 0 1104 0 -1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_39
timestamp 1608910539
transform 1 0 4692 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_27
timestamp 1608910539
transform 1 0 3588 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_62
timestamp 1608910539
transform 1 0 6808 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_59
timestamp 1608910539
transform 1 0 6532 0 -1 4752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_51
timestamp 1608910539
transform 1 0 5796 0 -1 4752
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608910539
transform 1 0 6716 0 -1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_74
timestamp 1608910539
transform 1 0 7912 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_98
timestamp 1608910539
transform 1 0 10120 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_86
timestamp 1608910539
transform 1 0 9016 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_123
timestamp 1608910539
transform 1 0 12420 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_110
timestamp 1608910539
transform 1 0 11224 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608910539
transform 1 0 12328 0 -1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_135
timestamp 1608910539
transform 1 0 13524 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_159
timestamp 1608910539
transform 1 0 15732 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_147
timestamp 1608910539
transform 1 0 14628 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_184
timestamp 1608910539
transform 1 0 18032 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_171
timestamp 1608910539
transform 1 0 16836 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608910539
transform 1 0 17940 0 -1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_208
timestamp 1608910539
transform 1 0 20240 0 -1 4752
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_196
timestamp 1608910539
transform 1 0 19136 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_222
timestamp 1608910539
transform 1 0 21528 0 -1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_218
timestamp 1608910539
transform 1 0 21160 0 -1 4752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608910539
transform -1 0 21896 0 -1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _87_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 20792 0 -1 4752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1608910539
transform 1 0 2484 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1608910539
transform 1 0 1380 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608910539
transform 1 0 1104 0 1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_32
timestamp 1608910539
transform 1 0 4048 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_27
timestamp 1608910539
transform 1 0 3588 0 1 4752
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608910539
transform 1 0 3956 0 1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_56
timestamp 1608910539
transform 1 0 6256 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_44
timestamp 1608910539
transform 1 0 5152 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_80
timestamp 1608910539
transform 1 0 8464 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_68
timestamp 1608910539
transform 1 0 7360 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1608910539
transform 1 0 9660 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608910539
transform 1 0 9568 0 1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_117
timestamp 1608910539
transform 1 0 11868 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_105
timestamp 1608910539
transform 1 0 10764 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_141
timestamp 1608910539
transform 1 0 14076 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_129
timestamp 1608910539
transform 1 0 12972 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_166
timestamp 1608910539
transform 1 0 16376 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_154
timestamp 1608910539
transform 1 0 15272 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608910539
transform 1 0 15180 0 1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_178
timestamp 1608910539
transform 1 0 17480 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_202
timestamp 1608910539
transform 1 0 19688 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_190
timestamp 1608910539
transform 1 0 18584 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_220
timestamp 1608910539
transform 1 0 21344 0 1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_215
timestamp 1608910539
transform 1 0 20884 0 1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1608910539
transform 1 0 21160 0 1 4752
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608910539
transform 1 0 20792 0 1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608910539
transform -1 0 21896 0 1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1608910539
transform 1 0 2484 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1608910539
transform 1 0 1380 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1608910539
transform 1 0 2484 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1608910539
transform 1 0 1380 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608910539
transform 1 0 1104 0 1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608910539
transform 1 0 1104 0 -1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_32
timestamp 1608910539
transform 1 0 4048 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1608910539
transform 1 0 3588 0 1 5840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_39
timestamp 1608910539
transform 1 0 4692 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_27
timestamp 1608910539
transform 1 0 3588 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608910539
transform 1 0 3956 0 1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_56
timestamp 1608910539
transform 1 0 6256 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_44
timestamp 1608910539
transform 1 0 5152 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_62
timestamp 1608910539
transform 1 0 6808 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_59
timestamp 1608910539
transform 1 0 6532 0 -1 5840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_51
timestamp 1608910539
transform 1 0 5796 0 -1 5840
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608910539
transform 1 0 6716 0 -1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_80
timestamp 1608910539
transform 1 0 8464 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_68
timestamp 1608910539
transform 1 0 7360 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_74
timestamp 1608910539
transform 1 0 7912 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1608910539
transform 1 0 9660 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_98
timestamp 1608910539
transform 1 0 10120 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_86
timestamp 1608910539
transform 1 0 9016 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608910539
transform 1 0 9568 0 1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_117
timestamp 1608910539
transform 1 0 11868 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_105
timestamp 1608910539
transform 1 0 10764 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_123
timestamp 1608910539
transform 1 0 12420 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_110
timestamp 1608910539
transform 1 0 11224 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608910539
transform 1 0 12328 0 -1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_141
timestamp 1608910539
transform 1 0 14076 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_129
timestamp 1608910539
transform 1 0 12972 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_135
timestamp 1608910539
transform 1 0 13524 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_166
timestamp 1608910539
transform 1 0 16376 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_154
timestamp 1608910539
transform 1 0 15272 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_159
timestamp 1608910539
transform 1 0 15732 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_147
timestamp 1608910539
transform 1 0 14628 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608910539
transform 1 0 15180 0 1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_178
timestamp 1608910539
transform 1 0 17480 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_184
timestamp 1608910539
transform 1 0 18032 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_171
timestamp 1608910539
transform 1 0 16836 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608910539
transform 1 0 17940 0 -1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_202
timestamp 1608910539
transform 1 0 19688 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_190
timestamp 1608910539
transform 1 0 18584 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_208
timestamp 1608910539
transform 1 0 20240 0 -1 5840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_196
timestamp 1608910539
transform 1 0 19136 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_219
timestamp 1608910539
transform 1 0 21252 0 1 5840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_222
timestamp 1608910539
transform 1 0 21528 0 -1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_218
timestamp 1608910539
transform 1 0 21160 0 -1 5840
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608910539
transform 1 0 20792 0 1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608910539
transform -1 0 21896 0 1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608910539
transform -1 0 21896 0 -1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1608910539
transform 1 0 20884 0 1 5840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1608910539
transform 1 0 20792 0 -1 5840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1608910539
transform 1 0 2484 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1608910539
transform 1 0 1380 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608910539
transform 1 0 1104 0 -1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_39
timestamp 1608910539
transform 1 0 4692 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_27
timestamp 1608910539
transform 1 0 3588 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_62
timestamp 1608910539
transform 1 0 6808 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_59
timestamp 1608910539
transform 1 0 6532 0 -1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_51
timestamp 1608910539
transform 1 0 5796 0 -1 6928
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608910539
transform 1 0 6716 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_77
timestamp 1608910539
transform 1 0 8188 0 -1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_74
timestamp 1608910539
transform 1 0 7912 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608910539
transform 1 0 8004 0 -1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 8372 0 -1 6928
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_8_95
timestamp 1608910539
transform 1 0 9844 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_125
timestamp 1608910539
transform 1 0 12604 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_120
timestamp 1608910539
transform 1 0 12144 0 -1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_109
timestamp 1608910539
transform 1 0 11132 0 -1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 10948 0 -1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 12420 0 -1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608910539
transform 1 0 12328 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 11316 0 -1 6928
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_141
timestamp 1608910539
transform 1 0 14076 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_137
timestamp 1608910539
transform 1 0 13708 0 -1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1608910539
transform 1 0 14168 0 -1 6928
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_8_155
timestamp 1608910539
transform 1 0 15364 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1608910539
transform 1 0 14996 0 -1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 15180 0 -1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_187
timestamp 1608910539
transform 1 0 18308 0 -1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_179
timestamp 1608910539
transform 1 0 17572 0 -1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_167
timestamp 1608910539
transform 1 0 16468 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608910539
transform 1 0 17940 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _35_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 18032 0 -1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_203
timestamp 1608910539
transform 1 0 19780 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_191
timestamp 1608910539
transform 1 0 18676 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 18492 0 -1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_221
timestamp 1608910539
transform 1 0 21436 0 -1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1608910539
transform 1 0 20884 0 -1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1608910539
transform 1 0 21252 0 -1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608910539
transform -1 0 21896 0 -1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1608910539
transform 1 0 2484 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1608910539
transform 1 0 1380 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608910539
transform 1 0 1104 0 1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_32
timestamp 1608910539
transform 1 0 4048 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_27
timestamp 1608910539
transform 1 0 3588 0 1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608910539
transform 1 0 3956 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_56
timestamp 1608910539
transform 1 0 6256 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_44
timestamp 1608910539
transform 1 0 5152 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_80
timestamp 1608910539
transform 1 0 8464 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_68
timestamp 1608910539
transform 1 0 7360 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_93
timestamp 1608910539
transform 1 0 9660 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608910539
transform 1 0 9568 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9844 0 1 6928
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_9_111
timestamp 1608910539
transform 1 0 11316 0 1 6928
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 11868 0 1 6928
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_140
timestamp 1608910539
transform 1 0 13984 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_137
timestamp 1608910539
transform 1 0 13708 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_133
timestamp 1608910539
transform 1 0 13340 0 1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 13800 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1608910539
transform 1 0 14168 0 1 6928
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_154
timestamp 1608910539
transform 1 0 15272 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_151
timestamp 1608910539
transform 1 0 14996 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608910539
transform 1 0 15180 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15364 0 1 6928
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_171
timestamp 1608910539
transform 1 0 16836 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 17020 0 1 6928
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_9_204
timestamp 1608910539
transform 1 0 19872 0 1 6928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_200
timestamp 1608910539
transform 1 0 19504 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_189
timestamp 1608910539
transform 1 0 18492 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 19688 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1608910539
transform 1 0 18676 0 1 6928
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_219
timestamp 1608910539
transform 1 0 21252 0 1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_212
timestamp 1608910539
transform 1 0 20608 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1608910539
transform 1 0 20424 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608910539
transform 1 0 20792 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608910539
transform -1 0 21896 0 1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1608910539
transform 1 0 20884 0 1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1608910539
transform 1 0 2484 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1608910539
transform 1 0 1380 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608910539
transform 1 0 1104 0 -1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_39
timestamp 1608910539
transform 1 0 4692 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_27
timestamp 1608910539
transform 1 0 3588 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_62
timestamp 1608910539
transform 1 0 6808 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_59
timestamp 1608910539
transform 1 0 6532 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_51
timestamp 1608910539
transform 1 0 5796 0 -1 8016
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608910539
transform 1 0 6716 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_74
timestamp 1608910539
transform 1 0 7912 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_98
timestamp 1608910539
transform 1 0 10120 0 -1 8016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_86
timestamp 1608910539
transform 1 0 9016 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1608910539
transform 1 0 10672 0 -1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_123
timestamp 1608910539
transform 1 0 12420 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_118
timestamp 1608910539
transform 1 0 11960 0 -1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_107
timestamp 1608910539
transform 1 0 10948 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608910539
transform 1 0 12328 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 11132 0 -1 8016
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_135
timestamp 1608910539
transform 1 0 13524 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 13616 0 -1 8016
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_10_157
timestamp 1608910539
transform 1 0 15548 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_152
timestamp 1608910539
transform 1 0 15088 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1608910539
transform 1 0 15272 0 -1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_184
timestamp 1608910539
transform 1 0 18032 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_181
timestamp 1608910539
transform 1 0 17756 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_169
timestamp 1608910539
transform 1 0 16652 0 -1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608910539
transform 1 0 17940 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1608910539
transform 1 0 16928 0 -1 8016
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 18216 0 -1 8016
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_10_202
timestamp 1608910539
transform 1 0 19688 0 -1 8016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_222
timestamp 1608910539
transform 1 0 21528 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_218
timestamp 1608910539
transform 1 0 21160 0 -1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_212
timestamp 1608910539
transform 1 0 20608 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1608910539
transform 1 0 20424 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608910539
transform -1 0 21896 0 -1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1608910539
transform 1 0 20792 0 -1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1608910539
transform 1 0 2484 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1608910539
transform 1 0 1380 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608910539
transform 1 0 1104 0 1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_32
timestamp 1608910539
transform 1 0 4048 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_27
timestamp 1608910539
transform 1 0 3588 0 1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608910539
transform 1 0 3956 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_56
timestamp 1608910539
transform 1 0 6256 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_44
timestamp 1608910539
transform 1 0 5152 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_80
timestamp 1608910539
transform 1 0 8464 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_68
timestamp 1608910539
transform 1 0 7360 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1608910539
transform 1 0 9660 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608910539
transform 1 0 9568 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_114
timestamp 1608910539
transform 1 0 11592 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_105
timestamp 1608910539
transform 1 0 10764 0 1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 11040 0 1 8016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_140
timestamp 1608910539
transform 1 0 13984 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_126
timestamp 1608910539
transform 1 0 12696 0 1 8016
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 13432 0 1 8016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_154
timestamp 1608910539
transform 1 0 15272 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_152
timestamp 1608910539
transform 1 0 15088 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608910539
transform 1 0 15180 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 16376 0 1 8016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1608910539
transform 1 0 18032 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_172
timestamp 1608910539
transform 1 0 16928 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_208
timestamp 1608910539
transform 1 0 20240 0 1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1608910539
transform 1 0 19136 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_219
timestamp 1608910539
transform 1 0 21252 0 1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_212
timestamp 1608910539
transform 1 0 20608 0 1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1608910539
transform 1 0 20424 0 1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608910539
transform 1 0 20792 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608910539
transform -1 0 21896 0 1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1608910539
transform 1 0 20884 0 1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1608910539
transform 1 0 2484 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1608910539
transform 1 0 1380 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608910539
transform 1 0 1104 0 -1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_39
timestamp 1608910539
transform 1 0 4692 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_27
timestamp 1608910539
transform 1 0 3588 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_62
timestamp 1608910539
transform 1 0 6808 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_59
timestamp 1608910539
transform 1 0 6532 0 -1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_51
timestamp 1608910539
transform 1 0 5796 0 -1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608910539
transform 1 0 6716 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_74
timestamp 1608910539
transform 1 0 7912 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_98
timestamp 1608910539
transform 1 0 10120 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_86
timestamp 1608910539
transform 1 0 9016 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_123
timestamp 1608910539
transform 1 0 12420 0 -1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_119
timestamp 1608910539
transform 1 0 12052 0 -1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_114
timestamp 1608910539
transform 1 0 11592 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_110
timestamp 1608910539
transform 1 0 11224 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608910539
transform 1 0 12328 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1608910539
transform 1 0 11684 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_136
timestamp 1608910539
transform 1 0 13616 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_131
timestamp 1608910539
transform 1 0 13156 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1608910539
transform 1 0 13248 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1608910539
transform 1 0 16376 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_158
timestamp 1608910539
transform 1 0 15640 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_154
timestamp 1608910539
transform 1 0 15272 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_148
timestamp 1608910539
transform 1 0 14720 0 -1 9104
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1608910539
transform 1 0 16008 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _42_
timestamp 1608910539
transform 1 0 15364 0 -1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_184
timestamp 1608910539
transform 1 0 18032 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_182
timestamp 1608910539
transform 1 0 17848 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_178
timestamp 1608910539
transform 1 0 17480 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608910539
transform 1 0 17940 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_208
timestamp 1608910539
transform 1 0 20240 0 -1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_204
timestamp 1608910539
transform 1 0 19872 0 -1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_196
timestamp 1608910539
transform 1 0 19136 0 -1 9104
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1608910539
transform 1 0 19688 0 -1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 20056 0 -1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_222
timestamp 1608910539
transform 1 0 21528 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_218
timestamp 1608910539
transform 1 0 21160 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_212
timestamp 1608910539
transform 1 0 20608 0 -1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1608910539
transform 1 0 20424 0 -1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608910539
transform -1 0 21896 0 -1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1608910539
transform 1 0 20792 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1608910539
transform 1 0 2484 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1608910539
transform 1 0 1380 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1608910539
transform 1 0 2484 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1608910539
transform 1 0 1380 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608910539
transform 1 0 1104 0 -1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608910539
transform 1 0 1104 0 1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_39
timestamp 1608910539
transform 1 0 4692 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_27
timestamp 1608910539
transform 1 0 3588 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_32
timestamp 1608910539
transform 1 0 4048 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_27
timestamp 1608910539
transform 1 0 3588 0 1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608910539
transform 1 0 3956 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_62
timestamp 1608910539
transform 1 0 6808 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_59
timestamp 1608910539
transform 1 0 6532 0 -1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_51
timestamp 1608910539
transform 1 0 5796 0 -1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_56
timestamp 1608910539
transform 1 0 6256 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_44
timestamp 1608910539
transform 1 0 5152 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1608910539
transform 1 0 6716 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_80
timestamp 1608910539
transform 1 0 8464 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_68
timestamp 1608910539
transform 1 0 7360 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 7912 0 -1 10192
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_14_102
timestamp 1608910539
transform 1 0 10488 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_90
timestamp 1608910539
transform 1 0 9384 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_97
timestamp 1608910539
transform 1 0 10028 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_93
timestamp 1608910539
transform 1 0 9660 0 1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608910539
transform 1 0 9568 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 10120 0 1 9104
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_14_123
timestamp 1608910539
transform 1 0 12420 0 -1 10192
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_114
timestamp 1608910539
transform 1 0 11592 0 -1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_114
timestamp 1608910539
transform 1 0 11592 0 1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1608910539
transform 1 0 12328 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 11776 0 1 9104
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_14_139
timestamp 1608910539
transform 1 0 13892 0 -1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_129
timestamp 1608910539
transform 1 0 12972 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_143
timestamp 1608910539
transform 1 0 14260 0 1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_132
timestamp 1608910539
transform 1 0 13248 0 1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1608910539
transform 1 0 13432 0 1 9104
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1608910539
transform 1 0 13064 0 -1 10192
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 14168 0 -1 10192
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_14_158
timestamp 1608910539
transform 1 0 15640 0 -1 10192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_163
timestamp 1608910539
transform 1 0 16100 0 1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_151
timestamp 1608910539
transform 1 0 14996 0 1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 16284 0 1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608910539
transform 1 0 15180 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1608910539
transform 1 0 15272 0 1 9104
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 16192 0 -1 10192
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_14_180
timestamp 1608910539
transform 1 0 17664 0 -1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_179
timestamp 1608910539
transform 1 0 17572 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_167
timestamp 1608910539
transform 1 0 16468 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1608910539
transform 1 0 17940 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 18032 0 -1 10192
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_14_200
timestamp 1608910539
transform 1 0 19504 0 -1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_207
timestamp 1608910539
transform 1 0 20148 0 1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1608910539
transform 1 0 19688 0 -1 10192
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 18676 0 1 9104
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_14_211
timestamp 1608910539
transform 1 0 20516 0 -1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_212
timestamp 1608910539
transform 1 0 20608 0 1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1608910539
transform 1 0 20424 0 1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_218
timestamp 1608910539
transform 1 0 21160 0 -1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608910539
transform 1 0 20792 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1608910539
transform 1 0 20792 0 -1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1608910539
transform 1 0 20884 0 1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_222
timestamp 1608910539
transform 1 0 21528 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_219
timestamp 1608910539
transform 1 0 21252 0 1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608910539
transform -1 0 21896 0 -1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608910539
transform -1 0 21896 0 1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1608910539
transform 1 0 2484 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1608910539
transform 1 0 1380 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608910539
transform 1 0 1104 0 1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_32
timestamp 1608910539
transform 1 0 4048 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_27
timestamp 1608910539
transform 1 0 3588 0 1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1608910539
transform 1 0 3956 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_56
timestamp 1608910539
transform 1 0 6256 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_44
timestamp 1608910539
transform 1 0 5152 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_74
timestamp 1608910539
transform 1 0 7912 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_68
timestamp 1608910539
transform 1 0 7360 0 1 10192
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8004 0 1 10192
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_15_101
timestamp 1608910539
transform 1 0 10396 0 1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_93
timestamp 1608910539
transform 1 0 9660 0 1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_84
timestamp 1608910539
transform 1 0 8832 0 1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1608910539
transform 1 0 9568 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1608910539
transform 1 0 10672 0 1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_122
timestamp 1608910539
transform 1 0 12328 0 1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_118
timestamp 1608910539
transform 1 0 11960 0 1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_107
timestamp 1608910539
transform 1 0 10948 0 1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 12512 0 1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 12144 0 1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1608910539
transform 1 0 11132 0 1 10192
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_144
timestamp 1608910539
transform 1 0 14352 0 1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_134
timestamp 1608910539
transform 1 0 13432 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_126
timestamp 1608910539
transform 1 0 12696 0 1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1608910539
transform 1 0 13524 0 1 10192
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_15_156
timestamp 1608910539
transform 1 0 15456 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_152
timestamp 1608910539
transform 1 0 15088 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_148
timestamp 1608910539
transform 1 0 14720 0 1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 15272 0 1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 14536 0 1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1608910539
transform 1 0 15180 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_180
timestamp 1608910539
transform 1 0 17664 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_168
timestamp 1608910539
transform 1 0 16560 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_206
timestamp 1608910539
transform 1 0 20056 0 1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_195
timestamp 1608910539
transform 1 0 19044 0 1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_192
timestamp 1608910539
transform 1 0 18768 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 18860 0 1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1608910539
transform 1 0 19228 0 1 10192
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1608910539
transform 1 0 20240 0 1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_219
timestamp 1608910539
transform 1 0 21252 0 1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_211
timestamp 1608910539
transform 1 0 20516 0 1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1608910539
transform 1 0 20792 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608910539
transform -1 0 21896 0 1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1608910539
transform 1 0 20884 0 1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1608910539
transform 1 0 2484 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1608910539
transform 1 0 1380 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608910539
transform 1 0 1104 0 -1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_39
timestamp 1608910539
transform 1 0 4692 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_27
timestamp 1608910539
transform 1 0 3588 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_62
timestamp 1608910539
transform 1 0 6808 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_59
timestamp 1608910539
transform 1 0 6532 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_51
timestamp 1608910539
transform 1 0 5796 0 -1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1608910539
transform 1 0 6716 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_74
timestamp 1608910539
transform 1 0 7912 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1608910539
transform 1 0 8096 0 -1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_101
timestamp 1608910539
transform 1 0 10396 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_93
timestamp 1608910539
transform 1 0 9660 0 -1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_89
timestamp 1608910539
transform 1 0 9292 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1608910539
transform 1 0 8924 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 9476 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 9108 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1608910539
transform 1 0 10488 0 -1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_16_123
timestamp 1608910539
transform 1 0 12420 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_119
timestamp 1608910539
transform 1 0 12052 0 -1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_111
timestamp 1608910539
transform 1 0 11316 0 -1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1608910539
transform 1 0 12328 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_138
timestamp 1608910539
transform 1 0 13800 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_right_track_0.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 13524 0 -1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_162
timestamp 1608910539
transform 1 0 16008 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_150
timestamp 1608910539
transform 1 0 14904 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_184
timestamp 1608910539
transform 1 0 18032 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_182
timestamp 1608910539
transform 1 0 17848 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_174
timestamp 1608910539
transform 1 0 17112 0 -1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1608910539
transform 1 0 17940 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_208
timestamp 1608910539
transform 1 0 20240 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_202
timestamp 1608910539
transform 1 0 19688 0 -1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__81__A
timestamp 1608910539
transform 1 0 20056 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 19136 0 -1 11280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_222
timestamp 1608910539
transform 1 0 21528 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_218
timestamp 1608910539
transform 1 0 21160 0 -1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_212
timestamp 1608910539
transform 1 0 20608 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__79__A
timestamp 1608910539
transform 1 0 20424 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608910539
transform -1 0 21896 0 -1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1608910539
transform 1 0 20792 0 -1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1608910539
transform 1 0 2484 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1608910539
transform 1 0 1380 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608910539
transform 1 0 1104 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_32
timestamp 1608910539
transform 1 0 4048 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_27
timestamp 1608910539
transform 1 0 3588 0 1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1608910539
transform 1 0 3956 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_56
timestamp 1608910539
transform 1 0 6256 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_44
timestamp 1608910539
transform 1 0 5152 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_73
timestamp 1608910539
transform 1 0 7820 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_68
timestamp 1608910539
transform 1 0 7360 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 7636 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8004 0 1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_88
timestamp 1608910539
transform 1 0 9200 0 1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_84
timestamp 1608910539
transform 1 0 8832 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9016 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1608910539
transform 1 0 9568 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 9660 0 1 11280
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_125
timestamp 1608910539
transform 1 0 12604 0 1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1608910539
transform 1 0 11500 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_109
timestamp 1608910539
transform 1 0 11132 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 11316 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_129
timestamp 1608910539
transform 1 0 12972 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 13064 0 1 11280
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_17_152
timestamp 1608910539
transform 1 0 15088 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_146
timestamp 1608910539
transform 1 0 14536 0 1 11280
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1608910539
transform 1 0 15180 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 15272 0 1 11280
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_183
timestamp 1608910539
transform 1 0 17940 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_178
timestamp 1608910539
transform 1 0 17480 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_170
timestamp 1608910539
transform 1 0 16744 0 1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1608910539
transform 1 0 18124 0 1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1608910539
transform 1 0 17664 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_204
timestamp 1608910539
transform 1 0 19872 0 1 11280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_200
timestamp 1608910539
transform 1 0 19504 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_194
timestamp 1608910539
transform 1 0 18952 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 19688 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1608910539
transform 1 0 19136 0 1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_219
timestamp 1608910539
transform 1 0 21252 0 1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_212
timestamp 1608910539
transform 1 0 20608 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__82__A
timestamp 1608910539
transform 1 0 20424 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1608910539
transform 1 0 20792 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608910539
transform -1 0 21896 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1608910539
transform 1 0 20884 0 1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1608910539
transform 1 0 2484 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1608910539
transform 1 0 1380 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608910539
transform 1 0 1104 0 -1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_39
timestamp 1608910539
transform 1 0 4692 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_27
timestamp 1608910539
transform 1 0 3588 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_62
timestamp 1608910539
transform 1 0 6808 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_59
timestamp 1608910539
transform 1 0 6532 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_51
timestamp 1608910539
transform 1 0 5796 0 -1 12368
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1608910539
transform 1 0 6716 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_74
timestamp 1608910539
transform 1 0 7912 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_98
timestamp 1608910539
transform 1 0 10120 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_86
timestamp 1608910539
transform 1 0 9016 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1608910539
transform 1 0 10304 0 -1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_123
timestamp 1608910539
transform 1 0 12420 0 -1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_118
timestamp 1608910539
transform 1 0 11960 0 -1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_109
timestamp 1608910539
transform 1 0 11132 0 -1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1608910539
transform 1 0 12328 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 11408 0 -1 12368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1608910539
transform 1 0 14076 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_130
timestamp 1608910539
transform 1 0 13064 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_127
timestamp 1608910539
transform 1 0 12788 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 12880 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 14260 0 -1 12368
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1608910539
transform 1 0 13248 0 -1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_156
timestamp 1608910539
transform 1 0 15456 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_153
timestamp 1608910539
transform 1 0 15180 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_149
timestamp 1608910539
transform 1 0 14812 0 -1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 15272 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 15640 0 -1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_18_182
timestamp 1608910539
transform 1 0 17848 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_178
timestamp 1608910539
transform 1 0 17480 0 -1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_167
timestamp 1608910539
transform 1 0 16468 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1608910539
transform 1 0 17940 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1608910539
transform 1 0 18032 0 -1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1608910539
transform 1 0 16652 0 -1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_202
timestamp 1608910539
transform 1 0 19688 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_198
timestamp 1608910539
transform 1 0 19320 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_193
timestamp 1608910539
transform 1 0 18860 0 -1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 19136 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__83__A
timestamp 1608910539
transform 1 0 19504 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 19872 0 -1 12368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_222
timestamp 1608910539
transform 1 0 21528 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_218
timestamp 1608910539
transform 1 0 21160 0 -1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_210
timestamp 1608910539
transform 1 0 20424 0 -1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608910539
transform -1 0 21896 0 -1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1608910539
transform 1 0 20792 0 -1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1608910539
transform 1 0 2484 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1608910539
transform 1 0 1380 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1608910539
transform 1 0 2484 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1608910539
transform 1 0 1380 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608910539
transform 1 0 1104 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608910539
transform 1 0 1104 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1608910539
transform 1 0 3588 0 -1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_32
timestamp 1608910539
transform 1 0 4048 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_27
timestamp 1608910539
transform 1 0 3588 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1608910539
transform 1 0 3956 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 3772 0 -1 13456
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_20_62
timestamp 1608910539
transform 1 0 6808 0 -1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_57
timestamp 1608910539
transform 1 0 6348 0 -1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_45
timestamp 1608910539
transform 1 0 5244 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_56
timestamp 1608910539
transform 1 0 6256 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_44
timestamp 1608910539
transform 1 0 5152 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1608910539
transform 1 0 6716 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_70
timestamp 1608910539
transform 1 0 7544 0 -1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_75
timestamp 1608910539
transform 1 0 8004 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_68
timestamp 1608910539
transform 1 0 7360 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_right_track_0.prog_clk
timestamp 1608910539
transform 1 0 7728 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 7728 0 -1 13456
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_20_92
timestamp 1608910539
transform 1 0 9568 0 -1 13456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_88
timestamp 1608910539
transform 1 0 9200 0 -1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_93
timestamp 1608910539
transform 1 0 9660 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_91
timestamp 1608910539
transform 1 0 9476 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_87
timestamp 1608910539
transform 1 0 9108 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9384 0 -1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1608910539
transform 1 0 9568 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_98
timestamp 1608910539
transform 1 0 10120 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1608910539
transform 1 0 9936 0 1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_right_track_0.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 10212 0 -1 13456
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_20_123
timestamp 1608910539
transform 1 0 12420 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_119
timestamp 1608910539
transform 1 0 12052 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_123
timestamp 1608910539
transform 1 0 12420 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_105
timestamp 1608910539
transform 1 0 10764 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1608910539
transform 1 0 12328 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1608910539
transform 1 0 12512 0 -1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 10948 0 1 12368
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1608910539
transform 1 0 12604 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_133
timestamp 1608910539
transform 1 0 13340 0 -1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_133
timestamp 1608910539
transform 1 0 13340 0 1 12368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_128
timestamp 1608910539
transform 1 0 12880 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 13524 0 -1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_right_track_0.prog_clk
timestamp 1608910539
transform 1 0 13064 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_137
timestamp 1608910539
transform 1 0 13708 0 -1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_143
timestamp 1608910539
transform 1 0 14260 0 1 12368
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 13892 0 -1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 14076 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1608910539
transform 1 0 14076 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_165
timestamp 1608910539
transform 1 0 16284 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_159
timestamp 1608910539
transform 1 0 15732 0 -1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_153
timestamp 1608910539
transform 1 0 15180 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_154
timestamp 1608910539
transform 1 0 15272 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_151
timestamp 1608910539
transform 1 0 14996 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 16100 0 -1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1608910539
transform 1 0 15180 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 15640 0 1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1608910539
transform 1 0 15456 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_171
timestamp 1608910539
transform 1 0 16836 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_167
timestamp 1608910539
transform 1 0 16468 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 16652 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1608910539
transform 1 0 17020 0 1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_184
timestamp 1608910539
transform 1 0 18032 0 -1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_177
timestamp 1608910539
transform 1 0 17388 0 -1 13456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_186
timestamp 1608910539
transform 1 0 18216 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_182
timestamp 1608910539
transform 1 0 17848 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 18032 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1608910539
transform 1 0 17940 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1608910539
transform 1 0 19228 0 -1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_196
timestamp 1608910539
transform 1 0 19136 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_190
timestamp 1608910539
transform 1 0 18584 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 18400 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 18952 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1608910539
transform 1 0 18400 0 -1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_207
timestamp 1608910539
transform 1 0 20148 0 -1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_202
timestamp 1608910539
transform 1 0 19688 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_206
timestamp 1608910539
transform 1 0 20056 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_200
timestamp 1608910539
transform 1 0 19504 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__85__A
timestamp 1608910539
transform 1 0 19320 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__84__A
timestamp 1608910539
transform 1 0 19964 0 -1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _85_
timestamp 1608910539
transform 1 0 19688 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1608910539
transform 1 0 19412 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1608910539
transform 1 0 20240 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_213
timestamp 1608910539
transform 1 0 20700 0 -1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_212
timestamp 1608910539
transform 1 0 20608 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1608910539
transform 1 0 20332 0 -1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1608910539
transform 1 0 20792 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _84_
timestamp 1608910539
transform 1 0 20884 0 -1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1608910539
transform 1 0 20884 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_219
timestamp 1608910539
transform 1 0 21252 0 -1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_219
timestamp 1608910539
transform 1 0 21252 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608910539
transform -1 0 21896 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608910539
transform -1 0 21896 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1608910539
transform 1 0 2484 0 1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1608910539
transform 1 0 1380 0 1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608910539
transform 1 0 1104 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1608910539
transform 1 0 4692 0 1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_36
timestamp 1608910539
transform 1 0 4416 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_32
timestamp 1608910539
transform 1 0 4048 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_27
timestamp 1608910539
transform 1 0 3588 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 4508 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1608910539
transform 1 0 3956 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 5796 0 1 13456
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_77
timestamp 1608910539
transform 1 0 8188 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_67
timestamp 1608910539
transform 1 0 7268 0 1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8004 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8372 0 1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_21_93
timestamp 1608910539
transform 1 0 9660 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_88
timestamp 1608910539
transform 1 0 9200 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1608910539
transform 1 0 9568 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 9936 0 1 13456
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_21_120
timestamp 1608910539
transform 1 0 12144 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_112
timestamp 1608910539
transform 1 0 11408 0 1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 12236 0 1 13456
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_137
timestamp 1608910539
transform 1 0 13708 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1608910539
transform 1 0 13892 0 1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_163
timestamp 1608910539
transform 1 0 16100 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_152
timestamp 1608910539
transform 1 0 15088 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_148
timestamp 1608910539
transform 1 0 14720 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1608910539
transform 1 0 15180 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 16284 0 1 13456
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1608910539
transform 1 0 15272 0 1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_175
timestamp 1608910539
transform 1 0 17204 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_171
timestamp 1608910539
transform 1 0 16836 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 17296 0 1 13456
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_21_207
timestamp 1608910539
transform 1 0 20148 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_203
timestamp 1608910539
transform 1 0 19780 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_192
timestamp 1608910539
transform 1 0 18768 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1608910539
transform 1 0 18952 0 1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _86_
timestamp 1608910539
transform 1 0 20240 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_219
timestamp 1608910539
transform 1 0 21252 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_212
timestamp 1608910539
transform 1 0 20608 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1608910539
transform 1 0 20792 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608910539
transform -1 0 21896 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1608910539
transform 1 0 20884 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_15
timestamp 1608910539
transform 1 0 2484 0 -1 14544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1608910539
transform 1 0 1380 0 -1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608910539
transform 1 0 1104 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_37
timestamp 1608910539
transform 1 0 4508 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1608910539
transform 1 0 4692 0 -1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 3036 0 -1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_22_60
timestamp 1608910539
transform 1 0 6624 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_52
timestamp 1608910539
transform 1 0 5888 0 -1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_48
timestamp 1608910539
transform 1 0 5520 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 5704 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1608910539
transform 1 0 6716 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 6808 0 -1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1608910539
transform 1 0 8648 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_78
timestamp 1608910539
transform 1 0 8280 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8464 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_101
timestamp 1608910539
transform 1 0 10396 0 -1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_93
timestamp 1608910539
transform 1 0 9660 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 9844 0 -1 14544
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8832 0 -1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_120
timestamp 1608910539
transform 1 0 12144 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_117
timestamp 1608910539
transform 1 0 11868 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_113
timestamp 1608910539
transform 1 0 11500 0 -1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 11960 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1608910539
transform 1 0 12328 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1608910539
transform 1 0 12420 0 -1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1608910539
transform 1 0 13800 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_132
timestamp 1608910539
transform 1 0 13248 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_right_track_0.prog_clk
timestamp 1608910539
transform 1 0 13524 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 13984 0 -1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_156
timestamp 1608910539
transform 1 0 15456 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1608910539
transform 1 0 15640 0 -1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_181
timestamp 1608910539
transform 1 0 17756 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_167
timestamp 1608910539
transform 1 0 16468 0 -1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 17572 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1608910539
transform 1 0 17940 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1608910539
transform 1 0 18032 0 -1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_203
timestamp 1608910539
transform 1 0 19780 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_197
timestamp 1608910539
transform 1 0 19228 0 -1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_193
timestamp 1608910539
transform 1 0 18860 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 19044 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__86__A
timestamp 1608910539
transform 1 0 19596 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 19964 0 -1 14544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_222
timestamp 1608910539
transform 1 0 21528 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_218
timestamp 1608910539
transform 1 0 21160 0 -1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_211
timestamp 1608910539
transform 1 0 20516 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608910539
transform -1 0 21896 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1608910539
transform 1 0 20792 0 -1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1608910539
transform 1 0 2484 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1608910539
transform 1 0 1380 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1608910539
transform 1 0 1104 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_32
timestamp 1608910539
transform 1 0 4048 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_27
timestamp 1608910539
transform 1 0 3588 0 1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1608910539
transform 1 0 3956 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1608910539
transform 1 0 4140 0 1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_23_59
timestamp 1608910539
transform 1 0 6532 0 1 14544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_47
timestamp 1608910539
transform 1 0 5428 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_42
timestamp 1608910539
transform 1 0 4968 0 1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1608910539
transform 1 0 5152 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_79
timestamp 1608910539
transform 1 0 8372 0 1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_74
timestamp 1608910539
transform 1 0 7912 0 1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_right_track_0.prog_clk
timestamp 1608910539
transform 1 0 8556 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1608910539
transform 1 0 7084 0 1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1608910539
transform 1 0 8096 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1608910539
transform 1 0 9660 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_84
timestamp 1608910539
transform 1 0 8832 0 1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1608910539
transform 1 0 9568 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_117
timestamp 1608910539
transform 1 0 11868 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_105
timestamp 1608910539
transform 1 0 10764 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_134
timestamp 1608910539
transform 1 0 13432 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_129
timestamp 1608910539
transform 1 0 12972 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 13248 0 1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_166
timestamp 1608910539
transform 1 0 16376 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_154
timestamp 1608910539
transform 1 0 15272 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_152
timestamp 1608910539
transform 1 0 15088 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_146
timestamp 1608910539
transform 1 0 14536 0 1 14544
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1608910539
transform 1 0 15180 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_178
timestamp 1608910539
transform 1 0 17480 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_202
timestamp 1608910539
transform 1 0 19688 0 1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_190
timestamp 1608910539
transform 1 0 18584 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 19872 0 1 14544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_219
timestamp 1608910539
transform 1 0 21252 0 1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_210
timestamp 1608910539
transform 1 0 20424 0 1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1608910539
transform 1 0 20792 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1608910539
transform -1 0 21896 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1608910539
transform 1 0 20884 0 1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1608910539
transform 1 0 1380 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1608910539
transform 1 0 1104 0 -1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 1748 0 -1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_24_35
timestamp 1608910539
transform 1 0 4324 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_23
timestamp 1608910539
transform 1 0 3220 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_62
timestamp 1608910539
transform 1 0 6808 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_59
timestamp 1608910539
transform 1 0 6532 0 -1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_47
timestamp 1608910539
transform 1 0 5428 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1608910539
transform 1 0 6716 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_79
timestamp 1608910539
transform 1 0 8372 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_75
timestamp 1608910539
transform 1 0 8004 0 -1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8188 0 -1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1608910539
transform 1 0 7176 0 -1 15632
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_24_103
timestamp 1608910539
transform 1 0 10580 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_91
timestamp 1608910539
transform 1 0 9476 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_123
timestamp 1608910539
transform 1 0 12420 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_121
timestamp 1608910539
transform 1 0 12236 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_115
timestamp 1608910539
transform 1 0 11684 0 -1 15632
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1608910539
transform 1 0 12328 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_135
timestamp 1608910539
transform 1 0 13524 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_159
timestamp 1608910539
transform 1 0 15732 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_147
timestamp 1608910539
transform 1 0 14628 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_171
timestamp 1608910539
transform 1 0 16836 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1608910539
transform 1 0 17940 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 18032 0 -1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_24_200
timestamp 1608910539
transform 1 0 19504 0 -1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 19780 0 -1 15632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_222
timestamp 1608910539
transform 1 0 21528 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_218
timestamp 1608910539
transform 1 0 21160 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_213
timestamp 1608910539
transform 1 0 20700 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_209
timestamp 1608910539
transform 1 0 20332 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1608910539
transform -1 0 21896 0 -1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1608910539
transform 1 0 20792 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_15
timestamp 1608910539
transform 1 0 2484 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1608910539
transform 1 0 1380 0 1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1608910539
transform 1 0 1104 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1608910539
transform 1 0 2760 0 1 15632
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_25_35
timestamp 1608910539
transform 1 0 4324 0 1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_32
timestamp 1608910539
transform 1 0 4048 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_27
timestamp 1608910539
transform 1 0 3588 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 4140 0 1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1608910539
transform 1 0 3956 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_60
timestamp 1608910539
transform 1 0 6624 0 1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_43
timestamp 1608910539
transform 1 0 5060 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 5152 0 1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_25_74
timestamp 1608910539
transform 1 0 7912 0 1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_68
timestamp 1608910539
transform 1 0 7360 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_right_track_0.prog_clk
timestamp 1608910539
transform 1 0 7636 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 8648 0 1 15632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_25_93
timestamp 1608910539
transform 1 0 9660 0 1 15632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_88
timestamp 1608910539
transform 1 0 9200 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1608910539
transform 1 0 9568 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 10212 0 1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_115
timestamp 1608910539
transform 1 0 11684 0 1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 11868 0 1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_133
timestamp 1608910539
transform 1 0 13340 0 1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 13524 0 1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_151
timestamp 1608910539
transform 1 0 14996 0 1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1608910539
transform 1 0 15180 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15272 0 1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_170
timestamp 1608910539
transform 1 0 16744 0 1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 16928 0 1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_25_205
timestamp 1608910539
transform 1 0 19964 0 1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_193
timestamp 1608910539
transform 1 0 18860 0 1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_188
timestamp 1608910539
transform 1 0 18400 0 1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1608910539
transform 1 0 18584 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_219
timestamp 1608910539
transform 1 0 21252 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_213
timestamp 1608910539
transform 1 0 20700 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1608910539
transform 1 0 20792 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1608910539
transform -1 0 21896 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1608910539
transform 1 0 20884 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1608910539
transform 1 0 1380 0 1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_15
timestamp 1608910539
transform 1 0 2484 0 -1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1608910539
transform 1 0 1380 0 -1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1608910539
transform 1 0 1104 0 1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1608910539
transform 1 0 1104 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 1748 0 1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_27_28
timestamp 1608910539
transform 1 0 3680 0 1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_23
timestamp 1608910539
transform 1 0 3220 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_31
timestamp 1608910539
transform 1 0 3956 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_21
timestamp 1608910539
transform 1 0 3036 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1608910539
transform 1 0 3956 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1608910539
transform 1 0 3128 0 -1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1608910539
transform 1 0 3404 0 1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_38
timestamp 1608910539
transform 1 0 4600 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_32
timestamp 1608910539
transform 1 0 4048 0 1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_35
timestamp 1608910539
transform 1 0 4324 0 -1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 4140 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 4692 0 -1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1608910539
transform 1 0 4324 0 1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4784 0 1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_27_60
timestamp 1608910539
transform 1 0 6624 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_56
timestamp 1608910539
transform 1 0 6256 0 1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_57
timestamp 1608910539
transform 1 0 6348 0 -1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_45
timestamp 1608910539
transform 1 0 5244 0 -1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 6716 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1608910539
transform 1 0 6716 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 6808 0 -1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_27_74
timestamp 1608910539
transform 1 0 7912 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_63
timestamp 1608910539
transform 1 0 6900 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_82
timestamp 1608910539
transform 1 0 8648 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_78
timestamp 1608910539
transform 1 0 8280 0 -1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8096 0 1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1608910539
transform 1 0 7084 0 1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 8740 0 -1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_27_93
timestamp 1608910539
transform 1 0 9660 0 1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_90
timestamp 1608910539
transform 1 0 9384 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_85
timestamp 1608910539
transform 1 0 8924 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1608910539
transform 1 0 9568 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _40_
timestamp 1608910539
transform 1 0 9108 0 1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_102
timestamp 1608910539
transform 1 0 10488 0 1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_99
timestamp 1608910539
transform 1 0 10212 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_99
timestamp 1608910539
transform 1 0 10212 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 10304 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10488 0 -1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1608910539
transform 1 0 11224 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_111
timestamp 1608910539
transform 1 0 11316 0 -1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 11040 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1608910539
transform 1 0 11408 0 1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_123
timestamp 1608910539
transform 1 0 12420 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_119
timestamp 1608910539
transform 1 0 12052 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_115
timestamp 1608910539
transform 1 0 11684 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 12604 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1608910539
transform 1 0 12328 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _41_
timestamp 1608910539
transform 1 0 11776 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_121
timestamp 1608910539
transform 1 0 12236 0 1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_145
timestamp 1608910539
transform 1 0 14444 0 1 16720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_133
timestamp 1608910539
transform 1 0 13340 0 1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_142
timestamp 1608910539
transform 1 0 14168 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1608910539
transform 1 0 13800 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_127
timestamp 1608910539
transform 1 0 12788 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 13984 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1608910539
transform 1 0 14352 0 -1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1608910539
transform 1 0 12972 0 -1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_27_161
timestamp 1608910539
transform 1 0 15916 0 1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_158
timestamp 1608910539
transform 1 0 15640 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_154
timestamp 1608910539
transform 1 0 15272 0 1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_158
timestamp 1608910539
transform 1 0 15640 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_153
timestamp 1608910539
transform 1 0 15180 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 15732 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1608910539
transform 1 0 15180 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1608910539
transform 1 0 15916 0 -1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1608910539
transform 1 0 15364 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_185
timestamp 1608910539
transform 1 0 18124 0 1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_173
timestamp 1608910539
transform 1 0 17020 0 1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_182
timestamp 1608910539
transform 1 0 17848 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_174
timestamp 1608910539
transform 1 0 17112 0 -1 16720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_170
timestamp 1608910539
transform 1 0 16744 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 16928 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1608910539
transform 1 0 17940 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1608910539
transform 1 0 18032 0 -1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_27_202
timestamp 1608910539
transform 1 0 19688 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_196
timestamp 1608910539
transform 1 0 19136 0 1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_189
timestamp 1608910539
transform 1 0 18492 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_208
timestamp 1608910539
transform 1 0 20240 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_201
timestamp 1608910539
transform 1 0 19596 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_193
timestamp 1608910539
transform 1 0 18860 0 -1 16720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 18584 0 1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 19780 0 1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 19688 0 -1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_213
timestamp 1608910539
transform 1 0 20700 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_209
timestamp 1608910539
transform 1 0 20332 0 1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1608910539
transform 1 0 20792 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 20424 0 -1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1608910539
transform 1 0 20884 0 1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_219
timestamp 1608910539
transform 1 0 21252 0 1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_222
timestamp 1608910539
transform 1 0 21528 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_216
timestamp 1608910539
transform 1 0 20976 0 -1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1608910539
transform -1 0 21896 0 1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1608910539
transform -1 0 21896 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1608910539
transform 1 0 2484 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1608910539
transform 1 0 1380 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1608910539
transform 1 0 1104 0 -1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_33
timestamp 1608910539
transform 1 0 4140 0 -1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_27
timestamp 1608910539
transform 1 0 3588 0 -1 17808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1608910539
transform 1 0 4232 0 -1 17808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_28_62
timestamp 1608910539
transform 1 0 6808 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_55
timestamp 1608910539
transform 1 0 6164 0 -1 17808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_43
timestamp 1608910539
transform 1 0 5060 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1608910539
transform 1 0 6716 0 -1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_76
timestamp 1608910539
transform 1 0 8096 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 7912 0 -1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_104
timestamp 1608910539
transform 1 0 10672 0 -1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_93
timestamp 1608910539
transform 1 0 9660 0 -1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_88
timestamp 1608910539
transform 1 0 9200 0 -1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9476 0 -1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1608910539
transform 1 0 9844 0 -1 17808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_28_123
timestamp 1608910539
transform 1 0 12420 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_120
timestamp 1608910539
transform 1 0 12144 0 -1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_108
timestamp 1608910539
transform 1 0 11040 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 10856 0 -1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1608910539
transform 1 0 12328 0 -1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_135
timestamp 1608910539
transform 1 0 13524 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_159
timestamp 1608910539
transform 1 0 15732 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_147
timestamp 1608910539
transform 1 0 14628 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_184
timestamp 1608910539
transform 1 0 18032 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_171
timestamp 1608910539
transform 1 0 16836 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1608910539
transform 1 0 17940 0 -1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_202
timestamp 1608910539
transform 1 0 19688 0 -1 17808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_196
timestamp 1608910539
transform 1 0 19136 0 -1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1608910539
transform 1 0 19320 0 -1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1608910539
transform 1 0 20240 0 -1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_222
timestamp 1608910539
transform 1 0 21528 0 -1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_218
timestamp 1608910539
transform 1 0 21160 0 -1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_212
timestamp 1608910539
transform 1 0 20608 0 -1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1608910539
transform -1 0 21896 0 -1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1608910539
transform 1 0 20792 0 -1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1608910539
transform 1 0 2484 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1608910539
transform 1 0 1380 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1608910539
transform 1 0 1104 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_32
timestamp 1608910539
transform 1 0 4048 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_27
timestamp 1608910539
transform 1 0 3588 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1608910539
transform 1 0 3956 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_56
timestamp 1608910539
transform 1 0 6256 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_44
timestamp 1608910539
transform 1 0 5152 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1608910539
transform 1 0 6624 0 1 17808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_29_77
timestamp 1608910539
transform 1 0 8188 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_73
timestamp 1608910539
transform 1 0 7820 0 1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_69
timestamp 1608910539
transform 1 0 7452 0 1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8004 0 1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 7636 0 1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_89
timestamp 1608910539
transform 1 0 9292 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1608910539
transform 1 0 9568 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 9660 0 1 17808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_29_125
timestamp 1608910539
transform 1 0 12604 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1608910539
transform 1 0 12144 0 1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_109
timestamp 1608910539
transform 1 0 11132 0 1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1608910539
transform 1 0 11316 0 1 17808
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1608910539
transform 1 0 12328 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_143
timestamp 1608910539
transform 1 0 14260 0 1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_132
timestamp 1608910539
transform 1 0 13248 0 1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_129
timestamp 1608910539
transform 1 0 12972 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 13064 0 1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1608910539
transform 1 0 13432 0 1 17808
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1608910539
transform 1 0 14444 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_154
timestamp 1608910539
transform 1 0 15272 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_152
timestamp 1608910539
transform 1 0 15088 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_148
timestamp 1608910539
transform 1 0 14720 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1608910539
transform 1 0 15180 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15548 0 1 17808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_29_173
timestamp 1608910539
transform 1 0 17020 0 1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 17204 0 1 17808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_29_200
timestamp 1608910539
transform 1 0 19504 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_196
timestamp 1608910539
transform 1 0 19136 0 1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_191
timestamp 1608910539
transform 1 0 18676 0 1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l2_in_0__S
timestamp 1608910539
transform 1 0 19320 0 1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1608910539
transform 1 0 18860 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_219
timestamp 1608910539
transform 1 0 21252 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_212
timestamp 1608910539
transform 1 0 20608 0 1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1608910539
transform 1 0 20792 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1608910539
transform -1 0 21896 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1608910539
transform 1 0 20884 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_11
timestamp 1608910539
transform 1 0 2116 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1608910539
transform 1 0 1380 0 -1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1608910539
transform 1 0 1104 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 2392 0 -1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_41
timestamp 1608910539
transform 1 0 4876 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_30
timestamp 1608910539
transform 1 0 3864 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1608910539
transform 1 0 4048 0 -1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_59
timestamp 1608910539
transform 1 0 6532 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_55
timestamp 1608910539
transform 1 0 6164 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_49
timestamp 1608910539
transform 1 0 5612 0 -1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_45
timestamp 1608910539
transform 1 0 5244 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 5428 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 5060 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1608910539
transform 1 0 6716 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1608910539
transform 1 0 6808 0 -1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1608910539
transform 1 0 6256 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_83
timestamp 1608910539
transform 1 0 8740 0 -1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_71
timestamp 1608910539
transform 1 0 7636 0 -1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_98
timestamp 1608910539
transform 1 0 10120 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_94
timestamp 1608910539
transform 1 0 9752 0 -1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1608910539
transform 1 0 9384 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_87
timestamp 1608910539
transform 1 0 9108 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9568 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9200 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 10212 0 -1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_120
timestamp 1608910539
transform 1 0 12144 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_115
timestamp 1608910539
transform 1 0 11684 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 11960 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1608910539
transform 1 0 12328 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1608910539
transform 1 0 12420 0 -1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_30_132
timestamp 1608910539
transform 1 0 13248 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 13524 0 -1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_165
timestamp 1608910539
transform 1 0 16284 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_151
timestamp 1608910539
transform 1 0 14996 0 -1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 16100 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_180
timestamp 1608910539
transform 1 0 17664 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_176
timestamp 1608910539
transform 1 0 17296 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 17480 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1608910539
transform 1 0 17940 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l2_in_0_
timestamp 1608910539
transform 1 0 18032 0 -1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l1_in_0_
timestamp 1608910539
transform 1 0 16468 0 -1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_202
timestamp 1608910539
transform 1 0 19688 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_193
timestamp 1608910539
transform 1 0 18860 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 19136 0 -1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 19872 0 -1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_222
timestamp 1608910539
transform 1 0 21528 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_218
timestamp 1608910539
transform 1 0 21160 0 -1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_210
timestamp 1608910539
transform 1 0 20424 0 -1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1608910539
transform -1 0 21896 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1608910539
transform 1 0 20792 0 -1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1608910539
transform 1 0 2484 0 1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1608910539
transform 1 0 1380 0 1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1608910539
transform 1 0 1104 0 1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_27
timestamp 1608910539
transform 1 0 3588 0 1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1608910539
transform 1 0 3956 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 4048 0 1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_31_54
timestamp 1608910539
transform 1 0 6072 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_48
timestamp 1608910539
transform 1 0 5520 0 1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 6164 0 1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_31_71
timestamp 1608910539
transform 1 0 7636 0 1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8372 0 1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_31_102
timestamp 1608910539
transform 1 0 10488 0 1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_88
timestamp 1608910539
transform 1 0 9200 0 1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1608910539
transform 1 0 9568 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1608910539
transform 1 0 9660 0 1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_124
timestamp 1608910539
transform 1 0 12512 0 1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 11040 0 1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_31_142
timestamp 1608910539
transform 1 0 14168 0 1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 12696 0 1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_31_150
timestamp 1608910539
transform 1 0 14904 0 1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1608910539
transform 1 0 15180 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 15272 0 1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_31_185
timestamp 1608910539
transform 1 0 18124 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_179
timestamp 1608910539
transform 1 0 17572 0 1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_31_170
timestamp 1608910539
transform 1 0 16744 0 1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 18216 0 1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 17020 0 1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_206
timestamp 1608910539
transform 1 0 20056 0 1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_198
timestamp 1608910539
transform 1 0 19320 0 1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 19504 0 1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1608910539
transform 1 0 20240 0 1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_219
timestamp 1608910539
transform 1 0 21252 0 1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_212
timestamp 1608910539
transform 1 0 20608 0 1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1608910539
transform 1 0 20792 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1608910539
transform -1 0 21896 0 1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1608910539
transform 1 0 20884 0 1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1608910539
transform 1 0 2484 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1608910539
transform 1 0 1380 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1608910539
transform 1 0 1104 0 -1 19984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_39
timestamp 1608910539
transform 1 0 4692 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_27
timestamp 1608910539
transform 1 0 3588 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 4784 0 -1 19984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_32_60
timestamp 1608910539
transform 1 0 6624 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_56
timestamp 1608910539
transform 1 0 6256 0 -1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1608910539
transform 1 0 6716 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 6808 0 -1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_74
timestamp 1608910539
transform 1 0 7912 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_68
timestamp 1608910539
transform 1 0 7360 0 -1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 8004 0 -1 19984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_32_96
timestamp 1608910539
transform 1 0 9936 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_91
timestamp 1608910539
transform 1 0 9476 0 -1 19984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1608910539
transform 1 0 9660 0 -1 19984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_123
timestamp 1608910539
transform 1 0 12420 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_120
timestamp 1608910539
transform 1 0 12144 0 -1 19984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_108
timestamp 1608910539
transform 1 0 11040 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1608910539
transform 1 0 12328 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_142
timestamp 1608910539
transform 1 0 14168 0 -1 19984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1608910539
transform 1 0 13892 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_135
timestamp 1608910539
transform 1 0 13524 0 -1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 13984 0 -1 19984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1608910539
transform 1 0 14352 0 -1 19984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_32_161
timestamp 1608910539
transform 1 0 15916 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_157
timestamp 1608910539
transform 1 0 15548 0 -1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_153
timestamp 1608910539
transform 1 0 15180 0 -1 19984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 15364 0 -1 19984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1608910539
transform 1 0 16008 0 -1 19984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_32_182
timestamp 1608910539
transform 1 0 17848 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_176
timestamp 1608910539
transform 1 0 17296 0 -1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_171
timestamp 1608910539
transform 1 0 16836 0 -1 19984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1608910539
transform 1 0 17940 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1608910539
transform 1 0 18032 0 -1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1608910539
transform 1 0 17020 0 -1 19984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_200
timestamp 1608910539
transform 1 0 19504 0 -1 19984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_196
timestamp 1608910539
transform 1 0 19136 0 -1 19984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_188
timestamp 1608910539
transform 1 0 18400 0 -1 19984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1608910539
transform 1 0 19320 0 -1 19984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 19780 0 -1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_222
timestamp 1608910539
transform 1 0 21528 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_218
timestamp 1608910539
transform 1 0 21160 0 -1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_213
timestamp 1608910539
transform 1 0 20700 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_209
timestamp 1608910539
transform 1 0 20332 0 -1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1608910539
transform -1 0 21896 0 -1 19984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1608910539
transform 1 0 20792 0 -1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1608910539
transform 1 0 2484 0 1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1608910539
transform 1 0 1380 0 1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1608910539
transform 1 0 1104 0 1 19984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_32
timestamp 1608910539
transform 1 0 4048 0 1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_27
timestamp 1608910539
transform 1 0 3588 0 1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1608910539
transform 1 0 3956 0 1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_56
timestamp 1608910539
transform 1 0 6256 0 1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_44
timestamp 1608910539
transform 1 0 5152 0 1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1608910539
transform 1 0 6808 0 1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_75
timestamp 1608910539
transform 1 0 8004 0 1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_63
timestamp 1608910539
transform 1 0 6900 0 1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_94
timestamp 1608910539
transform 1 0 9752 0 1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_87
timestamp 1608910539
transform 1 0 9108 0 1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1608910539
transform 1 0 9660 0 1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_125
timestamp 1608910539
transform 1 0 12604 0 1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_118
timestamp 1608910539
transform 1 0 11960 0 1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_106
timestamp 1608910539
transform 1 0 10856 0 1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1608910539
transform 1 0 12512 0 1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_137
timestamp 1608910539
transform 1 0 13708 0 1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_156
timestamp 1608910539
transform 1 0 15456 0 1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_149
timestamp 1608910539
transform 1 0 14812 0 1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1608910539
transform 1 0 15364 0 1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_187
timestamp 1608910539
transform 1 0 18308 0 1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_180
timestamp 1608910539
transform 1 0 17664 0 1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_168
timestamp 1608910539
transform 1 0 16560 0 1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1608910539
transform 1 0 18216 0 1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_199
timestamp 1608910539
transform 1 0 19412 0 1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1608910539
transform 1 0 19964 0 1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_222
timestamp 1608910539
transform 1 0 21528 0 1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_218
timestamp 1608910539
transform 1 0 21160 0 1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_215
timestamp 1608910539
transform 1 0 20884 0 1 19984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_209
timestamp 1608910539
transform 1 0 20332 0 1 19984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1608910539
transform 1 0 21068 0 1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1608910539
transform -1 0 21896 0 1 19984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1608910539
transform 1 0 20516 0 1 19984
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 5576 800 5696 6 ccff_head
port 0 nsew signal input
rlabel metal3 s 0 17000 800 17120 6 ccff_tail
port 1 nsew signal tristate
rlabel metal3 s 22200 4080 23000 4200 6 chanx_right_in[0]
port 2 nsew signal input
rlabel metal3 s 22200 8704 23000 8824 6 chanx_right_in[10]
port 3 nsew signal input
rlabel metal3 s 22200 9112 23000 9232 6 chanx_right_in[11]
port 4 nsew signal input
rlabel metal3 s 22200 9520 23000 9640 6 chanx_right_in[12]
port 5 nsew signal input
rlabel metal3 s 22200 10064 23000 10184 6 chanx_right_in[13]
port 6 nsew signal input
rlabel metal3 s 22200 10472 23000 10592 6 chanx_right_in[14]
port 7 nsew signal input
rlabel metal3 s 22200 11016 23000 11136 6 chanx_right_in[15]
port 8 nsew signal input
rlabel metal3 s 22200 11424 23000 11544 6 chanx_right_in[16]
port 9 nsew signal input
rlabel metal3 s 22200 11832 23000 11952 6 chanx_right_in[17]
port 10 nsew signal input
rlabel metal3 s 22200 12376 23000 12496 6 chanx_right_in[18]
port 11 nsew signal input
rlabel metal3 s 22200 12784 23000 12904 6 chanx_right_in[19]
port 12 nsew signal input
rlabel metal3 s 22200 4488 23000 4608 6 chanx_right_in[1]
port 13 nsew signal input
rlabel metal3 s 22200 5032 23000 5152 6 chanx_right_in[2]
port 14 nsew signal input
rlabel metal3 s 22200 5440 23000 5560 6 chanx_right_in[3]
port 15 nsew signal input
rlabel metal3 s 22200 5848 23000 5968 6 chanx_right_in[4]
port 16 nsew signal input
rlabel metal3 s 22200 6392 23000 6512 6 chanx_right_in[5]
port 17 nsew signal input
rlabel metal3 s 22200 6800 23000 6920 6 chanx_right_in[6]
port 18 nsew signal input
rlabel metal3 s 22200 7344 23000 7464 6 chanx_right_in[7]
port 19 nsew signal input
rlabel metal3 s 22200 7752 23000 7872 6 chanx_right_in[8]
port 20 nsew signal input
rlabel metal3 s 22200 8160 23000 8280 6 chanx_right_in[9]
port 21 nsew signal input
rlabel metal3 s 22200 13328 23000 13448 6 chanx_right_out[0]
port 22 nsew signal tristate
rlabel metal3 s 22200 17816 23000 17936 6 chanx_right_out[10]
port 23 nsew signal tristate
rlabel metal3 s 22200 18360 23000 18480 6 chanx_right_out[11]
port 24 nsew signal tristate
rlabel metal3 s 22200 18768 23000 18888 6 chanx_right_out[12]
port 25 nsew signal tristate
rlabel metal3 s 22200 19176 23000 19296 6 chanx_right_out[13]
port 26 nsew signal tristate
rlabel metal3 s 22200 19720 23000 19840 6 chanx_right_out[14]
port 27 nsew signal tristate
rlabel metal3 s 22200 20128 23000 20248 6 chanx_right_out[15]
port 28 nsew signal tristate
rlabel metal3 s 22200 20672 23000 20792 6 chanx_right_out[16]
port 29 nsew signal tristate
rlabel metal3 s 22200 21080 23000 21200 6 chanx_right_out[17]
port 30 nsew signal tristate
rlabel metal3 s 22200 21488 23000 21608 6 chanx_right_out[18]
port 31 nsew signal tristate
rlabel metal3 s 22200 22032 23000 22152 6 chanx_right_out[19]
port 32 nsew signal tristate
rlabel metal3 s 22200 13736 23000 13856 6 chanx_right_out[1]
port 33 nsew signal tristate
rlabel metal3 s 22200 14144 23000 14264 6 chanx_right_out[2]
port 34 nsew signal tristate
rlabel metal3 s 22200 14688 23000 14808 6 chanx_right_out[3]
port 35 nsew signal tristate
rlabel metal3 s 22200 15096 23000 15216 6 chanx_right_out[4]
port 36 nsew signal tristate
rlabel metal3 s 22200 15504 23000 15624 6 chanx_right_out[5]
port 37 nsew signal tristate
rlabel metal3 s 22200 16048 23000 16168 6 chanx_right_out[6]
port 38 nsew signal tristate
rlabel metal3 s 22200 16456 23000 16576 6 chanx_right_out[7]
port 39 nsew signal tristate
rlabel metal3 s 22200 17000 23000 17120 6 chanx_right_out[8]
port 40 nsew signal tristate
rlabel metal3 s 22200 17408 23000 17528 6 chanx_right_out[9]
port 41 nsew signal tristate
rlabel metal2 s 846 22056 902 22856 6 chany_top_in[0]
port 42 nsew signal input
rlabel metal2 s 6458 22056 6514 22856 6 chany_top_in[10]
port 43 nsew signal input
rlabel metal2 s 7010 22056 7066 22856 6 chany_top_in[11]
port 44 nsew signal input
rlabel metal2 s 7562 22056 7618 22856 6 chany_top_in[12]
port 45 nsew signal input
rlabel metal2 s 8114 22056 8170 22856 6 chany_top_in[13]
port 46 nsew signal input
rlabel metal2 s 8666 22056 8722 22856 6 chany_top_in[14]
port 47 nsew signal input
rlabel metal2 s 9218 22056 9274 22856 6 chany_top_in[15]
port 48 nsew signal input
rlabel metal2 s 9770 22056 9826 22856 6 chany_top_in[16]
port 49 nsew signal input
rlabel metal2 s 10322 22056 10378 22856 6 chany_top_in[17]
port 50 nsew signal input
rlabel metal2 s 10874 22056 10930 22856 6 chany_top_in[18]
port 51 nsew signal input
rlabel metal2 s 11426 22056 11482 22856 6 chany_top_in[19]
port 52 nsew signal input
rlabel metal2 s 1398 22056 1454 22856 6 chany_top_in[1]
port 53 nsew signal input
rlabel metal2 s 1950 22056 2006 22856 6 chany_top_in[2]
port 54 nsew signal input
rlabel metal2 s 2502 22056 2558 22856 6 chany_top_in[3]
port 55 nsew signal input
rlabel metal2 s 3054 22056 3110 22856 6 chany_top_in[4]
port 56 nsew signal input
rlabel metal2 s 3606 22056 3662 22856 6 chany_top_in[5]
port 57 nsew signal input
rlabel metal2 s 4158 22056 4214 22856 6 chany_top_in[6]
port 58 nsew signal input
rlabel metal2 s 4710 22056 4766 22856 6 chany_top_in[7]
port 59 nsew signal input
rlabel metal2 s 5262 22056 5318 22856 6 chany_top_in[8]
port 60 nsew signal input
rlabel metal2 s 5814 22056 5870 22856 6 chany_top_in[9]
port 61 nsew signal input
rlabel metal2 s 12070 22056 12126 22856 6 chany_top_out[0]
port 62 nsew signal tristate
rlabel metal2 s 17682 22056 17738 22856 6 chany_top_out[10]
port 63 nsew signal tristate
rlabel metal2 s 18234 22056 18290 22856 6 chany_top_out[11]
port 64 nsew signal tristate
rlabel metal2 s 18786 22056 18842 22856 6 chany_top_out[12]
port 65 nsew signal tristate
rlabel metal2 s 19338 22056 19394 22856 6 chany_top_out[13]
port 66 nsew signal tristate
rlabel metal2 s 19890 22056 19946 22856 6 chany_top_out[14]
port 67 nsew signal tristate
rlabel metal2 s 20442 22056 20498 22856 6 chany_top_out[15]
port 68 nsew signal tristate
rlabel metal2 s 20994 22056 21050 22856 6 chany_top_out[16]
port 69 nsew signal tristate
rlabel metal2 s 21546 22056 21602 22856 6 chany_top_out[17]
port 70 nsew signal tristate
rlabel metal2 s 22098 22056 22154 22856 6 chany_top_out[18]
port 71 nsew signal tristate
rlabel metal2 s 22650 22056 22706 22856 6 chany_top_out[19]
port 72 nsew signal tristate
rlabel metal2 s 12622 22056 12678 22856 6 chany_top_out[1]
port 73 nsew signal tristate
rlabel metal2 s 13174 22056 13230 22856 6 chany_top_out[2]
port 74 nsew signal tristate
rlabel metal2 s 13726 22056 13782 22856 6 chany_top_out[3]
port 75 nsew signal tristate
rlabel metal2 s 14278 22056 14334 22856 6 chany_top_out[4]
port 76 nsew signal tristate
rlabel metal2 s 14830 22056 14886 22856 6 chany_top_out[5]
port 77 nsew signal tristate
rlabel metal2 s 15382 22056 15438 22856 6 chany_top_out[6]
port 78 nsew signal tristate
rlabel metal2 s 15934 22056 15990 22856 6 chany_top_out[7]
port 79 nsew signal tristate
rlabel metal2 s 16486 22056 16542 22856 6 chany_top_out[8]
port 80 nsew signal tristate
rlabel metal2 s 17038 22056 17094 22856 6 chany_top_out[9]
port 81 nsew signal tristate
rlabel metal3 s 22200 22440 23000 22560 6 prog_clk_0_E_in
port 82 nsew signal input
rlabel metal3 s 22200 2176 23000 2296 6 right_bottom_grid_pin_11_
port 83 nsew signal input
rlabel metal3 s 22200 2720 23000 2840 6 right_bottom_grid_pin_13_
port 84 nsew signal input
rlabel metal3 s 22200 3128 23000 3248 6 right_bottom_grid_pin_15_
port 85 nsew signal input
rlabel metal3 s 22200 3672 23000 3792 6 right_bottom_grid_pin_17_
port 86 nsew signal input
rlabel metal3 s 22200 0 23000 120 6 right_bottom_grid_pin_1_
port 87 nsew signal input
rlabel metal3 s 22200 408 23000 528 6 right_bottom_grid_pin_3_
port 88 nsew signal input
rlabel metal3 s 22200 816 23000 936 6 right_bottom_grid_pin_5_
port 89 nsew signal input
rlabel metal3 s 22200 1360 23000 1480 6 right_bottom_grid_pin_7_
port 90 nsew signal input
rlabel metal3 s 22200 1768 23000 1888 6 right_bottom_grid_pin_9_
port 91 nsew signal input
rlabel metal2 s 294 22056 350 22856 6 top_left_grid_pin_1_
port 92 nsew signal input
rlabel metal4 s 18271 1984 18591 20576 6 VPWR
port 93 nsew power bidirectional
rlabel metal4 s 11340 1984 11660 20576 6 VPWR
port 94 nsew power bidirectional
rlabel metal4 s 4409 1984 4729 20576 6 VPWR
port 95 nsew power bidirectional
rlabel metal4 s 14805 1984 15125 20576 6 VGND
port 96 nsew ground bidirectional
rlabel metal4 s 7875 1984 8195 20576 6 VGND
port 97 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 23000 22856
<< end >>
