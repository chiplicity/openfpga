magic
tech sky130A
magscale 1 2
timestamp 1609018413
<< locali >>
rect 19291 13481 19383 13515
rect 19349 13379 19383 13481
rect 10609 13175 10643 13345
rect 5549 12699 5583 12869
rect 8309 12835 8343 12937
rect 7021 12087 7055 12393
rect 13277 11611 13311 11849
rect 13369 11543 13403 11781
rect 18889 11543 18923 11713
rect 3249 11135 3283 11305
rect 9321 9435 9355 9537
rect 9413 9367 9447 9605
rect 11621 8823 11655 9129
rect 11621 6171 11655 6341
rect 9413 5695 9447 5797
rect 3801 5015 3835 5321
rect 2973 3995 3007 4097
rect 13093 2839 13127 3077
<< viali >>
rect 1961 20553 1995 20587
rect 20729 20553 20763 20587
rect 2513 20485 2547 20519
rect 2973 20417 3007 20451
rect 1777 20349 1811 20383
rect 2329 20349 2363 20383
rect 3249 20349 3283 20383
rect 19809 20349 19843 20383
rect 20545 20349 20579 20383
rect 20177 20213 20211 20247
rect 21189 20213 21223 20247
rect 1961 20009 1995 20043
rect 20453 20009 20487 20043
rect 21097 20009 21131 20043
rect 1501 19873 1535 19907
rect 1777 19873 1811 19907
rect 2789 19873 2823 19907
rect 7941 19873 7975 19907
rect 8585 19873 8619 19907
rect 20269 19873 20303 19907
rect 20913 19873 20947 19907
rect 2973 19805 3007 19839
rect 8033 19805 8067 19839
rect 8217 19805 8251 19839
rect 2329 19669 2363 19703
rect 3617 19669 3651 19703
rect 7573 19669 7607 19703
rect 19901 19669 19935 19703
rect 1961 19465 1995 19499
rect 20453 19465 20487 19499
rect 7757 19329 7791 19363
rect 1777 19261 1811 19295
rect 2329 19261 2363 19295
rect 3157 19261 3191 19295
rect 7481 19261 7515 19295
rect 8125 19261 8159 19295
rect 8392 19261 8426 19295
rect 10057 19261 10091 19295
rect 10425 19261 10459 19295
rect 13277 19261 13311 19295
rect 18889 19261 18923 19295
rect 19165 19261 19199 19295
rect 19717 19261 19751 19295
rect 20269 19261 20303 19295
rect 20821 19261 20855 19295
rect 3424 19193 3458 19227
rect 10670 19193 10704 19227
rect 13522 19193 13556 19227
rect 2513 19125 2547 19159
rect 4537 19125 4571 19159
rect 7113 19125 7147 19159
rect 7573 19125 7607 19159
rect 9505 19125 9539 19159
rect 11805 19125 11839 19159
rect 14657 19125 14691 19159
rect 19349 19125 19383 19159
rect 19901 19125 19935 19159
rect 21005 19125 21039 19159
rect 1961 18921 1995 18955
rect 2513 18921 2547 18955
rect 3065 18921 3099 18955
rect 8585 18921 8619 18955
rect 21097 18921 21131 18955
rect 14565 18853 14599 18887
rect 20177 18853 20211 18887
rect 1777 18785 1811 18819
rect 2329 18785 2363 18819
rect 2881 18785 2915 18819
rect 4445 18785 4479 18819
rect 5437 18785 5471 18819
rect 7205 18785 7239 18819
rect 7472 18785 7506 18819
rect 12245 18785 12279 18819
rect 14657 18785 14691 18819
rect 15568 18785 15602 18819
rect 19901 18785 19935 18819
rect 20913 18785 20947 18819
rect 4537 18717 4571 18751
rect 4721 18717 4755 18751
rect 5181 18717 5215 18751
rect 11989 18717 12023 18751
rect 14749 18717 14783 18751
rect 15301 18717 15335 18751
rect 4077 18649 4111 18683
rect 13369 18649 13403 18683
rect 3525 18581 3559 18615
rect 6561 18581 6595 18615
rect 14197 18581 14231 18615
rect 16681 18581 16715 18615
rect 19533 18581 19567 18615
rect 1961 18377 1995 18411
rect 2605 18377 2639 18411
rect 4997 18377 5031 18411
rect 8125 18377 8159 18411
rect 20453 18377 20487 18411
rect 14473 18309 14507 18343
rect 3249 18241 3283 18275
rect 8677 18241 8711 18275
rect 10425 18241 10459 18275
rect 15025 18241 15059 18275
rect 15945 18241 15979 18275
rect 16037 18241 16071 18275
rect 1501 18173 1535 18207
rect 1777 18173 1811 18207
rect 3617 18173 3651 18207
rect 15853 18173 15887 18207
rect 19993 18173 20027 18207
rect 20269 18173 20303 18207
rect 20821 18173 20855 18207
rect 3884 18105 3918 18139
rect 10692 18105 10726 18139
rect 14933 18105 14967 18139
rect 17233 18105 17267 18139
rect 2973 18037 3007 18071
rect 3065 18037 3099 18071
rect 8493 18037 8527 18071
rect 8585 18037 8619 18071
rect 9229 18037 9263 18071
rect 11805 18037 11839 18071
rect 13093 18037 13127 18071
rect 14841 18037 14875 18071
rect 15485 18037 15519 18071
rect 19625 18037 19659 18071
rect 21005 18037 21039 18071
rect 1685 17833 1719 17867
rect 2973 17833 3007 17867
rect 4537 17833 4571 17867
rect 8401 17833 8435 17867
rect 12173 17833 12207 17867
rect 13369 17833 13403 17867
rect 15301 17833 15335 17867
rect 16773 17833 16807 17867
rect 3433 17765 3467 17799
rect 4077 17765 4111 17799
rect 6000 17765 6034 17799
rect 7941 17765 7975 17799
rect 8861 17765 8895 17799
rect 20085 17765 20119 17799
rect 1501 17697 1535 17731
rect 2053 17697 2087 17731
rect 3341 17697 3375 17731
rect 4905 17697 4939 17731
rect 7665 17697 7699 17731
rect 8769 17697 8803 17731
rect 9689 17697 9723 17731
rect 9956 17697 9990 17731
rect 13093 17697 13127 17731
rect 13737 17697 13771 17731
rect 14749 17697 14783 17731
rect 15669 17697 15703 17731
rect 17417 17697 17451 17731
rect 17684 17697 17718 17731
rect 19809 17697 19843 17731
rect 20913 17697 20947 17731
rect 2237 17629 2271 17663
rect 3525 17629 3559 17663
rect 4997 17629 5031 17663
rect 5089 17629 5123 17663
rect 5733 17629 5767 17663
rect 8953 17629 8987 17663
rect 11529 17629 11563 17663
rect 12265 17629 12299 17663
rect 12449 17629 12483 17663
rect 13829 17629 13863 17663
rect 13921 17629 13955 17663
rect 15761 17629 15795 17663
rect 15853 17629 15887 17663
rect 16865 17629 16899 17663
rect 17049 17629 17083 17663
rect 7113 17493 7147 17527
rect 11069 17493 11103 17527
rect 11805 17493 11839 17527
rect 14381 17493 14415 17527
rect 16405 17493 16439 17527
rect 18797 17493 18831 17527
rect 19533 17493 19567 17527
rect 21097 17493 21131 17527
rect 2513 17289 2547 17323
rect 3157 17289 3191 17323
rect 5089 17289 5123 17323
rect 7021 17289 7055 17323
rect 9045 17289 9079 17323
rect 13185 17289 13219 17323
rect 15117 17289 15151 17323
rect 1501 17221 1535 17255
rect 8125 17221 8159 17255
rect 3709 17153 3743 17187
rect 4169 17153 4203 17187
rect 5641 17153 5675 17187
rect 7573 17153 7607 17187
rect 9597 17153 9631 17187
rect 10885 17153 10919 17187
rect 11805 17153 11839 17187
rect 12449 17153 12483 17187
rect 13737 17153 13771 17187
rect 15669 17153 15703 17187
rect 16681 17153 16715 17187
rect 1777 17085 1811 17119
rect 2329 17085 2363 17119
rect 3617 17085 3651 17119
rect 7389 17085 7423 17119
rect 9413 17085 9447 17119
rect 10609 17085 10643 17119
rect 18153 17085 18187 17119
rect 19809 17085 19843 17119
rect 20821 17085 20855 17119
rect 4813 17017 4847 17051
rect 5457 17017 5491 17051
rect 7481 17017 7515 17051
rect 11621 17017 11655 17051
rect 11713 17017 11747 17051
rect 13553 17017 13587 17051
rect 15485 17017 15519 17051
rect 16497 17017 16531 17051
rect 17509 17017 17543 17051
rect 18420 17017 18454 17051
rect 20085 17017 20119 17051
rect 1961 16949 1995 16983
rect 3525 16949 3559 16983
rect 5549 16949 5583 16983
rect 8493 16949 8527 16983
rect 9505 16949 9539 16983
rect 10241 16949 10275 16983
rect 10701 16949 10735 16983
rect 11253 16949 11287 16983
rect 13645 16949 13679 16983
rect 15577 16949 15611 16983
rect 16129 16949 16163 16983
rect 16589 16949 16623 16983
rect 17233 16949 17267 16983
rect 19533 16949 19567 16983
rect 21005 16949 21039 16983
rect 5549 16745 5583 16779
rect 6009 16745 6043 16779
rect 7021 16745 7055 16779
rect 8033 16745 8067 16779
rect 10977 16745 11011 16779
rect 12449 16745 12483 16779
rect 13461 16745 13495 16779
rect 16221 16745 16255 16779
rect 17417 16745 17451 16779
rect 19533 16745 19567 16779
rect 21097 16745 21131 16779
rect 2973 16677 3007 16711
rect 5917 16677 5951 16711
rect 6561 16677 6595 16711
rect 7665 16677 7699 16711
rect 8493 16677 8527 16711
rect 12357 16677 12391 16711
rect 1777 16609 1811 16643
rect 2329 16609 2363 16643
rect 8401 16609 8435 16643
rect 10701 16609 10735 16643
rect 11345 16609 11379 16643
rect 13829 16609 13863 16643
rect 16589 16609 16623 16643
rect 17785 16609 17819 16643
rect 18521 16609 18555 16643
rect 19349 16609 19383 16643
rect 19901 16609 19935 16643
rect 20177 16609 20211 16643
rect 20913 16609 20947 16643
rect 6101 16541 6135 16575
rect 8677 16541 8711 16575
rect 11437 16541 11471 16575
rect 11621 16541 11655 16575
rect 12541 16541 12575 16575
rect 13921 16541 13955 16575
rect 14105 16541 14139 16575
rect 16681 16541 16715 16575
rect 16773 16541 16807 16575
rect 17877 16541 17911 16575
rect 17969 16541 18003 16575
rect 2513 16473 2547 16507
rect 3617 16473 3651 16507
rect 11989 16473 12023 16507
rect 13001 16473 13035 16507
rect 1961 16405 1995 16439
rect 3341 16405 3375 16439
rect 7297 16405 7331 16439
rect 9965 16405 9999 16439
rect 10333 16405 10367 16439
rect 14565 16405 14599 16439
rect 18981 16405 19015 16439
rect 3249 16201 3283 16235
rect 5825 16201 5859 16235
rect 7113 16201 7147 16235
rect 9873 16201 9907 16235
rect 17509 16201 17543 16235
rect 18521 16201 18555 16235
rect 1685 16133 1719 16167
rect 13277 16133 13311 16167
rect 2237 16065 2271 16099
rect 7757 16065 7791 16099
rect 20269 16065 20303 16099
rect 1501 15997 1535 16031
rect 2053 15997 2087 16031
rect 2881 15997 2915 16031
rect 4445 15997 4479 16031
rect 8125 15997 8159 16031
rect 8493 15997 8527 16031
rect 19993 15997 20027 16031
rect 20821 15997 20855 16031
rect 4712 15929 4746 15963
rect 7481 15929 7515 15963
rect 8760 15929 8794 15963
rect 6469 15861 6503 15895
rect 7573 15861 7607 15895
rect 11805 15861 11839 15895
rect 17049 15861 17083 15895
rect 19717 15861 19751 15895
rect 21005 15861 21039 15895
rect 1961 15657 1995 15691
rect 5457 15657 5491 15691
rect 8309 15657 8343 15691
rect 13829 15657 13863 15691
rect 14933 15657 14967 15691
rect 19073 15657 19107 15691
rect 20453 15657 20487 15691
rect 21097 15657 21131 15691
rect 6184 15589 6218 15623
rect 11612 15589 11646 15623
rect 15844 15589 15878 15623
rect 1777 15521 1811 15555
rect 3065 15521 3099 15555
rect 4077 15521 4111 15555
rect 4333 15521 4367 15555
rect 5917 15521 5951 15555
rect 8493 15521 8527 15555
rect 11345 15521 11379 15555
rect 14197 15521 14231 15555
rect 15577 15521 15611 15555
rect 17693 15521 17727 15555
rect 17960 15521 17994 15555
rect 20269 15521 20303 15555
rect 20913 15521 20947 15555
rect 3157 15453 3191 15487
rect 3341 15453 3375 15487
rect 14289 15453 14323 15487
rect 14473 15453 14507 15487
rect 19349 15453 19383 15487
rect 2697 15385 2731 15419
rect 7573 15385 7607 15419
rect 12725 15385 12759 15419
rect 2421 15317 2455 15351
rect 7297 15317 7331 15351
rect 16957 15317 16991 15351
rect 19901 15317 19935 15351
rect 6285 15113 6319 15147
rect 11529 15113 11563 15147
rect 12725 15113 12759 15147
rect 16957 15045 16991 15079
rect 8493 14977 8527 15011
rect 10149 14977 10183 15011
rect 13185 14977 13219 15011
rect 15485 14977 15519 15011
rect 17601 14977 17635 15011
rect 19349 14977 19383 15011
rect 20361 14977 20395 15011
rect 1777 14909 1811 14943
rect 2513 14909 2547 14943
rect 6469 14909 6503 14943
rect 6837 14909 6871 14943
rect 10405 14909 10439 14943
rect 12909 14909 12943 14943
rect 15301 14909 15335 14943
rect 20177 14909 20211 14943
rect 20821 14909 20855 14943
rect 2780 14841 2814 14875
rect 7104 14841 7138 14875
rect 8738 14841 8772 14875
rect 13452 14841 13486 14875
rect 17325 14841 17359 14875
rect 19165 14841 19199 14875
rect 1961 14773 1995 14807
rect 3893 14773 3927 14807
rect 8217 14773 8251 14807
rect 9873 14773 9907 14807
rect 14565 14773 14599 14807
rect 14841 14773 14875 14807
rect 15209 14773 15243 14807
rect 17417 14773 17451 14807
rect 18797 14773 18831 14807
rect 19257 14773 19291 14807
rect 19809 14773 19843 14807
rect 20269 14773 20303 14807
rect 21005 14773 21039 14807
rect 2329 14569 2363 14603
rect 4077 14569 4111 14603
rect 5825 14569 5859 14603
rect 6285 14569 6319 14603
rect 6837 14569 6871 14603
rect 7941 14569 7975 14603
rect 13645 14569 13679 14603
rect 14657 14569 14691 14603
rect 19441 14569 19475 14603
rect 1869 14501 1903 14535
rect 7205 14501 7239 14535
rect 12256 14501 12290 14535
rect 14013 14501 14047 14535
rect 19073 14501 19107 14535
rect 19809 14501 19843 14535
rect 21189 14501 21223 14535
rect 1593 14433 1627 14467
rect 2697 14433 2731 14467
rect 4445 14433 4479 14467
rect 6193 14433 6227 14467
rect 9689 14433 9723 14467
rect 9956 14433 9990 14467
rect 11989 14433 12023 14467
rect 16017 14433 16051 14467
rect 17684 14433 17718 14467
rect 20913 14433 20947 14467
rect 2789 14365 2823 14399
rect 2973 14365 3007 14399
rect 4537 14365 4571 14399
rect 4629 14365 4663 14399
rect 6469 14365 6503 14399
rect 7297 14365 7331 14399
rect 7481 14365 7515 14399
rect 14105 14365 14139 14399
rect 14289 14365 14323 14399
rect 15761 14365 15795 14399
rect 17417 14365 17451 14399
rect 19901 14365 19935 14399
rect 19993 14365 20027 14399
rect 13369 14297 13403 14331
rect 17141 14297 17175 14331
rect 5181 14229 5215 14263
rect 11069 14229 11103 14263
rect 18797 14229 18831 14263
rect 20453 14229 20487 14263
rect 1869 14025 1903 14059
rect 2237 14025 2271 14059
rect 4077 14025 4111 14059
rect 7113 14025 7147 14059
rect 8309 14025 8343 14059
rect 11345 14025 11379 14059
rect 15853 14025 15887 14059
rect 18521 14025 18555 14059
rect 19901 14025 19935 14059
rect 21097 14025 21131 14059
rect 13829 13957 13863 13991
rect 18153 13957 18187 13991
rect 18889 13957 18923 13991
rect 2789 13889 2823 13923
rect 4629 13889 4663 13923
rect 5641 13889 5675 13923
rect 7665 13889 7699 13923
rect 8861 13889 8895 13923
rect 9873 13889 9907 13923
rect 11989 13889 12023 13923
rect 14381 13889 14415 13923
rect 16497 13889 16531 13923
rect 19441 13889 19475 13923
rect 20361 13889 20395 13923
rect 20453 13889 20487 13923
rect 1685 13821 1719 13855
rect 7573 13821 7607 13855
rect 10609 13821 10643 13855
rect 11069 13821 11103 13855
rect 11713 13821 11747 13855
rect 14289 13821 14323 13855
rect 15577 13821 15611 13855
rect 20913 13821 20947 13855
rect 2605 13753 2639 13787
rect 3249 13753 3283 13787
rect 4445 13753 4479 13787
rect 5457 13753 5491 13787
rect 6193 13753 6227 13787
rect 11805 13753 11839 13787
rect 19257 13753 19291 13787
rect 2697 13685 2731 13719
rect 4537 13685 4571 13719
rect 5089 13685 5123 13719
rect 5549 13685 5583 13719
rect 7481 13685 7515 13719
rect 8677 13685 8711 13719
rect 8769 13685 8803 13719
rect 9321 13685 9355 13719
rect 9689 13685 9723 13719
rect 9781 13685 9815 13719
rect 14197 13685 14231 13719
rect 15393 13685 15427 13719
rect 16221 13685 16255 13719
rect 16313 13685 16347 13719
rect 17233 13685 17267 13719
rect 19349 13685 19383 13719
rect 20269 13685 20303 13719
rect 2421 13481 2455 13515
rect 4445 13481 4479 13515
rect 4813 13481 4847 13515
rect 6745 13481 6779 13515
rect 7757 13481 7791 13515
rect 9689 13481 9723 13515
rect 11161 13481 11195 13515
rect 15301 13481 15335 13515
rect 16313 13481 16347 13515
rect 16773 13481 16807 13515
rect 19257 13481 19291 13515
rect 19441 13481 19475 13515
rect 2789 13413 2823 13447
rect 5273 13413 5307 13447
rect 6285 13413 6319 13447
rect 12633 13413 12667 13447
rect 15669 13413 15703 13447
rect 17325 13413 17359 13447
rect 19809 13413 19843 13447
rect 1777 13345 1811 13379
rect 2881 13345 2915 13379
rect 5181 13345 5215 13379
rect 7113 13345 7147 13379
rect 7941 13345 7975 13379
rect 8309 13345 8343 13379
rect 10057 13345 10091 13379
rect 10609 13345 10643 13379
rect 10701 13345 10735 13379
rect 11529 13345 11563 13379
rect 12541 13345 12575 13379
rect 14105 13345 14139 13379
rect 16681 13345 16715 13379
rect 18797 13345 18831 13379
rect 19349 13345 19383 13379
rect 20453 13345 20487 13379
rect 20913 13345 20947 13379
rect 3065 13277 3099 13311
rect 5365 13277 5399 13311
rect 7205 13277 7239 13311
rect 7389 13277 7423 13311
rect 10149 13277 10183 13311
rect 10241 13277 10275 13311
rect 5917 13209 5951 13243
rect 11621 13277 11655 13311
rect 11805 13277 11839 13311
rect 12725 13277 12759 13311
rect 15761 13277 15795 13311
rect 15945 13277 15979 13311
rect 16865 13277 16899 13311
rect 18153 13277 18187 13311
rect 18889 13277 18923 13311
rect 19073 13277 19107 13311
rect 19901 13277 19935 13311
rect 19993 13277 20027 13311
rect 21097 13277 21131 13311
rect 13921 13209 13955 13243
rect 17785 13209 17819 13243
rect 2145 13141 2179 13175
rect 3433 13141 3467 13175
rect 10609 13141 10643 13175
rect 12173 13141 12207 13175
rect 18429 13141 18463 13175
rect 2237 12937 2271 12971
rect 3617 12937 3651 12971
rect 7389 12937 7423 12971
rect 8309 12937 8343 12971
rect 9137 12937 9171 12971
rect 15669 12937 15703 12971
rect 18337 12937 18371 12971
rect 19349 12937 19383 12971
rect 5549 12869 5583 12903
rect 2881 12801 2915 12835
rect 4169 12801 4203 12835
rect 5181 12801 5215 12835
rect 11161 12869 11195 12903
rect 11437 12869 11471 12903
rect 16589 12869 16623 12903
rect 7113 12801 7147 12835
rect 7849 12801 7883 12835
rect 8033 12801 8067 12835
rect 8309 12801 8343 12835
rect 9781 12801 9815 12835
rect 10793 12801 10827 12835
rect 13737 12801 13771 12835
rect 17417 12801 17451 12835
rect 18797 12801 18831 12835
rect 18889 12801 18923 12835
rect 19901 12801 19935 12835
rect 21097 12801 21131 12835
rect 7757 12733 7791 12767
rect 8493 12733 8527 12767
rect 14289 12733 14323 12767
rect 16129 12733 16163 12767
rect 18705 12733 18739 12767
rect 21005 12733 21039 12767
rect 3985 12665 4019 12699
rect 4997 12665 5031 12699
rect 5089 12665 5123 12699
rect 5549 12665 5583 12699
rect 5641 12665 5675 12699
rect 13553 12665 13587 12699
rect 13645 12665 13679 12699
rect 14534 12665 14568 12699
rect 17233 12665 17267 12699
rect 19809 12665 19843 12699
rect 2605 12597 2639 12631
rect 2697 12597 2731 12631
rect 4077 12597 4111 12631
rect 4629 12597 4663 12631
rect 9505 12597 9539 12631
rect 9597 12597 9631 12631
rect 10149 12597 10183 12631
rect 12449 12597 12483 12631
rect 13185 12597 13219 12631
rect 16865 12597 16899 12631
rect 17325 12597 17359 12631
rect 19717 12597 19751 12631
rect 20545 12597 20579 12631
rect 20913 12597 20947 12631
rect 2421 12393 2455 12427
rect 4721 12393 4755 12427
rect 7021 12393 7055 12427
rect 7205 12393 7239 12427
rect 9689 12393 9723 12427
rect 12449 12393 12483 12427
rect 14197 12393 14231 12427
rect 15301 12393 15335 12427
rect 17785 12393 17819 12427
rect 18061 12393 18095 12427
rect 18521 12393 18555 12427
rect 19349 12393 19383 12427
rect 21097 12393 21131 12427
rect 1777 12257 1811 12291
rect 2789 12257 2823 12291
rect 5089 12257 5123 12291
rect 5181 12257 5215 12291
rect 2881 12189 2915 12223
rect 3065 12189 3099 12223
rect 4445 12189 4479 12223
rect 5365 12189 5399 12223
rect 6745 12189 6779 12223
rect 2145 12121 2179 12155
rect 14841 12325 14875 12359
rect 15761 12325 15795 12359
rect 16672 12325 16706 12359
rect 20453 12325 20487 12359
rect 7573 12257 7607 12291
rect 7665 12257 7699 12291
rect 8309 12257 8343 12291
rect 10057 12257 10091 12291
rect 11069 12257 11103 12291
rect 11325 12257 11359 12291
rect 13073 12257 13107 12291
rect 15669 12257 15703 12291
rect 16405 12257 16439 12291
rect 18429 12257 18463 12291
rect 19717 12257 19751 12291
rect 20913 12257 20947 12291
rect 7757 12189 7791 12223
rect 10149 12189 10183 12223
rect 10241 12189 10275 12223
rect 12817 12189 12851 12223
rect 15853 12189 15887 12223
rect 18613 12189 18647 12223
rect 19809 12189 19843 12223
rect 19993 12189 20027 12223
rect 9137 12121 9171 12155
rect 6469 12053 6503 12087
rect 7021 12053 7055 12087
rect 8769 12053 8803 12087
rect 10793 12053 10827 12087
rect 14473 12053 14507 12087
rect 1869 11849 1903 11883
rect 3617 11849 3651 11883
rect 6837 11849 6871 11883
rect 8493 11849 8527 11883
rect 9505 11849 9539 11883
rect 10517 11849 10551 11883
rect 12449 11849 12483 11883
rect 13277 11849 13311 11883
rect 5825 11713 5859 11747
rect 6193 11713 6227 11747
rect 7297 11713 7331 11747
rect 7481 11713 7515 11747
rect 9137 11713 9171 11747
rect 10057 11713 10091 11747
rect 11161 11713 11195 11747
rect 13093 11713 13127 11747
rect 1685 11645 1719 11679
rect 2237 11645 2271 11679
rect 2504 11645 2538 11679
rect 7205 11645 7239 11679
rect 12817 11645 12851 11679
rect 8217 11577 8251 11611
rect 8953 11577 8987 11611
rect 10885 11577 10919 11611
rect 11621 11577 11655 11611
rect 12909 11577 12943 11611
rect 13277 11577 13311 11611
rect 13369 11781 13403 11815
rect 13921 11713 13955 11747
rect 14105 11713 14139 11747
rect 17601 11713 17635 11747
rect 18613 11713 18647 11747
rect 18889 11713 18923 11747
rect 13829 11645 13863 11679
rect 17325 11645 17359 11679
rect 18429 11645 18463 11679
rect 19993 11645 20027 11679
rect 20260 11577 20294 11611
rect 4353 11509 4387 11543
rect 8861 11509 8895 11543
rect 9873 11509 9907 11543
rect 9965 11509 9999 11543
rect 10977 11509 11011 11543
rect 11897 11509 11931 11543
rect 13369 11509 13403 11543
rect 13461 11509 13495 11543
rect 18061 11509 18095 11543
rect 18521 11509 18555 11543
rect 18889 11509 18923 11543
rect 19073 11509 19107 11543
rect 19625 11509 19659 11543
rect 21373 11509 21407 11543
rect 2421 11305 2455 11339
rect 2789 11305 2823 11339
rect 3249 11305 3283 11339
rect 5733 11305 5767 11339
rect 6929 11305 6963 11339
rect 9689 11305 9723 11339
rect 13921 11305 13955 11339
rect 17693 11305 17727 11339
rect 18981 11305 19015 11339
rect 21281 11305 21315 11339
rect 1961 11237 1995 11271
rect 1685 11169 1719 11203
rect 10793 11237 10827 11271
rect 13185 11237 13219 11271
rect 15546 11237 15580 11271
rect 4620 11169 4654 11203
rect 6285 11169 6319 11203
rect 7021 11169 7055 11203
rect 7941 11169 7975 11203
rect 8769 11169 8803 11203
rect 12357 11169 12391 11203
rect 15301 11169 15335 11203
rect 18061 11169 18095 11203
rect 20177 11169 20211 11203
rect 2881 11101 2915 11135
rect 3065 11101 3099 11135
rect 3249 11101 3283 11135
rect 4353 11101 4387 11135
rect 7205 11101 7239 11135
rect 8033 11101 8067 11135
rect 8125 11101 8159 11135
rect 13277 11101 13311 11135
rect 13461 11101 13495 11135
rect 18153 11101 18187 11135
rect 18337 11101 18371 11135
rect 19901 11101 19935 11135
rect 3525 11033 3559 11067
rect 8585 11033 8619 11067
rect 9229 11033 9263 11067
rect 10333 11033 10367 11067
rect 16681 11033 16715 11067
rect 19257 11033 19291 11067
rect 20913 11033 20947 11067
rect 6561 10965 6595 10999
rect 7573 10965 7607 10999
rect 12817 10965 12851 10999
rect 1593 10761 1627 10795
rect 2789 10761 2823 10795
rect 5273 10761 5307 10795
rect 9137 10761 9171 10795
rect 12541 10761 12575 10795
rect 20637 10761 20671 10795
rect 8677 10693 8711 10727
rect 9505 10693 9539 10727
rect 13093 10693 13127 10727
rect 18061 10693 18095 10727
rect 6377 10625 6411 10659
rect 9965 10625 9999 10659
rect 10149 10625 10183 10659
rect 14657 10625 14691 10659
rect 18613 10625 18647 10659
rect 19257 10625 19291 10659
rect 1869 10557 1903 10591
rect 2145 10557 2179 10591
rect 2605 10557 2639 10591
rect 3893 10557 3927 10591
rect 4160 10557 4194 10591
rect 6193 10557 6227 10591
rect 7021 10557 7055 10591
rect 7288 10557 7322 10591
rect 13277 10557 13311 10591
rect 18521 10557 18555 10591
rect 6101 10489 6135 10523
rect 9873 10489 9907 10523
rect 10517 10489 10551 10523
rect 14473 10489 14507 10523
rect 18429 10489 18463 10523
rect 19502 10489 19536 10523
rect 5733 10421 5767 10455
rect 8401 10421 8435 10455
rect 14013 10421 14047 10455
rect 14381 10421 14415 10455
rect 17141 10421 17175 10455
rect 17509 10421 17543 10455
rect 2329 10217 2363 10251
rect 4905 10217 4939 10251
rect 5365 10217 5399 10251
rect 5917 10217 5951 10251
rect 6285 10217 6319 10251
rect 6929 10217 6963 10251
rect 7941 10217 7975 10251
rect 15301 10217 15335 10251
rect 19533 10217 19567 10251
rect 14841 10149 14875 10183
rect 15761 10149 15795 10183
rect 18420 10149 18454 10183
rect 20269 10149 20303 10183
rect 21005 10149 21039 10183
rect 2697 10081 2731 10115
rect 5273 10081 5307 10115
rect 7297 10081 7331 10115
rect 7389 10081 7423 10115
rect 9689 10081 9723 10115
rect 9956 10081 9990 10115
rect 11601 10081 11635 10115
rect 13257 10081 13291 10115
rect 15669 10081 15703 10115
rect 16497 10081 16531 10115
rect 16764 10081 16798 10115
rect 18153 10081 18187 10115
rect 20177 10081 20211 10115
rect 2789 10013 2823 10047
rect 2973 10013 3007 10047
rect 5457 10013 5491 10047
rect 6377 10013 6411 10047
rect 6561 10013 6595 10047
rect 7481 10013 7515 10047
rect 11345 10013 11379 10047
rect 13001 10013 13035 10047
rect 15853 10013 15887 10047
rect 20453 10013 20487 10047
rect 11069 9945 11103 9979
rect 17877 9945 17911 9979
rect 8493 9877 8527 9911
rect 12725 9877 12759 9911
rect 14381 9877 14415 9911
rect 19809 9877 19843 9911
rect 6837 9673 6871 9707
rect 9413 9605 9447 9639
rect 16773 9605 16807 9639
rect 18061 9605 18095 9639
rect 7389 9537 7423 9571
rect 9321 9537 9355 9571
rect 2053 9469 2087 9503
rect 8033 9469 8067 9503
rect 8861 9469 8895 9503
rect 2320 9401 2354 9435
rect 9229 9401 9263 9435
rect 9321 9401 9355 9435
rect 10149 9537 10183 9571
rect 11161 9537 11195 9571
rect 15209 9537 15243 9571
rect 16221 9537 16255 9571
rect 18613 9537 18647 9571
rect 19625 9537 19659 9571
rect 10977 9469 11011 9503
rect 13093 9469 13127 9503
rect 13360 9469 13394 9503
rect 14933 9469 14967 9503
rect 17601 9469 17635 9503
rect 18429 9469 18463 9503
rect 19892 9469 19926 9503
rect 9873 9401 9907 9435
rect 16037 9401 16071 9435
rect 18521 9401 18555 9435
rect 3433 9333 3467 9367
rect 6469 9333 6503 9367
rect 7205 9333 7239 9367
rect 7297 9333 7331 9367
rect 7849 9333 7883 9367
rect 8401 9333 8435 9367
rect 9413 9333 9447 9367
rect 9505 9333 9539 9367
rect 9965 9333 9999 9367
rect 10517 9333 10551 9367
rect 10885 9333 10919 9367
rect 14473 9333 14507 9367
rect 14749 9333 14783 9367
rect 15669 9333 15703 9367
rect 16129 9333 16163 9367
rect 17141 9333 17175 9367
rect 21005 9333 21039 9367
rect 2237 9129 2271 9163
rect 3617 9129 3651 9163
rect 5457 9129 5491 9163
rect 7113 9129 7147 9163
rect 7389 9129 7423 9163
rect 8769 9129 8803 9163
rect 9689 9129 9723 9163
rect 10149 9129 10183 9163
rect 11621 9129 11655 9163
rect 14565 9129 14599 9163
rect 14657 9129 14691 9163
rect 20269 9129 20303 9163
rect 20913 9129 20947 9163
rect 4322 9061 4356 9095
rect 5978 9061 6012 9095
rect 2605 8993 2639 9027
rect 7757 8993 7791 9027
rect 10057 8993 10091 9027
rect 11161 8993 11195 9027
rect 2697 8925 2731 8959
rect 2881 8925 2915 8959
rect 4077 8925 4111 8959
rect 5733 8925 5767 8959
rect 7849 8925 7883 8959
rect 7941 8925 7975 8959
rect 8861 8925 8895 8959
rect 9045 8925 9079 8959
rect 10241 8925 10275 8959
rect 11253 8925 11287 8959
rect 11345 8925 11379 8959
rect 10793 8857 10827 8891
rect 12265 9061 12299 9095
rect 11805 8993 11839 9027
rect 13921 8993 13955 9027
rect 15945 8993 15979 9027
rect 20177 8993 20211 9027
rect 14749 8925 14783 8959
rect 20453 8925 20487 8959
rect 8401 8789 8435 8823
rect 11621 8789 11655 8823
rect 12633 8789 12667 8823
rect 13737 8789 13771 8823
rect 14197 8789 14231 8823
rect 15761 8789 15795 8823
rect 19441 8789 19475 8823
rect 19809 8789 19843 8823
rect 3249 8585 3283 8619
rect 5733 8585 5767 8619
rect 6837 8585 6871 8619
rect 8217 8585 8251 8619
rect 10149 8585 10183 8619
rect 10609 8585 10643 8619
rect 16865 8585 16899 8619
rect 17601 8585 17635 8619
rect 3893 8517 3927 8551
rect 7849 8517 7883 8551
rect 10977 8517 11011 8551
rect 17141 8517 17175 8551
rect 19349 8517 19383 8551
rect 4537 8449 4571 8483
rect 6377 8449 6411 8483
rect 7297 8449 7331 8483
rect 7481 8449 7515 8483
rect 8769 8449 8803 8483
rect 11529 8449 11563 8483
rect 13277 8449 13311 8483
rect 14473 8449 14507 8483
rect 14657 8449 14691 8483
rect 18613 8449 18647 8483
rect 19809 8449 19843 8483
rect 19993 8449 20027 8483
rect 1869 8381 1903 8415
rect 4353 8381 4387 8415
rect 5917 8381 5951 8415
rect 9036 8381 9070 8415
rect 11437 8381 11471 8415
rect 13185 8381 13219 8415
rect 14381 8381 14415 8415
rect 15485 8381 15519 8415
rect 18521 8381 18555 8415
rect 19717 8381 19751 8415
rect 2136 8313 2170 8347
rect 13093 8313 13127 8347
rect 15752 8313 15786 8347
rect 3525 8245 3559 8279
rect 4261 8245 4295 8279
rect 7205 8245 7239 8279
rect 11345 8245 11379 8279
rect 12725 8245 12759 8279
rect 14013 8245 14047 8279
rect 18061 8245 18095 8279
rect 18429 8245 18463 8279
rect 1685 8041 1719 8075
rect 2421 8041 2455 8075
rect 4077 8041 4111 8075
rect 4445 8041 4479 8075
rect 8033 8041 8067 8075
rect 11253 8041 11287 8075
rect 12173 8041 12207 8075
rect 14473 8041 14507 8075
rect 16037 8041 16071 8075
rect 17969 8041 18003 8075
rect 18245 8041 18279 8075
rect 4537 7973 4571 8007
rect 12992 7973 13026 8007
rect 19064 7973 19098 8007
rect 2789 7905 2823 7939
rect 5457 7905 5491 7939
rect 8217 7905 8251 7939
rect 12081 7905 12115 7939
rect 12725 7905 12759 7939
rect 15945 7905 15979 7939
rect 16856 7905 16890 7939
rect 18797 7905 18831 7939
rect 2881 7837 2915 7871
rect 3065 7837 3099 7871
rect 3433 7837 3467 7871
rect 4629 7837 4663 7871
rect 5549 7837 5583 7871
rect 5733 7837 5767 7871
rect 10885 7837 10919 7871
rect 12265 7837 12299 7871
rect 16221 7837 16255 7871
rect 16589 7837 16623 7871
rect 8493 7769 8527 7803
rect 2053 7701 2087 7735
rect 5089 7701 5123 7735
rect 7665 7701 7699 7735
rect 10425 7701 10459 7735
rect 11713 7701 11747 7735
rect 14105 7701 14139 7735
rect 14841 7701 14875 7735
rect 15577 7701 15611 7735
rect 20177 7701 20211 7735
rect 2421 7497 2455 7531
rect 4261 7497 4295 7531
rect 5273 7497 5307 7531
rect 9229 7497 9263 7531
rect 9689 7497 9723 7531
rect 21097 7497 21131 7531
rect 2973 7361 3007 7395
rect 4721 7361 4755 7395
rect 4905 7361 4939 7395
rect 5825 7361 5859 7395
rect 7849 7361 7883 7395
rect 17049 7361 17083 7395
rect 17141 7361 17175 7395
rect 19441 7361 19475 7395
rect 2789 7293 2823 7327
rect 5641 7293 5675 7327
rect 10701 7293 10735 7327
rect 10968 7293 11002 7327
rect 14013 7293 14047 7327
rect 14280 7293 14314 7327
rect 16957 7293 16991 7327
rect 19708 7293 19742 7327
rect 3801 7225 3835 7259
rect 4629 7225 4663 7259
rect 8094 7225 8128 7259
rect 1409 7157 1443 7191
rect 2053 7157 2087 7191
rect 2881 7157 2915 7191
rect 5733 7157 5767 7191
rect 6285 7157 6319 7191
rect 12081 7157 12115 7191
rect 15393 7157 15427 7191
rect 16589 7157 16623 7191
rect 19165 7157 19199 7191
rect 20821 7157 20855 7191
rect 2053 6953 2087 6987
rect 4169 6953 4203 6987
rect 5825 6953 5859 6987
rect 7757 6953 7791 6987
rect 8953 6953 8987 6987
rect 9689 6953 9723 6987
rect 12357 6953 12391 6987
rect 16773 6953 16807 6987
rect 19993 6953 20027 6987
rect 12265 6885 12299 6919
rect 14013 6885 14047 6919
rect 18981 6885 19015 6919
rect 1961 6817 1995 6851
rect 4445 6817 4479 6851
rect 4712 6817 4746 6851
rect 6633 6817 6667 6851
rect 8033 6817 8067 6851
rect 9045 6817 9079 6851
rect 10508 6817 10542 6851
rect 15660 6817 15694 6851
rect 20085 6817 20119 6851
rect 20913 6817 20947 6851
rect 2237 6749 2271 6783
rect 6377 6749 6411 6783
rect 9229 6749 9263 6783
rect 10241 6749 10275 6783
rect 12449 6749 12483 6783
rect 14473 6749 14507 6783
rect 15393 6749 15427 6783
rect 17049 6749 17083 6783
rect 19073 6749 19107 6783
rect 19257 6749 19291 6783
rect 20177 6749 20211 6783
rect 19625 6681 19659 6715
rect 1593 6613 1627 6647
rect 2697 6613 2731 6647
rect 8585 6613 8619 6647
rect 11621 6613 11655 6647
rect 11897 6613 11931 6647
rect 18613 6613 18647 6647
rect 9597 6409 9631 6443
rect 9873 6409 9907 6443
rect 11897 6409 11931 6443
rect 18153 6409 18187 6443
rect 18981 6409 19015 6443
rect 4997 6341 5031 6375
rect 11621 6341 11655 6375
rect 13185 6341 13219 6375
rect 2145 6273 2179 6307
rect 3065 6273 3099 6307
rect 6285 6273 6319 6307
rect 7389 6273 7423 6307
rect 8217 6273 8251 6307
rect 10333 6273 10367 6307
rect 10425 6273 10459 6307
rect 1869 6205 1903 6239
rect 7205 6205 7239 6239
rect 7941 6205 7975 6239
rect 13645 6273 13679 6307
rect 13829 6273 13863 6307
rect 14749 6273 14783 6307
rect 16221 6273 16255 6307
rect 16405 6273 16439 6307
rect 17325 6273 17359 6307
rect 19625 6273 19659 6307
rect 15393 6205 15427 6239
rect 16129 6205 16163 6239
rect 17141 6205 17175 6239
rect 17233 6205 17267 6239
rect 19993 6205 20027 6239
rect 20260 6205 20294 6239
rect 2881 6137 2915 6171
rect 8484 6137 8518 6171
rect 11621 6137 11655 6171
rect 12909 6137 12943 6171
rect 13553 6137 13587 6171
rect 1501 6069 1535 6103
rect 1961 6069 1995 6103
rect 2513 6069 2547 6103
rect 2973 6069 3007 6103
rect 3617 6069 3651 6103
rect 5457 6069 5491 6103
rect 5733 6069 5767 6103
rect 6101 6069 6135 6103
rect 6193 6069 6227 6103
rect 6837 6069 6871 6103
rect 7297 6069 7331 6103
rect 10241 6069 10275 6103
rect 11437 6069 11471 6103
rect 14197 6069 14231 6103
rect 14565 6069 14599 6103
rect 14657 6069 14691 6103
rect 15761 6069 15795 6103
rect 16773 6069 16807 6103
rect 18705 6069 18739 6103
rect 19349 6069 19383 6103
rect 19441 6069 19475 6103
rect 21373 6069 21407 6103
rect 1869 5865 1903 5899
rect 6193 5865 6227 5899
rect 7573 5865 7607 5899
rect 8585 5865 8619 5899
rect 14565 5865 14599 5899
rect 16497 5865 16531 5899
rect 17233 5865 17267 5899
rect 18245 5865 18279 5899
rect 19625 5865 19659 5899
rect 20085 5865 20119 5899
rect 2596 5797 2630 5831
rect 7665 5797 7699 5831
rect 9413 5797 9447 5831
rect 11069 5797 11103 5831
rect 4333 5729 4367 5763
rect 6561 5729 6595 5763
rect 8953 5729 8987 5763
rect 10333 5729 10367 5763
rect 10977 5729 11011 5763
rect 11989 5729 12023 5763
rect 12909 5729 12943 5763
rect 13176 5729 13210 5763
rect 16589 5729 16623 5763
rect 18337 5729 18371 5763
rect 19349 5729 19383 5763
rect 19993 5729 20027 5763
rect 2329 5661 2363 5695
rect 4077 5661 4111 5695
rect 6653 5661 6687 5695
rect 6837 5661 6871 5695
rect 7757 5661 7791 5695
rect 9045 5661 9079 5695
rect 9229 5661 9263 5695
rect 9413 5661 9447 5695
rect 11253 5661 11287 5695
rect 12081 5661 12115 5695
rect 12173 5661 12207 5695
rect 16773 5661 16807 5695
rect 18429 5661 18463 5695
rect 20269 5661 20303 5695
rect 5457 5593 5491 5627
rect 7205 5593 7239 5627
rect 15301 5593 15335 5627
rect 17877 5593 17911 5627
rect 3709 5525 3743 5559
rect 5917 5525 5951 5559
rect 8309 5525 8343 5559
rect 9689 5525 9723 5559
rect 10609 5525 10643 5559
rect 11621 5525 11655 5559
rect 14289 5525 14323 5559
rect 16129 5525 16163 5559
rect 18981 5525 19015 5559
rect 21281 5525 21315 5559
rect 3801 5321 3835 5355
rect 13829 5321 13863 5355
rect 16129 5321 16163 5355
rect 16497 5321 16531 5355
rect 19717 5321 19751 5355
rect 1501 5253 1535 5287
rect 2145 5185 2179 5219
rect 3065 5185 3099 5219
rect 1869 5117 1903 5151
rect 2881 5049 2915 5083
rect 2973 5049 3007 5083
rect 5273 5253 5307 5287
rect 3985 5185 4019 5219
rect 6101 5185 6135 5219
rect 10425 5185 10459 5219
rect 14657 5185 14691 5219
rect 15669 5185 15703 5219
rect 18061 5185 18095 5219
rect 20177 5185 20211 5219
rect 20269 5185 20303 5219
rect 5917 5117 5951 5151
rect 10692 5117 10726 5151
rect 12449 5117 12483 5151
rect 14473 5117 14507 5151
rect 15485 5117 15519 5151
rect 20085 5117 20119 5151
rect 20821 5117 20855 5151
rect 7573 5049 7607 5083
rect 12694 5049 12728 5083
rect 14565 5049 14599 5083
rect 18328 5049 18362 5083
rect 1961 4981 1995 5015
rect 2513 4981 2547 5015
rect 3525 4981 3559 5015
rect 3801 4981 3835 5015
rect 5549 4981 5583 5015
rect 6009 4981 6043 5015
rect 11805 4981 11839 5015
rect 14105 4981 14139 5015
rect 15117 4981 15151 5015
rect 15577 4981 15611 5015
rect 19441 4981 19475 5015
rect 21005 4981 21039 5015
rect 2237 4777 2271 4811
rect 2697 4777 2731 4811
rect 4169 4777 4203 4811
rect 5181 4777 5215 4811
rect 6285 4777 6319 4811
rect 7021 4777 7055 4811
rect 8309 4777 8343 4811
rect 8401 4777 8435 4811
rect 11345 4777 11379 4811
rect 11989 4777 12023 4811
rect 17141 4777 17175 4811
rect 20361 4777 20395 4811
rect 6377 4709 6411 4743
rect 7665 4709 7699 4743
rect 11437 4709 11471 4743
rect 18972 4709 19006 4743
rect 2605 4641 2639 4675
rect 14749 4641 14783 4675
rect 16028 4641 16062 4675
rect 18705 4641 18739 4675
rect 20913 4641 20947 4675
rect 2881 4573 2915 4607
rect 5273 4573 5307 4607
rect 5457 4573 5491 4607
rect 6469 4573 6503 4607
rect 8585 4573 8619 4607
rect 8953 4573 8987 4607
rect 11621 4573 11655 4607
rect 15761 4573 15795 4607
rect 4445 4505 4479 4539
rect 20085 4505 20119 4539
rect 3341 4437 3375 4471
rect 4813 4437 4847 4471
rect 5917 4437 5951 4471
rect 7941 4437 7975 4471
rect 10977 4437 11011 4471
rect 15393 4437 15427 4471
rect 21097 4437 21131 4471
rect 2881 4233 2915 4267
rect 3157 4233 3191 4267
rect 6837 4233 6871 4267
rect 19349 4233 19383 4267
rect 14933 4165 14967 4199
rect 2973 4097 3007 4131
rect 3709 4097 3743 4131
rect 5365 4097 5399 4131
rect 5457 4097 5491 4131
rect 6009 4097 6043 4131
rect 7849 4097 7883 4131
rect 8033 4097 8067 4131
rect 13553 4097 13587 4131
rect 15853 4097 15887 4131
rect 16773 4097 16807 4131
rect 18981 4097 19015 4131
rect 19625 4097 19659 4131
rect 1501 4029 1535 4063
rect 1768 4029 1802 4063
rect 5273 4029 5307 4063
rect 8401 4029 8435 4063
rect 13820 4029 13854 4063
rect 15669 4029 15703 4063
rect 16681 4029 16715 4063
rect 19892 4029 19926 4063
rect 2973 3961 3007 3995
rect 3525 3961 3559 3995
rect 3617 3961 3651 3995
rect 8668 3961 8702 3995
rect 16589 3961 16623 3995
rect 17233 3961 17267 3995
rect 18613 3961 18647 3995
rect 4905 3893 4939 3927
rect 7389 3893 7423 3927
rect 7757 3893 7791 3927
rect 9781 3893 9815 3927
rect 15209 3893 15243 3927
rect 15577 3893 15611 3927
rect 16221 3893 16255 3927
rect 21005 3893 21039 3927
rect 21373 3893 21407 3927
rect 3065 3689 3099 3723
rect 5273 3689 5307 3723
rect 5733 3689 5767 3723
rect 8217 3689 8251 3723
rect 8585 3689 8619 3723
rect 10701 3689 10735 3723
rect 11253 3689 11287 3723
rect 16681 3689 16715 3723
rect 20545 3689 20579 3723
rect 5641 3621 5675 3655
rect 9229 3621 9263 3655
rect 15568 3621 15602 3655
rect 1685 3553 1719 3587
rect 1941 3553 1975 3587
rect 6377 3553 6411 3587
rect 6644 3553 6678 3587
rect 9965 3553 9999 3587
rect 10609 3553 10643 3587
rect 11713 3553 11747 3587
rect 12449 3553 12483 3587
rect 13185 3553 13219 3587
rect 13737 3553 13771 3587
rect 15301 3553 15335 3587
rect 17141 3553 17175 3587
rect 18061 3553 18095 3587
rect 18889 3553 18923 3587
rect 19901 3553 19935 3587
rect 20913 3553 20947 3587
rect 5825 3485 5859 3519
rect 8677 3485 8711 3519
rect 8861 3485 8895 3519
rect 10885 3485 10919 3519
rect 11989 3485 12023 3519
rect 12725 3485 12759 3519
rect 17325 3485 17359 3519
rect 19165 3485 19199 3519
rect 3341 3349 3375 3383
rect 7757 3349 7791 3383
rect 10241 3349 10275 3383
rect 13369 3349 13403 3383
rect 13921 3349 13955 3383
rect 18245 3349 18279 3383
rect 20085 3349 20119 3383
rect 21097 3349 21131 3383
rect 5825 3145 5859 3179
rect 9505 3145 9539 3179
rect 4169 3077 4203 3111
rect 7757 3077 7791 3111
rect 13093 3077 13127 3111
rect 4445 3009 4479 3043
rect 8125 3009 8159 3043
rect 9965 3009 9999 3043
rect 10701 3009 10735 3043
rect 10793 3009 10827 3043
rect 2789 2941 2823 2975
rect 4712 2941 4746 2975
rect 6193 2941 6227 2975
rect 6837 2941 6871 2975
rect 7113 2941 7147 2975
rect 11253 2941 11287 2975
rect 12449 2941 12483 2975
rect 3056 2873 3090 2907
rect 8392 2873 8426 2907
rect 11529 2873 11563 2907
rect 12725 2873 12759 2907
rect 15945 3009 15979 3043
rect 16129 3009 16163 3043
rect 18245 3009 18279 3043
rect 20821 3009 20855 3043
rect 13185 2941 13219 2975
rect 13921 2941 13955 2975
rect 14657 2941 14691 2975
rect 16497 2941 16531 2975
rect 17233 2941 17267 2975
rect 18061 2941 18095 2975
rect 18797 2941 18831 2975
rect 19533 2941 19567 2975
rect 20361 2941 20395 2975
rect 14197 2873 14231 2907
rect 15853 2873 15887 2907
rect 16773 2873 16807 2907
rect 17509 2873 17543 2907
rect 19073 2873 19107 2907
rect 10241 2805 10275 2839
rect 10609 2805 10643 2839
rect 13093 2805 13127 2839
rect 13369 2805 13403 2839
rect 14841 2805 14875 2839
rect 15485 2805 15519 2839
rect 19717 2805 19751 2839
rect 5089 2601 5123 2635
rect 5181 2601 5215 2635
rect 5825 2601 5859 2635
rect 9045 2601 9079 2635
rect 9137 2601 9171 2635
rect 9781 2601 9815 2635
rect 10149 2601 10183 2635
rect 19073 2601 19107 2635
rect 6193 2533 6227 2567
rect 6929 2533 6963 2567
rect 12909 2533 12943 2567
rect 2789 2465 2823 2499
rect 10241 2465 10275 2499
rect 11805 2465 11839 2499
rect 12633 2465 12667 2499
rect 13369 2465 13403 2499
rect 13921 2465 13955 2499
rect 14749 2465 14783 2499
rect 16129 2465 16163 2499
rect 16681 2465 16715 2499
rect 17233 2465 17267 2499
rect 18521 2465 18555 2499
rect 19441 2465 19475 2499
rect 19993 2465 20027 2499
rect 20545 2465 20579 2499
rect 21189 2465 21223 2499
rect 3065 2397 3099 2431
rect 5273 2397 5307 2431
rect 6285 2397 6319 2431
rect 6469 2397 6503 2431
rect 9321 2397 9355 2431
rect 10333 2397 10367 2431
rect 8677 2329 8711 2363
rect 14105 2329 14139 2363
rect 20177 2329 20211 2363
rect 4721 2261 4755 2295
rect 11989 2261 12023 2295
rect 13553 2261 13587 2295
rect 14933 2261 14967 2295
rect 16313 2261 16347 2295
rect 16865 2261 16899 2295
rect 17417 2261 17451 2295
rect 18705 2261 18739 2295
rect 19625 2261 19659 2295
rect 20729 2261 20763 2295
<< metal1 >>
rect 1104 20698 21896 20720
rect 1104 20646 4447 20698
rect 4499 20646 4511 20698
rect 4563 20646 4575 20698
rect 4627 20646 4639 20698
rect 4691 20646 11378 20698
rect 11430 20646 11442 20698
rect 11494 20646 11506 20698
rect 11558 20646 11570 20698
rect 11622 20646 18308 20698
rect 18360 20646 18372 20698
rect 18424 20646 18436 20698
rect 18488 20646 18500 20698
rect 18552 20646 21896 20698
rect 1104 20624 21896 20646
rect 1949 20587 2007 20593
rect 1949 20553 1961 20587
rect 1995 20584 2007 20587
rect 2774 20584 2780 20596
rect 1995 20556 2780 20584
rect 1995 20553 2007 20556
rect 1949 20547 2007 20553
rect 2774 20544 2780 20556
rect 2832 20544 2838 20596
rect 20622 20544 20628 20596
rect 20680 20584 20686 20596
rect 20717 20587 20775 20593
rect 20717 20584 20729 20587
rect 20680 20556 20729 20584
rect 20680 20544 20686 20556
rect 20717 20553 20729 20556
rect 20763 20553 20775 20587
rect 20717 20547 20775 20553
rect 2501 20519 2559 20525
rect 2501 20485 2513 20519
rect 2547 20516 2559 20519
rect 2866 20516 2872 20528
rect 2547 20488 2872 20516
rect 2547 20485 2559 20488
rect 2501 20479 2559 20485
rect 2866 20476 2872 20488
rect 2924 20476 2930 20528
rect 2961 20451 3019 20457
rect 2961 20448 2973 20451
rect 1780 20420 2973 20448
rect 1780 20389 1808 20420
rect 2961 20417 2973 20420
rect 3007 20448 3019 20451
rect 7650 20448 7656 20460
rect 3007 20420 7656 20448
rect 3007 20417 3019 20420
rect 2961 20411 3019 20417
rect 7650 20408 7656 20420
rect 7708 20408 7714 20460
rect 1765 20383 1823 20389
rect 1765 20349 1777 20383
rect 1811 20349 1823 20383
rect 1765 20343 1823 20349
rect 2317 20383 2375 20389
rect 2317 20349 2329 20383
rect 2363 20380 2375 20383
rect 3237 20383 3295 20389
rect 3237 20380 3249 20383
rect 2363 20352 3249 20380
rect 2363 20349 2375 20352
rect 2317 20343 2375 20349
rect 3237 20349 3249 20352
rect 3283 20380 3295 20383
rect 10042 20380 10048 20392
rect 3283 20352 10048 20380
rect 3283 20349 3295 20352
rect 3237 20343 3295 20349
rect 10042 20340 10048 20352
rect 10100 20340 10106 20392
rect 19797 20383 19855 20389
rect 19797 20349 19809 20383
rect 19843 20380 19855 20383
rect 19978 20380 19984 20392
rect 19843 20352 19984 20380
rect 19843 20349 19855 20352
rect 19797 20343 19855 20349
rect 19978 20340 19984 20352
rect 20036 20380 20042 20392
rect 20533 20383 20591 20389
rect 20533 20380 20545 20383
rect 20036 20352 20545 20380
rect 20036 20340 20042 20352
rect 20533 20349 20545 20352
rect 20579 20349 20591 20383
rect 20533 20343 20591 20349
rect 20165 20247 20223 20253
rect 20165 20213 20177 20247
rect 20211 20244 20223 20247
rect 20254 20244 20260 20256
rect 20211 20216 20260 20244
rect 20211 20213 20223 20216
rect 20165 20207 20223 20213
rect 20254 20204 20260 20216
rect 20312 20204 20318 20256
rect 20806 20204 20812 20256
rect 20864 20244 20870 20256
rect 21177 20247 21235 20253
rect 21177 20244 21189 20247
rect 20864 20216 21189 20244
rect 20864 20204 20870 20216
rect 21177 20213 21189 20216
rect 21223 20213 21235 20247
rect 21177 20207 21235 20213
rect 1104 20154 21896 20176
rect 1104 20102 7912 20154
rect 7964 20102 7976 20154
rect 8028 20102 8040 20154
rect 8092 20102 8104 20154
rect 8156 20102 14843 20154
rect 14895 20102 14907 20154
rect 14959 20102 14971 20154
rect 15023 20102 15035 20154
rect 15087 20102 21896 20154
rect 1104 20080 21896 20102
rect 1946 20040 1952 20052
rect 1907 20012 1952 20040
rect 1946 20000 1952 20012
rect 2004 20000 2010 20052
rect 20438 20040 20444 20052
rect 20399 20012 20444 20040
rect 20438 20000 20444 20012
rect 20496 20000 20502 20052
rect 21082 20040 21088 20052
rect 21043 20012 21088 20040
rect 21082 20000 21088 20012
rect 21140 20000 21146 20052
rect 1489 19907 1547 19913
rect 1489 19873 1501 19907
rect 1535 19904 1547 19907
rect 1765 19907 1823 19913
rect 1765 19904 1777 19907
rect 1535 19876 1777 19904
rect 1535 19873 1547 19876
rect 1489 19867 1547 19873
rect 1765 19873 1777 19876
rect 1811 19873 1823 19907
rect 1765 19867 1823 19873
rect 2777 19907 2835 19913
rect 2777 19873 2789 19907
rect 2823 19904 2835 19907
rect 6822 19904 6828 19916
rect 2823 19876 6828 19904
rect 2823 19873 2835 19876
rect 2777 19867 2835 19873
rect 1780 19768 1808 19867
rect 6822 19864 6828 19876
rect 6880 19864 6886 19916
rect 7929 19907 7987 19913
rect 7929 19873 7941 19907
rect 7975 19904 7987 19907
rect 8573 19907 8631 19913
rect 8573 19904 8585 19907
rect 7975 19876 8585 19904
rect 7975 19873 7987 19876
rect 7929 19867 7987 19873
rect 8573 19873 8585 19876
rect 8619 19873 8631 19907
rect 8573 19867 8631 19873
rect 20162 19864 20168 19916
rect 20220 19904 20226 19916
rect 20257 19907 20315 19913
rect 20257 19904 20269 19907
rect 20220 19876 20269 19904
rect 20220 19864 20226 19876
rect 20257 19873 20269 19876
rect 20303 19873 20315 19907
rect 20257 19867 20315 19873
rect 20806 19864 20812 19916
rect 20864 19904 20870 19916
rect 20901 19907 20959 19913
rect 20901 19904 20913 19907
rect 20864 19876 20913 19904
rect 20864 19864 20870 19876
rect 20901 19873 20913 19876
rect 20947 19873 20959 19907
rect 20901 19867 20959 19873
rect 2866 19796 2872 19848
rect 2924 19836 2930 19848
rect 2961 19839 3019 19845
rect 2961 19836 2973 19839
rect 2924 19808 2973 19836
rect 2924 19796 2930 19808
rect 2961 19805 2973 19808
rect 3007 19805 3019 19839
rect 2961 19799 3019 19805
rect 7098 19796 7104 19848
rect 7156 19836 7162 19848
rect 8021 19839 8079 19845
rect 8021 19836 8033 19839
rect 7156 19808 8033 19836
rect 7156 19796 7162 19808
rect 8021 19805 8033 19808
rect 8067 19805 8079 19839
rect 8021 19799 8079 19805
rect 8205 19839 8263 19845
rect 8205 19805 8217 19839
rect 8251 19836 8263 19839
rect 8386 19836 8392 19848
rect 8251 19808 8392 19836
rect 8251 19805 8263 19808
rect 8205 19799 8263 19805
rect 8386 19796 8392 19808
rect 8444 19796 8450 19848
rect 5902 19768 5908 19780
rect 1780 19740 5908 19768
rect 5902 19728 5908 19740
rect 5960 19728 5966 19780
rect 2038 19660 2044 19712
rect 2096 19700 2102 19712
rect 2317 19703 2375 19709
rect 2317 19700 2329 19703
rect 2096 19672 2329 19700
rect 2096 19660 2102 19672
rect 2317 19669 2329 19672
rect 2363 19669 2375 19703
rect 3602 19700 3608 19712
rect 3563 19672 3608 19700
rect 2317 19663 2375 19669
rect 3602 19660 3608 19672
rect 3660 19660 3666 19712
rect 7558 19700 7564 19712
rect 7519 19672 7564 19700
rect 7558 19660 7564 19672
rect 7616 19660 7622 19712
rect 19886 19700 19892 19712
rect 19847 19672 19892 19700
rect 19886 19660 19892 19672
rect 19944 19660 19950 19712
rect 1104 19610 21896 19632
rect 1104 19558 4447 19610
rect 4499 19558 4511 19610
rect 4563 19558 4575 19610
rect 4627 19558 4639 19610
rect 4691 19558 11378 19610
rect 11430 19558 11442 19610
rect 11494 19558 11506 19610
rect 11558 19558 11570 19610
rect 11622 19558 18308 19610
rect 18360 19558 18372 19610
rect 18424 19558 18436 19610
rect 18488 19558 18500 19610
rect 18552 19558 21896 19610
rect 1104 19536 21896 19558
rect 1946 19496 1952 19508
rect 1907 19468 1952 19496
rect 1946 19456 1952 19468
rect 2004 19456 2010 19508
rect 9490 19496 9496 19508
rect 8128 19468 9496 19496
rect 7745 19363 7803 19369
rect 7745 19329 7757 19363
rect 7791 19360 7803 19363
rect 8128 19360 8156 19468
rect 9490 19456 9496 19468
rect 9548 19456 9554 19508
rect 20438 19496 20444 19508
rect 20399 19468 20444 19496
rect 20438 19456 20444 19468
rect 20496 19456 20502 19508
rect 7791 19332 8156 19360
rect 7791 19329 7803 19332
rect 7745 19323 7803 19329
rect 19886 19320 19892 19372
rect 19944 19360 19950 19372
rect 19944 19332 20392 19360
rect 19944 19320 19950 19332
rect 1765 19295 1823 19301
rect 1765 19261 1777 19295
rect 1811 19292 1823 19295
rect 2038 19292 2044 19304
rect 1811 19264 2044 19292
rect 1811 19261 1823 19264
rect 1765 19255 1823 19261
rect 2038 19252 2044 19264
rect 2096 19252 2102 19304
rect 2317 19295 2375 19301
rect 2317 19261 2329 19295
rect 2363 19261 2375 19295
rect 3142 19292 3148 19304
rect 3103 19264 3148 19292
rect 2317 19255 2375 19261
rect 2332 19224 2360 19255
rect 3142 19252 3148 19264
rect 3200 19252 3206 19304
rect 7469 19295 7527 19301
rect 7469 19261 7481 19295
rect 7515 19292 7527 19295
rect 7558 19292 7564 19304
rect 7515 19264 7564 19292
rect 7515 19261 7527 19264
rect 7469 19255 7527 19261
rect 7558 19252 7564 19264
rect 7616 19252 7622 19304
rect 8110 19292 8116 19304
rect 8071 19264 8116 19292
rect 8110 19252 8116 19264
rect 8168 19252 8174 19304
rect 8386 19301 8392 19304
rect 8380 19292 8392 19301
rect 8347 19264 8392 19292
rect 8380 19255 8392 19264
rect 8386 19252 8392 19255
rect 8444 19252 8450 19304
rect 10045 19295 10103 19301
rect 10045 19292 10057 19295
rect 8864 19264 10057 19292
rect 3412 19227 3470 19233
rect 2332 19196 3096 19224
rect 2501 19159 2559 19165
rect 2501 19125 2513 19159
rect 2547 19156 2559 19159
rect 2958 19156 2964 19168
rect 2547 19128 2964 19156
rect 2547 19125 2559 19128
rect 2501 19119 2559 19125
rect 2958 19116 2964 19128
rect 3016 19116 3022 19168
rect 3068 19156 3096 19196
rect 3412 19193 3424 19227
rect 3458 19224 3470 19227
rect 3510 19224 3516 19236
rect 3458 19196 3516 19224
rect 3458 19193 3470 19196
rect 3412 19187 3470 19193
rect 3510 19184 3516 19196
rect 3568 19184 3574 19236
rect 5718 19184 5724 19236
rect 5776 19224 5782 19236
rect 5776 19196 8156 19224
rect 5776 19184 5782 19196
rect 3602 19156 3608 19168
rect 3068 19128 3608 19156
rect 3602 19116 3608 19128
rect 3660 19116 3666 19168
rect 4525 19159 4583 19165
rect 4525 19125 4537 19159
rect 4571 19156 4583 19159
rect 5074 19156 5080 19168
rect 4571 19128 5080 19156
rect 4571 19125 4583 19128
rect 4525 19119 4583 19125
rect 5074 19116 5080 19128
rect 5132 19116 5138 19168
rect 6822 19116 6828 19168
rect 6880 19156 6886 19168
rect 7101 19159 7159 19165
rect 7101 19156 7113 19159
rect 6880 19128 7113 19156
rect 6880 19116 6886 19128
rect 7101 19125 7113 19128
rect 7147 19125 7159 19159
rect 7558 19156 7564 19168
rect 7519 19128 7564 19156
rect 7101 19119 7159 19125
rect 7558 19116 7564 19128
rect 7616 19116 7622 19168
rect 8128 19156 8156 19196
rect 8864 19156 8892 19264
rect 10045 19261 10057 19264
rect 10091 19261 10103 19295
rect 10410 19292 10416 19304
rect 10371 19264 10416 19292
rect 10045 19255 10103 19261
rect 10060 19224 10088 19255
rect 10410 19252 10416 19264
rect 10468 19252 10474 19304
rect 11974 19252 11980 19304
rect 12032 19292 12038 19304
rect 13265 19295 13323 19301
rect 13265 19292 13277 19295
rect 12032 19264 13277 19292
rect 12032 19252 12038 19264
rect 13265 19261 13277 19264
rect 13311 19261 13323 19295
rect 18874 19292 18880 19304
rect 18787 19264 18880 19292
rect 13265 19255 13323 19261
rect 18874 19252 18880 19264
rect 18932 19292 18938 19304
rect 19153 19295 19211 19301
rect 19153 19292 19165 19295
rect 18932 19264 19165 19292
rect 18932 19252 18938 19264
rect 19153 19261 19165 19264
rect 19199 19261 19211 19295
rect 19153 19255 19211 19261
rect 19334 19252 19340 19304
rect 19392 19292 19398 19304
rect 19705 19295 19763 19301
rect 19705 19292 19717 19295
rect 19392 19264 19717 19292
rect 19392 19252 19398 19264
rect 19705 19261 19717 19264
rect 19751 19261 19763 19295
rect 20254 19292 20260 19304
rect 20215 19264 20260 19292
rect 19705 19255 19763 19261
rect 20254 19252 20260 19264
rect 20312 19252 20318 19304
rect 20364 19292 20392 19332
rect 20809 19295 20867 19301
rect 20809 19292 20821 19295
rect 20364 19264 20821 19292
rect 20809 19261 20821 19264
rect 20855 19261 20867 19295
rect 20809 19255 20867 19261
rect 10658 19227 10716 19233
rect 10658 19224 10670 19227
rect 10060 19196 10670 19224
rect 10658 19193 10670 19196
rect 10704 19193 10716 19227
rect 10658 19187 10716 19193
rect 13354 19184 13360 19236
rect 13412 19224 13418 19236
rect 13510 19227 13568 19233
rect 13510 19224 13522 19227
rect 13412 19196 13522 19224
rect 13412 19184 13418 19196
rect 13510 19193 13522 19196
rect 13556 19193 13568 19227
rect 13510 19187 13568 19193
rect 19242 19184 19248 19236
rect 19300 19224 19306 19236
rect 19300 19196 19932 19224
rect 19300 19184 19306 19196
rect 9490 19156 9496 19168
rect 8128 19128 8892 19156
rect 9451 19128 9496 19156
rect 9490 19116 9496 19128
rect 9548 19116 9554 19168
rect 11790 19156 11796 19168
rect 11751 19128 11796 19156
rect 11790 19116 11796 19128
rect 11848 19116 11854 19168
rect 14645 19159 14703 19165
rect 14645 19125 14657 19159
rect 14691 19156 14703 19159
rect 14734 19156 14740 19168
rect 14691 19128 14740 19156
rect 14691 19125 14703 19128
rect 14645 19119 14703 19125
rect 14734 19116 14740 19128
rect 14792 19156 14798 19168
rect 15562 19156 15568 19168
rect 14792 19128 15568 19156
rect 14792 19116 14798 19128
rect 15562 19116 15568 19128
rect 15620 19116 15626 19168
rect 19150 19116 19156 19168
rect 19208 19156 19214 19168
rect 19904 19165 19932 19196
rect 19337 19159 19395 19165
rect 19337 19156 19349 19159
rect 19208 19128 19349 19156
rect 19208 19116 19214 19128
rect 19337 19125 19349 19128
rect 19383 19125 19395 19159
rect 19337 19119 19395 19125
rect 19889 19159 19947 19165
rect 19889 19125 19901 19159
rect 19935 19125 19947 19159
rect 20990 19156 20996 19168
rect 20951 19128 20996 19156
rect 19889 19119 19947 19125
rect 20990 19116 20996 19128
rect 21048 19116 21054 19168
rect 1104 19066 21896 19088
rect 1104 19014 7912 19066
rect 7964 19014 7976 19066
rect 8028 19014 8040 19066
rect 8092 19014 8104 19066
rect 8156 19014 14843 19066
rect 14895 19014 14907 19066
rect 14959 19014 14971 19066
rect 15023 19014 15035 19066
rect 15087 19014 21896 19066
rect 1104 18992 21896 19014
rect 1946 18952 1952 18964
rect 1907 18924 1952 18952
rect 1946 18912 1952 18924
rect 2004 18912 2010 18964
rect 2501 18955 2559 18961
rect 2501 18921 2513 18955
rect 2547 18952 2559 18955
rect 2774 18952 2780 18964
rect 2547 18924 2780 18952
rect 2547 18921 2559 18924
rect 2501 18915 2559 18921
rect 2774 18912 2780 18924
rect 2832 18912 2838 18964
rect 3050 18952 3056 18964
rect 3011 18924 3056 18952
rect 3050 18912 3056 18924
rect 3108 18912 3114 18964
rect 3602 18912 3608 18964
rect 3660 18952 3666 18964
rect 5442 18952 5448 18964
rect 3660 18924 5448 18952
rect 3660 18912 3666 18924
rect 5442 18912 5448 18924
rect 5500 18912 5506 18964
rect 8386 18912 8392 18964
rect 8444 18952 8450 18964
rect 8573 18955 8631 18961
rect 8573 18952 8585 18955
rect 8444 18924 8585 18952
rect 8444 18912 8450 18924
rect 8573 18921 8585 18924
rect 8619 18921 8631 18955
rect 8573 18915 8631 18921
rect 9490 18912 9496 18964
rect 9548 18952 9554 18964
rect 17218 18952 17224 18964
rect 9548 18924 17224 18952
rect 9548 18912 9554 18924
rect 17218 18912 17224 18924
rect 17276 18912 17282 18964
rect 21082 18952 21088 18964
rect 21043 18924 21088 18952
rect 21082 18912 21088 18924
rect 21140 18912 21146 18964
rect 6178 18884 6184 18896
rect 1780 18856 6184 18884
rect 1780 18825 1808 18856
rect 6178 18844 6184 18856
rect 6236 18844 6242 18896
rect 8202 18884 8208 18896
rect 7208 18856 8208 18884
rect 1765 18819 1823 18825
rect 1765 18785 1777 18819
rect 1811 18785 1823 18819
rect 1765 18779 1823 18785
rect 2317 18819 2375 18825
rect 2317 18785 2329 18819
rect 2363 18785 2375 18819
rect 2866 18816 2872 18828
rect 2827 18788 2872 18816
rect 2317 18779 2375 18785
rect 2332 18748 2360 18779
rect 2866 18776 2872 18788
rect 2924 18776 2930 18828
rect 3602 18776 3608 18828
rect 3660 18816 3666 18828
rect 4433 18819 4491 18825
rect 4433 18816 4445 18819
rect 3660 18788 4445 18816
rect 3660 18776 3666 18788
rect 4433 18785 4445 18788
rect 4479 18785 4491 18819
rect 4982 18816 4988 18828
rect 4433 18779 4491 18785
rect 4724 18788 4988 18816
rect 2332 18720 2811 18748
rect 2783 18612 2811 18720
rect 3142 18708 3148 18760
rect 3200 18748 3206 18760
rect 3200 18720 4292 18748
rect 3200 18708 3206 18720
rect 3234 18640 3240 18692
rect 3292 18680 3298 18692
rect 4065 18683 4123 18689
rect 4065 18680 4077 18683
rect 3292 18652 4077 18680
rect 3292 18640 3298 18652
rect 4065 18649 4077 18652
rect 4111 18649 4123 18683
rect 4264 18680 4292 18720
rect 4338 18708 4344 18760
rect 4396 18748 4402 18760
rect 4724 18757 4752 18788
rect 4982 18776 4988 18788
rect 5040 18816 5046 18828
rect 7208 18825 7236 18856
rect 8202 18844 8208 18856
rect 8260 18884 8266 18896
rect 10410 18884 10416 18896
rect 8260 18856 10416 18884
rect 8260 18844 8266 18856
rect 10410 18844 10416 18856
rect 10468 18844 10474 18896
rect 14553 18887 14611 18893
rect 14553 18853 14565 18887
rect 14599 18884 14611 18887
rect 15286 18884 15292 18896
rect 14599 18856 15292 18884
rect 14599 18853 14611 18856
rect 14553 18847 14611 18853
rect 15286 18844 15292 18856
rect 15344 18844 15350 18896
rect 17402 18884 17408 18896
rect 15396 18856 17408 18884
rect 5425 18819 5483 18825
rect 5425 18816 5437 18819
rect 5040 18788 5437 18816
rect 5040 18776 5046 18788
rect 5425 18785 5437 18788
rect 5471 18785 5483 18819
rect 5425 18779 5483 18785
rect 7193 18819 7251 18825
rect 7193 18785 7205 18819
rect 7239 18785 7251 18819
rect 7193 18779 7251 18785
rect 7460 18819 7518 18825
rect 7460 18785 7472 18819
rect 7506 18816 7518 18819
rect 8938 18816 8944 18828
rect 7506 18788 8944 18816
rect 7506 18785 7518 18788
rect 7460 18779 7518 18785
rect 8938 18776 8944 18788
rect 8996 18776 9002 18828
rect 11790 18776 11796 18828
rect 11848 18816 11854 18828
rect 12233 18819 12291 18825
rect 12233 18816 12245 18819
rect 11848 18788 12245 18816
rect 11848 18776 11854 18788
rect 12233 18785 12245 18788
rect 12279 18816 12291 18819
rect 14642 18816 14648 18828
rect 12279 18788 14504 18816
rect 14603 18788 14648 18816
rect 12279 18785 12291 18788
rect 12233 18779 12291 18785
rect 4525 18751 4583 18757
rect 4525 18748 4537 18751
rect 4396 18720 4537 18748
rect 4396 18708 4402 18720
rect 4525 18717 4537 18720
rect 4571 18717 4583 18751
rect 4525 18711 4583 18717
rect 4709 18751 4767 18757
rect 4709 18717 4721 18751
rect 4755 18717 4767 18751
rect 4709 18711 4767 18717
rect 5169 18751 5227 18757
rect 5169 18717 5181 18751
rect 5215 18717 5227 18751
rect 11974 18748 11980 18760
rect 11935 18720 11980 18748
rect 5169 18711 5227 18717
rect 5184 18680 5212 18711
rect 11974 18708 11980 18720
rect 12032 18708 12038 18760
rect 13354 18680 13360 18692
rect 4264 18652 5212 18680
rect 13315 18652 13360 18680
rect 4065 18643 4123 18649
rect 3513 18615 3571 18621
rect 3513 18612 3525 18615
rect 2783 18584 3525 18612
rect 3513 18581 3525 18584
rect 3559 18612 3571 18615
rect 3694 18612 3700 18624
rect 3559 18584 3700 18612
rect 3559 18581 3571 18584
rect 3513 18575 3571 18581
rect 3694 18572 3700 18584
rect 3752 18572 3758 18624
rect 5184 18612 5212 18652
rect 13354 18640 13360 18652
rect 13412 18640 13418 18692
rect 14476 18680 14504 18788
rect 14642 18776 14648 18788
rect 14700 18776 14706 18828
rect 14734 18748 14740 18760
rect 14695 18720 14740 18748
rect 14734 18708 14740 18720
rect 14792 18708 14798 18760
rect 15289 18751 15347 18757
rect 15289 18717 15301 18751
rect 15335 18748 15347 18751
rect 15396 18748 15424 18856
rect 17402 18844 17408 18856
rect 17460 18844 17466 18896
rect 20162 18884 20168 18896
rect 20123 18856 20168 18884
rect 20162 18844 20168 18856
rect 20220 18844 20226 18896
rect 15562 18825 15568 18828
rect 15556 18816 15568 18825
rect 15523 18788 15568 18816
rect 15556 18779 15568 18788
rect 15562 18776 15568 18779
rect 15620 18776 15626 18828
rect 19889 18819 19947 18825
rect 19889 18785 19901 18819
rect 19935 18785 19947 18819
rect 19889 18779 19947 18785
rect 15335 18720 15424 18748
rect 19904 18748 19932 18779
rect 20070 18776 20076 18828
rect 20128 18816 20134 18828
rect 20901 18819 20959 18825
rect 20901 18816 20913 18819
rect 20128 18788 20913 18816
rect 20128 18776 20134 18788
rect 20901 18785 20913 18788
rect 20947 18785 20959 18819
rect 20901 18779 20959 18785
rect 20346 18748 20352 18760
rect 19904 18720 20352 18748
rect 15335 18717 15347 18720
rect 15289 18711 15347 18717
rect 20346 18708 20352 18720
rect 20404 18708 20410 18760
rect 15194 18680 15200 18692
rect 14476 18652 15200 18680
rect 15194 18640 15200 18652
rect 15252 18640 15258 18692
rect 5534 18612 5540 18624
rect 5184 18584 5540 18612
rect 5534 18572 5540 18584
rect 5592 18572 5598 18624
rect 6549 18615 6607 18621
rect 6549 18581 6561 18615
rect 6595 18612 6607 18615
rect 6914 18612 6920 18624
rect 6595 18584 6920 18612
rect 6595 18581 6607 18584
rect 6549 18575 6607 18581
rect 6914 18572 6920 18584
rect 6972 18572 6978 18624
rect 14182 18612 14188 18624
rect 14143 18584 14188 18612
rect 14182 18572 14188 18584
rect 14240 18572 14246 18624
rect 16022 18572 16028 18624
rect 16080 18612 16086 18624
rect 16669 18615 16727 18621
rect 16669 18612 16681 18615
rect 16080 18584 16681 18612
rect 16080 18572 16086 18584
rect 16669 18581 16681 18584
rect 16715 18581 16727 18615
rect 16669 18575 16727 18581
rect 19334 18572 19340 18624
rect 19392 18612 19398 18624
rect 19521 18615 19579 18621
rect 19521 18612 19533 18615
rect 19392 18584 19533 18612
rect 19392 18572 19398 18584
rect 19521 18581 19533 18584
rect 19567 18581 19579 18615
rect 19521 18575 19579 18581
rect 1104 18522 21896 18544
rect 1104 18470 4447 18522
rect 4499 18470 4511 18522
rect 4563 18470 4575 18522
rect 4627 18470 4639 18522
rect 4691 18470 11378 18522
rect 11430 18470 11442 18522
rect 11494 18470 11506 18522
rect 11558 18470 11570 18522
rect 11622 18470 18308 18522
rect 18360 18470 18372 18522
rect 18424 18470 18436 18522
rect 18488 18470 18500 18522
rect 18552 18470 21896 18522
rect 1104 18448 21896 18470
rect 1946 18408 1952 18420
rect 1907 18380 1952 18408
rect 1946 18368 1952 18380
rect 2004 18368 2010 18420
rect 2593 18411 2651 18417
rect 2593 18377 2605 18411
rect 2639 18408 2651 18411
rect 3602 18408 3608 18420
rect 2639 18380 3608 18408
rect 2639 18377 2651 18380
rect 2593 18371 2651 18377
rect 3602 18368 3608 18380
rect 3660 18368 3666 18420
rect 4982 18408 4988 18420
rect 4943 18380 4988 18408
rect 4982 18368 4988 18380
rect 5040 18368 5046 18420
rect 7558 18368 7564 18420
rect 7616 18408 7622 18420
rect 8113 18411 8171 18417
rect 8113 18408 8125 18411
rect 7616 18380 8125 18408
rect 7616 18368 7622 18380
rect 8113 18377 8125 18380
rect 8159 18377 8171 18411
rect 20438 18408 20444 18420
rect 20399 18380 20444 18408
rect 8113 18371 8171 18377
rect 20438 18368 20444 18380
rect 20496 18368 20502 18420
rect 14461 18343 14519 18349
rect 14461 18309 14473 18343
rect 14507 18340 14519 18343
rect 14507 18312 15976 18340
rect 14507 18309 14519 18312
rect 14461 18303 14519 18309
rect 3237 18275 3295 18281
rect 3237 18241 3249 18275
rect 3283 18272 3295 18275
rect 3283 18244 3740 18272
rect 3283 18241 3295 18244
rect 3237 18235 3295 18241
rect 1489 18207 1547 18213
rect 1489 18173 1501 18207
rect 1535 18204 1547 18207
rect 1765 18207 1823 18213
rect 1765 18204 1777 18207
rect 1535 18176 1777 18204
rect 1535 18173 1547 18176
rect 1489 18167 1547 18173
rect 1765 18173 1777 18176
rect 1811 18173 1823 18207
rect 1765 18167 1823 18173
rect 1780 18136 1808 18167
rect 3142 18164 3148 18216
rect 3200 18204 3206 18216
rect 3605 18207 3663 18213
rect 3605 18204 3617 18207
rect 3200 18176 3617 18204
rect 3200 18164 3206 18176
rect 3605 18173 3617 18176
rect 3651 18173 3663 18207
rect 3605 18167 3663 18173
rect 3712 18136 3740 18244
rect 8386 18232 8392 18284
rect 8444 18272 8450 18284
rect 8665 18275 8723 18281
rect 8665 18272 8677 18275
rect 8444 18244 8677 18272
rect 8444 18232 8450 18244
rect 8665 18241 8677 18244
rect 8711 18241 8723 18275
rect 10410 18272 10416 18284
rect 10371 18244 10416 18272
rect 8665 18235 8723 18241
rect 10410 18232 10416 18244
rect 10468 18232 10474 18284
rect 14734 18232 14740 18284
rect 14792 18272 14798 18284
rect 15948 18281 15976 18312
rect 15013 18275 15071 18281
rect 15013 18272 15025 18275
rect 14792 18244 15025 18272
rect 14792 18232 14798 18244
rect 15013 18241 15025 18244
rect 15059 18241 15071 18275
rect 15013 18235 15071 18241
rect 15933 18275 15991 18281
rect 15933 18241 15945 18275
rect 15979 18241 15991 18275
rect 15933 18235 15991 18241
rect 16022 18232 16028 18284
rect 16080 18272 16086 18284
rect 16080 18244 16125 18272
rect 16080 18232 16086 18244
rect 14182 18164 14188 18216
rect 14240 18204 14246 18216
rect 15841 18207 15899 18213
rect 15841 18204 15853 18207
rect 14240 18176 15853 18204
rect 14240 18164 14246 18176
rect 15841 18173 15853 18176
rect 15887 18173 15899 18207
rect 15841 18167 15899 18173
rect 19981 18207 20039 18213
rect 19981 18173 19993 18207
rect 20027 18204 20039 18207
rect 20257 18207 20315 18213
rect 20257 18204 20269 18207
rect 20027 18176 20269 18204
rect 20027 18173 20039 18176
rect 19981 18167 20039 18173
rect 20257 18173 20269 18176
rect 20303 18204 20315 18207
rect 20530 18204 20536 18216
rect 20303 18176 20536 18204
rect 20303 18173 20315 18176
rect 20257 18167 20315 18173
rect 20530 18164 20536 18176
rect 20588 18164 20594 18216
rect 20809 18207 20867 18213
rect 20809 18173 20821 18207
rect 20855 18173 20867 18207
rect 20809 18167 20867 18173
rect 3872 18139 3930 18145
rect 3872 18136 3884 18139
rect 1780 18108 3648 18136
rect 3712 18108 3884 18136
rect 2958 18068 2964 18080
rect 2919 18040 2964 18068
rect 2958 18028 2964 18040
rect 3016 18028 3022 18080
rect 3050 18028 3056 18080
rect 3108 18068 3114 18080
rect 3620 18068 3648 18108
rect 3872 18105 3884 18108
rect 3918 18136 3930 18139
rect 5074 18136 5080 18148
rect 3918 18108 5080 18136
rect 3918 18105 3930 18108
rect 3872 18099 3930 18105
rect 5074 18096 5080 18108
rect 5132 18096 5138 18148
rect 5902 18096 5908 18148
rect 5960 18136 5966 18148
rect 9582 18136 9588 18148
rect 5960 18108 9588 18136
rect 5960 18096 5966 18108
rect 9582 18096 9588 18108
rect 9640 18096 9646 18148
rect 10680 18139 10738 18145
rect 10680 18105 10692 18139
rect 10726 18136 10738 18139
rect 10962 18136 10968 18148
rect 10726 18108 10968 18136
rect 10726 18105 10738 18108
rect 10680 18099 10738 18105
rect 10962 18096 10968 18108
rect 11020 18096 11026 18148
rect 14734 18096 14740 18148
rect 14792 18136 14798 18148
rect 14921 18139 14979 18145
rect 14921 18136 14933 18139
rect 14792 18108 14933 18136
rect 14792 18096 14798 18108
rect 14921 18105 14933 18108
rect 14967 18105 14979 18139
rect 14921 18099 14979 18105
rect 17034 18096 17040 18148
rect 17092 18136 17098 18148
rect 17221 18139 17279 18145
rect 17221 18136 17233 18139
rect 17092 18108 17233 18136
rect 17092 18096 17098 18108
rect 17221 18105 17233 18108
rect 17267 18105 17279 18139
rect 20824 18136 20852 18167
rect 17221 18099 17279 18105
rect 19812 18108 20852 18136
rect 19812 18080 19840 18108
rect 8202 18068 8208 18080
rect 3108 18040 3153 18068
rect 3620 18040 8208 18068
rect 3108 18028 3114 18040
rect 8202 18028 8208 18040
rect 8260 18028 8266 18080
rect 8478 18068 8484 18080
rect 8439 18040 8484 18068
rect 8478 18028 8484 18040
rect 8536 18028 8542 18080
rect 8570 18028 8576 18080
rect 8628 18068 8634 18080
rect 9214 18068 9220 18080
rect 8628 18040 8673 18068
rect 9175 18040 9220 18068
rect 8628 18028 8634 18040
rect 9214 18028 9220 18040
rect 9272 18068 9278 18080
rect 10502 18068 10508 18080
rect 9272 18040 10508 18068
rect 9272 18028 9278 18040
rect 10502 18028 10508 18040
rect 10560 18028 10566 18080
rect 11793 18071 11851 18077
rect 11793 18037 11805 18071
rect 11839 18068 11851 18071
rect 12158 18068 12164 18080
rect 11839 18040 12164 18068
rect 11839 18037 11851 18040
rect 11793 18031 11851 18037
rect 12158 18028 12164 18040
rect 12216 18028 12222 18080
rect 13081 18071 13139 18077
rect 13081 18037 13093 18071
rect 13127 18068 13139 18071
rect 13538 18068 13544 18080
rect 13127 18040 13544 18068
rect 13127 18037 13139 18040
rect 13081 18031 13139 18037
rect 13538 18028 13544 18040
rect 13596 18028 13602 18080
rect 13814 18028 13820 18080
rect 13872 18068 13878 18080
rect 14829 18071 14887 18077
rect 14829 18068 14841 18071
rect 13872 18040 14841 18068
rect 13872 18028 13878 18040
rect 14829 18037 14841 18040
rect 14875 18037 14887 18071
rect 14829 18031 14887 18037
rect 15473 18071 15531 18077
rect 15473 18037 15485 18071
rect 15519 18068 15531 18071
rect 17126 18068 17132 18080
rect 15519 18040 17132 18068
rect 15519 18037 15531 18040
rect 15473 18031 15531 18037
rect 17126 18028 17132 18040
rect 17184 18028 17190 18080
rect 19613 18071 19671 18077
rect 19613 18037 19625 18071
rect 19659 18068 19671 18071
rect 19794 18068 19800 18080
rect 19659 18040 19800 18068
rect 19659 18037 19671 18040
rect 19613 18031 19671 18037
rect 19794 18028 19800 18040
rect 19852 18028 19858 18080
rect 20990 18068 20996 18080
rect 20951 18040 20996 18068
rect 20990 18028 20996 18040
rect 21048 18028 21054 18080
rect 1104 17978 21896 18000
rect 1104 17926 7912 17978
rect 7964 17926 7976 17978
rect 8028 17926 8040 17978
rect 8092 17926 8104 17978
rect 8156 17926 14843 17978
rect 14895 17926 14907 17978
rect 14959 17926 14971 17978
rect 15023 17926 15035 17978
rect 15087 17926 21896 17978
rect 1104 17904 21896 17926
rect 1670 17864 1676 17876
rect 1631 17836 1676 17864
rect 1670 17824 1676 17836
rect 1728 17824 1734 17876
rect 2958 17864 2964 17876
rect 2919 17836 2964 17864
rect 2958 17824 2964 17836
rect 3016 17824 3022 17876
rect 4338 17824 4344 17876
rect 4396 17864 4402 17876
rect 4525 17867 4583 17873
rect 4525 17864 4537 17867
rect 4396 17836 4537 17864
rect 4396 17824 4402 17836
rect 4525 17833 4537 17836
rect 4571 17833 4583 17867
rect 4525 17827 4583 17833
rect 8389 17867 8447 17873
rect 8389 17833 8401 17867
rect 8435 17864 8447 17867
rect 8570 17864 8576 17876
rect 8435 17836 8576 17864
rect 8435 17833 8447 17836
rect 8389 17827 8447 17833
rect 8570 17824 8576 17836
rect 8628 17824 8634 17876
rect 12161 17867 12219 17873
rect 12161 17833 12173 17867
rect 12207 17864 12219 17867
rect 12434 17864 12440 17876
rect 12207 17836 12440 17864
rect 12207 17833 12219 17836
rect 12161 17827 12219 17833
rect 12434 17824 12440 17836
rect 12492 17824 12498 17876
rect 13357 17867 13415 17873
rect 13357 17833 13369 17867
rect 13403 17864 13415 17867
rect 14642 17864 14648 17876
rect 13403 17836 14648 17864
rect 13403 17833 13415 17836
rect 13357 17827 13415 17833
rect 14642 17824 14648 17836
rect 14700 17824 14706 17876
rect 15286 17864 15292 17876
rect 15247 17836 15292 17864
rect 15286 17824 15292 17836
rect 15344 17824 15350 17876
rect 16761 17867 16819 17873
rect 16761 17833 16773 17867
rect 16807 17864 16819 17867
rect 17034 17864 17040 17876
rect 16807 17836 17040 17864
rect 16807 17833 16819 17836
rect 16761 17827 16819 17833
rect 17034 17824 17040 17836
rect 17092 17824 17098 17876
rect 17494 17824 17500 17876
rect 17552 17864 17558 17876
rect 19886 17864 19892 17876
rect 17552 17836 19892 17864
rect 17552 17824 17558 17836
rect 19886 17824 19892 17836
rect 19944 17824 19950 17876
rect 3418 17796 3424 17808
rect 3379 17768 3424 17796
rect 3418 17756 3424 17768
rect 3476 17796 3482 17808
rect 4065 17799 4123 17805
rect 4065 17796 4077 17799
rect 3476 17768 4077 17796
rect 3476 17756 3482 17768
rect 4065 17765 4077 17768
rect 4111 17765 4123 17799
rect 4065 17759 4123 17765
rect 5988 17799 6046 17805
rect 5988 17765 6000 17799
rect 6034 17796 6046 17799
rect 6086 17796 6092 17808
rect 6034 17768 6092 17796
rect 6034 17765 6046 17768
rect 5988 17759 6046 17765
rect 6086 17756 6092 17768
rect 6144 17756 6150 17808
rect 6178 17756 6184 17808
rect 6236 17796 6242 17808
rect 7929 17799 7987 17805
rect 7929 17796 7941 17799
rect 6236 17768 7941 17796
rect 6236 17756 6242 17768
rect 7929 17765 7941 17768
rect 7975 17765 7987 17799
rect 7929 17759 7987 17765
rect 8202 17756 8208 17808
rect 8260 17796 8266 17808
rect 8849 17799 8907 17805
rect 8849 17796 8861 17799
rect 8260 17768 8861 17796
rect 8260 17756 8266 17768
rect 8849 17765 8861 17768
rect 8895 17796 8907 17799
rect 9214 17796 9220 17808
rect 8895 17768 9220 17796
rect 8895 17765 8907 17768
rect 8849 17759 8907 17765
rect 9214 17756 9220 17768
rect 9272 17756 9278 17808
rect 10410 17796 10416 17808
rect 9692 17768 10416 17796
rect 9692 17740 9720 17768
rect 10410 17756 10416 17768
rect 10468 17756 10474 17808
rect 10502 17756 10508 17808
rect 10560 17796 10566 17808
rect 11882 17796 11888 17808
rect 10560 17768 11888 17796
rect 10560 17756 10566 17768
rect 11882 17756 11888 17768
rect 11940 17756 11946 17808
rect 11992 17768 12480 17796
rect 1486 17728 1492 17740
rect 1447 17700 1492 17728
rect 1486 17688 1492 17700
rect 1544 17688 1550 17740
rect 2041 17731 2099 17737
rect 2041 17697 2053 17731
rect 2087 17728 2099 17731
rect 3234 17728 3240 17740
rect 2087 17700 3240 17728
rect 2087 17697 2099 17700
rect 2041 17691 2099 17697
rect 3234 17688 3240 17700
rect 3292 17688 3298 17740
rect 3329 17731 3387 17737
rect 3329 17697 3341 17731
rect 3375 17728 3387 17731
rect 4154 17728 4160 17740
rect 3375 17700 4160 17728
rect 3375 17697 3387 17700
rect 3329 17691 3387 17697
rect 4154 17688 4160 17700
rect 4212 17688 4218 17740
rect 4893 17731 4951 17737
rect 4893 17697 4905 17731
rect 4939 17728 4951 17731
rect 7006 17728 7012 17740
rect 4939 17700 7012 17728
rect 4939 17697 4951 17700
rect 4893 17691 4951 17697
rect 7006 17688 7012 17700
rect 7064 17688 7070 17740
rect 7653 17731 7711 17737
rect 7653 17697 7665 17731
rect 7699 17728 7711 17731
rect 8294 17728 8300 17740
rect 7699 17700 8300 17728
rect 7699 17697 7711 17700
rect 7653 17691 7711 17697
rect 8294 17688 8300 17700
rect 8352 17688 8358 17740
rect 8754 17728 8760 17740
rect 8715 17700 8760 17728
rect 8754 17688 8760 17700
rect 8812 17688 8818 17740
rect 9674 17728 9680 17740
rect 9587 17700 9680 17728
rect 9674 17688 9680 17700
rect 9732 17688 9738 17740
rect 9766 17688 9772 17740
rect 9824 17728 9830 17740
rect 9944 17731 10002 17737
rect 9944 17728 9956 17731
rect 9824 17700 9956 17728
rect 9824 17688 9830 17700
rect 9944 17697 9956 17700
rect 9990 17728 10002 17731
rect 11698 17728 11704 17740
rect 9990 17700 11704 17728
rect 9990 17697 10002 17700
rect 9944 17691 10002 17697
rect 11698 17688 11704 17700
rect 11756 17728 11762 17740
rect 11992 17728 12020 17768
rect 11756 17700 12020 17728
rect 11756 17688 11762 17700
rect 1762 17620 1768 17672
rect 1820 17660 1826 17672
rect 2225 17663 2283 17669
rect 2225 17660 2237 17663
rect 1820 17632 2237 17660
rect 1820 17620 1826 17632
rect 2225 17629 2237 17632
rect 2271 17629 2283 17663
rect 3510 17660 3516 17672
rect 3471 17632 3516 17660
rect 2225 17623 2283 17629
rect 3510 17620 3516 17632
rect 3568 17620 3574 17672
rect 4982 17660 4988 17672
rect 4943 17632 4988 17660
rect 4982 17620 4988 17632
rect 5040 17620 5046 17672
rect 5074 17620 5080 17672
rect 5132 17660 5138 17672
rect 5132 17632 5177 17660
rect 5132 17620 5138 17632
rect 5534 17620 5540 17672
rect 5592 17660 5598 17672
rect 5721 17663 5779 17669
rect 5721 17660 5733 17663
rect 5592 17632 5733 17660
rect 5592 17620 5598 17632
rect 5721 17629 5733 17632
rect 5767 17629 5779 17663
rect 5721 17623 5779 17629
rect 8938 17620 8944 17672
rect 8996 17660 9002 17672
rect 8996 17632 9041 17660
rect 8996 17620 9002 17632
rect 10686 17620 10692 17672
rect 10744 17660 10750 17672
rect 11517 17663 11575 17669
rect 11517 17660 11529 17663
rect 10744 17632 11529 17660
rect 10744 17620 10750 17632
rect 11517 17629 11529 17632
rect 11563 17660 11575 17663
rect 12250 17660 12256 17672
rect 11563 17632 12256 17660
rect 11563 17629 11575 17632
rect 11517 17623 11575 17629
rect 12250 17620 12256 17632
rect 12308 17620 12314 17672
rect 12452 17669 12480 17768
rect 13446 17756 13452 17808
rect 13504 17796 13510 17808
rect 13504 17768 13952 17796
rect 13504 17756 13510 17768
rect 13081 17731 13139 17737
rect 13081 17697 13093 17731
rect 13127 17728 13139 17731
rect 13262 17728 13268 17740
rect 13127 17700 13268 17728
rect 13127 17697 13139 17700
rect 13081 17691 13139 17697
rect 13262 17688 13268 17700
rect 13320 17688 13326 17740
rect 13722 17728 13728 17740
rect 13683 17700 13728 17728
rect 13722 17688 13728 17700
rect 13780 17688 13786 17740
rect 12437 17663 12495 17669
rect 12437 17629 12449 17663
rect 12483 17660 12495 17663
rect 12483 17632 13216 17660
rect 12483 17629 12495 17632
rect 12437 17623 12495 17629
rect 9490 17592 9496 17604
rect 7024 17564 9496 17592
rect 3602 17484 3608 17536
rect 3660 17524 3666 17536
rect 7024 17524 7052 17564
rect 9490 17552 9496 17564
rect 9548 17552 9554 17604
rect 3660 17496 7052 17524
rect 7101 17527 7159 17533
rect 3660 17484 3666 17496
rect 7101 17493 7113 17527
rect 7147 17524 7159 17527
rect 7190 17524 7196 17536
rect 7147 17496 7196 17524
rect 7147 17493 7159 17496
rect 7101 17487 7159 17493
rect 7190 17484 7196 17496
rect 7248 17484 7254 17536
rect 10962 17484 10968 17536
rect 11020 17524 11026 17536
rect 11057 17527 11115 17533
rect 11057 17524 11069 17527
rect 11020 17496 11069 17524
rect 11020 17484 11026 17496
rect 11057 17493 11069 17496
rect 11103 17493 11115 17527
rect 11057 17487 11115 17493
rect 11146 17484 11152 17536
rect 11204 17524 11210 17536
rect 11793 17527 11851 17533
rect 11793 17524 11805 17527
rect 11204 17496 11805 17524
rect 11204 17484 11210 17496
rect 11793 17493 11805 17496
rect 11839 17493 11851 17527
rect 13188 17524 13216 17632
rect 13630 17620 13636 17672
rect 13688 17660 13694 17672
rect 13924 17669 13952 17768
rect 13998 17756 14004 17808
rect 14056 17796 14062 17808
rect 20070 17796 20076 17808
rect 14056 17768 19564 17796
rect 20031 17768 20076 17796
rect 14056 17756 14062 17768
rect 14737 17731 14795 17737
rect 14737 17697 14749 17731
rect 14783 17728 14795 17731
rect 15657 17731 15715 17737
rect 15657 17728 15669 17731
rect 14783 17700 15669 17728
rect 14783 17697 14795 17700
rect 14737 17691 14795 17697
rect 15657 17697 15669 17700
rect 15703 17697 15715 17731
rect 17402 17728 17408 17740
rect 15657 17691 15715 17697
rect 15764 17700 17264 17728
rect 17363 17700 17408 17728
rect 13817 17663 13875 17669
rect 13817 17660 13829 17663
rect 13688 17632 13829 17660
rect 13688 17620 13694 17632
rect 13817 17629 13829 17632
rect 13863 17629 13875 17663
rect 13817 17623 13875 17629
rect 13909 17663 13967 17669
rect 13909 17629 13921 17663
rect 13955 17629 13967 17663
rect 13909 17623 13967 17629
rect 14274 17620 14280 17672
rect 14332 17660 14338 17672
rect 15764 17669 15792 17700
rect 15749 17663 15807 17669
rect 15749 17660 15761 17663
rect 14332 17632 15761 17660
rect 14332 17620 14338 17632
rect 15749 17629 15761 17632
rect 15795 17629 15807 17663
rect 15749 17623 15807 17629
rect 15838 17620 15844 17672
rect 15896 17660 15902 17672
rect 16850 17660 16856 17672
rect 15896 17632 15941 17660
rect 16811 17632 16856 17660
rect 15896 17620 15902 17632
rect 16850 17620 16856 17632
rect 16908 17620 16914 17672
rect 17037 17663 17095 17669
rect 17037 17629 17049 17663
rect 17083 17660 17095 17663
rect 17236 17660 17264 17700
rect 17402 17688 17408 17700
rect 17460 17688 17466 17740
rect 17494 17688 17500 17740
rect 17552 17688 17558 17740
rect 17678 17737 17684 17740
rect 17672 17691 17684 17737
rect 17736 17728 17742 17740
rect 17736 17700 17772 17728
rect 17678 17688 17684 17691
rect 17736 17688 17742 17700
rect 17954 17688 17960 17740
rect 18012 17728 18018 17740
rect 19334 17728 19340 17740
rect 18012 17700 19340 17728
rect 18012 17688 18018 17700
rect 19334 17688 19340 17700
rect 19392 17688 19398 17740
rect 17512 17660 17540 17688
rect 17083 17632 17172 17660
rect 17236 17632 17540 17660
rect 17083 17629 17095 17632
rect 17037 17623 17095 17629
rect 17144 17592 17172 17632
rect 13740 17564 17172 17592
rect 13740 17524 13768 17564
rect 13188 17496 13768 17524
rect 11793 17487 11851 17493
rect 14274 17484 14280 17536
rect 14332 17524 14338 17536
rect 14369 17527 14427 17533
rect 14369 17524 14381 17527
rect 14332 17496 14381 17524
rect 14332 17484 14338 17496
rect 14369 17493 14381 17496
rect 14415 17493 14427 17527
rect 16390 17524 16396 17536
rect 16351 17496 16396 17524
rect 14369 17487 14427 17493
rect 16390 17484 16396 17496
rect 16448 17484 16454 17536
rect 17144 17524 17172 17564
rect 19536 17533 19564 17768
rect 20070 17756 20076 17768
rect 20128 17756 20134 17808
rect 19610 17688 19616 17740
rect 19668 17728 19674 17740
rect 19797 17731 19855 17737
rect 19797 17728 19809 17731
rect 19668 17700 19809 17728
rect 19668 17688 19674 17700
rect 19797 17697 19809 17700
rect 19843 17697 19855 17731
rect 19797 17691 19855 17697
rect 20254 17688 20260 17740
rect 20312 17728 20318 17740
rect 20901 17731 20959 17737
rect 20901 17728 20913 17731
rect 20312 17700 20913 17728
rect 20312 17688 20318 17700
rect 20901 17697 20913 17700
rect 20947 17697 20959 17731
rect 20901 17691 20959 17697
rect 18785 17527 18843 17533
rect 18785 17524 18797 17527
rect 17144 17496 18797 17524
rect 18785 17493 18797 17496
rect 18831 17493 18843 17527
rect 18785 17487 18843 17493
rect 19521 17527 19579 17533
rect 19521 17493 19533 17527
rect 19567 17524 19579 17527
rect 19886 17524 19892 17536
rect 19567 17496 19892 17524
rect 19567 17493 19579 17496
rect 19521 17487 19579 17493
rect 19886 17484 19892 17496
rect 19944 17484 19950 17536
rect 21082 17524 21088 17536
rect 21043 17496 21088 17524
rect 21082 17484 21088 17496
rect 21140 17484 21146 17536
rect 1104 17434 21896 17456
rect 1104 17382 4447 17434
rect 4499 17382 4511 17434
rect 4563 17382 4575 17434
rect 4627 17382 4639 17434
rect 4691 17382 11378 17434
rect 11430 17382 11442 17434
rect 11494 17382 11506 17434
rect 11558 17382 11570 17434
rect 11622 17382 18308 17434
rect 18360 17382 18372 17434
rect 18424 17382 18436 17434
rect 18488 17382 18500 17434
rect 18552 17382 21896 17434
rect 1104 17360 21896 17382
rect 2501 17323 2559 17329
rect 2501 17289 2513 17323
rect 2547 17320 2559 17323
rect 2774 17320 2780 17332
rect 2547 17292 2780 17320
rect 2547 17289 2559 17292
rect 2501 17283 2559 17289
rect 2774 17280 2780 17292
rect 2832 17280 2838 17332
rect 3050 17280 3056 17332
rect 3108 17320 3114 17332
rect 3145 17323 3203 17329
rect 3145 17320 3157 17323
rect 3108 17292 3157 17320
rect 3108 17280 3114 17292
rect 3145 17289 3157 17292
rect 3191 17289 3203 17323
rect 3145 17283 3203 17289
rect 4982 17280 4988 17332
rect 5040 17320 5046 17332
rect 5077 17323 5135 17329
rect 5077 17320 5089 17323
rect 5040 17292 5089 17320
rect 5040 17280 5046 17292
rect 5077 17289 5089 17292
rect 5123 17289 5135 17323
rect 7006 17320 7012 17332
rect 6967 17292 7012 17320
rect 5077 17283 5135 17289
rect 7006 17280 7012 17292
rect 7064 17280 7070 17332
rect 8478 17280 8484 17332
rect 8536 17320 8542 17332
rect 9033 17323 9091 17329
rect 9033 17320 9045 17323
rect 8536 17292 9045 17320
rect 8536 17280 8542 17292
rect 9033 17289 9045 17292
rect 9079 17289 9091 17323
rect 9033 17283 9091 17289
rect 9490 17280 9496 17332
rect 9548 17320 9554 17332
rect 10134 17320 10140 17332
rect 9548 17292 10140 17320
rect 9548 17280 9554 17292
rect 10134 17280 10140 17292
rect 10192 17280 10198 17332
rect 13173 17323 13231 17329
rect 13173 17289 13185 17323
rect 13219 17320 13231 17323
rect 13814 17320 13820 17332
rect 13219 17292 13820 17320
rect 13219 17289 13231 17292
rect 13173 17283 13231 17289
rect 13814 17280 13820 17292
rect 13872 17280 13878 17332
rect 14734 17280 14740 17332
rect 14792 17320 14798 17332
rect 15105 17323 15163 17329
rect 15105 17320 15117 17323
rect 14792 17292 15117 17320
rect 14792 17280 14798 17292
rect 15105 17289 15117 17292
rect 15151 17289 15163 17323
rect 19702 17320 19708 17332
rect 15105 17283 15163 17289
rect 15212 17292 19708 17320
rect 1486 17252 1492 17264
rect 1399 17224 1492 17252
rect 1486 17212 1492 17224
rect 1544 17252 1550 17264
rect 3602 17252 3608 17264
rect 1544 17224 3608 17252
rect 1544 17212 1550 17224
rect 3602 17212 3608 17224
rect 3660 17212 3666 17264
rect 8113 17255 8171 17261
rect 3712 17224 5672 17252
rect 3510 17144 3516 17196
rect 3568 17184 3574 17196
rect 3712 17193 3740 17224
rect 3697 17187 3755 17193
rect 3697 17184 3709 17187
rect 3568 17156 3709 17184
rect 3568 17144 3574 17156
rect 3697 17153 3709 17156
rect 3743 17153 3755 17187
rect 4154 17184 4160 17196
rect 4115 17156 4160 17184
rect 3697 17147 3755 17153
rect 4154 17144 4160 17156
rect 4212 17144 4218 17196
rect 5644 17193 5672 17224
rect 8113 17221 8125 17255
rect 8159 17252 8171 17255
rect 10778 17252 10784 17264
rect 8159 17224 10784 17252
rect 8159 17221 8171 17224
rect 8113 17215 8171 17221
rect 5629 17187 5687 17193
rect 5629 17153 5641 17187
rect 5675 17184 5687 17187
rect 7190 17184 7196 17196
rect 5675 17156 7196 17184
rect 5675 17153 5687 17156
rect 5629 17147 5687 17153
rect 7190 17144 7196 17156
rect 7248 17184 7254 17196
rect 7561 17187 7619 17193
rect 7561 17184 7573 17187
rect 7248 17156 7573 17184
rect 7248 17144 7254 17156
rect 7561 17153 7573 17156
rect 7607 17153 7619 17187
rect 7561 17147 7619 17153
rect 1765 17119 1823 17125
rect 1765 17085 1777 17119
rect 1811 17116 1823 17119
rect 2222 17116 2228 17128
rect 1811 17088 2228 17116
rect 1811 17085 1823 17088
rect 1765 17079 1823 17085
rect 2222 17076 2228 17088
rect 2280 17076 2286 17128
rect 2314 17076 2320 17128
rect 2372 17116 2378 17128
rect 2372 17088 2417 17116
rect 2372 17076 2378 17088
rect 3326 17076 3332 17128
rect 3384 17116 3390 17128
rect 3605 17119 3663 17125
rect 3605 17116 3617 17119
rect 3384 17088 3617 17116
rect 3384 17076 3390 17088
rect 3605 17085 3617 17088
rect 3651 17085 3663 17119
rect 3605 17079 3663 17085
rect 7377 17119 7435 17125
rect 7377 17085 7389 17119
rect 7423 17116 7435 17119
rect 8128 17116 8156 17215
rect 10778 17212 10784 17224
rect 10836 17212 10842 17264
rect 15212 17252 15240 17292
rect 19702 17280 19708 17292
rect 19760 17280 19766 17332
rect 12912 17224 15240 17252
rect 8386 17144 8392 17196
rect 8444 17184 8450 17196
rect 8938 17184 8944 17196
rect 8444 17156 8944 17184
rect 8444 17144 8450 17156
rect 8938 17144 8944 17156
rect 8996 17184 9002 17196
rect 9585 17187 9643 17193
rect 9585 17184 9597 17187
rect 8996 17156 9597 17184
rect 8996 17144 9002 17156
rect 9585 17153 9597 17156
rect 9631 17153 9643 17187
rect 9585 17147 9643 17153
rect 10873 17187 10931 17193
rect 10873 17153 10885 17187
rect 10919 17184 10931 17187
rect 10962 17184 10968 17196
rect 10919 17156 10968 17184
rect 10919 17153 10931 17156
rect 10873 17147 10931 17153
rect 10962 17144 10968 17156
rect 11020 17184 11026 17196
rect 11793 17187 11851 17193
rect 11793 17184 11805 17187
rect 11020 17156 11805 17184
rect 11020 17144 11026 17156
rect 11793 17153 11805 17156
rect 11839 17153 11851 17187
rect 12434 17184 12440 17196
rect 12395 17156 12440 17184
rect 11793 17147 11851 17153
rect 12434 17144 12440 17156
rect 12492 17144 12498 17196
rect 7423 17088 8156 17116
rect 9401 17119 9459 17125
rect 7423 17085 7435 17088
rect 7377 17079 7435 17085
rect 9401 17085 9413 17119
rect 9447 17116 9459 17119
rect 10318 17116 10324 17128
rect 9447 17088 10324 17116
rect 9447 17085 9459 17088
rect 9401 17079 9459 17085
rect 10318 17076 10324 17088
rect 10376 17076 10382 17128
rect 10597 17119 10655 17125
rect 10597 17085 10609 17119
rect 10643 17116 10655 17119
rect 11146 17116 11152 17128
rect 10643 17088 11152 17116
rect 10643 17085 10655 17088
rect 10597 17079 10655 17085
rect 11146 17076 11152 17088
rect 11204 17076 11210 17128
rect 12066 17076 12072 17128
rect 12124 17116 12130 17128
rect 12912 17116 12940 17224
rect 17494 17212 17500 17264
rect 17552 17252 17558 17264
rect 17954 17252 17960 17264
rect 17552 17224 17960 17252
rect 17552 17212 17558 17224
rect 17954 17212 17960 17224
rect 18012 17212 18018 17264
rect 13446 17144 13452 17196
rect 13504 17184 13510 17196
rect 13725 17187 13783 17193
rect 13725 17184 13737 17187
rect 13504 17156 13737 17184
rect 13504 17144 13510 17156
rect 13725 17153 13737 17156
rect 13771 17184 13783 17187
rect 15657 17187 15715 17193
rect 15657 17184 15669 17187
rect 13771 17156 15669 17184
rect 13771 17153 13783 17156
rect 13725 17147 13783 17153
rect 15657 17153 15669 17156
rect 15703 17184 15715 17187
rect 15838 17184 15844 17196
rect 15703 17156 15844 17184
rect 15703 17153 15715 17156
rect 15657 17147 15715 17153
rect 15838 17144 15844 17156
rect 15896 17144 15902 17196
rect 16482 17144 16488 17196
rect 16540 17184 16546 17196
rect 16669 17187 16727 17193
rect 16669 17184 16681 17187
rect 16540 17156 16681 17184
rect 16540 17144 16546 17156
rect 16669 17153 16681 17156
rect 16715 17153 16727 17187
rect 16669 17147 16727 17153
rect 17126 17144 17132 17196
rect 17184 17184 17190 17196
rect 17184 17156 18276 17184
rect 17184 17144 17190 17156
rect 16390 17116 16396 17128
rect 12124 17088 12940 17116
rect 13004 17088 16396 17116
rect 12124 17076 12130 17088
rect 4801 17051 4859 17057
rect 4801 17017 4813 17051
rect 4847 17048 4859 17051
rect 5350 17048 5356 17060
rect 4847 17020 5356 17048
rect 4847 17017 4859 17020
rect 4801 17011 4859 17017
rect 5350 17008 5356 17020
rect 5408 17048 5414 17060
rect 5445 17051 5503 17057
rect 5445 17048 5457 17051
rect 5408 17020 5457 17048
rect 5408 17008 5414 17020
rect 5445 17017 5457 17020
rect 5491 17048 5503 17051
rect 6822 17048 6828 17060
rect 5491 17020 6828 17048
rect 5491 17017 5503 17020
rect 5445 17011 5503 17017
rect 6822 17008 6828 17020
rect 6880 17008 6886 17060
rect 7282 17008 7288 17060
rect 7340 17048 7346 17060
rect 7469 17051 7527 17057
rect 7469 17048 7481 17051
rect 7340 17020 7481 17048
rect 7340 17008 7346 17020
rect 7469 17017 7481 17020
rect 7515 17017 7527 17051
rect 7469 17011 7527 17017
rect 8202 17008 8208 17060
rect 8260 17048 8266 17060
rect 11609 17051 11667 17057
rect 11609 17048 11621 17051
rect 8260 17020 11621 17048
rect 8260 17008 8266 17020
rect 11609 17017 11621 17020
rect 11655 17017 11667 17051
rect 11609 17011 11667 17017
rect 11701 17051 11759 17057
rect 11701 17017 11713 17051
rect 11747 17048 11759 17051
rect 13004 17048 13032 17088
rect 16390 17076 16396 17088
rect 16448 17076 16454 17128
rect 17402 17076 17408 17128
rect 17460 17116 17466 17128
rect 17770 17116 17776 17128
rect 17460 17088 17776 17116
rect 17460 17076 17466 17088
rect 17770 17076 17776 17088
rect 17828 17116 17834 17128
rect 18141 17119 18199 17125
rect 18141 17116 18153 17119
rect 17828 17088 18153 17116
rect 17828 17076 17834 17088
rect 18141 17085 18153 17088
rect 18187 17085 18199 17119
rect 18248 17116 18276 17156
rect 19797 17119 19855 17125
rect 19797 17116 19809 17119
rect 18248 17088 19809 17116
rect 18141 17079 18199 17085
rect 19797 17085 19809 17088
rect 19843 17085 19855 17119
rect 19797 17079 19855 17085
rect 19886 17076 19892 17128
rect 19944 17116 19950 17128
rect 20809 17119 20867 17125
rect 20809 17116 20821 17119
rect 19944 17088 20821 17116
rect 19944 17076 19950 17088
rect 20809 17085 20821 17088
rect 20855 17085 20867 17119
rect 20809 17079 20867 17085
rect 13541 17051 13599 17057
rect 13541 17048 13553 17051
rect 11747 17020 13032 17048
rect 13096 17020 13553 17048
rect 11747 17017 11759 17020
rect 11701 17011 11759 17017
rect 1946 16980 1952 16992
rect 1907 16952 1952 16980
rect 1946 16940 1952 16952
rect 2004 16940 2010 16992
rect 3510 16980 3516 16992
rect 3471 16952 3516 16980
rect 3510 16940 3516 16952
rect 3568 16940 3574 16992
rect 5534 16980 5540 16992
rect 5495 16952 5540 16980
rect 5534 16940 5540 16952
rect 5592 16940 5598 16992
rect 8481 16983 8539 16989
rect 8481 16949 8493 16983
rect 8527 16980 8539 16983
rect 8754 16980 8760 16992
rect 8527 16952 8760 16980
rect 8527 16949 8539 16952
rect 8481 16943 8539 16949
rect 8754 16940 8760 16952
rect 8812 16980 8818 16992
rect 9306 16980 9312 16992
rect 8812 16952 9312 16980
rect 8812 16940 8818 16952
rect 9306 16940 9312 16952
rect 9364 16940 9370 16992
rect 9493 16983 9551 16989
rect 9493 16949 9505 16983
rect 9539 16980 9551 16983
rect 9950 16980 9956 16992
rect 9539 16952 9956 16980
rect 9539 16949 9551 16952
rect 9493 16943 9551 16949
rect 9950 16940 9956 16952
rect 10008 16940 10014 16992
rect 10226 16980 10232 16992
rect 10187 16952 10232 16980
rect 10226 16940 10232 16952
rect 10284 16940 10290 16992
rect 10689 16983 10747 16989
rect 10689 16949 10701 16983
rect 10735 16980 10747 16983
rect 10962 16980 10968 16992
rect 10735 16952 10968 16980
rect 10735 16949 10747 16952
rect 10689 16943 10747 16949
rect 10962 16940 10968 16952
rect 11020 16940 11026 16992
rect 11238 16980 11244 16992
rect 11199 16952 11244 16980
rect 11238 16940 11244 16952
rect 11296 16940 11302 16992
rect 12986 16940 12992 16992
rect 13044 16980 13050 16992
rect 13096 16980 13124 17020
rect 13541 17017 13553 17020
rect 13587 17017 13599 17051
rect 13541 17011 13599 17017
rect 15473 17051 15531 17057
rect 15473 17017 15485 17051
rect 15519 17048 15531 17051
rect 16485 17051 16543 17057
rect 15519 17020 16160 17048
rect 15519 17017 15531 17020
rect 15473 17011 15531 17017
rect 13044 16952 13124 16980
rect 13044 16940 13050 16952
rect 13446 16940 13452 16992
rect 13504 16980 13510 16992
rect 13633 16983 13691 16989
rect 13633 16980 13645 16983
rect 13504 16952 13645 16980
rect 13504 16940 13510 16952
rect 13633 16949 13645 16952
rect 13679 16949 13691 16983
rect 15562 16980 15568 16992
rect 15523 16952 15568 16980
rect 13633 16943 13691 16949
rect 15562 16940 15568 16952
rect 15620 16940 15626 16992
rect 16132 16989 16160 17020
rect 16485 17017 16497 17051
rect 16531 17048 16543 17051
rect 17497 17051 17555 17057
rect 17497 17048 17509 17051
rect 16531 17020 17509 17048
rect 16531 17017 16543 17020
rect 16485 17011 16543 17017
rect 17497 17017 17509 17020
rect 17543 17048 17555 17051
rect 18046 17048 18052 17060
rect 17543 17020 18052 17048
rect 17543 17017 17555 17020
rect 17497 17011 17555 17017
rect 18046 17008 18052 17020
rect 18104 17008 18110 17060
rect 18408 17051 18466 17057
rect 18408 17017 18420 17051
rect 18454 17048 18466 17051
rect 19058 17048 19064 17060
rect 18454 17020 19064 17048
rect 18454 17017 18466 17020
rect 18408 17011 18466 17017
rect 19058 17008 19064 17020
rect 19116 17008 19122 17060
rect 20073 17051 20131 17057
rect 20073 17017 20085 17051
rect 20119 17048 20131 17051
rect 20898 17048 20904 17060
rect 20119 17020 20904 17048
rect 20119 17017 20131 17020
rect 20073 17011 20131 17017
rect 20898 17008 20904 17020
rect 20956 17008 20962 17060
rect 16117 16983 16175 16989
rect 16117 16949 16129 16983
rect 16163 16949 16175 16983
rect 16117 16943 16175 16949
rect 16577 16983 16635 16989
rect 16577 16949 16589 16983
rect 16623 16980 16635 16983
rect 17218 16980 17224 16992
rect 16623 16952 17224 16980
rect 16623 16949 16635 16952
rect 16577 16943 16635 16949
rect 17218 16940 17224 16952
rect 17276 16940 17282 16992
rect 17678 16940 17684 16992
rect 17736 16980 17742 16992
rect 19521 16983 19579 16989
rect 19521 16980 19533 16983
rect 17736 16952 19533 16980
rect 17736 16940 17742 16952
rect 19521 16949 19533 16952
rect 19567 16949 19579 16983
rect 19521 16943 19579 16949
rect 20622 16940 20628 16992
rect 20680 16980 20686 16992
rect 20993 16983 21051 16989
rect 20993 16980 21005 16983
rect 20680 16952 21005 16980
rect 20680 16940 20686 16952
rect 20993 16949 21005 16952
rect 21039 16949 21051 16983
rect 20993 16943 21051 16949
rect 1104 16890 21896 16912
rect 1104 16838 7912 16890
rect 7964 16838 7976 16890
rect 8028 16838 8040 16890
rect 8092 16838 8104 16890
rect 8156 16838 14843 16890
rect 14895 16838 14907 16890
rect 14959 16838 14971 16890
rect 15023 16838 15035 16890
rect 15087 16838 21896 16890
rect 1104 16816 21896 16838
rect 5534 16776 5540 16788
rect 5495 16748 5540 16776
rect 5534 16736 5540 16748
rect 5592 16736 5598 16788
rect 5997 16779 6055 16785
rect 5997 16776 6009 16779
rect 5644 16748 6009 16776
rect 2961 16711 3019 16717
rect 2961 16677 2973 16711
rect 3007 16708 3019 16711
rect 5644 16708 5672 16748
rect 5997 16745 6009 16748
rect 6043 16776 6055 16779
rect 7009 16779 7067 16785
rect 7009 16776 7021 16779
rect 6043 16748 7021 16776
rect 6043 16745 6055 16748
rect 5997 16739 6055 16745
rect 7009 16745 7021 16748
rect 7055 16776 7067 16779
rect 7558 16776 7564 16788
rect 7055 16748 7564 16776
rect 7055 16745 7067 16748
rect 7009 16739 7067 16745
rect 7558 16736 7564 16748
rect 7616 16736 7622 16788
rect 8021 16779 8079 16785
rect 8021 16745 8033 16779
rect 8067 16776 8079 16779
rect 8202 16776 8208 16788
rect 8067 16748 8208 16776
rect 8067 16745 8079 16748
rect 8021 16739 8079 16745
rect 8202 16736 8208 16748
rect 8260 16736 8266 16788
rect 10962 16776 10968 16788
rect 10923 16748 10968 16776
rect 10962 16736 10968 16748
rect 11020 16736 11026 16788
rect 11238 16736 11244 16788
rect 11296 16776 11302 16788
rect 12437 16779 12495 16785
rect 12437 16776 12449 16779
rect 11296 16748 12449 16776
rect 11296 16736 11302 16748
rect 12437 16745 12449 16748
rect 12483 16745 12495 16779
rect 13446 16776 13452 16788
rect 13407 16748 13452 16776
rect 12437 16739 12495 16745
rect 13446 16736 13452 16748
rect 13504 16736 13510 16788
rect 15562 16736 15568 16788
rect 15620 16776 15626 16788
rect 16209 16779 16267 16785
rect 16209 16776 16221 16779
rect 15620 16748 16221 16776
rect 15620 16736 15626 16748
rect 16209 16745 16221 16748
rect 16255 16745 16267 16779
rect 16209 16739 16267 16745
rect 16850 16736 16856 16788
rect 16908 16776 16914 16788
rect 17405 16779 17463 16785
rect 17405 16776 17417 16779
rect 16908 16748 17417 16776
rect 16908 16736 16914 16748
rect 17405 16745 17417 16748
rect 17451 16745 17463 16779
rect 17405 16739 17463 16745
rect 19242 16736 19248 16788
rect 19300 16776 19306 16788
rect 19521 16779 19579 16785
rect 19521 16776 19533 16779
rect 19300 16748 19533 16776
rect 19300 16736 19306 16748
rect 19521 16745 19533 16748
rect 19567 16745 19579 16779
rect 19521 16739 19579 16745
rect 21085 16779 21143 16785
rect 21085 16745 21097 16779
rect 21131 16776 21143 16779
rect 21266 16776 21272 16788
rect 21131 16748 21272 16776
rect 21131 16745 21143 16748
rect 21085 16739 21143 16745
rect 21266 16736 21272 16748
rect 21324 16736 21330 16788
rect 5902 16708 5908 16720
rect 3007 16680 5672 16708
rect 5863 16680 5908 16708
rect 3007 16677 3019 16680
rect 2961 16671 3019 16677
rect 1762 16640 1768 16652
rect 1723 16612 1768 16640
rect 1762 16600 1768 16612
rect 1820 16600 1826 16652
rect 2317 16643 2375 16649
rect 2317 16609 2329 16643
rect 2363 16640 2375 16643
rect 2976 16640 3004 16671
rect 5902 16668 5908 16680
rect 5960 16708 5966 16720
rect 6549 16711 6607 16717
rect 6549 16708 6561 16711
rect 5960 16680 6561 16708
rect 5960 16668 5966 16680
rect 6549 16677 6561 16680
rect 6595 16677 6607 16711
rect 6549 16671 6607 16677
rect 6822 16668 6828 16720
rect 6880 16708 6886 16720
rect 7653 16711 7711 16717
rect 7653 16708 7665 16711
rect 6880 16680 7665 16708
rect 6880 16668 6886 16680
rect 7653 16677 7665 16680
rect 7699 16708 7711 16711
rect 8481 16711 8539 16717
rect 8481 16708 8493 16711
rect 7699 16680 8493 16708
rect 7699 16677 7711 16680
rect 7653 16671 7711 16677
rect 8481 16677 8493 16680
rect 8527 16677 8539 16711
rect 8481 16671 8539 16677
rect 10226 16668 10232 16720
rect 10284 16708 10290 16720
rect 12345 16711 12403 16717
rect 12345 16708 12357 16711
rect 10284 16680 12357 16708
rect 10284 16668 10290 16680
rect 12345 16677 12357 16680
rect 12391 16677 12403 16711
rect 12345 16671 12403 16677
rect 17880 16680 18552 16708
rect 2363 16612 3004 16640
rect 2363 16609 2375 16612
rect 2317 16603 2375 16609
rect 7282 16600 7288 16652
rect 7340 16640 7346 16652
rect 8389 16643 8447 16649
rect 8389 16640 8401 16643
rect 7340 16612 8401 16640
rect 7340 16600 7346 16612
rect 8389 16609 8401 16612
rect 8435 16609 8447 16643
rect 8389 16603 8447 16609
rect 10502 16600 10508 16652
rect 10560 16640 10566 16652
rect 10689 16643 10747 16649
rect 10689 16640 10701 16643
rect 10560 16612 10701 16640
rect 10560 16600 10566 16612
rect 10689 16609 10701 16612
rect 10735 16640 10747 16643
rect 11333 16643 11391 16649
rect 11333 16640 11345 16643
rect 10735 16612 11345 16640
rect 10735 16609 10747 16612
rect 10689 16603 10747 16609
rect 11333 16609 11345 16612
rect 11379 16640 11391 16643
rect 12066 16640 12072 16652
rect 11379 16612 11928 16640
rect 11379 16609 11391 16612
rect 11333 16603 11391 16609
rect 6086 16572 6092 16584
rect 6047 16544 6092 16572
rect 6086 16532 6092 16544
rect 6144 16532 6150 16584
rect 8665 16575 8723 16581
rect 8665 16541 8677 16575
rect 8711 16572 8723 16575
rect 9766 16572 9772 16584
rect 8711 16544 9772 16572
rect 8711 16541 8723 16544
rect 8665 16535 8723 16541
rect 9766 16532 9772 16544
rect 9824 16532 9830 16584
rect 10870 16532 10876 16584
rect 10928 16572 10934 16584
rect 11425 16575 11483 16581
rect 11425 16572 11437 16575
rect 10928 16544 11437 16572
rect 10928 16532 10934 16544
rect 11425 16541 11437 16544
rect 11471 16541 11483 16575
rect 11425 16535 11483 16541
rect 11609 16575 11667 16581
rect 11609 16541 11621 16575
rect 11655 16572 11667 16575
rect 11698 16572 11704 16584
rect 11655 16544 11704 16572
rect 11655 16541 11667 16544
rect 11609 16535 11667 16541
rect 11698 16532 11704 16544
rect 11756 16532 11762 16584
rect 2498 16504 2504 16516
rect 2459 16476 2504 16504
rect 2498 16464 2504 16476
rect 2556 16464 2562 16516
rect 3510 16464 3516 16516
rect 3568 16504 3574 16516
rect 3605 16507 3663 16513
rect 3605 16504 3617 16507
rect 3568 16476 3617 16504
rect 3568 16464 3574 16476
rect 3605 16473 3617 16476
rect 3651 16473 3663 16507
rect 3605 16467 3663 16473
rect 3694 16464 3700 16516
rect 3752 16504 3758 16516
rect 9030 16504 9036 16516
rect 3752 16476 9036 16504
rect 3752 16464 3758 16476
rect 9030 16464 9036 16476
rect 9088 16464 9094 16516
rect 1854 16396 1860 16448
rect 1912 16436 1918 16448
rect 1949 16439 2007 16445
rect 1949 16436 1961 16439
rect 1912 16408 1961 16436
rect 1912 16396 1918 16408
rect 1949 16405 1961 16408
rect 1995 16405 2007 16439
rect 1949 16399 2007 16405
rect 2314 16396 2320 16448
rect 2372 16436 2378 16448
rect 3329 16439 3387 16445
rect 3329 16436 3341 16439
rect 2372 16408 3341 16436
rect 2372 16396 2378 16408
rect 3329 16405 3341 16408
rect 3375 16436 3387 16439
rect 5994 16436 6000 16448
rect 3375 16408 6000 16436
rect 3375 16405 3387 16408
rect 3329 16399 3387 16405
rect 5994 16396 6000 16408
rect 6052 16396 6058 16448
rect 7282 16436 7288 16448
rect 7243 16408 7288 16436
rect 7282 16396 7288 16408
rect 7340 16396 7346 16448
rect 9950 16436 9956 16448
rect 9911 16408 9956 16436
rect 9950 16396 9956 16408
rect 10008 16396 10014 16448
rect 10318 16436 10324 16448
rect 10279 16408 10324 16436
rect 10318 16396 10324 16408
rect 10376 16396 10382 16448
rect 11900 16436 11928 16612
rect 11992 16612 12072 16640
rect 11992 16513 12020 16612
rect 12066 16600 12072 16612
rect 12124 16600 12130 16652
rect 13814 16640 13820 16652
rect 13775 16612 13820 16640
rect 13814 16600 13820 16612
rect 13872 16600 13878 16652
rect 16577 16643 16635 16649
rect 16577 16609 16589 16643
rect 16623 16640 16635 16643
rect 16850 16640 16856 16652
rect 16623 16612 16856 16640
rect 16623 16609 16635 16612
rect 16577 16603 16635 16609
rect 16850 16600 16856 16612
rect 16908 16600 16914 16652
rect 17218 16600 17224 16652
rect 17276 16640 17282 16652
rect 17773 16643 17831 16649
rect 17773 16640 17785 16643
rect 17276 16612 17785 16640
rect 17276 16600 17282 16612
rect 17773 16609 17785 16612
rect 17819 16640 17831 16643
rect 17880 16640 17908 16680
rect 18524 16649 18552 16680
rect 17819 16612 17908 16640
rect 18509 16643 18567 16649
rect 17819 16609 17831 16612
rect 17773 16603 17831 16609
rect 18509 16609 18521 16643
rect 18555 16640 18567 16643
rect 18555 16612 18920 16640
rect 18555 16609 18567 16612
rect 18509 16603 18567 16609
rect 12158 16532 12164 16584
rect 12216 16572 12222 16584
rect 12529 16575 12587 16581
rect 12529 16572 12541 16575
rect 12216 16544 12541 16572
rect 12216 16532 12222 16544
rect 12529 16541 12541 16544
rect 12575 16541 12587 16575
rect 12529 16535 12587 16541
rect 13909 16575 13967 16581
rect 13909 16541 13921 16575
rect 13955 16541 13967 16575
rect 13909 16535 13967 16541
rect 14093 16575 14151 16581
rect 14093 16541 14105 16575
rect 14139 16572 14151 16575
rect 15194 16572 15200 16584
rect 14139 16544 15200 16572
rect 14139 16541 14151 16544
rect 14093 16535 14151 16541
rect 11977 16507 12035 16513
rect 11977 16473 11989 16507
rect 12023 16473 12035 16507
rect 12986 16504 12992 16516
rect 12947 16476 12992 16504
rect 11977 16467 12035 16473
rect 12986 16464 12992 16476
rect 13044 16464 13050 16516
rect 13924 16504 13952 16535
rect 15194 16532 15200 16544
rect 15252 16532 15258 16584
rect 16666 16572 16672 16584
rect 16627 16544 16672 16572
rect 16666 16532 16672 16544
rect 16724 16532 16730 16584
rect 16761 16575 16819 16581
rect 16761 16541 16773 16575
rect 16807 16541 16819 16575
rect 17862 16572 17868 16584
rect 17823 16544 17868 16572
rect 16761 16535 16819 16541
rect 15212 16504 15240 16532
rect 16482 16504 16488 16516
rect 13924 16476 14596 16504
rect 15212 16476 16488 16504
rect 13998 16436 14004 16448
rect 11900 16408 14004 16436
rect 13998 16396 14004 16408
rect 14056 16396 14062 16448
rect 14568 16445 14596 16476
rect 16482 16464 16488 16476
rect 16540 16504 16546 16516
rect 16776 16504 16804 16535
rect 17862 16532 17868 16544
rect 17920 16532 17926 16584
rect 17957 16575 18015 16581
rect 17957 16541 17969 16575
rect 18003 16541 18015 16575
rect 18892 16572 18920 16612
rect 18966 16600 18972 16652
rect 19024 16640 19030 16652
rect 19337 16643 19395 16649
rect 19337 16640 19349 16643
rect 19024 16612 19349 16640
rect 19024 16600 19030 16612
rect 19337 16609 19349 16612
rect 19383 16609 19395 16643
rect 19518 16640 19524 16652
rect 19337 16603 19395 16609
rect 19444 16612 19524 16640
rect 19444 16572 19472 16612
rect 19518 16600 19524 16612
rect 19576 16600 19582 16652
rect 19702 16600 19708 16652
rect 19760 16640 19766 16652
rect 19889 16643 19947 16649
rect 19889 16640 19901 16643
rect 19760 16612 19901 16640
rect 19760 16600 19766 16612
rect 19889 16609 19901 16612
rect 19935 16609 19947 16643
rect 19889 16603 19947 16609
rect 20165 16643 20223 16649
rect 20165 16609 20177 16643
rect 20211 16640 20223 16643
rect 20714 16640 20720 16652
rect 20211 16612 20720 16640
rect 20211 16609 20223 16612
rect 20165 16603 20223 16609
rect 20714 16600 20720 16612
rect 20772 16600 20778 16652
rect 20898 16640 20904 16652
rect 20859 16612 20904 16640
rect 20898 16600 20904 16612
rect 20956 16600 20962 16652
rect 18892 16544 19472 16572
rect 17957 16535 18015 16541
rect 16540 16476 16804 16504
rect 16540 16464 16546 16476
rect 17678 16464 17684 16516
rect 17736 16504 17742 16516
rect 17972 16504 18000 16535
rect 17736 16476 18000 16504
rect 17736 16464 17742 16476
rect 14553 16439 14611 16445
rect 14553 16405 14565 16439
rect 14599 16436 14611 16439
rect 17034 16436 17040 16448
rect 14599 16408 17040 16436
rect 14599 16405 14611 16408
rect 14553 16399 14611 16405
rect 17034 16396 17040 16408
rect 17092 16396 17098 16448
rect 18966 16436 18972 16448
rect 18927 16408 18972 16436
rect 18966 16396 18972 16408
rect 19024 16396 19030 16448
rect 1104 16346 21896 16368
rect 1104 16294 4447 16346
rect 4499 16294 4511 16346
rect 4563 16294 4575 16346
rect 4627 16294 4639 16346
rect 4691 16294 11378 16346
rect 11430 16294 11442 16346
rect 11494 16294 11506 16346
rect 11558 16294 11570 16346
rect 11622 16294 18308 16346
rect 18360 16294 18372 16346
rect 18424 16294 18436 16346
rect 18488 16294 18500 16346
rect 18552 16294 21896 16346
rect 1104 16272 21896 16294
rect 3237 16235 3295 16241
rect 3237 16201 3249 16235
rect 3283 16232 3295 16235
rect 3326 16232 3332 16244
rect 3283 16204 3332 16232
rect 3283 16201 3295 16204
rect 3237 16195 3295 16201
rect 3326 16192 3332 16204
rect 3384 16232 3390 16244
rect 4246 16232 4252 16244
rect 3384 16204 4252 16232
rect 3384 16192 3390 16204
rect 4246 16192 4252 16204
rect 4304 16192 4310 16244
rect 5813 16235 5871 16241
rect 5813 16201 5825 16235
rect 5859 16232 5871 16235
rect 6086 16232 6092 16244
rect 5859 16204 6092 16232
rect 5859 16201 5871 16204
rect 5813 16195 5871 16201
rect 6086 16192 6092 16204
rect 6144 16192 6150 16244
rect 7098 16232 7104 16244
rect 7059 16204 7104 16232
rect 7098 16192 7104 16204
rect 7156 16192 7162 16244
rect 8386 16192 8392 16244
rect 8444 16232 8450 16244
rect 9861 16235 9919 16241
rect 9861 16232 9873 16235
rect 8444 16204 9873 16232
rect 8444 16192 8450 16204
rect 9861 16201 9873 16204
rect 9907 16201 9919 16235
rect 9861 16195 9919 16201
rect 10318 16192 10324 16244
rect 10376 16232 10382 16244
rect 13538 16232 13544 16244
rect 10376 16204 13544 16232
rect 10376 16192 10382 16204
rect 13538 16192 13544 16204
rect 13596 16192 13602 16244
rect 16666 16192 16672 16244
rect 16724 16232 16730 16244
rect 17497 16235 17555 16241
rect 17497 16232 17509 16235
rect 16724 16204 17509 16232
rect 16724 16192 16730 16204
rect 17497 16201 17509 16204
rect 17543 16232 17555 16235
rect 17954 16232 17960 16244
rect 17543 16204 17960 16232
rect 17543 16201 17555 16204
rect 17497 16195 17555 16201
rect 17954 16192 17960 16204
rect 18012 16232 18018 16244
rect 18138 16232 18144 16244
rect 18012 16204 18144 16232
rect 18012 16192 18018 16204
rect 18138 16192 18144 16204
rect 18196 16232 18202 16244
rect 18509 16235 18567 16241
rect 18509 16232 18521 16235
rect 18196 16204 18521 16232
rect 18196 16192 18202 16204
rect 18509 16201 18521 16204
rect 18555 16232 18567 16235
rect 18690 16232 18696 16244
rect 18555 16204 18696 16232
rect 18555 16201 18567 16204
rect 18509 16195 18567 16201
rect 18690 16192 18696 16204
rect 18748 16192 18754 16244
rect 1670 16164 1676 16176
rect 1631 16136 1676 16164
rect 1670 16124 1676 16136
rect 1728 16124 1734 16176
rect 1780 16136 2912 16164
rect 1489 16031 1547 16037
rect 1489 15997 1501 16031
rect 1535 16028 1547 16031
rect 1780 16028 1808 16136
rect 2222 16096 2228 16108
rect 2183 16068 2228 16096
rect 2222 16056 2228 16068
rect 2280 16056 2286 16108
rect 2884 16037 2912 16136
rect 9490 16124 9496 16176
rect 9548 16164 9554 16176
rect 13265 16167 13323 16173
rect 13265 16164 13277 16167
rect 9548 16136 13277 16164
rect 9548 16124 9554 16136
rect 13265 16133 13277 16136
rect 13311 16164 13323 16167
rect 13814 16164 13820 16176
rect 13311 16136 13820 16164
rect 13311 16133 13323 16136
rect 13265 16127 13323 16133
rect 13814 16124 13820 16136
rect 13872 16124 13878 16176
rect 7745 16099 7803 16105
rect 7745 16065 7757 16099
rect 7791 16096 7803 16099
rect 8386 16096 8392 16108
rect 7791 16068 8392 16096
rect 7791 16065 7803 16068
rect 7745 16059 7803 16065
rect 8386 16056 8392 16068
rect 8444 16056 8450 16108
rect 11698 16056 11704 16108
rect 11756 16096 11762 16108
rect 18966 16096 18972 16108
rect 11756 16068 18972 16096
rect 11756 16056 11762 16068
rect 18966 16056 18972 16068
rect 19024 16056 19030 16108
rect 20254 16096 20260 16108
rect 20215 16068 20260 16096
rect 20254 16056 20260 16068
rect 20312 16056 20318 16108
rect 1535 16000 1808 16028
rect 2041 16031 2099 16037
rect 1535 15997 1547 16000
rect 1489 15991 1547 15997
rect 2041 15997 2053 16031
rect 2087 15997 2099 16031
rect 2041 15991 2099 15997
rect 2869 16031 2927 16037
rect 2869 15997 2881 16031
rect 2915 16028 2927 16031
rect 4338 16028 4344 16040
rect 2915 16000 4344 16028
rect 2915 15997 2927 16000
rect 2869 15991 2927 15997
rect 2056 15960 2084 15991
rect 4338 15988 4344 16000
rect 4396 15988 4402 16040
rect 4430 15988 4436 16040
rect 4488 16028 4494 16040
rect 5626 16028 5632 16040
rect 4488 16000 5632 16028
rect 4488 15988 4494 16000
rect 5626 15988 5632 16000
rect 5684 15988 5690 16040
rect 7282 15988 7288 16040
rect 7340 16028 7346 16040
rect 8113 16031 8171 16037
rect 8113 16028 8125 16031
rect 7340 16000 8125 16028
rect 7340 15988 7346 16000
rect 8113 15997 8125 16000
rect 8159 15997 8171 16031
rect 8478 16028 8484 16040
rect 8391 16000 8484 16028
rect 8113 15991 8171 15997
rect 8478 15988 8484 16000
rect 8536 16028 8542 16040
rect 9674 16028 9680 16040
rect 8536 16000 9680 16028
rect 8536 15988 8542 16000
rect 9674 15988 9680 16000
rect 9732 15988 9738 16040
rect 13814 15988 13820 16040
rect 13872 16028 13878 16040
rect 19981 16031 20039 16037
rect 19981 16028 19993 16031
rect 13872 16000 19993 16028
rect 13872 15988 13878 16000
rect 19981 15997 19993 16000
rect 20027 15997 20039 16031
rect 19981 15991 20039 15997
rect 20714 15988 20720 16040
rect 20772 16028 20778 16040
rect 20809 16031 20867 16037
rect 20809 16028 20821 16031
rect 20772 16000 20821 16028
rect 20772 15988 20778 16000
rect 20809 15997 20821 16000
rect 20855 15997 20867 16031
rect 20809 15991 20867 15997
rect 4706 15969 4712 15972
rect 4700 15960 4712 15969
rect 2056 15932 4292 15960
rect 4667 15932 4712 15960
rect 4264 15892 4292 15932
rect 4700 15923 4712 15932
rect 4706 15920 4712 15923
rect 4764 15920 4770 15972
rect 7374 15920 7380 15972
rect 7432 15960 7438 15972
rect 7469 15963 7527 15969
rect 7469 15960 7481 15963
rect 7432 15932 7481 15960
rect 7432 15920 7438 15932
rect 7469 15929 7481 15932
rect 7515 15929 7527 15963
rect 7469 15923 7527 15929
rect 8748 15963 8806 15969
rect 8748 15929 8760 15963
rect 8794 15960 8806 15963
rect 8846 15960 8852 15972
rect 8794 15932 8852 15960
rect 8794 15929 8806 15932
rect 8748 15923 8806 15929
rect 8846 15920 8852 15932
rect 8904 15920 8910 15972
rect 9858 15920 9864 15972
rect 9916 15960 9922 15972
rect 16390 15960 16396 15972
rect 9916 15932 16396 15960
rect 9916 15920 9922 15932
rect 16390 15920 16396 15932
rect 16448 15920 16454 15972
rect 5810 15892 5816 15904
rect 4264 15864 5816 15892
rect 5810 15852 5816 15864
rect 5868 15852 5874 15904
rect 6457 15895 6515 15901
rect 6457 15861 6469 15895
rect 6503 15892 6515 15895
rect 6638 15892 6644 15904
rect 6503 15864 6644 15892
rect 6503 15861 6515 15864
rect 6457 15855 6515 15861
rect 6638 15852 6644 15864
rect 6696 15892 6702 15904
rect 7561 15895 7619 15901
rect 7561 15892 7573 15895
rect 6696 15864 7573 15892
rect 6696 15852 6702 15864
rect 7561 15861 7573 15864
rect 7607 15861 7619 15895
rect 7561 15855 7619 15861
rect 10870 15852 10876 15904
rect 10928 15892 10934 15904
rect 11793 15895 11851 15901
rect 11793 15892 11805 15895
rect 10928 15864 11805 15892
rect 10928 15852 10934 15864
rect 11793 15861 11805 15864
rect 11839 15861 11851 15895
rect 11793 15855 11851 15861
rect 16850 15852 16856 15904
rect 16908 15892 16914 15904
rect 17037 15895 17095 15901
rect 17037 15892 17049 15895
rect 16908 15864 17049 15892
rect 16908 15852 16914 15864
rect 17037 15861 17049 15864
rect 17083 15861 17095 15895
rect 19702 15892 19708 15904
rect 19663 15864 19708 15892
rect 17037 15855 17095 15861
rect 19702 15852 19708 15864
rect 19760 15852 19766 15904
rect 20622 15852 20628 15904
rect 20680 15892 20686 15904
rect 20993 15895 21051 15901
rect 20993 15892 21005 15895
rect 20680 15864 21005 15892
rect 20680 15852 20686 15864
rect 20993 15861 21005 15864
rect 21039 15861 21051 15895
rect 20993 15855 21051 15861
rect 1104 15802 21896 15824
rect 1104 15750 7912 15802
rect 7964 15750 7976 15802
rect 8028 15750 8040 15802
rect 8092 15750 8104 15802
rect 8156 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 15035 15802
rect 15087 15750 21896 15802
rect 1104 15728 21896 15750
rect 1946 15688 1952 15700
rect 1907 15660 1952 15688
rect 1946 15648 1952 15660
rect 2004 15648 2010 15700
rect 4706 15688 4712 15700
rect 3344 15660 4712 15688
rect 1765 15555 1823 15561
rect 1765 15521 1777 15555
rect 1811 15552 1823 15555
rect 2406 15552 2412 15564
rect 1811 15524 2412 15552
rect 1811 15521 1823 15524
rect 1765 15515 1823 15521
rect 2406 15512 2412 15524
rect 2464 15512 2470 15564
rect 3050 15552 3056 15564
rect 3011 15524 3056 15552
rect 3050 15512 3056 15524
rect 3108 15512 3114 15564
rect 2314 15444 2320 15496
rect 2372 15484 2378 15496
rect 3142 15484 3148 15496
rect 2372 15456 3004 15484
rect 3103 15456 3148 15484
rect 2372 15444 2378 15456
rect 1578 15376 1584 15428
rect 1636 15416 1642 15428
rect 2685 15419 2743 15425
rect 2685 15416 2697 15419
rect 1636 15388 2697 15416
rect 1636 15376 1642 15388
rect 2685 15385 2697 15388
rect 2731 15385 2743 15419
rect 2976 15416 3004 15456
rect 3142 15444 3148 15456
rect 3200 15444 3206 15496
rect 3344 15493 3372 15660
rect 4706 15648 4712 15660
rect 4764 15688 4770 15700
rect 5445 15691 5503 15697
rect 5445 15688 5457 15691
rect 4764 15660 5457 15688
rect 4764 15648 4770 15660
rect 5445 15657 5457 15660
rect 5491 15657 5503 15691
rect 5445 15651 5503 15657
rect 6914 15648 6920 15700
rect 6972 15648 6978 15700
rect 8297 15691 8355 15697
rect 8297 15657 8309 15691
rect 8343 15688 8355 15691
rect 8478 15688 8484 15700
rect 8343 15660 8484 15688
rect 8343 15657 8355 15660
rect 8297 15651 8355 15657
rect 8478 15648 8484 15660
rect 8536 15648 8542 15700
rect 13814 15688 13820 15700
rect 13775 15660 13820 15688
rect 13814 15648 13820 15660
rect 13872 15648 13878 15700
rect 14921 15691 14979 15697
rect 14921 15657 14933 15691
rect 14967 15688 14979 15691
rect 15378 15688 15384 15700
rect 14967 15660 15384 15688
rect 14967 15657 14979 15660
rect 14921 15651 14979 15657
rect 15378 15648 15384 15660
rect 15436 15688 15442 15700
rect 18874 15688 18880 15700
rect 15436 15660 18880 15688
rect 15436 15648 15442 15660
rect 18874 15648 18880 15660
rect 18932 15648 18938 15700
rect 19058 15688 19064 15700
rect 19019 15660 19064 15688
rect 19058 15648 19064 15660
rect 19116 15648 19122 15700
rect 20438 15688 20444 15700
rect 20399 15660 20444 15688
rect 20438 15648 20444 15660
rect 20496 15648 20502 15700
rect 21082 15688 21088 15700
rect 21043 15660 21088 15688
rect 21082 15648 21088 15660
rect 21140 15648 21146 15700
rect 4430 15620 4436 15632
rect 4080 15592 4436 15620
rect 4080 15561 4108 15592
rect 4430 15580 4436 15592
rect 4488 15580 4494 15632
rect 6172 15623 6230 15629
rect 6172 15589 6184 15623
rect 6218 15620 6230 15623
rect 6932 15620 6960 15648
rect 6218 15592 6960 15620
rect 11600 15623 11658 15629
rect 6218 15589 6230 15592
rect 6172 15583 6230 15589
rect 11600 15589 11612 15623
rect 11646 15620 11658 15623
rect 12158 15620 12164 15632
rect 11646 15592 12164 15620
rect 11646 15589 11658 15592
rect 11600 15583 11658 15589
rect 12158 15580 12164 15592
rect 12216 15580 12222 15632
rect 15832 15623 15890 15629
rect 15832 15589 15844 15623
rect 15878 15620 15890 15623
rect 16022 15620 16028 15632
rect 15878 15592 16028 15620
rect 15878 15589 15890 15592
rect 15832 15583 15890 15589
rect 16022 15580 16028 15592
rect 16080 15580 16086 15632
rect 4065 15555 4123 15561
rect 4065 15521 4077 15555
rect 4111 15521 4123 15555
rect 4065 15515 4123 15521
rect 3329 15487 3387 15493
rect 3329 15453 3341 15487
rect 3375 15453 3387 15487
rect 3329 15447 3387 15453
rect 4080 15416 4108 15515
rect 4154 15512 4160 15564
rect 4212 15552 4218 15564
rect 4321 15555 4379 15561
rect 4321 15552 4333 15555
rect 4212 15524 4333 15552
rect 4212 15512 4218 15524
rect 4321 15521 4333 15524
rect 4367 15521 4379 15555
rect 4321 15515 4379 15521
rect 5626 15512 5632 15564
rect 5684 15552 5690 15564
rect 5905 15555 5963 15561
rect 5905 15552 5917 15555
rect 5684 15524 5917 15552
rect 5684 15512 5690 15524
rect 5905 15521 5917 15524
rect 5951 15521 5963 15555
rect 5905 15515 5963 15521
rect 6914 15512 6920 15564
rect 6972 15552 6978 15564
rect 8481 15555 8539 15561
rect 8481 15552 8493 15555
rect 6972 15524 8493 15552
rect 6972 15512 6978 15524
rect 8481 15521 8493 15524
rect 8527 15521 8539 15555
rect 8481 15515 8539 15521
rect 11333 15555 11391 15561
rect 11333 15521 11345 15555
rect 11379 15552 11391 15555
rect 11974 15552 11980 15564
rect 11379 15524 11980 15552
rect 11379 15521 11391 15524
rect 11333 15515 11391 15521
rect 11974 15512 11980 15524
rect 12032 15512 12038 15564
rect 14182 15552 14188 15564
rect 14143 15524 14188 15552
rect 14182 15512 14188 15524
rect 14240 15512 14246 15564
rect 15565 15555 15623 15561
rect 15565 15521 15577 15555
rect 15611 15552 15623 15555
rect 15654 15552 15660 15564
rect 15611 15524 15660 15552
rect 15611 15521 15623 15524
rect 15565 15515 15623 15521
rect 15654 15512 15660 15524
rect 15712 15552 15718 15564
rect 17681 15555 17739 15561
rect 17681 15552 17693 15555
rect 15712 15524 17693 15552
rect 15712 15512 15718 15524
rect 17681 15521 17693 15524
rect 17727 15552 17739 15555
rect 17770 15552 17776 15564
rect 17727 15524 17776 15552
rect 17727 15521 17739 15524
rect 17681 15515 17739 15521
rect 17770 15512 17776 15524
rect 17828 15512 17834 15564
rect 17954 15561 17960 15564
rect 17948 15552 17960 15561
rect 17915 15524 17960 15552
rect 17948 15515 17960 15524
rect 17954 15512 17960 15515
rect 18012 15512 18018 15564
rect 19702 15512 19708 15564
rect 19760 15552 19766 15564
rect 20257 15555 20315 15561
rect 20257 15552 20269 15555
rect 19760 15524 20269 15552
rect 19760 15512 19766 15524
rect 20257 15521 20269 15524
rect 20303 15552 20315 15555
rect 20438 15552 20444 15564
rect 20303 15524 20444 15552
rect 20303 15521 20315 15524
rect 20257 15515 20315 15521
rect 20438 15512 20444 15524
rect 20496 15512 20502 15564
rect 20901 15555 20959 15561
rect 20901 15521 20913 15555
rect 20947 15521 20959 15555
rect 20901 15515 20959 15521
rect 13814 15444 13820 15496
rect 13872 15484 13878 15496
rect 14277 15487 14335 15493
rect 14277 15484 14289 15487
rect 13872 15456 14289 15484
rect 13872 15444 13878 15456
rect 14277 15453 14289 15456
rect 14323 15453 14335 15487
rect 14277 15447 14335 15453
rect 14461 15487 14519 15493
rect 14461 15453 14473 15487
rect 14507 15484 14519 15487
rect 14550 15484 14556 15496
rect 14507 15456 14556 15484
rect 14507 15453 14519 15456
rect 14461 15447 14519 15453
rect 14550 15444 14556 15456
rect 14608 15444 14614 15496
rect 19334 15484 19340 15496
rect 19295 15456 19340 15484
rect 19334 15444 19340 15456
rect 19392 15444 19398 15496
rect 20916 15484 20944 15515
rect 19904 15456 20944 15484
rect 7374 15416 7380 15428
rect 2976 15388 4108 15416
rect 6840 15388 7380 15416
rect 2685 15379 2743 15385
rect 6840 15360 6868 15388
rect 7374 15376 7380 15388
rect 7432 15416 7438 15428
rect 7561 15419 7619 15425
rect 7561 15416 7573 15419
rect 7432 15388 7573 15416
rect 7432 15376 7438 15388
rect 7561 15385 7573 15388
rect 7607 15385 7619 15419
rect 7561 15379 7619 15385
rect 12342 15376 12348 15428
rect 12400 15416 12406 15428
rect 12713 15419 12771 15425
rect 12713 15416 12725 15419
rect 12400 15388 12725 15416
rect 12400 15376 12406 15388
rect 12713 15385 12725 15388
rect 12759 15416 12771 15419
rect 15194 15416 15200 15428
rect 12759 15388 15200 15416
rect 12759 15385 12771 15388
rect 12713 15379 12771 15385
rect 15194 15376 15200 15388
rect 15252 15376 15258 15428
rect 19904 15360 19932 15456
rect 2406 15348 2412 15360
rect 2367 15320 2412 15348
rect 2406 15308 2412 15320
rect 2464 15308 2470 15360
rect 6822 15308 6828 15360
rect 6880 15308 6886 15360
rect 7285 15351 7343 15357
rect 7285 15317 7297 15351
rect 7331 15348 7343 15351
rect 7466 15348 7472 15360
rect 7331 15320 7472 15348
rect 7331 15317 7343 15320
rect 7285 15311 7343 15317
rect 7466 15308 7472 15320
rect 7524 15308 7530 15360
rect 16942 15348 16948 15360
rect 16903 15320 16948 15348
rect 16942 15308 16948 15320
rect 17000 15308 17006 15360
rect 19886 15348 19892 15360
rect 19847 15320 19892 15348
rect 19886 15308 19892 15320
rect 19944 15308 19950 15360
rect 1104 15258 21896 15280
rect 1104 15206 4447 15258
rect 4499 15206 4511 15258
rect 4563 15206 4575 15258
rect 4627 15206 4639 15258
rect 4691 15206 11378 15258
rect 11430 15206 11442 15258
rect 11494 15206 11506 15258
rect 11558 15206 11570 15258
rect 11622 15206 18308 15258
rect 18360 15206 18372 15258
rect 18424 15206 18436 15258
rect 18488 15206 18500 15258
rect 18552 15206 21896 15258
rect 1104 15184 21896 15206
rect 5626 15104 5632 15156
rect 5684 15144 5690 15156
rect 6273 15147 6331 15153
rect 6273 15144 6285 15147
rect 5684 15116 6285 15144
rect 5684 15104 5690 15116
rect 6273 15113 6285 15116
rect 6319 15113 6331 15147
rect 6273 15107 6331 15113
rect 8846 15104 8852 15156
rect 8904 15144 8910 15156
rect 11517 15147 11575 15153
rect 11517 15144 11529 15147
rect 8904 15116 11529 15144
rect 8904 15104 8910 15116
rect 11517 15113 11529 15116
rect 11563 15113 11575 15147
rect 11517 15107 11575 15113
rect 11974 15104 11980 15156
rect 12032 15144 12038 15156
rect 12713 15147 12771 15153
rect 12713 15144 12725 15147
rect 12032 15116 12725 15144
rect 12032 15104 12038 15116
rect 12713 15113 12725 15116
rect 12759 15113 12771 15147
rect 12713 15107 12771 15113
rect 12728 15020 12756 15107
rect 16945 15079 17003 15085
rect 16945 15045 16957 15079
rect 16991 15045 17003 15079
rect 16945 15039 17003 15045
rect 8478 15008 8484 15020
rect 8439 14980 8484 15008
rect 8478 14968 8484 14980
rect 8536 14968 8542 15020
rect 9674 14968 9680 15020
rect 9732 15008 9738 15020
rect 10137 15011 10195 15017
rect 10137 15008 10149 15011
rect 9732 14980 10149 15008
rect 9732 14968 9738 14980
rect 10137 14977 10149 14980
rect 10183 14977 10195 15011
rect 12710 15008 12716 15020
rect 12623 14980 12716 15008
rect 10137 14971 10195 14977
rect 12710 14968 12716 14980
rect 12768 15008 12774 15020
rect 13173 15011 13231 15017
rect 13173 15008 13185 15011
rect 12768 14980 13185 15008
rect 12768 14968 12774 14980
rect 13173 14977 13185 14980
rect 13219 14977 13231 15011
rect 13173 14971 13231 14977
rect 15194 14968 15200 15020
rect 15252 15008 15258 15020
rect 15473 15011 15531 15017
rect 15473 15008 15485 15011
rect 15252 14980 15485 15008
rect 15252 14968 15258 14980
rect 15473 14977 15485 14980
rect 15519 15008 15531 15011
rect 15930 15008 15936 15020
rect 15519 14980 15936 15008
rect 15519 14977 15531 14980
rect 15473 14971 15531 14977
rect 15930 14968 15936 14980
rect 15988 14968 15994 15020
rect 1762 14940 1768 14952
rect 1723 14912 1768 14940
rect 1762 14900 1768 14912
rect 1820 14900 1826 14952
rect 2314 14900 2320 14952
rect 2372 14940 2378 14952
rect 2501 14943 2559 14949
rect 2501 14940 2513 14943
rect 2372 14912 2513 14940
rect 2372 14900 2378 14912
rect 2501 14909 2513 14912
rect 2547 14909 2559 14943
rect 2501 14903 2559 14909
rect 6457 14943 6515 14949
rect 6457 14909 6469 14943
rect 6503 14909 6515 14943
rect 6457 14903 6515 14909
rect 6825 14943 6883 14949
rect 6825 14909 6837 14943
rect 6871 14940 6883 14943
rect 8496 14940 8524 14968
rect 6871 14912 8524 14940
rect 6871 14909 6883 14912
rect 6825 14903 6883 14909
rect 2774 14881 2780 14884
rect 2768 14835 2780 14881
rect 2832 14872 2838 14884
rect 6472 14872 6500 14903
rect 9858 14900 9864 14952
rect 9916 14940 9922 14952
rect 10393 14943 10451 14949
rect 10393 14940 10405 14943
rect 9916 14912 10405 14940
rect 9916 14900 9922 14912
rect 10393 14909 10405 14912
rect 10439 14909 10451 14943
rect 10393 14903 10451 14909
rect 12897 14943 12955 14949
rect 12897 14909 12909 14943
rect 12943 14909 12955 14943
rect 12897 14903 12955 14909
rect 15289 14943 15347 14949
rect 15289 14909 15301 14943
rect 15335 14940 15347 14943
rect 15378 14940 15384 14952
rect 15335 14912 15384 14940
rect 15335 14909 15347 14912
rect 15289 14903 15347 14909
rect 6914 14872 6920 14884
rect 2832 14844 2868 14872
rect 6472 14844 6920 14872
rect 2774 14832 2780 14835
rect 2832 14832 2838 14844
rect 6914 14832 6920 14844
rect 6972 14832 6978 14884
rect 7092 14875 7150 14881
rect 7092 14841 7104 14875
rect 7138 14872 7150 14875
rect 7466 14872 7472 14884
rect 7138 14844 7472 14872
rect 7138 14841 7150 14844
rect 7092 14835 7150 14841
rect 7466 14832 7472 14844
rect 7524 14832 7530 14884
rect 8726 14875 8784 14881
rect 8726 14872 8738 14875
rect 8220 14844 8738 14872
rect 1946 14804 1952 14816
rect 1907 14776 1952 14804
rect 1946 14764 1952 14776
rect 2004 14764 2010 14816
rect 3878 14804 3884 14816
rect 3839 14776 3884 14804
rect 3878 14764 3884 14776
rect 3936 14804 3942 14816
rect 4154 14804 4160 14816
rect 3936 14776 4160 14804
rect 3936 14764 3942 14776
rect 4154 14764 4160 14776
rect 4212 14764 4218 14816
rect 6454 14764 6460 14816
rect 6512 14804 6518 14816
rect 8220 14813 8248 14844
rect 8726 14841 8738 14844
rect 8772 14841 8784 14875
rect 8726 14835 8784 14841
rect 8205 14807 8263 14813
rect 8205 14804 8217 14807
rect 6512 14776 8217 14804
rect 6512 14764 6518 14776
rect 8205 14773 8217 14776
rect 8251 14773 8263 14807
rect 8205 14767 8263 14773
rect 9861 14807 9919 14813
rect 9861 14773 9873 14807
rect 9907 14804 9919 14807
rect 10226 14804 10232 14816
rect 9907 14776 10232 14804
rect 9907 14773 9919 14776
rect 9861 14767 9919 14773
rect 10226 14764 10232 14776
rect 10284 14764 10290 14816
rect 12912 14804 12940 14903
rect 15378 14900 15384 14912
rect 15436 14900 15442 14952
rect 16960 14940 16988 15039
rect 19058 15036 19064 15088
rect 19116 15076 19122 15088
rect 19116 15048 20392 15076
rect 19116 15036 19122 15048
rect 17589 15011 17647 15017
rect 17589 14977 17601 15011
rect 17635 15008 17647 15011
rect 17954 15008 17960 15020
rect 17635 14980 17960 15008
rect 17635 14977 17647 14980
rect 17589 14971 17647 14977
rect 17954 14968 17960 14980
rect 18012 15008 18018 15020
rect 18782 15008 18788 15020
rect 18012 14980 18788 15008
rect 18012 14968 18018 14980
rect 18782 14968 18788 14980
rect 18840 14968 18846 15020
rect 19242 14968 19248 15020
rect 19300 15008 19306 15020
rect 20364 15017 20392 15048
rect 19337 15011 19395 15017
rect 19337 15008 19349 15011
rect 19300 14980 19349 15008
rect 19300 14968 19306 14980
rect 19337 14977 19349 14980
rect 19383 14977 19395 15011
rect 19337 14971 19395 14977
rect 20349 15011 20407 15017
rect 20349 14977 20361 15011
rect 20395 14977 20407 15011
rect 20349 14971 20407 14977
rect 20165 14943 20223 14949
rect 20165 14940 20177 14943
rect 16960 14912 20177 14940
rect 20165 14909 20177 14912
rect 20211 14909 20223 14943
rect 20806 14940 20812 14952
rect 20767 14912 20812 14940
rect 20165 14903 20223 14909
rect 20806 14900 20812 14912
rect 20864 14900 20870 14952
rect 13446 14881 13452 14884
rect 13440 14872 13452 14881
rect 13407 14844 13452 14872
rect 13440 14835 13452 14844
rect 13446 14832 13452 14835
rect 13504 14832 13510 14884
rect 17313 14875 17371 14881
rect 17313 14841 17325 14875
rect 17359 14872 17371 14875
rect 19153 14875 19211 14881
rect 17359 14844 18828 14872
rect 17359 14841 17371 14844
rect 17313 14835 17371 14841
rect 13906 14804 13912 14816
rect 12912 14776 13912 14804
rect 13906 14764 13912 14776
rect 13964 14764 13970 14816
rect 14550 14804 14556 14816
rect 14511 14776 14556 14804
rect 14550 14764 14556 14776
rect 14608 14764 14614 14816
rect 14734 14764 14740 14816
rect 14792 14804 14798 14816
rect 14829 14807 14887 14813
rect 14829 14804 14841 14807
rect 14792 14776 14841 14804
rect 14792 14764 14798 14776
rect 14829 14773 14841 14776
rect 14875 14773 14887 14807
rect 15194 14804 15200 14816
rect 15155 14776 15200 14804
rect 14829 14767 14887 14773
rect 15194 14764 15200 14776
rect 15252 14764 15258 14816
rect 15838 14764 15844 14816
rect 15896 14804 15902 14816
rect 18800 14813 18828 14844
rect 19153 14841 19165 14875
rect 19199 14872 19211 14875
rect 19334 14872 19340 14884
rect 19199 14844 19340 14872
rect 19199 14841 19211 14844
rect 19153 14835 19211 14841
rect 19334 14832 19340 14844
rect 19392 14832 19398 14884
rect 17405 14807 17463 14813
rect 17405 14804 17417 14807
rect 15896 14776 17417 14804
rect 15896 14764 15902 14776
rect 17405 14773 17417 14776
rect 17451 14773 17463 14807
rect 17405 14767 17463 14773
rect 18785 14807 18843 14813
rect 18785 14773 18797 14807
rect 18831 14773 18843 14807
rect 18785 14767 18843 14773
rect 19245 14807 19303 14813
rect 19245 14773 19257 14807
rect 19291 14804 19303 14807
rect 19426 14804 19432 14816
rect 19291 14776 19432 14804
rect 19291 14773 19303 14776
rect 19245 14767 19303 14773
rect 19426 14764 19432 14776
rect 19484 14764 19490 14816
rect 19797 14807 19855 14813
rect 19797 14773 19809 14807
rect 19843 14804 19855 14807
rect 20070 14804 20076 14816
rect 19843 14776 20076 14804
rect 19843 14773 19855 14776
rect 19797 14767 19855 14773
rect 20070 14764 20076 14776
rect 20128 14764 20134 14816
rect 20254 14804 20260 14816
rect 20215 14776 20260 14804
rect 20254 14764 20260 14776
rect 20312 14764 20318 14816
rect 20990 14804 20996 14816
rect 20951 14776 20996 14804
rect 20990 14764 20996 14776
rect 21048 14764 21054 14816
rect 1104 14714 21896 14736
rect 1104 14662 7912 14714
rect 7964 14662 7976 14714
rect 8028 14662 8040 14714
rect 8092 14662 8104 14714
rect 8156 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 15035 14714
rect 15087 14662 21896 14714
rect 1104 14640 21896 14662
rect 2317 14603 2375 14609
rect 2317 14569 2329 14603
rect 2363 14600 2375 14603
rect 3050 14600 3056 14612
rect 2363 14572 3056 14600
rect 2363 14569 2375 14572
rect 2317 14563 2375 14569
rect 3050 14560 3056 14572
rect 3108 14560 3114 14612
rect 3142 14560 3148 14612
rect 3200 14600 3206 14612
rect 4065 14603 4123 14609
rect 4065 14600 4077 14603
rect 3200 14572 4077 14600
rect 3200 14560 3206 14572
rect 4065 14569 4077 14572
rect 4111 14569 4123 14603
rect 5810 14600 5816 14612
rect 5771 14572 5816 14600
rect 4065 14563 4123 14569
rect 5810 14560 5816 14572
rect 5868 14560 5874 14612
rect 6273 14603 6331 14609
rect 6273 14569 6285 14603
rect 6319 14600 6331 14603
rect 6825 14603 6883 14609
rect 6825 14600 6837 14603
rect 6319 14572 6837 14600
rect 6319 14569 6331 14572
rect 6273 14563 6331 14569
rect 6825 14569 6837 14572
rect 6871 14569 6883 14603
rect 6825 14563 6883 14569
rect 7650 14560 7656 14612
rect 7708 14600 7714 14612
rect 7929 14603 7987 14609
rect 7929 14600 7941 14603
rect 7708 14572 7941 14600
rect 7708 14560 7714 14572
rect 7929 14569 7941 14572
rect 7975 14569 7987 14603
rect 7929 14563 7987 14569
rect 13633 14603 13691 14609
rect 13633 14569 13645 14603
rect 13679 14600 13691 14603
rect 14182 14600 14188 14612
rect 13679 14572 14188 14600
rect 13679 14569 13691 14572
rect 13633 14563 13691 14569
rect 14182 14560 14188 14572
rect 14240 14560 14246 14612
rect 14645 14603 14703 14609
rect 14645 14569 14657 14603
rect 14691 14600 14703 14603
rect 15194 14600 15200 14612
rect 14691 14572 15200 14600
rect 14691 14569 14703 14572
rect 14645 14563 14703 14569
rect 15194 14560 15200 14572
rect 15252 14560 15258 14612
rect 19426 14600 19432 14612
rect 19387 14572 19432 14600
rect 19426 14560 19432 14572
rect 19484 14560 19490 14612
rect 1762 14492 1768 14544
rect 1820 14532 1826 14544
rect 1857 14535 1915 14541
rect 1857 14532 1869 14535
rect 1820 14504 1869 14532
rect 1820 14492 1826 14504
rect 1857 14501 1869 14504
rect 1903 14501 1915 14535
rect 1857 14495 1915 14501
rect 7193 14535 7251 14541
rect 7193 14501 7205 14535
rect 7239 14532 7251 14535
rect 7374 14532 7380 14544
rect 7239 14504 7380 14532
rect 7239 14501 7251 14504
rect 7193 14495 7251 14501
rect 7374 14492 7380 14504
rect 7432 14492 7438 14544
rect 12244 14535 12302 14541
rect 12244 14501 12256 14535
rect 12290 14532 12302 14535
rect 12342 14532 12348 14544
rect 12290 14504 12348 14532
rect 12290 14501 12302 14504
rect 12244 14495 12302 14501
rect 12342 14492 12348 14504
rect 12400 14492 12406 14544
rect 14001 14535 14059 14541
rect 14001 14501 14013 14535
rect 14047 14532 14059 14535
rect 14734 14532 14740 14544
rect 14047 14504 14740 14532
rect 14047 14501 14059 14504
rect 14001 14495 14059 14501
rect 14734 14492 14740 14504
rect 14792 14492 14798 14544
rect 17954 14492 17960 14544
rect 18012 14532 18018 14544
rect 19061 14535 19119 14541
rect 19061 14532 19073 14535
rect 18012 14504 19073 14532
rect 18012 14492 18018 14504
rect 19061 14501 19073 14504
rect 19107 14532 19119 14535
rect 19797 14535 19855 14541
rect 19797 14532 19809 14535
rect 19107 14504 19809 14532
rect 19107 14501 19119 14504
rect 19061 14495 19119 14501
rect 19797 14501 19809 14504
rect 19843 14532 19855 14535
rect 20714 14532 20720 14544
rect 19843 14504 20720 14532
rect 19843 14501 19855 14504
rect 19797 14495 19855 14501
rect 20714 14492 20720 14504
rect 20772 14492 20778 14544
rect 20806 14492 20812 14544
rect 20864 14532 20870 14544
rect 21177 14535 21235 14541
rect 21177 14532 21189 14535
rect 20864 14504 21189 14532
rect 20864 14492 20870 14504
rect 21177 14501 21189 14504
rect 21223 14501 21235 14535
rect 21177 14495 21235 14501
rect 1578 14464 1584 14476
rect 1539 14436 1584 14464
rect 1578 14424 1584 14436
rect 1636 14424 1642 14476
rect 2222 14424 2228 14476
rect 2280 14464 2286 14476
rect 2685 14467 2743 14473
rect 2685 14464 2697 14467
rect 2280 14436 2697 14464
rect 2280 14424 2286 14436
rect 2685 14433 2697 14436
rect 2731 14433 2743 14467
rect 2685 14427 2743 14433
rect 4154 14424 4160 14476
rect 4212 14464 4218 14476
rect 4433 14467 4491 14473
rect 4433 14464 4445 14467
rect 4212 14436 4445 14464
rect 4212 14424 4218 14436
rect 4433 14433 4445 14436
rect 4479 14433 4491 14467
rect 6178 14464 6184 14476
rect 6139 14436 6184 14464
rect 4433 14427 4491 14433
rect 6178 14424 6184 14436
rect 6236 14424 6242 14476
rect 9674 14464 9680 14476
rect 9635 14436 9680 14464
rect 9674 14424 9680 14436
rect 9732 14424 9738 14476
rect 9944 14467 10002 14473
rect 9944 14433 9956 14467
rect 9990 14464 10002 14467
rect 10226 14464 10232 14476
rect 9990 14436 10232 14464
rect 9990 14433 10002 14436
rect 9944 14427 10002 14433
rect 10226 14424 10232 14436
rect 10284 14424 10290 14476
rect 11974 14464 11980 14476
rect 11935 14436 11980 14464
rect 11974 14424 11980 14436
rect 12032 14424 12038 14476
rect 15194 14424 15200 14476
rect 15252 14464 15258 14476
rect 15378 14464 15384 14476
rect 15252 14436 15384 14464
rect 15252 14424 15258 14436
rect 15378 14424 15384 14436
rect 15436 14424 15442 14476
rect 15654 14424 15660 14476
rect 15712 14464 15718 14476
rect 16005 14467 16063 14473
rect 16005 14464 16017 14467
rect 15712 14436 16017 14464
rect 15712 14424 15718 14436
rect 16005 14433 16017 14436
rect 16051 14433 16063 14467
rect 17672 14467 17730 14473
rect 17672 14464 17684 14467
rect 16005 14427 16063 14433
rect 17144 14436 17684 14464
rect 2498 14356 2504 14408
rect 2556 14396 2562 14408
rect 2777 14399 2835 14405
rect 2777 14396 2789 14399
rect 2556 14368 2789 14396
rect 2556 14356 2562 14368
rect 2777 14365 2789 14368
rect 2823 14365 2835 14399
rect 2777 14359 2835 14365
rect 2961 14399 3019 14405
rect 2961 14365 2973 14399
rect 3007 14396 3019 14399
rect 3878 14396 3884 14408
rect 3007 14368 3884 14396
rect 3007 14365 3019 14368
rect 2961 14359 3019 14365
rect 3878 14356 3884 14368
rect 3936 14356 3942 14408
rect 4062 14356 4068 14408
rect 4120 14396 4126 14408
rect 4525 14399 4583 14405
rect 4525 14396 4537 14399
rect 4120 14368 4537 14396
rect 4120 14356 4126 14368
rect 4525 14365 4537 14368
rect 4571 14365 4583 14399
rect 4525 14359 4583 14365
rect 4617 14399 4675 14405
rect 4617 14365 4629 14399
rect 4663 14365 4675 14399
rect 6454 14396 6460 14408
rect 6415 14368 6460 14396
rect 4617 14359 4675 14365
rect 3896 14328 3924 14356
rect 4632 14328 4660 14359
rect 6454 14356 6460 14368
rect 6512 14356 6518 14408
rect 7098 14356 7104 14408
rect 7156 14396 7162 14408
rect 7285 14399 7343 14405
rect 7285 14396 7297 14399
rect 7156 14368 7297 14396
rect 7156 14356 7162 14368
rect 7285 14365 7297 14368
rect 7331 14365 7343 14399
rect 7466 14396 7472 14408
rect 7427 14368 7472 14396
rect 7285 14359 7343 14365
rect 7466 14356 7472 14368
rect 7524 14356 7530 14408
rect 14090 14396 14096 14408
rect 14051 14368 14096 14396
rect 14090 14356 14096 14368
rect 14148 14356 14154 14408
rect 14277 14399 14335 14405
rect 14277 14365 14289 14399
rect 14323 14396 14335 14399
rect 14366 14396 14372 14408
rect 14323 14368 14372 14396
rect 14323 14365 14335 14368
rect 14277 14359 14335 14365
rect 3896 14300 4660 14328
rect 13357 14331 13415 14337
rect 13357 14297 13369 14331
rect 13403 14328 13415 14331
rect 13446 14328 13452 14340
rect 13403 14300 13452 14328
rect 13403 14297 13415 14300
rect 13357 14291 13415 14297
rect 13446 14288 13452 14300
rect 13504 14328 13510 14340
rect 14292 14328 14320 14359
rect 14366 14356 14372 14368
rect 14424 14356 14430 14408
rect 15746 14396 15752 14408
rect 15707 14368 15752 14396
rect 15746 14356 15752 14368
rect 15804 14356 15810 14408
rect 13504 14300 14320 14328
rect 13504 14288 13510 14300
rect 16758 14288 16764 14340
rect 16816 14328 16822 14340
rect 17144 14337 17172 14436
rect 17672 14433 17684 14436
rect 17718 14464 17730 14467
rect 19242 14464 19248 14476
rect 17718 14436 19248 14464
rect 17718 14433 17730 14436
rect 17672 14427 17730 14433
rect 19242 14424 19248 14436
rect 19300 14424 19306 14476
rect 19702 14424 19708 14476
rect 19760 14464 19766 14476
rect 19760 14436 20024 14464
rect 19760 14424 19766 14436
rect 19996 14405 20024 14436
rect 20070 14424 20076 14476
rect 20128 14464 20134 14476
rect 20901 14467 20959 14473
rect 20901 14464 20913 14467
rect 20128 14436 20913 14464
rect 20128 14424 20134 14436
rect 20901 14433 20913 14436
rect 20947 14433 20959 14467
rect 20901 14427 20959 14433
rect 17405 14399 17463 14405
rect 17405 14365 17417 14399
rect 17451 14365 17463 14399
rect 17405 14359 17463 14365
rect 19889 14399 19947 14405
rect 19889 14365 19901 14399
rect 19935 14365 19947 14399
rect 19889 14359 19947 14365
rect 19981 14399 20039 14405
rect 19981 14365 19993 14399
rect 20027 14365 20039 14399
rect 19981 14359 20039 14365
rect 17129 14331 17187 14337
rect 17129 14328 17141 14331
rect 16816 14300 17141 14328
rect 16816 14288 16822 14300
rect 17129 14297 17141 14300
rect 17175 14297 17187 14331
rect 17129 14291 17187 14297
rect 5169 14263 5227 14269
rect 5169 14229 5181 14263
rect 5215 14260 5227 14263
rect 5258 14260 5264 14272
rect 5215 14232 5264 14260
rect 5215 14229 5227 14232
rect 5169 14223 5227 14229
rect 5258 14220 5264 14232
rect 5316 14220 5322 14272
rect 9858 14220 9864 14272
rect 9916 14260 9922 14272
rect 11057 14263 11115 14269
rect 11057 14260 11069 14263
rect 9916 14232 11069 14260
rect 9916 14220 9922 14232
rect 11057 14229 11069 14232
rect 11103 14229 11115 14263
rect 11057 14223 11115 14229
rect 15746 14220 15752 14272
rect 15804 14260 15810 14272
rect 17420 14260 17448 14359
rect 19904 14328 19932 14359
rect 19904 14300 20208 14328
rect 20180 14272 20208 14300
rect 18782 14260 18788 14272
rect 15804 14232 17448 14260
rect 18743 14232 18788 14260
rect 15804 14220 15810 14232
rect 18782 14220 18788 14232
rect 18840 14220 18846 14272
rect 20162 14220 20168 14272
rect 20220 14260 20226 14272
rect 20438 14260 20444 14272
rect 20220 14232 20444 14260
rect 20220 14220 20226 14232
rect 20438 14220 20444 14232
rect 20496 14220 20502 14272
rect 1104 14170 21896 14192
rect 1104 14118 4447 14170
rect 4499 14118 4511 14170
rect 4563 14118 4575 14170
rect 4627 14118 4639 14170
rect 4691 14118 11378 14170
rect 11430 14118 11442 14170
rect 11494 14118 11506 14170
rect 11558 14118 11570 14170
rect 11622 14118 18308 14170
rect 18360 14118 18372 14170
rect 18424 14118 18436 14170
rect 18488 14118 18500 14170
rect 18552 14118 21896 14170
rect 1104 14096 21896 14118
rect 1854 14056 1860 14068
rect 1815 14028 1860 14056
rect 1854 14016 1860 14028
rect 1912 14016 1918 14068
rect 2222 14056 2228 14068
rect 2183 14028 2228 14056
rect 2222 14016 2228 14028
rect 2280 14016 2286 14068
rect 4062 14056 4068 14068
rect 4023 14028 4068 14056
rect 4062 14016 4068 14028
rect 4120 14016 4126 14068
rect 7098 14056 7104 14068
rect 7059 14028 7104 14056
rect 7098 14016 7104 14028
rect 7156 14016 7162 14068
rect 8294 14056 8300 14068
rect 8255 14028 8300 14056
rect 8294 14016 8300 14028
rect 8352 14016 8358 14068
rect 11333 14059 11391 14065
rect 11333 14025 11345 14059
rect 11379 14056 11391 14059
rect 14090 14056 14096 14068
rect 11379 14028 14096 14056
rect 11379 14025 11391 14028
rect 11333 14019 11391 14025
rect 14090 14016 14096 14028
rect 14148 14016 14154 14068
rect 15838 14056 15844 14068
rect 15799 14028 15844 14056
rect 15838 14016 15844 14028
rect 15896 14016 15902 14068
rect 18046 14016 18052 14068
rect 18104 14056 18110 14068
rect 18509 14059 18567 14065
rect 18509 14056 18521 14059
rect 18104 14028 18521 14056
rect 18104 14016 18110 14028
rect 18509 14025 18521 14028
rect 18555 14025 18567 14059
rect 18509 14019 18567 14025
rect 19889 14059 19947 14065
rect 19889 14025 19901 14059
rect 19935 14056 19947 14059
rect 20254 14056 20260 14068
rect 19935 14028 20260 14056
rect 19935 14025 19947 14028
rect 19889 14019 19947 14025
rect 20254 14016 20260 14028
rect 20312 14016 20318 14068
rect 21082 14056 21088 14068
rect 21043 14028 21088 14056
rect 21082 14016 21088 14028
rect 21140 14016 21146 14068
rect 13814 13988 13820 14000
rect 13775 13960 13820 13988
rect 13814 13948 13820 13960
rect 13872 13948 13878 14000
rect 13906 13948 13912 14000
rect 13964 13988 13970 14000
rect 18138 13988 18144 14000
rect 13964 13960 15608 13988
rect 18099 13960 18144 13988
rect 13964 13948 13970 13960
rect 2774 13880 2780 13932
rect 2832 13920 2838 13932
rect 2958 13920 2964 13932
rect 2832 13892 2964 13920
rect 2832 13880 2838 13892
rect 2958 13880 2964 13892
rect 3016 13920 3022 13932
rect 4617 13923 4675 13929
rect 4617 13920 4629 13923
rect 3016 13892 4629 13920
rect 3016 13880 3022 13892
rect 4617 13889 4629 13892
rect 4663 13889 4675 13923
rect 4617 13883 4675 13889
rect 5166 13880 5172 13932
rect 5224 13920 5230 13932
rect 5629 13923 5687 13929
rect 5629 13920 5641 13923
rect 5224 13892 5641 13920
rect 5224 13880 5230 13892
rect 5629 13889 5641 13892
rect 5675 13889 5687 13923
rect 5629 13883 5687 13889
rect 5994 13880 6000 13932
rect 6052 13920 6058 13932
rect 6052 13892 6960 13920
rect 6052 13880 6058 13892
rect 1673 13855 1731 13861
rect 1673 13821 1685 13855
rect 1719 13852 1731 13855
rect 2130 13852 2136 13864
rect 1719 13824 2136 13852
rect 1719 13821 1731 13824
rect 1673 13815 1731 13821
rect 2130 13812 2136 13824
rect 2188 13812 2194 13864
rect 6932 13852 6960 13892
rect 7006 13880 7012 13932
rect 7064 13920 7070 13932
rect 7653 13923 7711 13929
rect 7653 13920 7665 13923
rect 7064 13892 7665 13920
rect 7064 13880 7070 13892
rect 7653 13889 7665 13892
rect 7699 13920 7711 13923
rect 8202 13920 8208 13932
rect 7699 13892 8208 13920
rect 7699 13889 7711 13892
rect 7653 13883 7711 13889
rect 8202 13880 8208 13892
rect 8260 13880 8266 13932
rect 8846 13920 8852 13932
rect 8807 13892 8852 13920
rect 8846 13880 8852 13892
rect 8904 13880 8910 13932
rect 9858 13920 9864 13932
rect 9819 13892 9864 13920
rect 9858 13880 9864 13892
rect 9916 13880 9922 13932
rect 10318 13880 10324 13932
rect 10376 13920 10382 13932
rect 10376 13892 11100 13920
rect 10376 13880 10382 13892
rect 7561 13855 7619 13861
rect 7561 13852 7573 13855
rect 6932 13824 7573 13852
rect 7561 13821 7573 13824
rect 7607 13852 7619 13855
rect 8294 13852 8300 13864
rect 7607 13824 8300 13852
rect 7607 13821 7619 13824
rect 7561 13815 7619 13821
rect 8294 13812 8300 13824
rect 8352 13812 8358 13864
rect 10410 13812 10416 13864
rect 10468 13852 10474 13864
rect 11072 13861 11100 13892
rect 11790 13880 11796 13932
rect 11848 13920 11854 13932
rect 11977 13923 12035 13929
rect 11977 13920 11989 13923
rect 11848 13892 11989 13920
rect 11848 13880 11854 13892
rect 11977 13889 11989 13892
rect 12023 13920 12035 13923
rect 12342 13920 12348 13932
rect 12023 13892 12348 13920
rect 12023 13889 12035 13892
rect 11977 13883 12035 13889
rect 12342 13880 12348 13892
rect 12400 13880 12406 13932
rect 14366 13920 14372 13932
rect 14327 13892 14372 13920
rect 14366 13880 14372 13892
rect 14424 13880 14430 13932
rect 10597 13855 10655 13861
rect 10597 13852 10609 13855
rect 10468 13824 10609 13852
rect 10468 13812 10474 13824
rect 10597 13821 10609 13824
rect 10643 13821 10655 13855
rect 10597 13815 10655 13821
rect 11057 13855 11115 13861
rect 11057 13821 11069 13855
rect 11103 13852 11115 13855
rect 11698 13852 11704 13864
rect 11103 13824 11704 13852
rect 11103 13821 11115 13824
rect 11057 13815 11115 13821
rect 2593 13787 2651 13793
rect 2593 13753 2605 13787
rect 2639 13784 2651 13787
rect 3237 13787 3295 13793
rect 3237 13784 3249 13787
rect 2639 13756 3249 13784
rect 2639 13753 2651 13756
rect 2593 13747 2651 13753
rect 3237 13753 3249 13756
rect 3283 13753 3295 13787
rect 3237 13747 3295 13753
rect 4433 13787 4491 13793
rect 4433 13753 4445 13787
rect 4479 13784 4491 13787
rect 5445 13787 5503 13793
rect 4479 13756 5120 13784
rect 4479 13753 4491 13756
rect 4433 13747 4491 13753
rect 2682 13716 2688 13728
rect 2643 13688 2688 13716
rect 2682 13676 2688 13688
rect 2740 13676 2746 13728
rect 4522 13676 4528 13728
rect 4580 13716 4586 13728
rect 5092 13725 5120 13756
rect 5445 13753 5457 13787
rect 5491 13784 5503 13787
rect 6181 13787 6239 13793
rect 6181 13784 6193 13787
rect 5491 13756 6193 13784
rect 5491 13753 5503 13756
rect 5445 13747 5503 13753
rect 6181 13753 6193 13756
rect 6227 13784 6239 13787
rect 6362 13784 6368 13796
rect 6227 13756 6368 13784
rect 6227 13753 6239 13756
rect 6181 13747 6239 13753
rect 6362 13744 6368 13756
rect 6420 13744 6426 13796
rect 10612 13784 10640 13815
rect 11698 13812 11704 13824
rect 11756 13812 11762 13864
rect 14277 13855 14335 13861
rect 14277 13821 14289 13855
rect 14323 13852 14335 13855
rect 15286 13852 15292 13864
rect 14323 13824 15292 13852
rect 14323 13821 14335 13824
rect 14277 13815 14335 13821
rect 15286 13812 15292 13824
rect 15344 13812 15350 13864
rect 15580 13861 15608 13960
rect 18138 13948 18144 13960
rect 18196 13948 18202 14000
rect 18877 13991 18935 13997
rect 18877 13957 18889 13991
rect 18923 13988 18935 13991
rect 18923 13960 20392 13988
rect 18923 13957 18935 13960
rect 18877 13951 18935 13957
rect 16485 13923 16543 13929
rect 16485 13889 16497 13923
rect 16531 13920 16543 13923
rect 16758 13920 16764 13932
rect 16531 13892 16764 13920
rect 16531 13889 16543 13892
rect 16485 13883 16543 13889
rect 16758 13880 16764 13892
rect 16816 13880 16822 13932
rect 18156 13920 18184 13948
rect 18966 13920 18972 13932
rect 18156 13892 18972 13920
rect 18966 13880 18972 13892
rect 19024 13880 19030 13932
rect 19242 13880 19248 13932
rect 19300 13920 19306 13932
rect 20364 13929 20392 13960
rect 19429 13923 19487 13929
rect 19429 13920 19441 13923
rect 19300 13892 19441 13920
rect 19300 13880 19306 13892
rect 19429 13889 19441 13892
rect 19475 13889 19487 13923
rect 19429 13883 19487 13889
rect 20349 13923 20407 13929
rect 20349 13889 20361 13923
rect 20395 13889 20407 13923
rect 20349 13883 20407 13889
rect 20441 13923 20499 13929
rect 20441 13889 20453 13923
rect 20487 13889 20499 13923
rect 20441 13883 20499 13889
rect 15565 13855 15623 13861
rect 15565 13821 15577 13855
rect 15611 13821 15623 13855
rect 15565 13815 15623 13821
rect 18782 13812 18788 13864
rect 18840 13852 18846 13864
rect 20456 13852 20484 13883
rect 18840 13824 20484 13852
rect 18840 13812 18846 13824
rect 20806 13812 20812 13864
rect 20864 13852 20870 13864
rect 20901 13855 20959 13861
rect 20901 13852 20913 13855
rect 20864 13824 20913 13852
rect 20864 13812 20870 13824
rect 20901 13821 20913 13824
rect 20947 13821 20959 13855
rect 20901 13815 20959 13821
rect 11793 13787 11851 13793
rect 11793 13784 11805 13787
rect 7392 13756 9996 13784
rect 10612 13756 11805 13784
rect 5077 13719 5135 13725
rect 4580 13688 4625 13716
rect 4580 13676 4586 13688
rect 5077 13685 5089 13719
rect 5123 13685 5135 13719
rect 5077 13679 5135 13685
rect 5258 13676 5264 13728
rect 5316 13716 5322 13728
rect 5537 13719 5595 13725
rect 5537 13716 5549 13719
rect 5316 13688 5549 13716
rect 5316 13676 5322 13688
rect 5537 13685 5549 13688
rect 5583 13716 5595 13719
rect 7392 13716 7420 13756
rect 5583 13688 7420 13716
rect 7469 13719 7527 13725
rect 5583 13685 5595 13688
rect 5537 13679 5595 13685
rect 7469 13685 7481 13719
rect 7515 13716 7527 13719
rect 7650 13716 7656 13728
rect 7515 13688 7656 13716
rect 7515 13685 7527 13688
rect 7469 13679 7527 13685
rect 7650 13676 7656 13688
rect 7708 13676 7714 13728
rect 8662 13716 8668 13728
rect 8623 13688 8668 13716
rect 8662 13676 8668 13688
rect 8720 13676 8726 13728
rect 8757 13719 8815 13725
rect 8757 13685 8769 13719
rect 8803 13716 8815 13719
rect 9309 13719 9367 13725
rect 9309 13716 9321 13719
rect 8803 13688 9321 13716
rect 8803 13685 8815 13688
rect 8757 13679 8815 13685
rect 9309 13685 9321 13688
rect 9355 13685 9367 13719
rect 9674 13716 9680 13728
rect 9635 13688 9680 13716
rect 9309 13679 9367 13685
rect 9674 13676 9680 13688
rect 9732 13676 9738 13728
rect 9766 13676 9772 13728
rect 9824 13716 9830 13728
rect 9968 13716 9996 13756
rect 11793 13753 11805 13756
rect 11839 13753 11851 13787
rect 11793 13747 11851 13753
rect 11882 13744 11888 13796
rect 11940 13784 11946 13796
rect 15470 13784 15476 13796
rect 11940 13756 15476 13784
rect 11940 13744 11946 13756
rect 15470 13744 15476 13756
rect 15528 13744 15534 13796
rect 19245 13787 19303 13793
rect 19245 13753 19257 13787
rect 19291 13784 19303 13787
rect 19426 13784 19432 13796
rect 19291 13756 19432 13784
rect 19291 13753 19303 13756
rect 19245 13747 19303 13753
rect 19426 13744 19432 13756
rect 19484 13744 19490 13796
rect 19978 13744 19984 13796
rect 20036 13784 20042 13796
rect 20438 13784 20444 13796
rect 20036 13756 20444 13784
rect 20036 13744 20042 13756
rect 20438 13744 20444 13756
rect 20496 13744 20502 13796
rect 11146 13716 11152 13728
rect 9824 13688 9869 13716
rect 9968 13688 11152 13716
rect 9824 13676 9830 13688
rect 11146 13676 11152 13688
rect 11204 13676 11210 13728
rect 14182 13716 14188 13728
rect 14143 13688 14188 13716
rect 14182 13676 14188 13688
rect 14240 13676 14246 13728
rect 15381 13719 15439 13725
rect 15381 13685 15393 13719
rect 15427 13716 15439 13719
rect 15838 13716 15844 13728
rect 15427 13688 15844 13716
rect 15427 13685 15439 13688
rect 15381 13679 15439 13685
rect 15838 13676 15844 13688
rect 15896 13676 15902 13728
rect 16206 13716 16212 13728
rect 16167 13688 16212 13716
rect 16206 13676 16212 13688
rect 16264 13676 16270 13728
rect 16298 13676 16304 13728
rect 16356 13716 16362 13728
rect 17218 13716 17224 13728
rect 16356 13688 16401 13716
rect 17179 13688 17224 13716
rect 16356 13676 16362 13688
rect 17218 13676 17224 13688
rect 17276 13676 17282 13728
rect 19334 13716 19340 13728
rect 19295 13688 19340 13716
rect 19334 13676 19340 13688
rect 19392 13676 19398 13728
rect 20254 13716 20260 13728
rect 20215 13688 20260 13716
rect 20254 13676 20260 13688
rect 20312 13676 20318 13728
rect 1104 13626 21896 13648
rect 1104 13574 7912 13626
rect 7964 13574 7976 13626
rect 8028 13574 8040 13626
rect 8092 13574 8104 13626
rect 8156 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 15035 13626
rect 15087 13574 21896 13626
rect 1104 13552 21896 13574
rect 2409 13515 2467 13521
rect 2409 13481 2421 13515
rect 2455 13512 2467 13515
rect 2682 13512 2688 13524
rect 2455 13484 2688 13512
rect 2455 13481 2467 13484
rect 2409 13475 2467 13481
rect 2682 13472 2688 13484
rect 2740 13472 2746 13524
rect 4246 13472 4252 13524
rect 4304 13512 4310 13524
rect 4433 13515 4491 13521
rect 4433 13512 4445 13515
rect 4304 13484 4445 13512
rect 4304 13472 4310 13484
rect 4433 13481 4445 13484
rect 4479 13481 4491 13515
rect 4433 13475 4491 13481
rect 4522 13472 4528 13524
rect 4580 13512 4586 13524
rect 4801 13515 4859 13521
rect 4801 13512 4813 13515
rect 4580 13484 4813 13512
rect 4580 13472 4586 13484
rect 4801 13481 4813 13484
rect 4847 13481 4859 13515
rect 4801 13475 4859 13481
rect 6178 13472 6184 13524
rect 6236 13512 6242 13524
rect 6733 13515 6791 13521
rect 6733 13512 6745 13515
rect 6236 13484 6745 13512
rect 6236 13472 6242 13484
rect 6733 13481 6745 13484
rect 6779 13481 6791 13515
rect 6733 13475 6791 13481
rect 6914 13472 6920 13524
rect 6972 13512 6978 13524
rect 7745 13515 7803 13521
rect 7745 13512 7757 13515
rect 6972 13484 7757 13512
rect 6972 13472 6978 13484
rect 7745 13481 7757 13484
rect 7791 13481 7803 13515
rect 7745 13475 7803 13481
rect 9677 13515 9735 13521
rect 9677 13481 9689 13515
rect 9723 13512 9735 13515
rect 9766 13512 9772 13524
rect 9723 13484 9772 13512
rect 9723 13481 9735 13484
rect 9677 13475 9735 13481
rect 9766 13472 9772 13484
rect 9824 13472 9830 13524
rect 11149 13515 11207 13521
rect 11149 13481 11161 13515
rect 11195 13512 11207 13515
rect 14182 13512 14188 13524
rect 11195 13484 14188 13512
rect 11195 13481 11207 13484
rect 11149 13475 11207 13481
rect 14182 13472 14188 13484
rect 14240 13472 14246 13524
rect 15286 13512 15292 13524
rect 15247 13484 15292 13512
rect 15286 13472 15292 13484
rect 15344 13472 15350 13524
rect 16298 13512 16304 13524
rect 16259 13484 16304 13512
rect 16298 13472 16304 13484
rect 16356 13472 16362 13524
rect 16761 13515 16819 13521
rect 16761 13481 16773 13515
rect 16807 13512 16819 13515
rect 17218 13512 17224 13524
rect 16807 13484 17224 13512
rect 16807 13481 16819 13484
rect 16761 13475 16819 13481
rect 17218 13472 17224 13484
rect 17276 13472 17282 13524
rect 19245 13515 19303 13521
rect 19245 13512 19257 13515
rect 17512 13484 19257 13512
rect 2777 13447 2835 13453
rect 2777 13413 2789 13447
rect 2823 13444 2835 13447
rect 3142 13444 3148 13456
rect 2823 13416 3148 13444
rect 2823 13413 2835 13416
rect 2777 13407 2835 13413
rect 3142 13404 3148 13416
rect 3200 13404 3206 13456
rect 1765 13379 1823 13385
rect 1765 13345 1777 13379
rect 1811 13376 1823 13379
rect 2869 13379 2927 13385
rect 2869 13376 2881 13379
rect 1811 13348 2881 13376
rect 1811 13345 1823 13348
rect 1765 13339 1823 13345
rect 2869 13345 2881 13348
rect 2915 13376 2927 13379
rect 3694 13376 3700 13388
rect 2915 13348 3700 13376
rect 2915 13345 2927 13348
rect 2869 13339 2927 13345
rect 3694 13336 3700 13348
rect 3752 13336 3758 13388
rect 4264 13376 4292 13472
rect 4338 13404 4344 13456
rect 4396 13444 4402 13456
rect 5074 13444 5080 13456
rect 4396 13416 5080 13444
rect 4396 13404 4402 13416
rect 5074 13404 5080 13416
rect 5132 13444 5138 13456
rect 5261 13447 5319 13453
rect 5261 13444 5273 13447
rect 5132 13416 5273 13444
rect 5132 13404 5138 13416
rect 5261 13413 5273 13416
rect 5307 13444 5319 13447
rect 6273 13447 6331 13453
rect 6273 13444 6285 13447
rect 5307 13416 6285 13444
rect 5307 13413 5319 13416
rect 5261 13407 5319 13413
rect 6273 13413 6285 13416
rect 6319 13413 6331 13447
rect 6273 13407 6331 13413
rect 6362 13404 6368 13456
rect 6420 13444 6426 13456
rect 7006 13444 7012 13456
rect 6420 13416 7012 13444
rect 6420 13404 6426 13416
rect 7006 13404 7012 13416
rect 7064 13444 7070 13456
rect 12618 13444 12624 13456
rect 7064 13416 11284 13444
rect 12579 13416 12624 13444
rect 7064 13404 7070 13416
rect 11256 13388 11284 13416
rect 12618 13404 12624 13416
rect 12676 13404 12682 13456
rect 13262 13404 13268 13456
rect 13320 13444 13326 13456
rect 15657 13447 15715 13453
rect 13320 13416 15608 13444
rect 13320 13404 13326 13416
rect 4982 13376 4988 13388
rect 4264 13348 4988 13376
rect 4982 13336 4988 13348
rect 5040 13336 5046 13388
rect 5169 13379 5227 13385
rect 5169 13345 5181 13379
rect 5215 13376 5227 13379
rect 5442 13376 5448 13388
rect 5215 13348 5448 13376
rect 5215 13345 5227 13348
rect 5169 13339 5227 13345
rect 5442 13336 5448 13348
rect 5500 13376 5506 13388
rect 7098 13376 7104 13388
rect 5500 13348 5948 13376
rect 7059 13348 7104 13376
rect 5500 13336 5506 13348
rect 3053 13311 3111 13317
rect 3053 13277 3065 13311
rect 3099 13277 3111 13311
rect 3053 13271 3111 13277
rect 3068 13240 3096 13271
rect 4798 13268 4804 13320
rect 4856 13308 4862 13320
rect 5258 13308 5264 13320
rect 4856 13280 5264 13308
rect 4856 13268 4862 13280
rect 5258 13268 5264 13280
rect 5316 13268 5322 13320
rect 5353 13311 5411 13317
rect 5353 13277 5365 13311
rect 5399 13277 5411 13311
rect 5353 13271 5411 13277
rect 5166 13240 5172 13252
rect 3068 13212 5172 13240
rect 5166 13200 5172 13212
rect 5224 13240 5230 13252
rect 5368 13240 5396 13271
rect 5920 13249 5948 13348
rect 7098 13336 7104 13348
rect 7156 13336 7162 13388
rect 7929 13379 7987 13385
rect 7929 13345 7941 13379
rect 7975 13376 7987 13379
rect 8202 13376 8208 13388
rect 7975 13348 8208 13376
rect 7975 13345 7987 13348
rect 7929 13339 7987 13345
rect 8202 13336 8208 13348
rect 8260 13336 8266 13388
rect 8294 13336 8300 13388
rect 8352 13376 8358 13388
rect 8754 13376 8760 13388
rect 8352 13348 8760 13376
rect 8352 13336 8358 13348
rect 8754 13336 8760 13348
rect 8812 13336 8818 13388
rect 10042 13376 10048 13388
rect 10003 13348 10048 13376
rect 10042 13336 10048 13348
rect 10100 13376 10106 13388
rect 10597 13379 10655 13385
rect 10597 13376 10609 13379
rect 10100 13348 10609 13376
rect 10100 13336 10106 13348
rect 10597 13345 10609 13348
rect 10643 13376 10655 13379
rect 10689 13379 10747 13385
rect 10689 13376 10701 13379
rect 10643 13348 10701 13376
rect 10643 13345 10655 13348
rect 10597 13339 10655 13345
rect 10689 13345 10701 13348
rect 10735 13345 10747 13379
rect 10689 13339 10747 13345
rect 11238 13336 11244 13388
rect 11296 13376 11302 13388
rect 11517 13379 11575 13385
rect 11517 13376 11529 13379
rect 11296 13348 11529 13376
rect 11296 13336 11302 13348
rect 11517 13345 11529 13348
rect 11563 13345 11575 13379
rect 11517 13339 11575 13345
rect 12529 13379 12587 13385
rect 12529 13345 12541 13379
rect 12575 13376 12587 13379
rect 12802 13376 12808 13388
rect 12575 13348 12808 13376
rect 12575 13345 12587 13348
rect 12529 13339 12587 13345
rect 12802 13336 12808 13348
rect 12860 13336 12866 13388
rect 14090 13376 14096 13388
rect 14051 13348 14096 13376
rect 14090 13336 14096 13348
rect 14148 13336 14154 13388
rect 15580 13376 15608 13416
rect 15657 13413 15669 13447
rect 15703 13444 15715 13447
rect 17313 13447 17371 13453
rect 17313 13444 17325 13447
rect 15703 13416 17325 13444
rect 15703 13413 15715 13416
rect 15657 13407 15715 13413
rect 17313 13413 17325 13416
rect 17359 13444 17371 13447
rect 17402 13444 17408 13456
rect 17359 13416 17408 13444
rect 17359 13413 17371 13416
rect 17313 13407 17371 13413
rect 17402 13404 17408 13416
rect 17460 13404 17466 13456
rect 16666 13376 16672 13388
rect 15580 13348 16528 13376
rect 16627 13348 16672 13376
rect 7190 13308 7196 13320
rect 7151 13280 7196 13308
rect 7190 13268 7196 13280
rect 7248 13268 7254 13320
rect 7377 13311 7435 13317
rect 7377 13277 7389 13311
rect 7423 13308 7435 13311
rect 7466 13308 7472 13320
rect 7423 13280 7472 13308
rect 7423 13277 7435 13280
rect 7377 13271 7435 13277
rect 7466 13268 7472 13280
rect 7524 13268 7530 13320
rect 10134 13308 10140 13320
rect 10095 13280 10140 13308
rect 10134 13268 10140 13280
rect 10192 13268 10198 13320
rect 10226 13268 10232 13320
rect 10284 13308 10290 13320
rect 10284 13280 10329 13308
rect 10284 13268 10290 13280
rect 11146 13268 11152 13320
rect 11204 13308 11210 13320
rect 11609 13311 11667 13317
rect 11609 13308 11621 13311
rect 11204 13280 11621 13308
rect 11204 13268 11210 13280
rect 11609 13277 11621 13280
rect 11655 13277 11667 13311
rect 11790 13308 11796 13320
rect 11751 13280 11796 13308
rect 11609 13271 11667 13277
rect 11790 13268 11796 13280
rect 11848 13268 11854 13320
rect 12713 13311 12771 13317
rect 12713 13277 12725 13311
rect 12759 13308 12771 13311
rect 12894 13308 12900 13320
rect 12759 13280 12900 13308
rect 12759 13277 12771 13280
rect 12713 13271 12771 13277
rect 12894 13268 12900 13280
rect 12952 13268 12958 13320
rect 15746 13308 15752 13320
rect 15707 13280 15752 13308
rect 15746 13268 15752 13280
rect 15804 13268 15810 13320
rect 15930 13308 15936 13320
rect 15891 13280 15936 13308
rect 15930 13268 15936 13280
rect 15988 13268 15994 13320
rect 16500 13308 16528 13348
rect 16666 13336 16672 13348
rect 16724 13336 16730 13388
rect 17512 13376 17540 13484
rect 19245 13481 19257 13484
rect 19291 13481 19303 13515
rect 19245 13475 19303 13481
rect 19334 13472 19340 13524
rect 19392 13512 19398 13524
rect 19429 13515 19487 13521
rect 19429 13512 19441 13515
rect 19392 13484 19441 13512
rect 19392 13472 19398 13484
rect 19429 13481 19441 13484
rect 19475 13481 19487 13515
rect 19429 13475 19487 13481
rect 19797 13447 19855 13453
rect 19797 13444 19809 13447
rect 16776 13348 17540 13376
rect 18616 13416 19809 13444
rect 16776 13308 16804 13348
rect 18616 13320 18644 13416
rect 19797 13413 19809 13416
rect 19843 13413 19855 13447
rect 20806 13444 20812 13456
rect 19797 13407 19855 13413
rect 20456 13416 20812 13444
rect 18782 13376 18788 13388
rect 18743 13348 18788 13376
rect 18782 13336 18788 13348
rect 18840 13336 18846 13388
rect 20456 13385 20484 13416
rect 20806 13404 20812 13416
rect 20864 13404 20870 13456
rect 19337 13379 19395 13385
rect 19337 13345 19349 13379
rect 19383 13376 19395 13379
rect 20441 13379 20499 13385
rect 20441 13376 20453 13379
rect 19383 13348 20453 13376
rect 19383 13345 19395 13348
rect 19337 13339 19395 13345
rect 20441 13345 20453 13348
rect 20487 13345 20499 13379
rect 20441 13339 20499 13345
rect 20714 13336 20720 13388
rect 20772 13376 20778 13388
rect 20901 13379 20959 13385
rect 20901 13376 20913 13379
rect 20772 13348 20913 13376
rect 20772 13336 20778 13348
rect 20901 13345 20913 13348
rect 20947 13345 20959 13379
rect 20901 13339 20959 13345
rect 16500 13280 16804 13308
rect 16853 13311 16911 13317
rect 16853 13277 16865 13311
rect 16899 13277 16911 13311
rect 16853 13271 16911 13277
rect 18141 13311 18199 13317
rect 18141 13277 18153 13311
rect 18187 13308 18199 13311
rect 18598 13308 18604 13320
rect 18187 13280 18604 13308
rect 18187 13277 18199 13280
rect 18141 13271 18199 13277
rect 5224 13212 5396 13240
rect 5905 13243 5963 13249
rect 5224 13200 5230 13212
rect 5905 13209 5917 13243
rect 5951 13240 5963 13243
rect 11882 13240 11888 13252
rect 5951 13212 11888 13240
rect 5951 13209 5963 13212
rect 5905 13203 5963 13209
rect 11882 13200 11888 13212
rect 11940 13200 11946 13252
rect 13906 13240 13912 13252
rect 11992 13212 13768 13240
rect 13867 13212 13912 13240
rect 2130 13172 2136 13184
rect 2091 13144 2136 13172
rect 2130 13132 2136 13144
rect 2188 13132 2194 13184
rect 3142 13132 3148 13184
rect 3200 13172 3206 13184
rect 3418 13172 3424 13184
rect 3200 13144 3424 13172
rect 3200 13132 3206 13144
rect 3418 13132 3424 13144
rect 3476 13132 3482 13184
rect 7650 13132 7656 13184
rect 7708 13172 7714 13184
rect 8294 13172 8300 13184
rect 7708 13144 8300 13172
rect 7708 13132 7714 13144
rect 8294 13132 8300 13144
rect 8352 13132 8358 13184
rect 10597 13175 10655 13181
rect 10597 13141 10609 13175
rect 10643 13172 10655 13175
rect 11992 13172 12020 13212
rect 10643 13144 12020 13172
rect 12161 13175 12219 13181
rect 10643 13141 10655 13144
rect 10597 13135 10655 13141
rect 12161 13141 12173 13175
rect 12207 13172 12219 13175
rect 13630 13172 13636 13184
rect 12207 13144 13636 13172
rect 12207 13141 12219 13144
rect 12161 13135 12219 13141
rect 13630 13132 13636 13144
rect 13688 13132 13694 13184
rect 13740 13172 13768 13212
rect 13906 13200 13912 13212
rect 13964 13200 13970 13252
rect 15562 13200 15568 13252
rect 15620 13240 15626 13252
rect 16482 13240 16488 13252
rect 15620 13212 16488 13240
rect 15620 13200 15626 13212
rect 16482 13200 16488 13212
rect 16540 13240 16546 13252
rect 16868 13240 16896 13271
rect 18598 13268 18604 13280
rect 18656 13268 18662 13320
rect 18874 13308 18880 13320
rect 18835 13280 18880 13308
rect 18874 13268 18880 13280
rect 18932 13268 18938 13320
rect 19061 13311 19119 13317
rect 19061 13277 19073 13311
rect 19107 13308 19119 13311
rect 19150 13308 19156 13320
rect 19107 13280 19156 13308
rect 19107 13277 19119 13280
rect 19061 13271 19119 13277
rect 19150 13268 19156 13280
rect 19208 13268 19214 13320
rect 19889 13311 19947 13317
rect 19889 13277 19901 13311
rect 19935 13277 19947 13311
rect 19889 13271 19947 13277
rect 16540 13212 16896 13240
rect 17773 13243 17831 13249
rect 16540 13200 16546 13212
rect 17773 13209 17785 13243
rect 17819 13240 17831 13243
rect 18690 13240 18696 13252
rect 17819 13212 18696 13240
rect 17819 13209 17831 13212
rect 17773 13203 17831 13209
rect 18690 13200 18696 13212
rect 18748 13200 18754 13252
rect 18966 13200 18972 13252
rect 19024 13240 19030 13252
rect 19904 13240 19932 13271
rect 19978 13268 19984 13320
rect 20036 13308 20042 13320
rect 21082 13308 21088 13320
rect 20036 13280 20081 13308
rect 21043 13280 21088 13308
rect 20036 13268 20042 13280
rect 21082 13268 21088 13280
rect 21140 13268 21146 13320
rect 19024 13212 19932 13240
rect 19024 13200 19030 13212
rect 18138 13172 18144 13184
rect 13740 13144 18144 13172
rect 18138 13132 18144 13144
rect 18196 13132 18202 13184
rect 18417 13175 18475 13181
rect 18417 13141 18429 13175
rect 18463 13172 18475 13175
rect 20254 13172 20260 13184
rect 18463 13144 20260 13172
rect 18463 13141 18475 13144
rect 18417 13135 18475 13141
rect 20254 13132 20260 13144
rect 20312 13132 20318 13184
rect 1104 13082 21896 13104
rect 1104 13030 4447 13082
rect 4499 13030 4511 13082
rect 4563 13030 4575 13082
rect 4627 13030 4639 13082
rect 4691 13030 11378 13082
rect 11430 13030 11442 13082
rect 11494 13030 11506 13082
rect 11558 13030 11570 13082
rect 11622 13030 18308 13082
rect 18360 13030 18372 13082
rect 18424 13030 18436 13082
rect 18488 13030 18500 13082
rect 18552 13030 21896 13082
rect 1104 13008 21896 13030
rect 2225 12971 2283 12977
rect 2225 12937 2237 12971
rect 2271 12968 2283 12971
rect 2498 12968 2504 12980
rect 2271 12940 2504 12968
rect 2271 12937 2283 12940
rect 2225 12931 2283 12937
rect 2498 12928 2504 12940
rect 2556 12928 2562 12980
rect 3605 12971 3663 12977
rect 3605 12937 3617 12971
rect 3651 12968 3663 12971
rect 4154 12968 4160 12980
rect 3651 12940 4160 12968
rect 3651 12937 3663 12940
rect 3605 12931 3663 12937
rect 4154 12928 4160 12940
rect 4212 12928 4218 12980
rect 7374 12968 7380 12980
rect 7335 12940 7380 12968
rect 7374 12928 7380 12940
rect 7432 12928 7438 12980
rect 8297 12971 8355 12977
rect 8297 12968 8309 12971
rect 7760 12940 8309 12968
rect 5537 12903 5595 12909
rect 5537 12869 5549 12903
rect 5583 12900 5595 12903
rect 7760 12900 7788 12940
rect 8297 12937 8309 12940
rect 8343 12937 8355 12971
rect 8297 12931 8355 12937
rect 8662 12928 8668 12980
rect 8720 12968 8726 12980
rect 9125 12971 9183 12977
rect 9125 12968 9137 12971
rect 8720 12940 9137 12968
rect 8720 12928 8726 12940
rect 9125 12937 9137 12940
rect 9171 12937 9183 12971
rect 15654 12968 15660 12980
rect 9125 12931 9183 12937
rect 9232 12940 13584 12968
rect 15615 12940 15660 12968
rect 9232 12900 9260 12940
rect 10410 12900 10416 12912
rect 5583 12872 7788 12900
rect 7852 12872 9260 12900
rect 9692 12872 10416 12900
rect 5583 12869 5595 12872
rect 5537 12863 5595 12869
rect 2869 12835 2927 12841
rect 2869 12801 2881 12835
rect 2915 12832 2927 12835
rect 2958 12832 2964 12844
rect 2915 12804 2964 12832
rect 2915 12801 2927 12804
rect 2869 12795 2927 12801
rect 2958 12792 2964 12804
rect 3016 12832 3022 12844
rect 3602 12832 3608 12844
rect 3016 12804 3608 12832
rect 3016 12792 3022 12804
rect 3602 12792 3608 12804
rect 3660 12832 3666 12844
rect 4157 12835 4215 12841
rect 4157 12832 4169 12835
rect 3660 12804 4169 12832
rect 3660 12792 3666 12804
rect 4157 12801 4169 12804
rect 4203 12801 4215 12835
rect 5166 12832 5172 12844
rect 5127 12804 5172 12832
rect 4157 12795 4215 12801
rect 5166 12792 5172 12804
rect 5224 12832 5230 12844
rect 5442 12832 5448 12844
rect 5224 12804 5448 12832
rect 5224 12792 5230 12804
rect 5442 12792 5448 12804
rect 5500 12792 5506 12844
rect 7101 12835 7159 12841
rect 7101 12801 7113 12835
rect 7147 12832 7159 12835
rect 7466 12832 7472 12844
rect 7147 12804 7472 12832
rect 7147 12801 7159 12804
rect 7101 12795 7159 12801
rect 7466 12792 7472 12804
rect 7524 12832 7530 12844
rect 7852 12841 7880 12872
rect 7837 12835 7895 12841
rect 7837 12832 7849 12835
rect 7524 12804 7849 12832
rect 7524 12792 7530 12804
rect 7837 12801 7849 12804
rect 7883 12801 7895 12835
rect 7837 12795 7895 12801
rect 8021 12835 8079 12841
rect 8021 12801 8033 12835
rect 8067 12832 8079 12835
rect 8110 12832 8116 12844
rect 8067 12804 8116 12832
rect 8067 12801 8079 12804
rect 8021 12795 8079 12801
rect 8110 12792 8116 12804
rect 8168 12792 8174 12844
rect 8297 12835 8355 12841
rect 8297 12801 8309 12835
rect 8343 12832 8355 12835
rect 9692 12832 9720 12872
rect 10410 12860 10416 12872
rect 10468 12860 10474 12912
rect 11146 12900 11152 12912
rect 11107 12872 11152 12900
rect 11146 12860 11152 12872
rect 11204 12860 11210 12912
rect 11238 12860 11244 12912
rect 11296 12900 11302 12912
rect 11425 12903 11483 12909
rect 11425 12900 11437 12903
rect 11296 12872 11437 12900
rect 11296 12860 11302 12872
rect 11425 12869 11437 12872
rect 11471 12869 11483 12903
rect 11425 12863 11483 12869
rect 12894 12860 12900 12912
rect 12952 12900 12958 12912
rect 13556 12900 13584 12940
rect 15654 12928 15660 12940
rect 15712 12928 15718 12980
rect 18325 12971 18383 12977
rect 18325 12937 18337 12971
rect 18371 12968 18383 12971
rect 18782 12968 18788 12980
rect 18371 12940 18788 12968
rect 18371 12937 18383 12940
rect 18325 12931 18383 12937
rect 18782 12928 18788 12940
rect 18840 12928 18846 12980
rect 18874 12928 18880 12980
rect 18932 12968 18938 12980
rect 19337 12971 19395 12977
rect 19337 12968 19349 12971
rect 18932 12940 19349 12968
rect 18932 12928 18938 12940
rect 19337 12937 19349 12940
rect 19383 12937 19395 12971
rect 19337 12931 19395 12937
rect 12952 12872 13216 12900
rect 13556 12872 14320 12900
rect 12952 12860 12958 12872
rect 8343 12804 9720 12832
rect 9769 12835 9827 12841
rect 8343 12801 8355 12804
rect 8297 12795 8355 12801
rect 9769 12801 9781 12835
rect 9815 12832 9827 12835
rect 9858 12832 9864 12844
rect 9815 12804 9864 12832
rect 9815 12801 9827 12804
rect 9769 12795 9827 12801
rect 9858 12792 9864 12804
rect 9916 12792 9922 12844
rect 10134 12792 10140 12844
rect 10192 12832 10198 12844
rect 10781 12835 10839 12841
rect 10781 12832 10793 12835
rect 10192 12804 10793 12832
rect 10192 12792 10198 12804
rect 10781 12801 10793 12804
rect 10827 12832 10839 12835
rect 13078 12832 13084 12844
rect 10827 12804 13084 12832
rect 10827 12801 10839 12804
rect 10781 12795 10839 12801
rect 13078 12792 13084 12804
rect 13136 12792 13142 12844
rect 13188 12832 13216 12872
rect 13725 12835 13783 12841
rect 13725 12832 13737 12835
rect 13188 12804 13737 12832
rect 13725 12801 13737 12804
rect 13771 12801 13783 12835
rect 14292 12832 14320 12872
rect 15746 12860 15752 12912
rect 15804 12900 15810 12912
rect 16577 12903 16635 12909
rect 16577 12900 16589 12903
rect 15804 12872 16589 12900
rect 15804 12860 15810 12872
rect 16577 12869 16589 12872
rect 16623 12900 16635 12903
rect 18598 12900 18604 12912
rect 16623 12872 18604 12900
rect 16623 12869 16635 12872
rect 16577 12863 16635 12869
rect 18598 12860 18604 12872
rect 18656 12860 18662 12912
rect 19150 12900 19156 12912
rect 18800 12872 19156 12900
rect 14292 12804 14412 12832
rect 13725 12795 13783 12801
rect 4062 12724 4068 12776
rect 4120 12764 4126 12776
rect 7745 12767 7803 12773
rect 4120 12736 5764 12764
rect 4120 12724 4126 12736
rect 3973 12699 4031 12705
rect 3973 12665 3985 12699
rect 4019 12696 4031 12699
rect 4706 12696 4712 12708
rect 4019 12668 4712 12696
rect 4019 12665 4031 12668
rect 3973 12659 4031 12665
rect 4706 12656 4712 12668
rect 4764 12656 4770 12708
rect 4982 12696 4988 12708
rect 4943 12668 4988 12696
rect 4982 12656 4988 12668
rect 5040 12656 5046 12708
rect 5077 12699 5135 12705
rect 5077 12665 5089 12699
rect 5123 12696 5135 12699
rect 5537 12699 5595 12705
rect 5537 12696 5549 12699
rect 5123 12668 5549 12696
rect 5123 12665 5135 12668
rect 5077 12659 5135 12665
rect 5537 12665 5549 12668
rect 5583 12696 5595 12699
rect 5629 12699 5687 12705
rect 5629 12696 5641 12699
rect 5583 12668 5641 12696
rect 5583 12665 5595 12668
rect 5537 12659 5595 12665
rect 5629 12665 5641 12668
rect 5675 12665 5687 12699
rect 5629 12659 5687 12665
rect 2590 12628 2596 12640
rect 2551 12600 2596 12628
rect 2590 12588 2596 12600
rect 2648 12588 2654 12640
rect 2682 12588 2688 12640
rect 2740 12628 2746 12640
rect 4065 12631 4123 12637
rect 2740 12600 2785 12628
rect 2740 12588 2746 12600
rect 4065 12597 4077 12631
rect 4111 12628 4123 12631
rect 4617 12631 4675 12637
rect 4617 12628 4629 12631
rect 4111 12600 4629 12628
rect 4111 12597 4123 12600
rect 4065 12591 4123 12597
rect 4617 12597 4629 12600
rect 4663 12597 4675 12631
rect 5736 12628 5764 12736
rect 7745 12733 7757 12767
rect 7791 12764 7803 12767
rect 8481 12767 8539 12773
rect 8481 12764 8493 12767
rect 7791 12736 8493 12764
rect 7791 12733 7803 12736
rect 7745 12727 7803 12733
rect 8481 12733 8493 12736
rect 8527 12764 8539 12767
rect 8570 12764 8576 12776
rect 8527 12736 8576 12764
rect 8527 12733 8539 12736
rect 8481 12727 8539 12733
rect 8570 12724 8576 12736
rect 8628 12764 8634 12776
rect 13354 12764 13360 12776
rect 8628 12736 13360 12764
rect 8628 12724 8634 12736
rect 13354 12724 13360 12736
rect 13412 12724 13418 12776
rect 13814 12724 13820 12776
rect 13872 12764 13878 12776
rect 14277 12767 14335 12773
rect 14277 12764 14289 12767
rect 13872 12736 14289 12764
rect 13872 12724 13878 12736
rect 14277 12733 14289 12736
rect 14323 12733 14335 12767
rect 14384 12764 14412 12804
rect 16482 12792 16488 12844
rect 16540 12832 16546 12844
rect 16540 12804 17080 12832
rect 16540 12792 16546 12804
rect 16117 12767 16175 12773
rect 16117 12764 16129 12767
rect 14384 12736 16129 12764
rect 14277 12727 14335 12733
rect 16117 12733 16129 12736
rect 16163 12764 16175 12767
rect 16666 12764 16672 12776
rect 16163 12736 16672 12764
rect 16163 12733 16175 12736
rect 16117 12727 16175 12733
rect 16666 12724 16672 12736
rect 16724 12724 16730 12776
rect 17052 12764 17080 12804
rect 17126 12792 17132 12844
rect 17184 12832 17190 12844
rect 17405 12835 17463 12841
rect 17405 12832 17417 12835
rect 17184 12804 17417 12832
rect 17184 12792 17190 12804
rect 17405 12801 17417 12804
rect 17451 12801 17463 12835
rect 17405 12795 17463 12801
rect 18046 12792 18052 12844
rect 18104 12832 18110 12844
rect 18800 12841 18828 12872
rect 19150 12860 19156 12872
rect 19208 12860 19214 12912
rect 18785 12835 18843 12841
rect 18785 12832 18797 12835
rect 18104 12804 18797 12832
rect 18104 12792 18110 12804
rect 18785 12801 18797 12804
rect 18831 12801 18843 12835
rect 18785 12795 18843 12801
rect 18877 12835 18935 12841
rect 18877 12801 18889 12835
rect 18923 12832 18935 12835
rect 19702 12832 19708 12844
rect 18923 12804 19708 12832
rect 18923 12801 18935 12804
rect 18877 12795 18935 12801
rect 18690 12764 18696 12776
rect 17052 12736 18552 12764
rect 18651 12736 18696 12764
rect 7650 12656 7656 12708
rect 7708 12696 7714 12708
rect 8110 12696 8116 12708
rect 7708 12668 8116 12696
rect 7708 12656 7714 12668
rect 8110 12656 8116 12668
rect 8168 12656 8174 12708
rect 10594 12696 10600 12708
rect 8220 12668 10600 12696
rect 8220 12628 8248 12668
rect 10594 12656 10600 12668
rect 10652 12656 10658 12708
rect 11882 12656 11888 12708
rect 11940 12696 11946 12708
rect 13541 12699 13599 12705
rect 13541 12696 13553 12699
rect 11940 12668 13553 12696
rect 11940 12656 11946 12668
rect 13541 12665 13553 12668
rect 13587 12665 13599 12699
rect 13541 12659 13599 12665
rect 13633 12699 13691 12705
rect 13633 12665 13645 12699
rect 13679 12696 13691 12699
rect 13679 12668 14136 12696
rect 13679 12665 13691 12668
rect 13633 12659 13691 12665
rect 5736 12600 8248 12628
rect 4617 12591 4675 12597
rect 8478 12588 8484 12640
rect 8536 12628 8542 12640
rect 9493 12631 9551 12637
rect 9493 12628 9505 12631
rect 8536 12600 9505 12628
rect 8536 12588 8542 12600
rect 9493 12597 9505 12600
rect 9539 12597 9551 12631
rect 9493 12591 9551 12597
rect 9585 12631 9643 12637
rect 9585 12597 9597 12631
rect 9631 12628 9643 12631
rect 9674 12628 9680 12640
rect 9631 12600 9680 12628
rect 9631 12597 9643 12600
rect 9585 12591 9643 12597
rect 9674 12588 9680 12600
rect 9732 12588 9738 12640
rect 9950 12588 9956 12640
rect 10008 12628 10014 12640
rect 10137 12631 10195 12637
rect 10137 12628 10149 12631
rect 10008 12600 10149 12628
rect 10008 12588 10014 12600
rect 10137 12597 10149 12600
rect 10183 12597 10195 12631
rect 10137 12591 10195 12597
rect 12434 12588 12440 12640
rect 12492 12628 12498 12640
rect 13173 12631 13231 12637
rect 12492 12600 12537 12628
rect 12492 12588 12498 12600
rect 13173 12597 13185 12631
rect 13219 12628 13231 12631
rect 13906 12628 13912 12640
rect 13219 12600 13912 12628
rect 13219 12597 13231 12600
rect 13173 12591 13231 12597
rect 13906 12588 13912 12600
rect 13964 12588 13970 12640
rect 14108 12628 14136 12668
rect 14182 12656 14188 12708
rect 14240 12696 14246 12708
rect 14522 12699 14580 12705
rect 14522 12696 14534 12699
rect 14240 12668 14534 12696
rect 14240 12656 14246 12668
rect 14522 12665 14534 12668
rect 14568 12665 14580 12699
rect 14522 12659 14580 12665
rect 17221 12699 17279 12705
rect 17221 12665 17233 12699
rect 17267 12696 17279 12699
rect 17678 12696 17684 12708
rect 17267 12668 17684 12696
rect 17267 12665 17279 12668
rect 17221 12659 17279 12665
rect 17678 12656 17684 12668
rect 17736 12656 17742 12708
rect 18524 12696 18552 12736
rect 18690 12724 18696 12736
rect 18748 12724 18754 12776
rect 18892 12764 18920 12795
rect 19702 12792 19708 12804
rect 19760 12832 19766 12844
rect 19889 12835 19947 12841
rect 19889 12832 19901 12835
rect 19760 12804 19901 12832
rect 19760 12792 19766 12804
rect 19889 12801 19901 12804
rect 19935 12832 19947 12835
rect 19978 12832 19984 12844
rect 19935 12804 19984 12832
rect 19935 12801 19947 12804
rect 19889 12795 19947 12801
rect 19978 12792 19984 12804
rect 20036 12792 20042 12844
rect 20254 12792 20260 12844
rect 20312 12832 20318 12844
rect 21085 12835 21143 12841
rect 21085 12832 21097 12835
rect 20312 12804 21097 12832
rect 20312 12792 20318 12804
rect 21085 12801 21097 12804
rect 21131 12801 21143 12835
rect 21085 12795 21143 12801
rect 20990 12764 20996 12776
rect 18800 12736 18920 12764
rect 19260 12736 20996 12764
rect 18800 12696 18828 12736
rect 18524 12668 18828 12696
rect 19260 12640 19288 12736
rect 20990 12724 20996 12736
rect 21048 12724 21054 12776
rect 19518 12656 19524 12708
rect 19576 12696 19582 12708
rect 19797 12699 19855 12705
rect 19797 12696 19809 12699
rect 19576 12668 19809 12696
rect 19576 12656 19582 12668
rect 19797 12665 19809 12668
rect 19843 12665 19855 12699
rect 19797 12659 19855 12665
rect 16853 12631 16911 12637
rect 16853 12628 16865 12631
rect 14108 12600 16865 12628
rect 16853 12597 16865 12600
rect 16899 12597 16911 12631
rect 16853 12591 16911 12597
rect 17313 12631 17371 12637
rect 17313 12597 17325 12631
rect 17359 12628 17371 12631
rect 18046 12628 18052 12640
rect 17359 12600 18052 12628
rect 17359 12597 17371 12600
rect 17313 12591 17371 12597
rect 18046 12588 18052 12600
rect 18104 12588 18110 12640
rect 18138 12588 18144 12640
rect 18196 12628 18202 12640
rect 19242 12628 19248 12640
rect 18196 12600 19248 12628
rect 18196 12588 18202 12600
rect 19242 12588 19248 12600
rect 19300 12588 19306 12640
rect 19334 12588 19340 12640
rect 19392 12628 19398 12640
rect 19705 12631 19763 12637
rect 19705 12628 19717 12631
rect 19392 12600 19717 12628
rect 19392 12588 19398 12600
rect 19705 12597 19717 12600
rect 19751 12597 19763 12631
rect 20530 12628 20536 12640
rect 20491 12600 20536 12628
rect 19705 12591 19763 12597
rect 20530 12588 20536 12600
rect 20588 12588 20594 12640
rect 20898 12628 20904 12640
rect 20859 12600 20904 12628
rect 20898 12588 20904 12600
rect 20956 12588 20962 12640
rect 1104 12538 21896 12560
rect 1104 12486 7912 12538
rect 7964 12486 7976 12538
rect 8028 12486 8040 12538
rect 8092 12486 8104 12538
rect 8156 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 15035 12538
rect 15087 12486 21896 12538
rect 1104 12464 21896 12486
rect 2409 12427 2467 12433
rect 2409 12393 2421 12427
rect 2455 12424 2467 12427
rect 2682 12424 2688 12436
rect 2455 12396 2688 12424
rect 2455 12393 2467 12396
rect 2409 12387 2467 12393
rect 2682 12384 2688 12396
rect 2740 12384 2746 12436
rect 4706 12424 4712 12436
rect 4667 12396 4712 12424
rect 4706 12384 4712 12396
rect 4764 12384 4770 12436
rect 7009 12427 7067 12433
rect 7009 12424 7021 12427
rect 5000 12396 7021 12424
rect 1765 12291 1823 12297
rect 1765 12257 1777 12291
rect 1811 12288 1823 12291
rect 2777 12291 2835 12297
rect 2777 12288 2789 12291
rect 1811 12260 2789 12288
rect 1811 12257 1823 12260
rect 1765 12251 1823 12257
rect 2777 12257 2789 12260
rect 2823 12288 2835 12291
rect 3326 12288 3332 12300
rect 2823 12260 3332 12288
rect 2823 12257 2835 12260
rect 2777 12251 2835 12257
rect 3326 12248 3332 12260
rect 3384 12248 3390 12300
rect 4338 12248 4344 12300
rect 4396 12288 4402 12300
rect 5000 12288 5028 12396
rect 7009 12393 7021 12396
rect 7055 12393 7067 12427
rect 7190 12424 7196 12436
rect 7151 12396 7196 12424
rect 7009 12387 7067 12393
rect 7190 12384 7196 12396
rect 7248 12384 7254 12436
rect 9674 12424 9680 12436
rect 9635 12396 9680 12424
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 10686 12424 10692 12436
rect 9784 12396 10692 12424
rect 5534 12316 5540 12368
rect 5592 12356 5598 12368
rect 9784 12356 9812 12396
rect 10686 12384 10692 12396
rect 10744 12384 10750 12436
rect 12437 12427 12495 12433
rect 12437 12393 12449 12427
rect 12483 12424 12495 12427
rect 12894 12424 12900 12436
rect 12483 12396 12900 12424
rect 12483 12393 12495 12396
rect 12437 12387 12495 12393
rect 12894 12384 12900 12396
rect 12952 12384 12958 12436
rect 13354 12384 13360 12436
rect 13412 12424 13418 12436
rect 14182 12424 14188 12436
rect 13412 12396 14044 12424
rect 14143 12396 14188 12424
rect 13412 12384 13418 12396
rect 10962 12356 10968 12368
rect 5592 12328 9812 12356
rect 9876 12328 10968 12356
rect 5592 12316 5598 12328
rect 5077 12291 5135 12297
rect 5077 12288 5089 12291
rect 4396 12260 5089 12288
rect 4396 12248 4402 12260
rect 5077 12257 5089 12260
rect 5123 12257 5135 12291
rect 5077 12251 5135 12257
rect 5169 12291 5227 12297
rect 5169 12257 5181 12291
rect 5215 12288 5227 12291
rect 6454 12288 6460 12300
rect 5215 12260 6460 12288
rect 5215 12257 5227 12260
rect 5169 12251 5227 12257
rect 2869 12223 2927 12229
rect 2869 12189 2881 12223
rect 2915 12220 2927 12223
rect 3053 12223 3111 12229
rect 2915 12192 3004 12220
rect 2915 12189 2927 12192
rect 2869 12183 2927 12189
rect 2133 12155 2191 12161
rect 2133 12121 2145 12155
rect 2179 12152 2191 12155
rect 2976 12152 3004 12192
rect 3053 12189 3065 12223
rect 3099 12189 3111 12223
rect 3053 12183 3111 12189
rect 4433 12223 4491 12229
rect 4433 12189 4445 12223
rect 4479 12220 4491 12223
rect 5184 12220 5212 12251
rect 6454 12248 6460 12260
rect 6512 12288 6518 12300
rect 7561 12291 7619 12297
rect 7561 12288 7573 12291
rect 6512 12260 7573 12288
rect 6512 12248 6518 12260
rect 7561 12257 7573 12260
rect 7607 12257 7619 12291
rect 7561 12251 7619 12257
rect 7653 12291 7711 12297
rect 7653 12257 7665 12291
rect 7699 12288 7711 12291
rect 8297 12291 8355 12297
rect 8297 12288 8309 12291
rect 7699 12260 8309 12288
rect 7699 12257 7711 12260
rect 7653 12251 7711 12257
rect 8297 12257 8309 12260
rect 8343 12288 8355 12291
rect 9876 12288 9904 12328
rect 10962 12316 10968 12328
rect 11020 12316 11026 12368
rect 12710 12356 12716 12368
rect 11072 12328 12716 12356
rect 11072 12297 11100 12328
rect 12710 12316 12716 12328
rect 12768 12356 12774 12368
rect 13814 12356 13820 12368
rect 12768 12328 13820 12356
rect 12768 12316 12774 12328
rect 13814 12316 13820 12328
rect 13872 12316 13878 12368
rect 14016 12356 14044 12396
rect 14182 12384 14188 12396
rect 14240 12384 14246 12436
rect 15289 12427 15347 12433
rect 15289 12393 15301 12427
rect 15335 12424 15347 12427
rect 16206 12424 16212 12436
rect 15335 12396 16212 12424
rect 15335 12393 15347 12396
rect 15289 12387 15347 12393
rect 16206 12384 16212 12396
rect 16264 12384 16270 12436
rect 16758 12384 16764 12436
rect 16816 12424 16822 12436
rect 17126 12424 17132 12436
rect 16816 12396 17132 12424
rect 16816 12384 16822 12396
rect 17126 12384 17132 12396
rect 17184 12424 17190 12436
rect 17773 12427 17831 12433
rect 17773 12424 17785 12427
rect 17184 12396 17785 12424
rect 17184 12384 17190 12396
rect 17773 12393 17785 12396
rect 17819 12393 17831 12427
rect 18046 12424 18052 12436
rect 18007 12396 18052 12424
rect 17773 12387 17831 12393
rect 18046 12384 18052 12396
rect 18104 12384 18110 12436
rect 18509 12427 18567 12433
rect 18509 12393 18521 12427
rect 18555 12424 18567 12427
rect 18598 12424 18604 12436
rect 18555 12396 18604 12424
rect 18555 12393 18567 12396
rect 18509 12387 18567 12393
rect 18598 12384 18604 12396
rect 18656 12424 18662 12436
rect 18966 12424 18972 12436
rect 18656 12396 18972 12424
rect 18656 12384 18662 12396
rect 18966 12384 18972 12396
rect 19024 12384 19030 12436
rect 19337 12427 19395 12433
rect 19337 12393 19349 12427
rect 19383 12424 19395 12427
rect 19426 12424 19432 12436
rect 19383 12396 19432 12424
rect 19383 12393 19395 12396
rect 19337 12387 19395 12393
rect 19426 12384 19432 12396
rect 19484 12384 19490 12436
rect 21085 12427 21143 12433
rect 21085 12393 21097 12427
rect 21131 12424 21143 12427
rect 21174 12424 21180 12436
rect 21131 12396 21180 12424
rect 21131 12393 21143 12396
rect 21085 12387 21143 12393
rect 21174 12384 21180 12396
rect 21232 12384 21238 12436
rect 14829 12359 14887 12365
rect 14829 12356 14841 12359
rect 14016 12328 14841 12356
rect 14829 12325 14841 12328
rect 14875 12356 14887 12359
rect 15749 12359 15807 12365
rect 15749 12356 15761 12359
rect 14875 12328 15761 12356
rect 14875 12325 14887 12328
rect 14829 12319 14887 12325
rect 15749 12325 15761 12328
rect 15795 12325 15807 12359
rect 15749 12319 15807 12325
rect 16660 12359 16718 12365
rect 16660 12325 16672 12359
rect 16706 12356 16718 12359
rect 16942 12356 16948 12368
rect 16706 12328 16948 12356
rect 16706 12325 16718 12328
rect 16660 12319 16718 12325
rect 16942 12316 16948 12328
rect 17000 12356 17006 12368
rect 17000 12328 18644 12356
rect 17000 12316 17006 12328
rect 8343 12260 9904 12288
rect 10045 12291 10103 12297
rect 8343 12257 8355 12260
rect 8297 12251 8355 12257
rect 10045 12257 10057 12291
rect 10091 12257 10103 12291
rect 10045 12251 10103 12257
rect 11057 12291 11115 12297
rect 11057 12257 11069 12291
rect 11103 12257 11115 12291
rect 11057 12251 11115 12257
rect 4479 12192 5212 12220
rect 5353 12223 5411 12229
rect 4479 12189 4491 12192
rect 4433 12183 4491 12189
rect 5353 12189 5365 12223
rect 5399 12220 5411 12223
rect 5442 12220 5448 12232
rect 5399 12192 5448 12220
rect 5399 12189 5411 12192
rect 5353 12183 5411 12189
rect 2179 12124 3004 12152
rect 3068 12152 3096 12183
rect 5368 12152 5396 12183
rect 5442 12180 5448 12192
rect 5500 12180 5506 12232
rect 6733 12223 6791 12229
rect 6733 12189 6745 12223
rect 6779 12220 6791 12223
rect 7190 12220 7196 12232
rect 6779 12192 7196 12220
rect 6779 12189 6791 12192
rect 6733 12183 6791 12189
rect 7190 12180 7196 12192
rect 7248 12180 7254 12232
rect 7742 12220 7748 12232
rect 7703 12192 7748 12220
rect 7742 12180 7748 12192
rect 7800 12180 7806 12232
rect 6638 12152 6644 12164
rect 3068 12124 5396 12152
rect 5440 12124 6644 12152
rect 2179 12121 2191 12124
rect 2133 12115 2191 12121
rect 2976 12084 3004 12124
rect 3786 12084 3792 12096
rect 2976 12056 3792 12084
rect 3786 12044 3792 12056
rect 3844 12084 3850 12096
rect 5440 12084 5468 12124
rect 6638 12112 6644 12124
rect 6696 12112 6702 12164
rect 9125 12155 9183 12161
rect 9125 12152 9137 12155
rect 6748 12124 9137 12152
rect 6748 12096 6776 12124
rect 9125 12121 9137 12124
rect 9171 12152 9183 12155
rect 9950 12152 9956 12164
rect 9171 12124 9956 12152
rect 9171 12121 9183 12124
rect 9125 12115 9183 12121
rect 9950 12112 9956 12124
rect 10008 12112 10014 12164
rect 6454 12084 6460 12096
rect 3844 12056 5468 12084
rect 6415 12056 6460 12084
rect 3844 12044 3850 12056
rect 6454 12044 6460 12056
rect 6512 12044 6518 12096
rect 6730 12044 6736 12096
rect 6788 12044 6794 12096
rect 7009 12087 7067 12093
rect 7009 12053 7021 12087
rect 7055 12084 7067 12087
rect 8757 12087 8815 12093
rect 8757 12084 8769 12087
rect 7055 12056 8769 12084
rect 7055 12053 7067 12056
rect 7009 12047 7067 12053
rect 8757 12053 8769 12056
rect 8803 12084 8815 12087
rect 10060 12084 10088 12251
rect 11146 12248 11152 12300
rect 11204 12288 11210 12300
rect 11313 12291 11371 12297
rect 11313 12288 11325 12291
rect 11204 12260 11325 12288
rect 11204 12248 11210 12260
rect 11313 12257 11325 12260
rect 11359 12257 11371 12291
rect 11313 12251 11371 12257
rect 11606 12248 11612 12300
rect 11664 12288 11670 12300
rect 11664 12260 12204 12288
rect 11664 12248 11670 12260
rect 10137 12223 10195 12229
rect 10137 12189 10149 12223
rect 10183 12189 10195 12223
rect 10137 12183 10195 12189
rect 8803 12056 10088 12084
rect 10152 12084 10180 12183
rect 10226 12180 10232 12232
rect 10284 12220 10290 12232
rect 10284 12192 10329 12220
rect 10284 12180 10290 12192
rect 12176 12164 12204 12260
rect 12894 12248 12900 12300
rect 12952 12288 12958 12300
rect 13061 12291 13119 12297
rect 13061 12288 13073 12291
rect 12952 12260 13073 12288
rect 12952 12248 12958 12260
rect 13061 12257 13073 12260
rect 13107 12257 13119 12291
rect 15657 12291 15715 12297
rect 15657 12288 15669 12291
rect 13061 12251 13119 12257
rect 14476 12260 15669 12288
rect 12805 12223 12863 12229
rect 12805 12189 12817 12223
rect 12851 12189 12863 12223
rect 12805 12183 12863 12189
rect 12158 12112 12164 12164
rect 12216 12152 12222 12164
rect 12216 12124 12388 12152
rect 12216 12112 12222 12124
rect 10781 12087 10839 12093
rect 10781 12084 10793 12087
rect 10152 12056 10793 12084
rect 8803 12053 8815 12056
rect 8757 12047 8815 12053
rect 10781 12053 10793 12056
rect 10827 12084 10839 12087
rect 12250 12084 12256 12096
rect 10827 12056 12256 12084
rect 10827 12053 10839 12056
rect 10781 12047 10839 12053
rect 12250 12044 12256 12056
rect 12308 12044 12314 12096
rect 12360 12084 12388 12124
rect 12710 12112 12716 12164
rect 12768 12152 12774 12164
rect 12820 12152 12848 12183
rect 12768 12124 12848 12152
rect 12768 12112 12774 12124
rect 14476 12093 14504 12260
rect 15657 12257 15669 12260
rect 15703 12257 15715 12291
rect 15657 12251 15715 12257
rect 15930 12248 15936 12300
rect 15988 12288 15994 12300
rect 16393 12291 16451 12297
rect 16393 12288 16405 12291
rect 15988 12260 16405 12288
rect 15988 12248 15994 12260
rect 16393 12257 16405 12260
rect 16439 12288 16451 12291
rect 18138 12288 18144 12300
rect 16439 12260 18144 12288
rect 16439 12257 16451 12260
rect 16393 12251 16451 12257
rect 18138 12248 18144 12260
rect 18196 12248 18202 12300
rect 18417 12291 18475 12297
rect 18417 12257 18429 12291
rect 18463 12257 18475 12291
rect 18417 12251 18475 12257
rect 15841 12223 15899 12229
rect 15841 12189 15853 12223
rect 15887 12189 15899 12223
rect 15841 12183 15899 12189
rect 15654 12112 15660 12164
rect 15712 12152 15718 12164
rect 15856 12152 15884 12183
rect 15712 12124 15884 12152
rect 18432 12152 18460 12251
rect 18616 12232 18644 12328
rect 19242 12316 19248 12368
rect 19300 12356 19306 12368
rect 20441 12359 20499 12365
rect 20441 12356 20453 12359
rect 19300 12328 20453 12356
rect 19300 12316 19306 12328
rect 20441 12325 20453 12328
rect 20487 12325 20499 12359
rect 20441 12319 20499 12325
rect 19705 12291 19763 12297
rect 19705 12288 19717 12291
rect 19260 12260 19717 12288
rect 18598 12220 18604 12232
rect 18559 12192 18604 12220
rect 18598 12180 18604 12192
rect 18656 12180 18662 12232
rect 19260 12164 19288 12260
rect 19705 12257 19717 12260
rect 19751 12257 19763 12291
rect 19705 12251 19763 12257
rect 20901 12291 20959 12297
rect 20901 12257 20913 12291
rect 20947 12288 20959 12291
rect 21082 12288 21088 12300
rect 20947 12260 21088 12288
rect 20947 12257 20959 12260
rect 20901 12251 20959 12257
rect 21082 12248 21088 12260
rect 21140 12248 21146 12300
rect 19797 12223 19855 12229
rect 19797 12189 19809 12223
rect 19843 12189 19855 12223
rect 19978 12220 19984 12232
rect 19939 12192 19984 12220
rect 19797 12183 19855 12189
rect 19242 12152 19248 12164
rect 18432 12124 19248 12152
rect 15712 12112 15718 12124
rect 19242 12112 19248 12124
rect 19300 12112 19306 12164
rect 19702 12112 19708 12164
rect 19760 12152 19766 12164
rect 19812 12152 19840 12183
rect 19978 12180 19984 12192
rect 20036 12180 20042 12232
rect 19760 12124 19840 12152
rect 19760 12112 19766 12124
rect 14461 12087 14519 12093
rect 14461 12084 14473 12087
rect 12360 12056 14473 12084
rect 14461 12053 14473 12056
rect 14507 12053 14519 12087
rect 14461 12047 14519 12053
rect 14642 12044 14648 12096
rect 14700 12084 14706 12096
rect 19886 12084 19892 12096
rect 14700 12056 19892 12084
rect 14700 12044 14706 12056
rect 19886 12044 19892 12056
rect 19944 12044 19950 12096
rect 20714 12044 20720 12096
rect 20772 12084 20778 12096
rect 20990 12084 20996 12096
rect 20772 12056 20996 12084
rect 20772 12044 20778 12056
rect 20990 12044 20996 12056
rect 21048 12044 21054 12096
rect 1104 11994 21896 12016
rect 1104 11942 4447 11994
rect 4499 11942 4511 11994
rect 4563 11942 4575 11994
rect 4627 11942 4639 11994
rect 4691 11942 11378 11994
rect 11430 11942 11442 11994
rect 11494 11942 11506 11994
rect 11558 11942 11570 11994
rect 11622 11942 18308 11994
rect 18360 11942 18372 11994
rect 18424 11942 18436 11994
rect 18488 11942 18500 11994
rect 18552 11942 21896 11994
rect 1104 11920 21896 11942
rect 1857 11883 1915 11889
rect 1857 11849 1869 11883
rect 1903 11880 1915 11883
rect 2866 11880 2872 11892
rect 1903 11852 2872 11880
rect 1903 11849 1915 11852
rect 1857 11843 1915 11849
rect 2866 11840 2872 11852
rect 2924 11840 2930 11892
rect 3602 11880 3608 11892
rect 3563 11852 3608 11880
rect 3602 11840 3608 11852
rect 3660 11840 3666 11892
rect 6825 11883 6883 11889
rect 6825 11849 6837 11883
rect 6871 11880 6883 11883
rect 7098 11880 7104 11892
rect 6871 11852 7104 11880
rect 6871 11849 6883 11852
rect 6825 11843 6883 11849
rect 7098 11840 7104 11852
rect 7156 11840 7162 11892
rect 8478 11880 8484 11892
rect 8439 11852 8484 11880
rect 8478 11840 8484 11852
rect 8536 11840 8542 11892
rect 9493 11883 9551 11889
rect 9493 11849 9505 11883
rect 9539 11880 9551 11883
rect 9766 11880 9772 11892
rect 9539 11852 9772 11880
rect 9539 11849 9551 11852
rect 9493 11843 9551 11849
rect 9766 11840 9772 11852
rect 9824 11840 9830 11892
rect 10505 11883 10563 11889
rect 10505 11849 10517 11883
rect 10551 11880 10563 11883
rect 11882 11880 11888 11892
rect 10551 11852 11888 11880
rect 10551 11849 10563 11852
rect 10505 11843 10563 11849
rect 11882 11840 11888 11852
rect 11940 11840 11946 11892
rect 12437 11883 12495 11889
rect 12437 11849 12449 11883
rect 12483 11880 12495 11883
rect 12618 11880 12624 11892
rect 12483 11852 12624 11880
rect 12483 11849 12495 11852
rect 12437 11843 12495 11849
rect 12618 11840 12624 11852
rect 12676 11840 12682 11892
rect 13265 11883 13323 11889
rect 13265 11849 13277 11883
rect 13311 11880 13323 11883
rect 14642 11880 14648 11892
rect 13311 11852 14648 11880
rect 13311 11849 13323 11852
rect 13265 11843 13323 11849
rect 14642 11840 14648 11852
rect 14700 11840 14706 11892
rect 14734 11840 14740 11892
rect 14792 11880 14798 11892
rect 20714 11880 20720 11892
rect 14792 11852 20720 11880
rect 14792 11840 14798 11852
rect 20714 11840 20720 11852
rect 20772 11840 20778 11892
rect 4062 11772 4068 11824
rect 4120 11812 4126 11824
rect 12526 11812 12532 11824
rect 4120 11784 12532 11812
rect 4120 11772 4126 11784
rect 12526 11772 12532 11784
rect 12584 11772 12590 11824
rect 13357 11815 13415 11821
rect 13357 11781 13369 11815
rect 13403 11812 13415 11815
rect 19058 11812 19064 11824
rect 13403 11784 19064 11812
rect 13403 11781 13415 11784
rect 13357 11775 13415 11781
rect 19058 11772 19064 11784
rect 19116 11772 19122 11824
rect 3510 11704 3516 11756
rect 3568 11744 3574 11756
rect 5813 11747 5871 11753
rect 5813 11744 5825 11747
rect 3568 11716 5825 11744
rect 3568 11704 3574 11716
rect 5813 11713 5825 11716
rect 5859 11744 5871 11747
rect 6181 11747 6239 11753
rect 6181 11744 6193 11747
rect 5859 11716 6193 11744
rect 5859 11713 5871 11716
rect 5813 11707 5871 11713
rect 6181 11713 6193 11716
rect 6227 11744 6239 11747
rect 6914 11744 6920 11756
rect 6227 11716 6920 11744
rect 6227 11713 6239 11716
rect 6181 11707 6239 11713
rect 6914 11704 6920 11716
rect 6972 11744 6978 11756
rect 7285 11747 7343 11753
rect 7285 11744 7297 11747
rect 6972 11716 7297 11744
rect 6972 11704 6978 11716
rect 7285 11713 7297 11716
rect 7331 11713 7343 11747
rect 7285 11707 7343 11713
rect 7469 11747 7527 11753
rect 7469 11713 7481 11747
rect 7515 11744 7527 11747
rect 7742 11744 7748 11756
rect 7515 11716 7748 11744
rect 7515 11713 7527 11716
rect 7469 11707 7527 11713
rect 7742 11704 7748 11716
rect 7800 11704 7806 11756
rect 9125 11747 9183 11753
rect 9125 11713 9137 11747
rect 9171 11744 9183 11747
rect 10045 11747 10103 11753
rect 10045 11744 10057 11747
rect 9171 11716 10057 11744
rect 9171 11713 9183 11716
rect 9125 11707 9183 11713
rect 10045 11713 10057 11716
rect 10091 11744 10103 11747
rect 10226 11744 10232 11756
rect 10091 11716 10232 11744
rect 10091 11713 10103 11716
rect 10045 11707 10103 11713
rect 10226 11704 10232 11716
rect 10284 11704 10290 11756
rect 11146 11744 11152 11756
rect 11059 11716 11152 11744
rect 11146 11704 11152 11716
rect 11204 11744 11210 11756
rect 13081 11747 13139 11753
rect 13081 11744 13093 11747
rect 11204 11716 13093 11744
rect 11204 11704 11210 11716
rect 13081 11713 13093 11716
rect 13127 11744 13139 11747
rect 13906 11744 13912 11756
rect 13127 11716 13676 11744
rect 13867 11716 13912 11744
rect 13127 11713 13139 11716
rect 13081 11707 13139 11713
rect 1673 11679 1731 11685
rect 1673 11645 1685 11679
rect 1719 11676 1731 11679
rect 1946 11676 1952 11688
rect 1719 11648 1952 11676
rect 1719 11645 1731 11648
rect 1673 11639 1731 11645
rect 1946 11636 1952 11648
rect 2004 11636 2010 11688
rect 2225 11679 2283 11685
rect 2225 11645 2237 11679
rect 2271 11676 2283 11679
rect 2314 11676 2320 11688
rect 2271 11648 2320 11676
rect 2271 11645 2283 11648
rect 2225 11639 2283 11645
rect 2314 11636 2320 11648
rect 2372 11636 2378 11688
rect 2492 11679 2550 11685
rect 2492 11645 2504 11679
rect 2538 11676 2550 11679
rect 3234 11676 3240 11688
rect 2538 11648 3240 11676
rect 2538 11645 2550 11648
rect 2492 11639 2550 11645
rect 3234 11636 3240 11648
rect 3292 11636 3298 11688
rect 3878 11636 3884 11688
rect 3936 11676 3942 11688
rect 5074 11676 5080 11688
rect 3936 11648 5080 11676
rect 3936 11636 3942 11648
rect 5074 11636 5080 11648
rect 5132 11636 5138 11688
rect 7190 11676 7196 11688
rect 7151 11648 7196 11676
rect 7190 11636 7196 11648
rect 7248 11636 7254 11688
rect 8294 11636 8300 11688
rect 8352 11676 8358 11688
rect 11974 11676 11980 11688
rect 8352 11648 11980 11676
rect 8352 11636 8358 11648
rect 11974 11636 11980 11648
rect 12032 11636 12038 11688
rect 12805 11679 12863 11685
rect 12805 11676 12817 11679
rect 12084 11648 12817 11676
rect 2866 11568 2872 11620
rect 2924 11608 2930 11620
rect 8205 11611 8263 11617
rect 8205 11608 8217 11611
rect 2924 11580 8217 11608
rect 2924 11568 2930 11580
rect 8205 11577 8217 11580
rect 8251 11608 8263 11611
rect 8941 11611 8999 11617
rect 8941 11608 8953 11611
rect 8251 11580 8953 11608
rect 8251 11577 8263 11580
rect 8205 11571 8263 11577
rect 8941 11577 8953 11580
rect 8987 11577 8999 11611
rect 10873 11611 10931 11617
rect 10873 11608 10885 11611
rect 8941 11571 8999 11577
rect 9876 11580 10885 11608
rect 3602 11500 3608 11552
rect 3660 11540 3666 11552
rect 4338 11540 4344 11552
rect 3660 11512 4344 11540
rect 3660 11500 3666 11512
rect 4338 11500 4344 11512
rect 4396 11500 4402 11552
rect 7098 11500 7104 11552
rect 7156 11540 7162 11552
rect 7558 11540 7564 11552
rect 7156 11512 7564 11540
rect 7156 11500 7162 11512
rect 7558 11500 7564 11512
rect 7616 11500 7622 11552
rect 8846 11540 8852 11552
rect 8807 11512 8852 11540
rect 8846 11500 8852 11512
rect 8904 11500 8910 11552
rect 9122 11500 9128 11552
rect 9180 11540 9186 11552
rect 9876 11549 9904 11580
rect 10873 11577 10885 11580
rect 10919 11577 10931 11611
rect 10873 11571 10931 11577
rect 11609 11611 11667 11617
rect 11609 11577 11621 11611
rect 11655 11608 11667 11611
rect 11790 11608 11796 11620
rect 11655 11580 11796 11608
rect 11655 11577 11667 11580
rect 11609 11571 11667 11577
rect 11790 11568 11796 11580
rect 11848 11608 11854 11620
rect 12084 11608 12112 11648
rect 12805 11645 12817 11648
rect 12851 11676 12863 11679
rect 12851 11648 13216 11676
rect 12851 11645 12863 11648
rect 12805 11639 12863 11645
rect 11848 11580 12112 11608
rect 11848 11568 11854 11580
rect 12158 11568 12164 11620
rect 12216 11608 12222 11620
rect 12342 11608 12348 11620
rect 12216 11580 12348 11608
rect 12216 11568 12222 11580
rect 12342 11568 12348 11580
rect 12400 11608 12406 11620
rect 12897 11611 12955 11617
rect 12897 11608 12909 11611
rect 12400 11580 12909 11608
rect 12400 11568 12406 11580
rect 12897 11577 12909 11580
rect 12943 11577 12955 11611
rect 13188 11608 13216 11648
rect 13648 11620 13676 11716
rect 13906 11704 13912 11716
rect 13964 11704 13970 11756
rect 14093 11747 14151 11753
rect 14093 11713 14105 11747
rect 14139 11744 14151 11747
rect 14182 11744 14188 11756
rect 14139 11716 14188 11744
rect 14139 11713 14151 11716
rect 14093 11707 14151 11713
rect 14182 11704 14188 11716
rect 14240 11704 14246 11756
rect 17402 11704 17408 11756
rect 17460 11744 17466 11756
rect 17589 11747 17647 11753
rect 17589 11744 17601 11747
rect 17460 11716 17601 11744
rect 17460 11704 17466 11716
rect 17589 11713 17601 11716
rect 17635 11744 17647 11747
rect 17954 11744 17960 11756
rect 17635 11716 17960 11744
rect 17635 11713 17647 11716
rect 17589 11707 17647 11713
rect 17954 11704 17960 11716
rect 18012 11704 18018 11756
rect 18230 11744 18236 11756
rect 18064 11716 18236 11744
rect 13722 11636 13728 11688
rect 13780 11676 13786 11688
rect 13817 11679 13875 11685
rect 13817 11676 13829 11679
rect 13780 11648 13829 11676
rect 13780 11636 13786 11648
rect 13817 11645 13829 11648
rect 13863 11645 13875 11679
rect 13817 11639 13875 11645
rect 17313 11679 17371 11685
rect 17313 11645 17325 11679
rect 17359 11676 17371 11679
rect 17770 11676 17776 11688
rect 17359 11648 17776 11676
rect 17359 11645 17371 11648
rect 17313 11639 17371 11645
rect 17770 11636 17776 11648
rect 17828 11636 17834 11688
rect 18064 11676 18092 11716
rect 18230 11704 18236 11716
rect 18288 11704 18294 11756
rect 18598 11744 18604 11756
rect 18559 11716 18604 11744
rect 18598 11704 18604 11716
rect 18656 11704 18662 11756
rect 18877 11747 18935 11753
rect 18877 11713 18889 11747
rect 18923 11744 18935 11747
rect 19334 11744 19340 11756
rect 18923 11716 19340 11744
rect 18923 11713 18935 11716
rect 18877 11707 18935 11713
rect 19334 11704 19340 11716
rect 19392 11744 19398 11756
rect 19886 11744 19892 11756
rect 19392 11716 19892 11744
rect 19392 11704 19398 11716
rect 19886 11704 19892 11716
rect 19944 11704 19950 11756
rect 18414 11676 18420 11688
rect 17972 11648 18092 11676
rect 18375 11648 18420 11676
rect 13265 11611 13323 11617
rect 13265 11608 13277 11611
rect 13188 11580 13277 11608
rect 12897 11571 12955 11577
rect 13265 11577 13277 11580
rect 13311 11577 13323 11611
rect 13630 11608 13636 11620
rect 13543 11580 13636 11608
rect 13265 11571 13323 11577
rect 13630 11568 13636 11580
rect 13688 11608 13694 11620
rect 16758 11608 16764 11620
rect 13688 11580 16764 11608
rect 13688 11568 13694 11580
rect 16758 11568 16764 11580
rect 16816 11568 16822 11620
rect 17972 11608 18000 11648
rect 18414 11636 18420 11648
rect 18472 11636 18478 11688
rect 18506 11636 18512 11688
rect 18564 11676 18570 11688
rect 19981 11679 20039 11685
rect 19981 11676 19993 11679
rect 18564 11648 19993 11676
rect 18564 11636 18570 11648
rect 19981 11645 19993 11648
rect 20027 11645 20039 11679
rect 20990 11676 20996 11688
rect 19981 11639 20039 11645
rect 20088 11648 20996 11676
rect 16868 11580 18000 11608
rect 9861 11543 9919 11549
rect 9861 11540 9873 11543
rect 9180 11512 9873 11540
rect 9180 11500 9186 11512
rect 9861 11509 9873 11512
rect 9907 11509 9919 11543
rect 9861 11503 9919 11509
rect 9950 11500 9956 11552
rect 10008 11540 10014 11552
rect 10965 11543 11023 11549
rect 10965 11540 10977 11543
rect 10008 11512 10977 11540
rect 10008 11500 10014 11512
rect 10965 11509 10977 11512
rect 11011 11509 11023 11543
rect 11882 11540 11888 11552
rect 11843 11512 11888 11540
rect 10965 11503 11023 11509
rect 11882 11500 11888 11512
rect 11940 11500 11946 11552
rect 11974 11500 11980 11552
rect 12032 11540 12038 11552
rect 13357 11543 13415 11549
rect 13357 11540 13369 11543
rect 12032 11512 13369 11540
rect 12032 11500 12038 11512
rect 13357 11509 13369 11512
rect 13403 11509 13415 11543
rect 13357 11503 13415 11509
rect 13449 11543 13507 11549
rect 13449 11509 13461 11543
rect 13495 11540 13507 11543
rect 16868 11540 16896 11580
rect 18230 11568 18236 11620
rect 18288 11608 18294 11620
rect 20088 11608 20116 11648
rect 20990 11636 20996 11648
rect 21048 11636 21054 11688
rect 20254 11617 20260 11620
rect 20248 11608 20260 11617
rect 18288 11580 20116 11608
rect 20167 11580 20260 11608
rect 18288 11568 18294 11580
rect 20248 11571 20260 11580
rect 20312 11608 20318 11620
rect 20622 11608 20628 11620
rect 20312 11580 20628 11608
rect 20254 11568 20260 11571
rect 20312 11568 20318 11580
rect 20622 11568 20628 11580
rect 20680 11568 20686 11620
rect 13495 11512 16896 11540
rect 13495 11509 13507 11512
rect 13449 11503 13507 11509
rect 17678 11500 17684 11552
rect 17736 11540 17742 11552
rect 18049 11543 18107 11549
rect 18049 11540 18061 11543
rect 17736 11512 18061 11540
rect 17736 11500 17742 11512
rect 18049 11509 18061 11512
rect 18095 11509 18107 11543
rect 18049 11503 18107 11509
rect 18138 11500 18144 11552
rect 18196 11540 18202 11552
rect 18509 11543 18567 11549
rect 18509 11540 18521 11543
rect 18196 11512 18521 11540
rect 18196 11500 18202 11512
rect 18509 11509 18521 11512
rect 18555 11540 18567 11543
rect 18877 11543 18935 11549
rect 18877 11540 18889 11543
rect 18555 11512 18889 11540
rect 18555 11509 18567 11512
rect 18509 11503 18567 11509
rect 18877 11509 18889 11512
rect 18923 11509 18935 11543
rect 18877 11503 18935 11509
rect 18966 11500 18972 11552
rect 19024 11540 19030 11552
rect 19061 11543 19119 11549
rect 19061 11540 19073 11543
rect 19024 11512 19073 11540
rect 19024 11500 19030 11512
rect 19061 11509 19073 11512
rect 19107 11509 19119 11543
rect 19061 11503 19119 11509
rect 19242 11500 19248 11552
rect 19300 11540 19306 11552
rect 19613 11543 19671 11549
rect 19613 11540 19625 11543
rect 19300 11512 19625 11540
rect 19300 11500 19306 11512
rect 19613 11509 19625 11512
rect 19659 11509 19671 11543
rect 21358 11540 21364 11552
rect 21319 11512 21364 11540
rect 19613 11503 19671 11509
rect 21358 11500 21364 11512
rect 21416 11500 21422 11552
rect 1104 11450 21896 11472
rect 1104 11398 7912 11450
rect 7964 11398 7976 11450
rect 8028 11398 8040 11450
rect 8092 11398 8104 11450
rect 8156 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 15035 11450
rect 15087 11398 21896 11450
rect 1104 11376 21896 11398
rect 2409 11339 2467 11345
rect 2409 11305 2421 11339
rect 2455 11336 2467 11339
rect 2590 11336 2596 11348
rect 2455 11308 2596 11336
rect 2455 11305 2467 11308
rect 2409 11299 2467 11305
rect 2590 11296 2596 11308
rect 2648 11296 2654 11348
rect 2777 11339 2835 11345
rect 2777 11305 2789 11339
rect 2823 11336 2835 11339
rect 2866 11336 2872 11348
rect 2823 11308 2872 11336
rect 2823 11305 2835 11308
rect 2777 11299 2835 11305
rect 2866 11296 2872 11308
rect 2924 11296 2930 11348
rect 3234 11336 3240 11348
rect 3147 11308 3240 11336
rect 3234 11296 3240 11308
rect 3292 11336 3298 11348
rect 5442 11336 5448 11348
rect 3292 11308 5448 11336
rect 3292 11296 3298 11308
rect 5442 11296 5448 11308
rect 5500 11336 5506 11348
rect 5721 11339 5779 11345
rect 5721 11336 5733 11339
rect 5500 11308 5733 11336
rect 5500 11296 5506 11308
rect 5721 11305 5733 11308
rect 5767 11305 5779 11339
rect 6914 11336 6920 11348
rect 6875 11308 6920 11336
rect 5721 11299 5779 11305
rect 6914 11296 6920 11308
rect 6972 11296 6978 11348
rect 8846 11296 8852 11348
rect 8904 11336 8910 11348
rect 9677 11339 9735 11345
rect 9677 11336 9689 11339
rect 8904 11308 9689 11336
rect 8904 11296 8910 11308
rect 9677 11305 9689 11308
rect 9723 11305 9735 11339
rect 13909 11339 13967 11345
rect 13909 11336 13921 11339
rect 9677 11299 9735 11305
rect 10796 11308 13921 11336
rect 1946 11268 1952 11280
rect 1907 11240 1952 11268
rect 1946 11228 1952 11240
rect 2004 11228 2010 11280
rect 4890 11268 4896 11280
rect 2700 11240 4896 11268
rect 1673 11203 1731 11209
rect 1673 11169 1685 11203
rect 1719 11200 1731 11203
rect 2700 11200 2728 11240
rect 4890 11228 4896 11240
rect 4948 11228 4954 11280
rect 5074 11228 5080 11280
rect 5132 11268 5138 11280
rect 10796 11277 10824 11308
rect 13909 11305 13921 11308
rect 13955 11336 13967 11339
rect 14734 11336 14740 11348
rect 13955 11308 14740 11336
rect 13955 11305 13967 11308
rect 13909 11299 13967 11305
rect 14734 11296 14740 11308
rect 14792 11296 14798 11348
rect 15194 11296 15200 11348
rect 15252 11336 15258 11348
rect 17586 11336 17592 11348
rect 15252 11308 17592 11336
rect 15252 11296 15258 11308
rect 17586 11296 17592 11308
rect 17644 11296 17650 11348
rect 17681 11339 17739 11345
rect 17681 11305 17693 11339
rect 17727 11305 17739 11339
rect 17681 11299 17739 11305
rect 18969 11339 19027 11345
rect 18969 11305 18981 11339
rect 19015 11336 19027 11339
rect 19058 11336 19064 11348
rect 19015 11308 19064 11336
rect 19015 11305 19027 11308
rect 18969 11299 19027 11305
rect 10781 11271 10839 11277
rect 5132 11240 8248 11268
rect 5132 11228 5138 11240
rect 2958 11200 2964 11212
rect 1719 11172 2728 11200
rect 2792 11172 2964 11200
rect 1719 11169 1731 11172
rect 1673 11163 1731 11169
rect 1578 11092 1584 11144
rect 1636 11132 1642 11144
rect 2792 11132 2820 11172
rect 2958 11160 2964 11172
rect 3016 11160 3022 11212
rect 4608 11203 4666 11209
rect 4608 11169 4620 11203
rect 4654 11200 4666 11203
rect 5166 11200 5172 11212
rect 4654 11172 5172 11200
rect 4654 11169 4666 11172
rect 4608 11163 4666 11169
rect 5166 11160 5172 11172
rect 5224 11160 5230 11212
rect 6273 11203 6331 11209
rect 6273 11169 6285 11203
rect 6319 11200 6331 11203
rect 6638 11200 6644 11212
rect 6319 11172 6644 11200
rect 6319 11169 6331 11172
rect 6273 11163 6331 11169
rect 6638 11160 6644 11172
rect 6696 11200 6702 11212
rect 7009 11203 7067 11209
rect 7009 11200 7021 11203
rect 6696 11172 7021 11200
rect 6696 11160 6702 11172
rect 7009 11169 7021 11172
rect 7055 11169 7067 11203
rect 7009 11163 7067 11169
rect 7107 11172 7319 11200
rect 1636 11104 2820 11132
rect 2869 11135 2927 11141
rect 1636 11092 1642 11104
rect 2869 11101 2881 11135
rect 2915 11101 2927 11135
rect 2869 11095 2927 11101
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11132 3111 11135
rect 3237 11135 3295 11141
rect 3237 11132 3249 11135
rect 3099 11104 3249 11132
rect 3099 11101 3111 11104
rect 3053 11095 3111 11101
rect 3237 11101 3249 11104
rect 3283 11101 3295 11135
rect 3237 11095 3295 11101
rect 2884 11064 2912 11095
rect 4154 11092 4160 11144
rect 4212 11132 4218 11144
rect 4341 11135 4399 11141
rect 4341 11132 4353 11135
rect 4212 11104 4353 11132
rect 4212 11092 4218 11104
rect 4341 11101 4353 11104
rect 4387 11101 4399 11135
rect 6822 11132 6828 11144
rect 4341 11095 4399 11101
rect 5736 11104 6828 11132
rect 3510 11064 3516 11076
rect 2884 11036 3516 11064
rect 3510 11024 3516 11036
rect 3568 11024 3574 11076
rect 3694 10956 3700 11008
rect 3752 10996 3758 11008
rect 5736 10996 5764 11104
rect 6822 11092 6828 11104
rect 6880 11132 6886 11144
rect 7107 11132 7135 11172
rect 6880 11104 7135 11132
rect 7193 11135 7251 11141
rect 6880 11092 6886 11104
rect 7193 11101 7205 11135
rect 7239 11101 7251 11135
rect 7291 11132 7319 11172
rect 7742 11160 7748 11212
rect 7800 11200 7806 11212
rect 7929 11203 7987 11209
rect 7929 11200 7941 11203
rect 7800 11172 7941 11200
rect 7800 11160 7806 11172
rect 7929 11169 7941 11172
rect 7975 11169 7987 11203
rect 7929 11163 7987 11169
rect 8018 11132 8024 11144
rect 7291 11104 8024 11132
rect 7193 11095 7251 11101
rect 7208 11064 7236 11095
rect 8018 11092 8024 11104
rect 8076 11092 8082 11144
rect 8113 11135 8171 11141
rect 8113 11101 8125 11135
rect 8159 11101 8171 11135
rect 8220 11132 8248 11240
rect 10781 11237 10793 11271
rect 10827 11237 10839 11271
rect 10781 11231 10839 11237
rect 13078 11228 13084 11280
rect 13136 11268 13142 11280
rect 13173 11271 13231 11277
rect 13173 11268 13185 11271
rect 13136 11240 13185 11268
rect 13136 11228 13142 11240
rect 13173 11237 13185 11240
rect 13219 11237 13231 11271
rect 13173 11231 13231 11237
rect 14550 11228 14556 11280
rect 14608 11268 14614 11280
rect 15534 11271 15592 11277
rect 15534 11268 15546 11271
rect 14608 11240 15546 11268
rect 14608 11228 14614 11240
rect 15534 11237 15546 11240
rect 15580 11237 15592 11271
rect 15534 11231 15592 11237
rect 8757 11203 8815 11209
rect 8757 11169 8769 11203
rect 8803 11200 8815 11203
rect 12345 11203 12403 11209
rect 12345 11200 12357 11203
rect 8803 11172 12357 11200
rect 8803 11169 8815 11172
rect 8757 11163 8815 11169
rect 12345 11169 12357 11172
rect 12391 11200 12403 11203
rect 12434 11200 12440 11212
rect 12391 11172 12440 11200
rect 12391 11169 12403 11172
rect 12345 11163 12403 11169
rect 12434 11160 12440 11172
rect 12492 11160 12498 11212
rect 12526 11160 12532 11212
rect 12584 11200 12590 11212
rect 15194 11200 15200 11212
rect 12584 11172 15200 11200
rect 12584 11160 12590 11172
rect 15194 11160 15200 11172
rect 15252 11160 15258 11212
rect 15289 11203 15347 11209
rect 15289 11169 15301 11203
rect 15335 11200 15347 11203
rect 15930 11200 15936 11212
rect 15335 11172 15936 11200
rect 15335 11169 15347 11172
rect 15289 11163 15347 11169
rect 15930 11160 15936 11172
rect 15988 11160 15994 11212
rect 13265 11135 13323 11141
rect 8220 11104 13216 11132
rect 8113 11095 8171 11101
rect 7282 11064 7288 11076
rect 7195 11036 7288 11064
rect 7282 11024 7288 11036
rect 7340 11064 7346 11076
rect 8128 11064 8156 11095
rect 7340 11036 8156 11064
rect 7340 11024 7346 11036
rect 8202 11024 8208 11076
rect 8260 11064 8266 11076
rect 8573 11067 8631 11073
rect 8573 11064 8585 11067
rect 8260 11036 8585 11064
rect 8260 11024 8266 11036
rect 8573 11033 8585 11036
rect 8619 11033 8631 11067
rect 8573 11027 8631 11033
rect 9122 11024 9128 11076
rect 9180 11064 9186 11076
rect 9217 11067 9275 11073
rect 9217 11064 9229 11067
rect 9180 11036 9229 11064
rect 9180 11024 9186 11036
rect 9217 11033 9229 11036
rect 9263 11064 9275 11067
rect 10321 11067 10379 11073
rect 10321 11064 10333 11067
rect 9263 11036 10333 11064
rect 9263 11033 9275 11036
rect 9217 11027 9275 11033
rect 10321 11033 10333 11036
rect 10367 11033 10379 11067
rect 13188 11064 13216 11104
rect 13265 11101 13277 11135
rect 13311 11132 13323 11135
rect 13354 11132 13360 11144
rect 13311 11104 13360 11132
rect 13311 11101 13323 11104
rect 13265 11095 13323 11101
rect 13354 11092 13360 11104
rect 13412 11092 13418 11144
rect 13449 11135 13507 11141
rect 13449 11101 13461 11135
rect 13495 11132 13507 11135
rect 13630 11132 13636 11144
rect 13495 11104 13636 11132
rect 13495 11101 13507 11104
rect 13449 11095 13507 11101
rect 13630 11092 13636 11104
rect 13688 11092 13694 11144
rect 17687 11132 17715 11299
rect 19058 11296 19064 11308
rect 19116 11296 19122 11348
rect 20898 11296 20904 11348
rect 20956 11336 20962 11348
rect 21269 11339 21327 11345
rect 21269 11336 21281 11339
rect 20956 11308 21281 11336
rect 20956 11296 20962 11308
rect 21269 11305 21281 11308
rect 21315 11305 21327 11339
rect 21269 11299 21327 11305
rect 18782 11228 18788 11280
rect 18840 11268 18846 11280
rect 19150 11268 19156 11280
rect 18840 11240 19156 11268
rect 18840 11228 18846 11240
rect 19150 11228 19156 11240
rect 19208 11228 19214 11280
rect 18046 11200 18052 11212
rect 18007 11172 18052 11200
rect 18046 11160 18052 11172
rect 18104 11160 18110 11212
rect 19702 11200 19708 11212
rect 18248 11172 19708 11200
rect 17954 11132 17960 11144
rect 17687 11104 17960 11132
rect 17954 11092 17960 11104
rect 18012 11092 18018 11144
rect 18138 11132 18144 11144
rect 18099 11104 18144 11132
rect 18138 11092 18144 11104
rect 18196 11092 18202 11144
rect 14642 11064 14648 11076
rect 13188 11036 14648 11064
rect 10321 11027 10379 11033
rect 14642 11024 14648 11036
rect 14700 11024 14706 11076
rect 16666 11064 16672 11076
rect 16627 11036 16672 11064
rect 16666 11024 16672 11036
rect 16724 11024 16730 11076
rect 16850 11024 16856 11076
rect 16908 11064 16914 11076
rect 18248 11064 18276 11172
rect 19702 11160 19708 11172
rect 19760 11200 19766 11212
rect 20165 11203 20223 11209
rect 20165 11200 20177 11203
rect 19760 11172 20177 11200
rect 19760 11160 19766 11172
rect 20165 11169 20177 11172
rect 20211 11169 20223 11203
rect 20165 11163 20223 11169
rect 18325 11135 18383 11141
rect 18325 11101 18337 11135
rect 18371 11132 18383 11135
rect 19150 11132 19156 11144
rect 18371 11104 19156 11132
rect 18371 11101 18383 11104
rect 18325 11095 18383 11101
rect 19150 11092 19156 11104
rect 19208 11092 19214 11144
rect 19886 11132 19892 11144
rect 19847 11104 19892 11132
rect 19886 11092 19892 11104
rect 19944 11092 19950 11144
rect 20254 11092 20260 11144
rect 20312 11132 20318 11144
rect 20438 11132 20444 11144
rect 20312 11104 20444 11132
rect 20312 11092 20318 11104
rect 20438 11092 20444 11104
rect 20496 11092 20502 11144
rect 19242 11064 19248 11076
rect 16908 11036 18276 11064
rect 19203 11036 19248 11064
rect 16908 11024 16914 11036
rect 19242 11024 19248 11036
rect 19300 11024 19306 11076
rect 19518 11024 19524 11076
rect 19576 11064 19582 11076
rect 20070 11064 20076 11076
rect 19576 11036 20076 11064
rect 19576 11024 19582 11036
rect 20070 11024 20076 11036
rect 20128 11064 20134 11076
rect 20901 11067 20959 11073
rect 20901 11064 20913 11067
rect 20128 11036 20913 11064
rect 20128 11024 20134 11036
rect 20901 11033 20913 11036
rect 20947 11033 20959 11067
rect 20901 11027 20959 11033
rect 6546 10996 6552 11008
rect 3752 10968 5764 10996
rect 6507 10968 6552 10996
rect 3752 10956 3758 10968
rect 6546 10956 6552 10968
rect 6604 10956 6610 11008
rect 6914 10956 6920 11008
rect 6972 10996 6978 11008
rect 7561 10999 7619 11005
rect 7561 10996 7573 10999
rect 6972 10968 7573 10996
rect 6972 10956 6978 10968
rect 7561 10965 7573 10968
rect 7607 10965 7619 10999
rect 12802 10996 12808 11008
rect 12763 10968 12808 10996
rect 7561 10959 7619 10965
rect 12802 10956 12808 10968
rect 12860 10956 12866 11008
rect 15470 10956 15476 11008
rect 15528 10996 15534 11008
rect 18874 10996 18880 11008
rect 15528 10968 18880 10996
rect 15528 10956 15534 10968
rect 18874 10956 18880 10968
rect 18932 10956 18938 11008
rect 1104 10906 21896 10928
rect 1104 10854 4447 10906
rect 4499 10854 4511 10906
rect 4563 10854 4575 10906
rect 4627 10854 4639 10906
rect 4691 10854 11378 10906
rect 11430 10854 11442 10906
rect 11494 10854 11506 10906
rect 11558 10854 11570 10906
rect 11622 10854 18308 10906
rect 18360 10854 18372 10906
rect 18424 10854 18436 10906
rect 18488 10854 18500 10906
rect 18552 10854 21896 10906
rect 1104 10832 21896 10854
rect 1578 10792 1584 10804
rect 1539 10764 1584 10792
rect 1578 10752 1584 10764
rect 1636 10752 1642 10804
rect 2774 10752 2780 10804
rect 2832 10792 2838 10804
rect 2832 10764 2877 10792
rect 2832 10752 2838 10764
rect 4062 10752 4068 10804
rect 4120 10792 4126 10804
rect 4120 10764 5120 10792
rect 4120 10752 4126 10764
rect 5092 10724 5120 10764
rect 5166 10752 5172 10804
rect 5224 10792 5230 10804
rect 5261 10795 5319 10801
rect 5261 10792 5273 10795
rect 5224 10764 5273 10792
rect 5224 10752 5230 10764
rect 5261 10761 5273 10764
rect 5307 10761 5319 10795
rect 9125 10795 9183 10801
rect 9125 10792 9137 10795
rect 5261 10755 5319 10761
rect 7024 10764 9137 10792
rect 7024 10724 7052 10764
rect 9125 10761 9137 10764
rect 9171 10761 9183 10795
rect 12526 10792 12532 10804
rect 12439 10764 12532 10792
rect 9125 10755 9183 10761
rect 5092 10696 7052 10724
rect 8018 10684 8024 10736
rect 8076 10724 8082 10736
rect 8665 10727 8723 10733
rect 8665 10724 8677 10727
rect 8076 10696 8677 10724
rect 8076 10684 8082 10696
rect 8665 10693 8677 10696
rect 8711 10693 8723 10727
rect 8665 10687 8723 10693
rect 6365 10659 6423 10665
rect 6365 10656 6377 10659
rect 6104 10628 6377 10656
rect 1854 10588 1860 10600
rect 1815 10560 1860 10588
rect 1854 10548 1860 10560
rect 1912 10548 1918 10600
rect 2133 10591 2191 10597
rect 2133 10557 2145 10591
rect 2179 10588 2191 10591
rect 2593 10591 2651 10597
rect 2593 10588 2605 10591
rect 2179 10560 2605 10588
rect 2179 10557 2191 10560
rect 2133 10551 2191 10557
rect 2593 10557 2605 10560
rect 2639 10557 2651 10591
rect 2593 10551 2651 10557
rect 3881 10591 3939 10597
rect 3881 10557 3893 10591
rect 3927 10557 3939 10591
rect 3881 10551 3939 10557
rect 4148 10591 4206 10597
rect 4148 10557 4160 10591
rect 4194 10588 4206 10591
rect 6104 10588 6132 10628
rect 6365 10625 6377 10628
rect 6411 10656 6423 10659
rect 6638 10656 6644 10668
rect 6411 10628 6644 10656
rect 6411 10625 6423 10628
rect 6365 10619 6423 10625
rect 6638 10616 6644 10628
rect 6696 10656 6702 10668
rect 9140 10656 9168 10755
rect 12526 10752 12532 10764
rect 12584 10792 12590 10804
rect 13354 10792 13360 10804
rect 12584 10764 13360 10792
rect 12584 10752 12590 10764
rect 13354 10752 13360 10764
rect 13412 10792 13418 10804
rect 16022 10792 16028 10804
rect 13412 10764 16028 10792
rect 13412 10752 13418 10764
rect 16022 10752 16028 10764
rect 16080 10792 16086 10804
rect 19978 10792 19984 10804
rect 16080 10764 19984 10792
rect 16080 10752 16086 10764
rect 19978 10752 19984 10764
rect 20036 10752 20042 10804
rect 20622 10792 20628 10804
rect 20583 10764 20628 10792
rect 20622 10752 20628 10764
rect 20680 10752 20686 10804
rect 9493 10727 9551 10733
rect 9493 10693 9505 10727
rect 9539 10724 9551 10727
rect 10778 10724 10784 10736
rect 9539 10696 10784 10724
rect 9539 10693 9551 10696
rect 9493 10687 9551 10693
rect 10778 10684 10784 10696
rect 10836 10684 10842 10736
rect 13081 10727 13139 10733
rect 13081 10693 13093 10727
rect 13127 10724 13139 10727
rect 14090 10724 14096 10736
rect 13127 10696 14096 10724
rect 13127 10693 13139 10696
rect 13081 10687 13139 10693
rect 14090 10684 14096 10696
rect 14148 10684 14154 10736
rect 18049 10727 18107 10733
rect 18049 10693 18061 10727
rect 18095 10693 18107 10727
rect 18049 10687 18107 10693
rect 18248 10696 19288 10724
rect 9953 10659 10011 10665
rect 9953 10656 9965 10659
rect 6696 10628 7135 10656
rect 9140 10628 9965 10656
rect 6696 10616 6702 10628
rect 4194 10560 6132 10588
rect 6181 10591 6239 10597
rect 4194 10557 4206 10560
rect 4148 10551 4206 10557
rect 6181 10557 6193 10591
rect 6227 10588 6239 10591
rect 6546 10588 6552 10600
rect 6227 10560 6552 10588
rect 6227 10557 6239 10560
rect 6181 10551 6239 10557
rect 3896 10452 3924 10551
rect 6546 10548 6552 10560
rect 6604 10548 6610 10600
rect 7009 10591 7067 10597
rect 7009 10557 7021 10591
rect 7055 10557 7067 10591
rect 7009 10551 7067 10557
rect 6089 10523 6147 10529
rect 6089 10489 6101 10523
rect 6135 10520 6147 10523
rect 6914 10520 6920 10532
rect 6135 10492 6920 10520
rect 6135 10489 6147 10492
rect 6089 10483 6147 10489
rect 6914 10480 6920 10492
rect 6972 10480 6978 10532
rect 4154 10452 4160 10464
rect 3896 10424 4160 10452
rect 4154 10412 4160 10424
rect 4212 10412 4218 10464
rect 5718 10452 5724 10464
rect 5679 10424 5724 10452
rect 5718 10412 5724 10424
rect 5776 10412 5782 10464
rect 7024 10452 7052 10551
rect 7107 10520 7135 10628
rect 9953 10625 9965 10628
rect 9999 10625 10011 10659
rect 10134 10656 10140 10668
rect 10095 10628 10140 10656
rect 9953 10619 10011 10625
rect 10134 10616 10140 10628
rect 10192 10616 10198 10668
rect 14645 10659 14703 10665
rect 14645 10625 14657 10659
rect 14691 10656 14703 10659
rect 14734 10656 14740 10668
rect 14691 10628 14740 10656
rect 14691 10625 14703 10628
rect 14645 10619 14703 10625
rect 14734 10616 14740 10628
rect 14792 10616 14798 10668
rect 18064 10656 18092 10687
rect 18138 10656 18144 10668
rect 18064 10628 18144 10656
rect 18138 10616 18144 10628
rect 18196 10616 18202 10668
rect 7282 10597 7288 10600
rect 7276 10588 7288 10597
rect 7243 10560 7288 10588
rect 7276 10551 7288 10560
rect 7282 10548 7288 10551
rect 7340 10548 7346 10600
rect 12434 10548 12440 10600
rect 12492 10588 12498 10600
rect 13265 10591 13323 10597
rect 13265 10588 13277 10591
rect 12492 10560 13277 10588
rect 12492 10548 12498 10560
rect 13265 10557 13277 10560
rect 13311 10557 13323 10591
rect 13265 10551 13323 10557
rect 14550 10548 14556 10600
rect 14608 10588 14614 10600
rect 17678 10588 17684 10600
rect 14608 10560 17684 10588
rect 14608 10548 14614 10560
rect 17678 10548 17684 10560
rect 17736 10548 17742 10600
rect 17862 10548 17868 10600
rect 17920 10588 17926 10600
rect 18248 10588 18276 10696
rect 18598 10656 18604 10668
rect 18559 10628 18604 10656
rect 18598 10616 18604 10628
rect 18656 10616 18662 10668
rect 19260 10665 19288 10696
rect 19245 10659 19303 10665
rect 19245 10625 19257 10659
rect 19291 10625 19303 10659
rect 19245 10619 19303 10625
rect 17920 10560 18276 10588
rect 18509 10591 18567 10597
rect 17920 10548 17926 10560
rect 18509 10557 18521 10591
rect 18555 10588 18567 10591
rect 19058 10588 19064 10600
rect 18555 10560 19064 10588
rect 18555 10557 18567 10560
rect 18509 10551 18567 10557
rect 19058 10548 19064 10560
rect 19116 10548 19122 10600
rect 9861 10523 9919 10529
rect 7107 10492 8432 10520
rect 8294 10452 8300 10464
rect 7024 10424 8300 10452
rect 8294 10412 8300 10424
rect 8352 10412 8358 10464
rect 8404 10461 8432 10492
rect 9861 10489 9873 10523
rect 9907 10520 9919 10523
rect 10505 10523 10563 10529
rect 10505 10520 10517 10523
rect 9907 10492 10517 10520
rect 9907 10489 9919 10492
rect 9861 10483 9919 10489
rect 10505 10489 10517 10492
rect 10551 10489 10563 10523
rect 10505 10483 10563 10489
rect 13814 10480 13820 10532
rect 13872 10520 13878 10532
rect 14461 10523 14519 10529
rect 14461 10520 14473 10523
rect 13872 10492 14473 10520
rect 13872 10480 13878 10492
rect 14461 10489 14473 10492
rect 14507 10489 14519 10523
rect 18417 10523 18475 10529
rect 18417 10520 18429 10523
rect 14461 10483 14519 10489
rect 17144 10492 18429 10520
rect 17144 10464 17172 10492
rect 18417 10489 18429 10492
rect 18463 10489 18475 10523
rect 18417 10483 18475 10489
rect 19150 10480 19156 10532
rect 19208 10520 19214 10532
rect 19490 10523 19548 10529
rect 19490 10520 19502 10523
rect 19208 10492 19502 10520
rect 19208 10480 19214 10492
rect 19490 10489 19502 10492
rect 19536 10489 19548 10523
rect 19490 10483 19548 10489
rect 8389 10455 8447 10461
rect 8389 10421 8401 10455
rect 8435 10421 8447 10455
rect 13998 10452 14004 10464
rect 13959 10424 14004 10452
rect 8389 10415 8447 10421
rect 13998 10412 14004 10424
rect 14056 10412 14062 10464
rect 14366 10452 14372 10464
rect 14327 10424 14372 10452
rect 14366 10412 14372 10424
rect 14424 10412 14430 10464
rect 17126 10452 17132 10464
rect 17087 10424 17132 10452
rect 17126 10412 17132 10424
rect 17184 10412 17190 10464
rect 17497 10455 17555 10461
rect 17497 10421 17509 10455
rect 17543 10452 17555 10455
rect 18138 10452 18144 10464
rect 17543 10424 18144 10452
rect 17543 10421 17555 10424
rect 17497 10415 17555 10421
rect 18138 10412 18144 10424
rect 18196 10412 18202 10464
rect 1104 10362 21896 10384
rect 1104 10310 7912 10362
rect 7964 10310 7976 10362
rect 8028 10310 8040 10362
rect 8092 10310 8104 10362
rect 8156 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 15035 10362
rect 15087 10310 21896 10362
rect 1104 10288 21896 10310
rect 1854 10208 1860 10260
rect 1912 10248 1918 10260
rect 2317 10251 2375 10257
rect 2317 10248 2329 10251
rect 1912 10220 2329 10248
rect 1912 10208 1918 10220
rect 2317 10217 2329 10220
rect 2363 10217 2375 10251
rect 4890 10248 4896 10260
rect 4851 10220 4896 10248
rect 2317 10211 2375 10217
rect 4890 10208 4896 10220
rect 4948 10208 4954 10260
rect 5353 10251 5411 10257
rect 5353 10217 5365 10251
rect 5399 10248 5411 10251
rect 5905 10251 5963 10257
rect 5905 10248 5917 10251
rect 5399 10220 5917 10248
rect 5399 10217 5411 10220
rect 5353 10211 5411 10217
rect 5905 10217 5917 10220
rect 5951 10217 5963 10251
rect 5905 10211 5963 10217
rect 6273 10251 6331 10257
rect 6273 10217 6285 10251
rect 6319 10248 6331 10251
rect 6917 10251 6975 10257
rect 6917 10248 6929 10251
rect 6319 10220 6929 10248
rect 6319 10217 6331 10220
rect 6273 10211 6331 10217
rect 6917 10217 6929 10220
rect 6963 10217 6975 10251
rect 6917 10211 6975 10217
rect 7742 10208 7748 10260
rect 7800 10248 7806 10260
rect 7929 10251 7987 10257
rect 7929 10248 7941 10251
rect 7800 10220 7941 10248
rect 7800 10208 7806 10220
rect 7929 10217 7941 10220
rect 7975 10217 7987 10251
rect 7929 10211 7987 10217
rect 14366 10208 14372 10260
rect 14424 10248 14430 10260
rect 15289 10251 15347 10257
rect 15289 10248 15301 10251
rect 14424 10220 15301 10248
rect 14424 10208 14430 10220
rect 15289 10217 15301 10220
rect 15335 10217 15347 10251
rect 15289 10211 15347 10217
rect 15764 10220 18736 10248
rect 4062 10140 4068 10192
rect 4120 10180 4126 10192
rect 14550 10180 14556 10192
rect 4120 10152 14556 10180
rect 4120 10140 4126 10152
rect 14550 10140 14556 10152
rect 14608 10140 14614 10192
rect 14642 10140 14648 10192
rect 14700 10180 14706 10192
rect 15764 10189 15792 10220
rect 14829 10183 14887 10189
rect 14829 10180 14841 10183
rect 14700 10152 14841 10180
rect 14700 10140 14706 10152
rect 14829 10149 14841 10152
rect 14875 10180 14887 10183
rect 15749 10183 15807 10189
rect 15749 10180 15761 10183
rect 14875 10152 15761 10180
rect 14875 10149 14887 10152
rect 14829 10143 14887 10149
rect 15749 10149 15761 10152
rect 15795 10149 15807 10183
rect 17862 10180 17868 10192
rect 15749 10143 15807 10149
rect 16592 10152 17868 10180
rect 16592 10124 16620 10152
rect 17862 10140 17868 10152
rect 17920 10180 17926 10192
rect 18408 10183 18466 10189
rect 18408 10180 18420 10183
rect 17920 10152 18184 10180
rect 17920 10140 17926 10152
rect 2682 10112 2688 10124
rect 2643 10084 2688 10112
rect 2682 10072 2688 10084
rect 2740 10072 2746 10124
rect 5261 10115 5319 10121
rect 5261 10081 5273 10115
rect 5307 10112 5319 10115
rect 5718 10112 5724 10124
rect 5307 10084 5724 10112
rect 5307 10081 5319 10084
rect 5261 10075 5319 10081
rect 5718 10072 5724 10084
rect 5776 10072 5782 10124
rect 6454 10072 6460 10124
rect 6512 10112 6518 10124
rect 7285 10115 7343 10121
rect 7285 10112 7297 10115
rect 6512 10084 7297 10112
rect 6512 10072 6518 10084
rect 7285 10081 7297 10084
rect 7331 10081 7343 10115
rect 7285 10075 7343 10081
rect 7377 10115 7435 10121
rect 7377 10081 7389 10115
rect 7423 10112 7435 10115
rect 7423 10084 7604 10112
rect 7423 10081 7435 10084
rect 7377 10075 7435 10081
rect 2774 10004 2780 10056
rect 2832 10044 2838 10056
rect 2961 10047 3019 10053
rect 2832 10016 2877 10044
rect 2832 10004 2838 10016
rect 2961 10013 2973 10047
rect 3007 10044 3019 10047
rect 3418 10044 3424 10056
rect 3007 10016 3424 10044
rect 3007 10013 3019 10016
rect 2961 10007 3019 10013
rect 3418 10004 3424 10016
rect 3476 10004 3482 10056
rect 5166 10004 5172 10056
rect 5224 10044 5230 10056
rect 5445 10047 5503 10053
rect 5445 10044 5457 10047
rect 5224 10016 5457 10044
rect 5224 10004 5230 10016
rect 5445 10013 5457 10016
rect 5491 10013 5503 10047
rect 6362 10044 6368 10056
rect 6323 10016 6368 10044
rect 5445 10007 5503 10013
rect 6362 10004 6368 10016
rect 6420 10004 6426 10056
rect 6549 10047 6607 10053
rect 6549 10013 6561 10047
rect 6595 10044 6607 10047
rect 6638 10044 6644 10056
rect 6595 10016 6644 10044
rect 6595 10013 6607 10016
rect 6549 10007 6607 10013
rect 6638 10004 6644 10016
rect 6696 10004 6702 10056
rect 7469 10047 7527 10053
rect 7469 10013 7481 10047
rect 7515 10013 7527 10047
rect 7469 10007 7527 10013
rect 2406 9936 2412 9988
rect 2464 9976 2470 9988
rect 6914 9976 6920 9988
rect 2464 9948 6920 9976
rect 2464 9936 2470 9948
rect 6914 9936 6920 9948
rect 6972 9936 6978 9988
rect 7282 9936 7288 9988
rect 7340 9976 7346 9988
rect 7484 9976 7512 10007
rect 7340 9948 7512 9976
rect 7340 9936 7346 9948
rect 7576 9908 7604 10084
rect 8294 10072 8300 10124
rect 8352 10112 8358 10124
rect 9677 10115 9735 10121
rect 9677 10112 9689 10115
rect 8352 10084 9689 10112
rect 8352 10072 8358 10084
rect 9677 10081 9689 10084
rect 9723 10081 9735 10115
rect 9677 10075 9735 10081
rect 9944 10115 10002 10121
rect 9944 10081 9956 10115
rect 9990 10112 10002 10115
rect 10226 10112 10232 10124
rect 9990 10084 10232 10112
rect 9990 10081 10002 10084
rect 9944 10075 10002 10081
rect 10226 10072 10232 10084
rect 10284 10072 10290 10124
rect 11238 10112 11244 10124
rect 11072 10084 11244 10112
rect 11072 9985 11100 10084
rect 11238 10072 11244 10084
rect 11296 10112 11302 10124
rect 11589 10115 11647 10121
rect 11589 10112 11601 10115
rect 11296 10084 11601 10112
rect 11296 10072 11302 10084
rect 11589 10081 11601 10084
rect 11635 10081 11647 10115
rect 11589 10075 11647 10081
rect 13078 10072 13084 10124
rect 13136 10112 13142 10124
rect 13245 10115 13303 10121
rect 13245 10112 13257 10115
rect 13136 10084 13257 10112
rect 13136 10072 13142 10084
rect 13245 10081 13257 10084
rect 13291 10112 13303 10115
rect 15654 10112 15660 10124
rect 13291 10084 15240 10112
rect 15615 10084 15660 10112
rect 13291 10081 13303 10084
rect 13245 10075 13303 10081
rect 11333 10047 11391 10053
rect 11333 10013 11345 10047
rect 11379 10013 11391 10047
rect 12986 10044 12992 10056
rect 11333 10007 11391 10013
rect 12452 10016 12992 10044
rect 11057 9979 11115 9985
rect 11057 9945 11069 9979
rect 11103 9945 11115 9979
rect 11057 9939 11115 9945
rect 8481 9911 8539 9917
rect 8481 9908 8493 9911
rect 7576 9880 8493 9908
rect 8481 9877 8493 9880
rect 8527 9908 8539 9911
rect 10962 9908 10968 9920
rect 8527 9880 10968 9908
rect 8527 9877 8539 9880
rect 8481 9871 8539 9877
rect 10962 9868 10968 9880
rect 11020 9868 11026 9920
rect 11348 9908 11376 10007
rect 12452 9908 12480 10016
rect 12986 10004 12992 10016
rect 13044 10004 13050 10056
rect 15212 9976 15240 10084
rect 15654 10072 15660 10084
rect 15712 10072 15718 10124
rect 16485 10115 16543 10121
rect 16485 10081 16497 10115
rect 16531 10112 16543 10115
rect 16574 10112 16580 10124
rect 16531 10084 16580 10112
rect 16531 10081 16543 10084
rect 16485 10075 16543 10081
rect 16574 10072 16580 10084
rect 16632 10072 16638 10124
rect 16758 10121 16764 10124
rect 16752 10075 16764 10121
rect 16816 10112 16822 10124
rect 18156 10121 18184 10152
rect 18248 10152 18420 10180
rect 18141 10115 18199 10121
rect 16816 10084 16852 10112
rect 16758 10072 16764 10075
rect 16816 10072 16822 10084
rect 18141 10081 18153 10115
rect 18187 10081 18199 10115
rect 18141 10075 18199 10081
rect 15841 10047 15899 10053
rect 15841 10013 15853 10047
rect 15887 10013 15899 10047
rect 18248 10044 18276 10152
rect 18408 10149 18420 10152
rect 18454 10180 18466 10183
rect 18598 10180 18604 10192
rect 18454 10152 18604 10180
rect 18454 10149 18466 10152
rect 18408 10143 18466 10149
rect 18598 10140 18604 10152
rect 18656 10140 18662 10192
rect 18708 10180 18736 10220
rect 19150 10208 19156 10260
rect 19208 10248 19214 10260
rect 19521 10251 19579 10257
rect 19521 10248 19533 10251
rect 19208 10220 19533 10248
rect 19208 10208 19214 10220
rect 19521 10217 19533 10220
rect 19567 10217 19579 10251
rect 19521 10211 19579 10217
rect 20254 10180 20260 10192
rect 18708 10152 20260 10180
rect 20254 10140 20260 10152
rect 20312 10180 20318 10192
rect 20993 10183 21051 10189
rect 20993 10180 21005 10183
rect 20312 10152 21005 10180
rect 20312 10140 20318 10152
rect 20993 10149 21005 10152
rect 21039 10149 21051 10183
rect 20993 10143 21051 10149
rect 20165 10115 20223 10121
rect 20165 10081 20177 10115
rect 20211 10112 20223 10115
rect 20898 10112 20904 10124
rect 20211 10084 20904 10112
rect 20211 10081 20223 10084
rect 20165 10075 20223 10081
rect 20898 10072 20904 10084
rect 20956 10072 20962 10124
rect 15841 10007 15899 10013
rect 17880 10016 18276 10044
rect 20441 10047 20499 10053
rect 15856 9976 15884 10007
rect 16206 9976 16212 9988
rect 15212 9948 16212 9976
rect 16206 9936 16212 9948
rect 16264 9936 16270 9988
rect 17880 9985 17908 10016
rect 20441 10013 20453 10047
rect 20487 10044 20499 10047
rect 20714 10044 20720 10056
rect 20487 10016 20720 10044
rect 20487 10013 20499 10016
rect 20441 10007 20499 10013
rect 20714 10004 20720 10016
rect 20772 10044 20778 10056
rect 21358 10044 21364 10056
rect 20772 10016 21364 10044
rect 20772 10004 20778 10016
rect 21358 10004 21364 10016
rect 21416 10004 21422 10056
rect 17865 9979 17923 9985
rect 17865 9945 17877 9979
rect 17911 9945 17923 9979
rect 17865 9939 17923 9945
rect 12710 9908 12716 9920
rect 11348 9880 12480 9908
rect 12671 9880 12716 9908
rect 12710 9868 12716 9880
rect 12768 9868 12774 9920
rect 14369 9911 14427 9917
rect 14369 9877 14381 9911
rect 14415 9908 14427 9911
rect 14734 9908 14740 9920
rect 14415 9880 14740 9908
rect 14415 9877 14427 9880
rect 14369 9871 14427 9877
rect 14734 9868 14740 9880
rect 14792 9868 14798 9920
rect 16224 9908 16252 9936
rect 16666 9908 16672 9920
rect 16224 9880 16672 9908
rect 16666 9868 16672 9880
rect 16724 9868 16730 9920
rect 19702 9868 19708 9920
rect 19760 9908 19766 9920
rect 19797 9911 19855 9917
rect 19797 9908 19809 9911
rect 19760 9880 19809 9908
rect 19760 9868 19766 9880
rect 19797 9877 19809 9880
rect 19843 9877 19855 9911
rect 19797 9871 19855 9877
rect 1104 9818 21896 9840
rect 1104 9766 4447 9818
rect 4499 9766 4511 9818
rect 4563 9766 4575 9818
rect 4627 9766 4639 9818
rect 4691 9766 11378 9818
rect 11430 9766 11442 9818
rect 11494 9766 11506 9818
rect 11558 9766 11570 9818
rect 11622 9766 18308 9818
rect 18360 9766 18372 9818
rect 18424 9766 18436 9818
rect 18488 9766 18500 9818
rect 18552 9766 21896 9818
rect 1104 9744 21896 9766
rect 4062 9664 4068 9716
rect 4120 9704 4126 9716
rect 4120 9676 6316 9704
rect 4120 9664 4126 9676
rect 6288 9636 6316 9676
rect 6362 9664 6368 9716
rect 6420 9704 6426 9716
rect 6825 9707 6883 9713
rect 6825 9704 6837 9707
rect 6420 9676 6837 9704
rect 6420 9664 6426 9676
rect 6825 9673 6837 9676
rect 6871 9673 6883 9707
rect 12526 9704 12532 9716
rect 6825 9667 6883 9673
rect 6932 9676 12532 9704
rect 6932 9636 6960 9676
rect 12526 9664 12532 9676
rect 12584 9664 12590 9716
rect 17862 9664 17868 9716
rect 17920 9704 17926 9716
rect 17920 9676 18736 9704
rect 17920 9664 17926 9676
rect 6288 9608 6960 9636
rect 9401 9639 9459 9645
rect 9401 9605 9413 9639
rect 9447 9636 9459 9639
rect 9490 9636 9496 9648
rect 9447 9608 9496 9636
rect 9447 9605 9459 9608
rect 9401 9599 9459 9605
rect 9490 9596 9496 9608
rect 9548 9596 9554 9648
rect 16761 9639 16819 9645
rect 16761 9605 16773 9639
rect 16807 9636 16819 9639
rect 16850 9636 16856 9648
rect 16807 9608 16856 9636
rect 16807 9605 16819 9608
rect 16761 9599 16819 9605
rect 16850 9596 16856 9608
rect 16908 9596 16914 9648
rect 18046 9636 18052 9648
rect 18007 9608 18052 9636
rect 18046 9596 18052 9608
rect 18104 9596 18110 9648
rect 7282 9528 7288 9580
rect 7340 9568 7346 9580
rect 7377 9571 7435 9577
rect 7377 9568 7389 9571
rect 7340 9540 7389 9568
rect 7340 9528 7346 9540
rect 7377 9537 7389 9540
rect 7423 9537 7435 9571
rect 7377 9531 7435 9537
rect 9309 9571 9367 9577
rect 9309 9537 9321 9571
rect 9355 9568 9367 9571
rect 9950 9568 9956 9580
rect 9355 9540 9956 9568
rect 9355 9537 9367 9540
rect 9309 9531 9367 9537
rect 9950 9528 9956 9540
rect 10008 9528 10014 9580
rect 10134 9568 10140 9580
rect 10095 9540 10140 9568
rect 10134 9528 10140 9540
rect 10192 9528 10198 9580
rect 11149 9571 11207 9577
rect 11149 9537 11161 9571
rect 11195 9568 11207 9571
rect 11238 9568 11244 9580
rect 11195 9540 11244 9568
rect 11195 9537 11207 9540
rect 11149 9531 11207 9537
rect 11238 9528 11244 9540
rect 11296 9528 11302 9580
rect 14090 9528 14096 9580
rect 14148 9568 14154 9580
rect 15197 9571 15255 9577
rect 14148 9540 14964 9568
rect 14148 9528 14154 9540
rect 2041 9503 2099 9509
rect 2041 9469 2053 9503
rect 2087 9500 2099 9503
rect 8021 9503 8079 9509
rect 2087 9472 2268 9500
rect 2087 9469 2099 9472
rect 2041 9463 2099 9469
rect 2240 9364 2268 9472
rect 8021 9469 8033 9503
rect 8067 9500 8079 9503
rect 8202 9500 8208 9512
rect 8067 9472 8208 9500
rect 8067 9469 8079 9472
rect 8021 9463 8079 9469
rect 8202 9460 8208 9472
rect 8260 9460 8266 9512
rect 8849 9503 8907 9509
rect 8849 9469 8861 9503
rect 8895 9500 8907 9503
rect 9582 9500 9588 9512
rect 8895 9472 9588 9500
rect 8895 9469 8907 9472
rect 8849 9463 8907 9469
rect 2308 9435 2366 9441
rect 2308 9401 2320 9435
rect 2354 9432 2366 9435
rect 2866 9432 2872 9444
rect 2354 9404 2872 9432
rect 2354 9401 2366 9404
rect 2308 9395 2366 9401
rect 2866 9392 2872 9404
rect 2924 9392 2930 9444
rect 3970 9392 3976 9444
rect 4028 9432 4034 9444
rect 8864 9432 8892 9463
rect 9582 9460 9588 9472
rect 9640 9460 9646 9512
rect 10965 9503 11023 9509
rect 10965 9500 10977 9503
rect 9692 9472 10977 9500
rect 4028 9404 8892 9432
rect 9217 9435 9275 9441
rect 4028 9392 4034 9404
rect 9217 9401 9229 9435
rect 9263 9432 9275 9435
rect 9309 9435 9367 9441
rect 9309 9432 9321 9435
rect 9263 9404 9321 9432
rect 9263 9401 9275 9404
rect 9217 9395 9275 9401
rect 9309 9401 9321 9404
rect 9355 9401 9367 9435
rect 9309 9395 9367 9401
rect 2498 9364 2504 9376
rect 2240 9336 2504 9364
rect 2498 9324 2504 9336
rect 2556 9324 2562 9376
rect 3418 9364 3424 9376
rect 3379 9336 3424 9364
rect 3418 9324 3424 9336
rect 3476 9324 3482 9376
rect 6454 9364 6460 9376
rect 6415 9336 6460 9364
rect 6454 9324 6460 9336
rect 6512 9324 6518 9376
rect 6822 9324 6828 9376
rect 6880 9364 6886 9376
rect 7193 9367 7251 9373
rect 7193 9364 7205 9367
rect 6880 9336 7205 9364
rect 6880 9324 6886 9336
rect 7193 9333 7205 9336
rect 7239 9333 7251 9367
rect 7193 9327 7251 9333
rect 7285 9367 7343 9373
rect 7285 9333 7297 9367
rect 7331 9364 7343 9367
rect 7374 9364 7380 9376
rect 7331 9336 7380 9364
rect 7331 9333 7343 9336
rect 7285 9327 7343 9333
rect 7374 9324 7380 9336
rect 7432 9324 7438 9376
rect 7837 9367 7895 9373
rect 7837 9333 7849 9367
rect 7883 9364 7895 9367
rect 8202 9364 8208 9376
rect 7883 9336 8208 9364
rect 7883 9333 7895 9336
rect 7837 9327 7895 9333
rect 8202 9324 8208 9336
rect 8260 9324 8266 9376
rect 8386 9364 8392 9376
rect 8347 9336 8392 9364
rect 8386 9324 8392 9336
rect 8444 9324 8450 9376
rect 9398 9364 9404 9376
rect 9359 9336 9404 9364
rect 9398 9324 9404 9336
rect 9456 9324 9462 9376
rect 9493 9367 9551 9373
rect 9493 9333 9505 9367
rect 9539 9364 9551 9367
rect 9692 9364 9720 9472
rect 10965 9469 10977 9472
rect 11011 9469 11023 9503
rect 10965 9463 11023 9469
rect 12986 9460 12992 9512
rect 13044 9500 13050 9512
rect 13081 9503 13139 9509
rect 13081 9500 13093 9503
rect 13044 9472 13093 9500
rect 13044 9460 13050 9472
rect 13081 9469 13093 9472
rect 13127 9469 13139 9503
rect 13081 9463 13139 9469
rect 13348 9503 13406 9509
rect 13348 9469 13360 9503
rect 13394 9500 13406 9503
rect 14734 9500 14740 9512
rect 13394 9472 14740 9500
rect 13394 9469 13406 9472
rect 13348 9463 13406 9469
rect 9766 9392 9772 9444
rect 9824 9432 9830 9444
rect 9861 9435 9919 9441
rect 9861 9432 9873 9435
rect 9824 9404 9873 9432
rect 9824 9392 9830 9404
rect 9861 9401 9873 9404
rect 9907 9432 9919 9435
rect 10318 9432 10324 9444
rect 9907 9404 10324 9432
rect 9907 9401 9919 9404
rect 9861 9395 9919 9401
rect 10318 9392 10324 9404
rect 10376 9392 10382 9444
rect 10520 9404 11468 9432
rect 9539 9336 9720 9364
rect 9539 9333 9551 9336
rect 9493 9327 9551 9333
rect 9950 9324 9956 9376
rect 10008 9364 10014 9376
rect 10520 9373 10548 9404
rect 10505 9367 10563 9373
rect 10008 9336 10053 9364
rect 10008 9324 10014 9336
rect 10505 9333 10517 9367
rect 10551 9333 10563 9367
rect 10505 9327 10563 9333
rect 10778 9324 10784 9376
rect 10836 9364 10842 9376
rect 10873 9367 10931 9373
rect 10873 9364 10885 9367
rect 10836 9336 10885 9364
rect 10836 9324 10842 9336
rect 10873 9333 10885 9336
rect 10919 9333 10931 9367
rect 11440 9364 11468 9404
rect 11790 9392 11796 9444
rect 11848 9432 11854 9444
rect 13096 9432 13124 9463
rect 14734 9460 14740 9472
rect 14792 9460 14798 9512
rect 14936 9509 14964 9540
rect 15197 9537 15209 9571
rect 15243 9568 15255 9571
rect 15654 9568 15660 9580
rect 15243 9540 15660 9568
rect 15243 9537 15255 9540
rect 15197 9531 15255 9537
rect 15654 9528 15660 9540
rect 15712 9528 15718 9580
rect 16206 9568 16212 9580
rect 16167 9540 16212 9568
rect 16206 9528 16212 9540
rect 16264 9528 16270 9580
rect 18322 9568 18328 9580
rect 16316 9540 18328 9568
rect 14921 9503 14979 9509
rect 14921 9469 14933 9503
rect 14967 9469 14979 9503
rect 16316 9500 16344 9540
rect 18322 9528 18328 9540
rect 18380 9528 18386 9580
rect 18598 9568 18604 9580
rect 18559 9540 18604 9568
rect 18598 9528 18604 9540
rect 18656 9528 18662 9580
rect 18708 9568 18736 9676
rect 19613 9571 19671 9577
rect 19613 9568 19625 9571
rect 18708 9540 19625 9568
rect 19613 9537 19625 9540
rect 19659 9537 19671 9571
rect 19613 9531 19671 9537
rect 17586 9500 17592 9512
rect 14921 9463 14979 9469
rect 15948 9472 16344 9500
rect 17547 9472 17592 9500
rect 13722 9432 13728 9444
rect 11848 9404 13032 9432
rect 13096 9404 13728 9432
rect 11848 9392 11854 9404
rect 12618 9364 12624 9376
rect 11440 9336 12624 9364
rect 10873 9327 10931 9333
rect 12618 9324 12624 9336
rect 12676 9324 12682 9376
rect 13004 9364 13032 9404
rect 13722 9392 13728 9404
rect 13780 9392 13786 9444
rect 15948 9432 15976 9472
rect 17586 9460 17592 9472
rect 17644 9460 17650 9512
rect 18138 9460 18144 9512
rect 18196 9500 18202 9512
rect 18417 9503 18475 9509
rect 18417 9500 18429 9503
rect 18196 9472 18429 9500
rect 18196 9460 18202 9472
rect 18417 9469 18429 9472
rect 18463 9469 18475 9503
rect 18417 9463 18475 9469
rect 19880 9503 19938 9509
rect 19880 9469 19892 9503
rect 19926 9500 19938 9503
rect 20714 9500 20720 9512
rect 19926 9472 20720 9500
rect 19926 9469 19938 9472
rect 19880 9463 19938 9469
rect 20714 9460 20720 9472
rect 20772 9460 20778 9512
rect 13832 9404 15976 9432
rect 16025 9435 16083 9441
rect 13832 9364 13860 9404
rect 16025 9401 16037 9435
rect 16071 9432 16083 9435
rect 17604 9432 17632 9460
rect 18509 9435 18567 9441
rect 18509 9432 18521 9435
rect 16071 9404 17172 9432
rect 17604 9404 18521 9432
rect 16071 9401 16083 9404
rect 16025 9395 16083 9401
rect 13004 9336 13860 9364
rect 14461 9367 14519 9373
rect 14461 9333 14473 9367
rect 14507 9364 14519 9367
rect 14550 9364 14556 9376
rect 14507 9336 14556 9364
rect 14507 9333 14519 9336
rect 14461 9327 14519 9333
rect 14550 9324 14556 9336
rect 14608 9324 14614 9376
rect 14737 9367 14795 9373
rect 14737 9333 14749 9367
rect 14783 9364 14795 9367
rect 15194 9364 15200 9376
rect 14783 9336 15200 9364
rect 14783 9333 14795 9336
rect 14737 9327 14795 9333
rect 15194 9324 15200 9336
rect 15252 9324 15258 9376
rect 15654 9364 15660 9376
rect 15615 9336 15660 9364
rect 15654 9324 15660 9336
rect 15712 9324 15718 9376
rect 16117 9367 16175 9373
rect 16117 9333 16129 9367
rect 16163 9364 16175 9367
rect 16850 9364 16856 9376
rect 16163 9336 16856 9364
rect 16163 9333 16175 9336
rect 16117 9327 16175 9333
rect 16850 9324 16856 9336
rect 16908 9324 16914 9376
rect 17144 9373 17172 9404
rect 18509 9401 18521 9404
rect 18555 9401 18567 9435
rect 18509 9395 18567 9401
rect 17129 9367 17187 9373
rect 17129 9333 17141 9367
rect 17175 9364 17187 9367
rect 18782 9364 18788 9376
rect 17175 9336 18788 9364
rect 17175 9333 17187 9336
rect 17129 9327 17187 9333
rect 18782 9324 18788 9336
rect 18840 9324 18846 9376
rect 19978 9324 19984 9376
rect 20036 9364 20042 9376
rect 20993 9367 21051 9373
rect 20993 9364 21005 9367
rect 20036 9336 21005 9364
rect 20036 9324 20042 9336
rect 20993 9333 21005 9336
rect 21039 9333 21051 9367
rect 20993 9327 21051 9333
rect 1104 9274 21896 9296
rect 1104 9222 7912 9274
rect 7964 9222 7976 9274
rect 8028 9222 8040 9274
rect 8092 9222 8104 9274
rect 8156 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 15035 9274
rect 15087 9222 21896 9274
rect 1104 9200 21896 9222
rect 2225 9163 2283 9169
rect 2225 9129 2237 9163
rect 2271 9160 2283 9163
rect 2682 9160 2688 9172
rect 2271 9132 2688 9160
rect 2271 9129 2283 9132
rect 2225 9123 2283 9129
rect 2682 9120 2688 9132
rect 2740 9120 2746 9172
rect 3605 9163 3663 9169
rect 3605 9129 3617 9163
rect 3651 9160 3663 9163
rect 4982 9160 4988 9172
rect 3651 9132 4988 9160
rect 3651 9129 3663 9132
rect 3605 9123 3663 9129
rect 4982 9120 4988 9132
rect 5040 9120 5046 9172
rect 5445 9163 5503 9169
rect 5445 9129 5457 9163
rect 5491 9129 5503 9163
rect 5445 9123 5503 9129
rect 7101 9163 7159 9169
rect 7101 9129 7113 9163
rect 7147 9160 7159 9163
rect 7190 9160 7196 9172
rect 7147 9132 7196 9160
rect 7147 9129 7159 9132
rect 7101 9123 7159 9129
rect 2498 9052 2504 9104
rect 2556 9092 2562 9104
rect 2556 9064 3372 9092
rect 2556 9052 2562 9064
rect 2590 9024 2596 9036
rect 2551 8996 2596 9024
rect 2590 8984 2596 8996
rect 2648 8984 2654 9036
rect 2682 8956 2688 8968
rect 2643 8928 2688 8956
rect 2682 8916 2688 8928
rect 2740 8916 2746 8968
rect 2866 8956 2872 8968
rect 2827 8928 2872 8956
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 3344 8956 3372 9064
rect 3418 9052 3424 9104
rect 3476 9092 3482 9104
rect 4310 9095 4368 9101
rect 4310 9092 4322 9095
rect 3476 9064 4322 9092
rect 3476 9052 3482 9064
rect 4310 9061 4322 9064
rect 4356 9061 4368 9095
rect 5460 9092 5488 9123
rect 7190 9120 7196 9132
rect 7248 9120 7254 9172
rect 7374 9160 7380 9172
rect 7335 9132 7380 9160
rect 7374 9120 7380 9132
rect 7432 9120 7438 9172
rect 7742 9120 7748 9172
rect 7800 9160 7806 9172
rect 8757 9163 8815 9169
rect 8757 9160 8769 9163
rect 7800 9132 8769 9160
rect 7800 9120 7806 9132
rect 8757 9129 8769 9132
rect 8803 9129 8815 9163
rect 8757 9123 8815 9129
rect 8846 9120 8852 9172
rect 8904 9160 8910 9172
rect 9306 9160 9312 9172
rect 8904 9132 9312 9160
rect 8904 9120 8910 9132
rect 9306 9120 9312 9132
rect 9364 9120 9370 9172
rect 9677 9163 9735 9169
rect 9677 9129 9689 9163
rect 9723 9160 9735 9163
rect 9950 9160 9956 9172
rect 9723 9132 9956 9160
rect 9723 9129 9735 9132
rect 9677 9123 9735 9129
rect 9950 9120 9956 9132
rect 10008 9120 10014 9172
rect 10137 9163 10195 9169
rect 10137 9129 10149 9163
rect 10183 9160 10195 9163
rect 10318 9160 10324 9172
rect 10183 9132 10324 9160
rect 10183 9129 10195 9132
rect 10137 9123 10195 9129
rect 10318 9120 10324 9132
rect 10376 9160 10382 9172
rect 11609 9163 11667 9169
rect 10376 9132 11560 9160
rect 10376 9120 10382 9132
rect 5966 9095 6024 9101
rect 5966 9092 5978 9095
rect 5460 9064 5978 9092
rect 4310 9055 4368 9061
rect 5966 9061 5978 9064
rect 6012 9092 6024 9095
rect 7466 9092 7472 9104
rect 6012 9064 7472 9092
rect 6012 9061 6024 9064
rect 5966 9055 6024 9061
rect 7466 9052 7472 9064
rect 7524 9092 7530 9104
rect 11532 9092 11560 9132
rect 11609 9129 11621 9163
rect 11655 9160 11667 9163
rect 14553 9163 14611 9169
rect 14553 9160 14565 9163
rect 11655 9132 14565 9160
rect 11655 9129 11667 9132
rect 11609 9123 11667 9129
rect 14553 9129 14565 9132
rect 14599 9129 14611 9163
rect 14553 9123 14611 9129
rect 14645 9163 14703 9169
rect 14645 9129 14657 9163
rect 14691 9160 14703 9163
rect 15654 9160 15660 9172
rect 14691 9132 15660 9160
rect 14691 9129 14703 9132
rect 14645 9123 14703 9129
rect 15654 9120 15660 9132
rect 15712 9120 15718 9172
rect 20257 9163 20315 9169
rect 20257 9129 20269 9163
rect 20303 9160 20315 9163
rect 20530 9160 20536 9172
rect 20303 9132 20536 9160
rect 20303 9129 20315 9132
rect 20257 9123 20315 9129
rect 20530 9120 20536 9132
rect 20588 9120 20594 9172
rect 20898 9160 20904 9172
rect 20859 9132 20904 9160
rect 20898 9120 20904 9132
rect 20956 9120 20962 9172
rect 12253 9095 12311 9101
rect 12253 9092 12265 9095
rect 7524 9064 7972 9092
rect 7524 9052 7530 9064
rect 4154 8984 4160 9036
rect 4212 8984 4218 9036
rect 6546 8984 6552 9036
rect 6604 9024 6610 9036
rect 7282 9024 7288 9036
rect 6604 8996 7288 9024
rect 6604 8984 6610 8996
rect 7282 8984 7288 8996
rect 7340 9024 7346 9036
rect 7745 9027 7803 9033
rect 7745 9024 7757 9027
rect 7340 8996 7757 9024
rect 7340 8984 7346 8996
rect 7745 8993 7757 8996
rect 7791 8993 7803 9027
rect 7745 8987 7803 8993
rect 4065 8959 4123 8965
rect 4065 8956 4077 8959
rect 3344 8928 4077 8956
rect 4065 8925 4077 8928
rect 4111 8956 4123 8959
rect 4172 8956 4200 8984
rect 4111 8928 4200 8956
rect 4111 8925 4123 8928
rect 4065 8919 4123 8925
rect 5442 8916 5448 8968
rect 5500 8956 5506 8968
rect 5721 8959 5779 8965
rect 5721 8956 5733 8959
rect 5500 8928 5733 8956
rect 5500 8916 5506 8928
rect 5721 8925 5733 8928
rect 5767 8925 5779 8959
rect 5721 8919 5779 8925
rect 6914 8916 6920 8968
rect 6972 8956 6978 8968
rect 7374 8956 7380 8968
rect 6972 8928 7380 8956
rect 6972 8916 6978 8928
rect 7374 8916 7380 8928
rect 7432 8956 7438 8968
rect 7944 8965 7972 9064
rect 9048 9064 10824 9092
rect 7837 8959 7895 8965
rect 7837 8956 7849 8959
rect 7432 8928 7849 8956
rect 7432 8916 7438 8928
rect 7837 8925 7849 8928
rect 7883 8925 7895 8959
rect 7837 8919 7895 8925
rect 7929 8959 7987 8965
rect 7929 8925 7941 8959
rect 7975 8925 7987 8959
rect 8386 8956 8392 8968
rect 7929 8919 7987 8925
rect 8312 8928 8392 8956
rect 7852 8888 7880 8919
rect 8312 8888 8340 8928
rect 8386 8916 8392 8928
rect 8444 8916 8450 8968
rect 8662 8916 8668 8968
rect 8720 8956 8726 8968
rect 9048 8965 9076 9064
rect 9490 8984 9496 9036
rect 9548 9024 9554 9036
rect 9858 9024 9864 9036
rect 9548 8996 9864 9024
rect 9548 8984 9554 8996
rect 9858 8984 9864 8996
rect 9916 8984 9922 9036
rect 10042 9024 10048 9036
rect 10003 8996 10048 9024
rect 10042 8984 10048 8996
rect 10100 8984 10106 9036
rect 10318 9024 10324 9036
rect 10152 8996 10324 9024
rect 8849 8959 8907 8965
rect 8849 8956 8861 8959
rect 8720 8928 8861 8956
rect 8720 8916 8726 8928
rect 8849 8925 8861 8928
rect 8895 8925 8907 8959
rect 8849 8919 8907 8925
rect 9033 8959 9091 8965
rect 9033 8925 9045 8959
rect 9079 8925 9091 8959
rect 10152 8956 10180 8996
rect 10318 8984 10324 8996
rect 10376 8984 10382 9036
rect 10796 9024 10824 9064
rect 10971 9064 11376 9092
rect 11532 9064 12265 9092
rect 10971 9024 10999 9064
rect 11146 9024 11152 9036
rect 10796 8996 10999 9024
rect 11107 8996 11152 9024
rect 11146 8984 11152 8996
rect 11204 8984 11210 9036
rect 9033 8919 9091 8925
rect 9232 8928 10180 8956
rect 10229 8959 10287 8965
rect 7852 8860 8340 8888
rect 8754 8848 8760 8900
rect 8812 8888 8818 8900
rect 9232 8888 9260 8928
rect 10229 8925 10241 8959
rect 10275 8925 10287 8959
rect 10229 8919 10287 8925
rect 8812 8860 9260 8888
rect 8812 8848 8818 8860
rect 9306 8848 9312 8900
rect 9364 8888 9370 8900
rect 10244 8888 10272 8919
rect 10962 8916 10968 8968
rect 11020 8956 11026 8968
rect 11348 8965 11376 9064
rect 12253 9061 12265 9064
rect 12299 9092 12311 9095
rect 19150 9092 19156 9104
rect 12299 9064 19156 9092
rect 12299 9061 12311 9064
rect 12253 9055 12311 9061
rect 19150 9052 19156 9064
rect 19208 9052 19214 9104
rect 20070 9052 20076 9104
rect 20128 9092 20134 9104
rect 21174 9092 21180 9104
rect 20128 9064 21180 9092
rect 20128 9052 20134 9064
rect 21174 9052 21180 9064
rect 21232 9052 21238 9104
rect 11422 8984 11428 9036
rect 11480 9024 11486 9036
rect 11790 9024 11796 9036
rect 11480 8996 11796 9024
rect 11480 8984 11486 8996
rect 11790 8984 11796 8996
rect 11848 8984 11854 9036
rect 13909 9027 13967 9033
rect 13909 8993 13921 9027
rect 13955 9024 13967 9027
rect 15194 9024 15200 9036
rect 13955 8996 15200 9024
rect 13955 8993 13967 8996
rect 13909 8987 13967 8993
rect 15194 8984 15200 8996
rect 15252 9024 15258 9036
rect 15933 9027 15991 9033
rect 15933 9024 15945 9027
rect 15252 8996 15945 9024
rect 15252 8984 15258 8996
rect 15933 8993 15945 8996
rect 15979 8993 15991 9027
rect 20165 9027 20223 9033
rect 20165 9024 20177 9027
rect 15933 8987 15991 8993
rect 19444 8996 20177 9024
rect 11241 8959 11299 8965
rect 11241 8956 11253 8959
rect 11020 8928 11253 8956
rect 11020 8916 11026 8928
rect 11241 8925 11253 8928
rect 11287 8925 11299 8959
rect 11241 8919 11299 8925
rect 11333 8959 11391 8965
rect 11333 8925 11345 8959
rect 11379 8956 11391 8959
rect 13078 8956 13084 8968
rect 11379 8928 13084 8956
rect 11379 8925 11391 8928
rect 11333 8919 11391 8925
rect 13078 8916 13084 8928
rect 13136 8916 13142 8968
rect 14734 8956 14740 8968
rect 14695 8928 14740 8956
rect 14734 8916 14740 8928
rect 14792 8916 14798 8968
rect 9364 8860 10272 8888
rect 10781 8891 10839 8897
rect 9364 8848 9370 8860
rect 10781 8857 10793 8891
rect 10827 8888 10839 8891
rect 13814 8888 13820 8900
rect 10827 8860 13820 8888
rect 10827 8857 10839 8860
rect 10781 8851 10839 8857
rect 13814 8848 13820 8860
rect 13872 8848 13878 8900
rect 16390 8848 16396 8900
rect 16448 8888 16454 8900
rect 19058 8888 19064 8900
rect 16448 8860 19064 8888
rect 16448 8848 16454 8860
rect 19058 8848 19064 8860
rect 19116 8848 19122 8900
rect 8389 8823 8447 8829
rect 8389 8789 8401 8823
rect 8435 8820 8447 8823
rect 11609 8823 11667 8829
rect 11609 8820 11621 8823
rect 8435 8792 11621 8820
rect 8435 8789 8447 8792
rect 8389 8783 8447 8789
rect 11609 8789 11621 8792
rect 11655 8789 11667 8823
rect 11609 8783 11667 8789
rect 12621 8823 12679 8829
rect 12621 8789 12633 8823
rect 12667 8820 12679 8823
rect 13078 8820 13084 8832
rect 12667 8792 13084 8820
rect 12667 8789 12679 8792
rect 12621 8783 12679 8789
rect 13078 8780 13084 8792
rect 13136 8780 13142 8832
rect 13722 8820 13728 8832
rect 13683 8792 13728 8820
rect 13722 8780 13728 8792
rect 13780 8780 13786 8832
rect 14185 8823 14243 8829
rect 14185 8789 14197 8823
rect 14231 8820 14243 8823
rect 14458 8820 14464 8832
rect 14231 8792 14464 8820
rect 14231 8789 14243 8792
rect 14185 8783 14243 8789
rect 14458 8780 14464 8792
rect 14516 8780 14522 8832
rect 15749 8823 15807 8829
rect 15749 8789 15761 8823
rect 15795 8820 15807 8823
rect 16574 8820 16580 8832
rect 15795 8792 16580 8820
rect 15795 8789 15807 8792
rect 15749 8783 15807 8789
rect 16574 8780 16580 8792
rect 16632 8780 16638 8832
rect 16666 8780 16672 8832
rect 16724 8820 16730 8832
rect 19444 8829 19472 8996
rect 20165 8993 20177 8996
rect 20211 8993 20223 9027
rect 20165 8987 20223 8993
rect 20441 8959 20499 8965
rect 20441 8925 20453 8959
rect 20487 8956 20499 8959
rect 20714 8956 20720 8968
rect 20487 8928 20720 8956
rect 20487 8925 20499 8928
rect 20441 8919 20499 8925
rect 20714 8916 20720 8928
rect 20772 8916 20778 8968
rect 19429 8823 19487 8829
rect 19429 8820 19441 8823
rect 16724 8792 19441 8820
rect 16724 8780 16730 8792
rect 19429 8789 19441 8792
rect 19475 8789 19487 8823
rect 19794 8820 19800 8832
rect 19755 8792 19800 8820
rect 19429 8783 19487 8789
rect 19794 8780 19800 8792
rect 19852 8780 19858 8832
rect 1104 8730 21896 8752
rect 1104 8678 4447 8730
rect 4499 8678 4511 8730
rect 4563 8678 4575 8730
rect 4627 8678 4639 8730
rect 4691 8678 11378 8730
rect 11430 8678 11442 8730
rect 11494 8678 11506 8730
rect 11558 8678 11570 8730
rect 11622 8678 18308 8730
rect 18360 8678 18372 8730
rect 18424 8678 18436 8730
rect 18488 8678 18500 8730
rect 18552 8678 21896 8730
rect 1104 8656 21896 8678
rect 2866 8576 2872 8628
rect 2924 8616 2930 8628
rect 3237 8619 3295 8625
rect 3237 8616 3249 8619
rect 2924 8588 3249 8616
rect 2924 8576 2930 8588
rect 3237 8585 3249 8588
rect 3283 8616 3295 8619
rect 3283 8588 4660 8616
rect 3283 8585 3295 8588
rect 3237 8579 3295 8585
rect 4632 8560 4660 8588
rect 4890 8576 4896 8628
rect 4948 8616 4954 8628
rect 5442 8616 5448 8628
rect 4948 8588 5448 8616
rect 4948 8576 4954 8588
rect 5442 8576 5448 8588
rect 5500 8616 5506 8628
rect 5721 8619 5779 8625
rect 5721 8616 5733 8619
rect 5500 8588 5733 8616
rect 5500 8576 5506 8588
rect 5721 8585 5733 8588
rect 5767 8585 5779 8619
rect 6822 8616 6828 8628
rect 6783 8588 6828 8616
rect 5721 8579 5779 8585
rect 6822 8576 6828 8588
rect 6880 8576 6886 8628
rect 7282 8576 7288 8628
rect 7340 8616 7346 8628
rect 8205 8619 8263 8625
rect 8205 8616 8217 8619
rect 7340 8588 8217 8616
rect 7340 8576 7346 8588
rect 8205 8585 8217 8588
rect 8251 8616 8263 8619
rect 9766 8616 9772 8628
rect 8251 8588 9772 8616
rect 8251 8585 8263 8588
rect 8205 8579 8263 8585
rect 9766 8576 9772 8588
rect 9824 8576 9830 8628
rect 10134 8616 10140 8628
rect 10095 8588 10140 8616
rect 10134 8576 10140 8588
rect 10192 8576 10198 8628
rect 10594 8616 10600 8628
rect 10555 8588 10600 8616
rect 10594 8576 10600 8588
rect 10652 8576 10658 8628
rect 11698 8576 11704 8628
rect 11756 8616 11762 8628
rect 16666 8616 16672 8628
rect 11756 8588 16672 8616
rect 11756 8576 11762 8588
rect 16666 8576 16672 8588
rect 16724 8576 16730 8628
rect 16758 8576 16764 8628
rect 16816 8616 16822 8628
rect 16853 8619 16911 8625
rect 16853 8616 16865 8619
rect 16816 8588 16865 8616
rect 16816 8576 16822 8588
rect 16853 8585 16865 8588
rect 16899 8585 16911 8619
rect 16853 8579 16911 8585
rect 17494 8576 17500 8628
rect 17552 8616 17558 8628
rect 17589 8619 17647 8625
rect 17589 8616 17601 8619
rect 17552 8588 17601 8616
rect 17552 8576 17558 8588
rect 17589 8585 17601 8588
rect 17635 8585 17647 8619
rect 17589 8579 17647 8585
rect 3881 8551 3939 8557
rect 3881 8517 3893 8551
rect 3927 8548 3939 8551
rect 4338 8548 4344 8560
rect 3927 8520 4344 8548
rect 3927 8517 3939 8520
rect 3881 8511 3939 8517
rect 4338 8508 4344 8520
rect 4396 8508 4402 8560
rect 4614 8508 4620 8560
rect 4672 8508 4678 8560
rect 7837 8551 7895 8557
rect 7837 8548 7849 8551
rect 7300 8520 7849 8548
rect 4525 8483 4583 8489
rect 4525 8449 4537 8483
rect 4571 8480 4583 8483
rect 5534 8480 5540 8492
rect 4571 8452 5540 8480
rect 4571 8449 4583 8452
rect 4525 8443 4583 8449
rect 5534 8440 5540 8452
rect 5592 8440 5598 8492
rect 6178 8440 6184 8492
rect 6236 8480 6242 8492
rect 7300 8489 7328 8520
rect 7837 8517 7849 8520
rect 7883 8548 7895 8551
rect 8662 8548 8668 8560
rect 7883 8520 8668 8548
rect 7883 8517 7895 8520
rect 7837 8511 7895 8517
rect 8662 8508 8668 8520
rect 8720 8508 8726 8560
rect 10965 8551 11023 8557
rect 10965 8517 10977 8551
rect 11011 8548 11023 8551
rect 11422 8548 11428 8560
rect 11011 8520 11428 8548
rect 11011 8517 11023 8520
rect 10965 8511 11023 8517
rect 11422 8508 11428 8520
rect 11480 8508 11486 8560
rect 16482 8508 16488 8560
rect 16540 8548 16546 8560
rect 17129 8551 17187 8557
rect 17129 8548 17141 8551
rect 16540 8520 17141 8548
rect 16540 8508 16546 8520
rect 17129 8517 17141 8520
rect 17175 8517 17187 8551
rect 17129 8511 17187 8517
rect 6365 8483 6423 8489
rect 6365 8480 6377 8483
rect 6236 8452 6377 8480
rect 6236 8440 6242 8452
rect 6365 8449 6377 8452
rect 6411 8480 6423 8483
rect 7285 8483 7343 8489
rect 7285 8480 7297 8483
rect 6411 8452 7297 8480
rect 6411 8449 6423 8452
rect 6365 8443 6423 8449
rect 7285 8449 7297 8452
rect 7331 8449 7343 8483
rect 7466 8480 7472 8492
rect 7427 8452 7472 8480
rect 7285 8443 7343 8449
rect 7466 8440 7472 8452
rect 7524 8440 7530 8492
rect 8294 8440 8300 8492
rect 8352 8480 8358 8492
rect 8757 8483 8815 8489
rect 8757 8480 8769 8483
rect 8352 8452 8769 8480
rect 8352 8440 8358 8452
rect 8757 8449 8769 8452
rect 8803 8449 8815 8483
rect 8757 8443 8815 8449
rect 11238 8440 11244 8492
rect 11296 8480 11302 8492
rect 11517 8483 11575 8489
rect 11517 8480 11529 8483
rect 11296 8452 11529 8480
rect 11296 8440 11302 8452
rect 11517 8449 11529 8452
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 12710 8440 12716 8492
rect 12768 8480 12774 8492
rect 12986 8480 12992 8492
rect 12768 8452 12992 8480
rect 12768 8440 12774 8452
rect 12986 8440 12992 8452
rect 13044 8480 13050 8492
rect 13265 8483 13323 8489
rect 13265 8480 13277 8483
rect 13044 8452 13277 8480
rect 13044 8440 13050 8452
rect 13265 8449 13277 8452
rect 13311 8449 13323 8483
rect 13265 8443 13323 8449
rect 14458 8440 14464 8492
rect 14516 8480 14522 8492
rect 14645 8483 14703 8489
rect 14516 8452 14561 8480
rect 14516 8440 14522 8452
rect 14645 8449 14657 8483
rect 14691 8480 14703 8483
rect 14826 8480 14832 8492
rect 14691 8452 14832 8480
rect 14691 8449 14703 8452
rect 14645 8443 14703 8449
rect 14826 8440 14832 8452
rect 14884 8440 14890 8492
rect 1857 8415 1915 8421
rect 1857 8381 1869 8415
rect 1903 8412 1915 8415
rect 2498 8412 2504 8424
rect 1903 8384 2504 8412
rect 1903 8381 1915 8384
rect 1857 8375 1915 8381
rect 2498 8372 2504 8384
rect 2556 8372 2562 8424
rect 4341 8415 4399 8421
rect 4341 8381 4353 8415
rect 4387 8412 4399 8415
rect 4982 8412 4988 8424
rect 4387 8384 4988 8412
rect 4387 8381 4399 8384
rect 4341 8375 4399 8381
rect 4982 8372 4988 8384
rect 5040 8372 5046 8424
rect 5905 8415 5963 8421
rect 5905 8381 5917 8415
rect 5951 8412 5963 8415
rect 8202 8412 8208 8424
rect 5951 8384 8208 8412
rect 5951 8381 5963 8384
rect 5905 8375 5963 8381
rect 8202 8372 8208 8384
rect 8260 8372 8266 8424
rect 9024 8415 9082 8421
rect 9024 8381 9036 8415
rect 9070 8412 9082 8415
rect 9306 8412 9312 8424
rect 9070 8384 9312 8412
rect 9070 8381 9082 8384
rect 9024 8375 9082 8381
rect 9306 8372 9312 8384
rect 9364 8372 9370 8424
rect 10594 8372 10600 8424
rect 10652 8412 10658 8424
rect 11425 8415 11483 8421
rect 11425 8412 11437 8415
rect 10652 8384 11437 8412
rect 10652 8372 10658 8384
rect 11425 8381 11437 8384
rect 11471 8381 11483 8415
rect 13170 8412 13176 8424
rect 13131 8384 13176 8412
rect 11425 8375 11483 8381
rect 13170 8372 13176 8384
rect 13228 8372 13234 8424
rect 13998 8372 14004 8424
rect 14056 8412 14062 8424
rect 14369 8415 14427 8421
rect 14369 8412 14381 8415
rect 14056 8384 14381 8412
rect 14056 8372 14062 8384
rect 14369 8381 14381 8384
rect 14415 8381 14427 8415
rect 14369 8375 14427 8381
rect 15473 8415 15531 8421
rect 15473 8381 15485 8415
rect 15519 8381 15531 8415
rect 17604 8412 17632 8579
rect 19337 8551 19395 8557
rect 19337 8517 19349 8551
rect 19383 8548 19395 8551
rect 19518 8548 19524 8560
rect 19383 8520 19524 8548
rect 19383 8517 19395 8520
rect 19337 8511 19395 8517
rect 19518 8508 19524 8520
rect 19576 8508 19582 8560
rect 18138 8440 18144 8492
rect 18196 8480 18202 8492
rect 18601 8483 18659 8489
rect 18601 8480 18613 8483
rect 18196 8452 18613 8480
rect 18196 8440 18202 8452
rect 18601 8449 18613 8452
rect 18647 8449 18659 8483
rect 19794 8480 19800 8492
rect 19755 8452 19800 8480
rect 18601 8443 18659 8449
rect 19794 8440 19800 8452
rect 19852 8440 19858 8492
rect 19978 8480 19984 8492
rect 19939 8452 19984 8480
rect 19978 8440 19984 8452
rect 20036 8440 20042 8492
rect 18509 8415 18567 8421
rect 18509 8412 18521 8415
rect 17604 8384 18521 8412
rect 15473 8375 15531 8381
rect 18509 8381 18521 8384
rect 18555 8381 18567 8415
rect 19702 8412 19708 8424
rect 19663 8384 19708 8412
rect 18509 8375 18567 8381
rect 2124 8347 2182 8353
rect 2124 8313 2136 8347
rect 2170 8344 2182 8347
rect 3050 8344 3056 8356
rect 2170 8316 3056 8344
rect 2170 8313 2182 8316
rect 2124 8307 2182 8313
rect 3050 8304 3056 8316
rect 3108 8304 3114 8356
rect 5074 8304 5080 8356
rect 5132 8344 5138 8356
rect 12526 8344 12532 8356
rect 5132 8316 12532 8344
rect 5132 8304 5138 8316
rect 12526 8304 12532 8316
rect 12584 8304 12590 8356
rect 13078 8344 13084 8356
rect 13039 8316 13084 8344
rect 13078 8304 13084 8316
rect 13136 8304 13142 8356
rect 13722 8304 13728 8356
rect 13780 8344 13786 8356
rect 15488 8344 15516 8375
rect 19702 8372 19708 8384
rect 19760 8372 19766 8424
rect 13780 8316 15516 8344
rect 15740 8347 15798 8353
rect 13780 8304 13786 8316
rect 15740 8313 15752 8347
rect 15786 8344 15798 8347
rect 16206 8344 16212 8356
rect 15786 8316 16212 8344
rect 15786 8313 15798 8316
rect 15740 8307 15798 8313
rect 16206 8304 16212 8316
rect 16264 8304 16270 8356
rect 16666 8304 16672 8356
rect 16724 8344 16730 8356
rect 19610 8344 19616 8356
rect 16724 8316 19616 8344
rect 16724 8304 16730 8316
rect 19610 8304 19616 8316
rect 19668 8304 19674 8356
rect 2314 8236 2320 8288
rect 2372 8276 2378 8288
rect 3513 8279 3571 8285
rect 3513 8276 3525 8279
rect 2372 8248 3525 8276
rect 2372 8236 2378 8248
rect 3513 8245 3525 8248
rect 3559 8276 3571 8279
rect 3602 8276 3608 8288
rect 3559 8248 3608 8276
rect 3559 8245 3571 8248
rect 3513 8239 3571 8245
rect 3602 8236 3608 8248
rect 3660 8276 3666 8288
rect 4249 8279 4307 8285
rect 4249 8276 4261 8279
rect 3660 8248 4261 8276
rect 3660 8236 3666 8248
rect 4249 8245 4261 8248
rect 4295 8245 4307 8279
rect 4249 8239 4307 8245
rect 6914 8236 6920 8288
rect 6972 8276 6978 8288
rect 7193 8279 7251 8285
rect 7193 8276 7205 8279
rect 6972 8248 7205 8276
rect 6972 8236 6978 8248
rect 7193 8245 7205 8248
rect 7239 8245 7251 8279
rect 11330 8276 11336 8288
rect 11291 8248 11336 8276
rect 7193 8239 7251 8245
rect 11330 8236 11336 8248
rect 11388 8236 11394 8288
rect 11422 8236 11428 8288
rect 11480 8276 11486 8288
rect 12250 8276 12256 8288
rect 11480 8248 12256 8276
rect 11480 8236 11486 8248
rect 12250 8236 12256 8248
rect 12308 8236 12314 8288
rect 12710 8276 12716 8288
rect 12671 8248 12716 8276
rect 12710 8236 12716 8248
rect 12768 8236 12774 8288
rect 14001 8279 14059 8285
rect 14001 8245 14013 8279
rect 14047 8276 14059 8279
rect 14182 8276 14188 8288
rect 14047 8248 14188 8276
rect 14047 8245 14059 8248
rect 14001 8239 14059 8245
rect 14182 8236 14188 8248
rect 14240 8236 14246 8288
rect 14642 8236 14648 8288
rect 14700 8276 14706 8288
rect 17770 8276 17776 8288
rect 14700 8248 17776 8276
rect 14700 8236 14706 8248
rect 17770 8236 17776 8248
rect 17828 8236 17834 8288
rect 18046 8276 18052 8288
rect 18007 8248 18052 8276
rect 18046 8236 18052 8248
rect 18104 8236 18110 8288
rect 18414 8276 18420 8288
rect 18375 8248 18420 8276
rect 18414 8236 18420 8248
rect 18472 8236 18478 8288
rect 1104 8186 21896 8208
rect 1104 8134 7912 8186
rect 7964 8134 7976 8186
rect 8028 8134 8040 8186
rect 8092 8134 8104 8186
rect 8156 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 15035 8186
rect 15087 8134 21896 8186
rect 1104 8112 21896 8134
rect 1578 8032 1584 8084
rect 1636 8072 1642 8084
rect 1673 8075 1731 8081
rect 1673 8072 1685 8075
rect 1636 8044 1685 8072
rect 1636 8032 1642 8044
rect 1673 8041 1685 8044
rect 1719 8041 1731 8075
rect 1673 8035 1731 8041
rect 2409 8075 2467 8081
rect 2409 8041 2421 8075
rect 2455 8072 2467 8075
rect 2682 8072 2688 8084
rect 2455 8044 2688 8072
rect 2455 8041 2467 8044
rect 2409 8035 2467 8041
rect 1688 7948 1716 8035
rect 2682 8032 2688 8044
rect 2740 8032 2746 8084
rect 2774 8032 2780 8084
rect 2832 8072 2838 8084
rect 4065 8075 4123 8081
rect 4065 8072 4077 8075
rect 2832 8044 4077 8072
rect 2832 8032 2838 8044
rect 4065 8041 4077 8044
rect 4111 8041 4123 8075
rect 4065 8035 4123 8041
rect 4338 8032 4344 8084
rect 4396 8072 4402 8084
rect 4433 8075 4491 8081
rect 4433 8072 4445 8075
rect 4396 8044 4445 8072
rect 4396 8032 4402 8044
rect 4433 8041 4445 8044
rect 4479 8041 4491 8075
rect 4433 8035 4491 8041
rect 8021 8075 8079 8081
rect 8021 8041 8033 8075
rect 8067 8072 8079 8075
rect 8294 8072 8300 8084
rect 8067 8044 8300 8072
rect 8067 8041 8079 8044
rect 8021 8035 8079 8041
rect 8294 8032 8300 8044
rect 8352 8032 8358 8084
rect 11241 8075 11299 8081
rect 11241 8041 11253 8075
rect 11287 8072 11299 8075
rect 11330 8072 11336 8084
rect 11287 8044 11336 8072
rect 11287 8041 11299 8044
rect 11241 8035 11299 8041
rect 11330 8032 11336 8044
rect 11388 8032 11394 8084
rect 12161 8075 12219 8081
rect 12161 8041 12173 8075
rect 12207 8072 12219 8075
rect 12710 8072 12716 8084
rect 12207 8044 12716 8072
rect 12207 8041 12219 8044
rect 12161 8035 12219 8041
rect 12710 8032 12716 8044
rect 12768 8032 12774 8084
rect 13170 8032 13176 8084
rect 13228 8072 13234 8084
rect 14461 8075 14519 8081
rect 14461 8072 14473 8075
rect 13228 8044 14473 8072
rect 13228 8032 13234 8044
rect 14461 8041 14473 8044
rect 14507 8072 14519 8075
rect 14642 8072 14648 8084
rect 14507 8044 14648 8072
rect 14507 8041 14519 8044
rect 14461 8035 14519 8041
rect 14642 8032 14648 8044
rect 14700 8032 14706 8084
rect 16025 8075 16083 8081
rect 16025 8041 16037 8075
rect 16071 8072 16083 8075
rect 16482 8072 16488 8084
rect 16071 8044 16488 8072
rect 16071 8041 16083 8044
rect 16025 8035 16083 8041
rect 16482 8032 16488 8044
rect 16540 8032 16546 8084
rect 16574 8032 16580 8084
rect 16632 8072 16638 8084
rect 17862 8072 17868 8084
rect 16632 8044 17868 8072
rect 16632 8032 16638 8044
rect 17862 8032 17868 8044
rect 17920 8032 17926 8084
rect 17957 8075 18015 8081
rect 17957 8041 17969 8075
rect 18003 8072 18015 8075
rect 18138 8072 18144 8084
rect 18003 8044 18144 8072
rect 18003 8041 18015 8044
rect 17957 8035 18015 8041
rect 4525 8007 4583 8013
rect 4525 7973 4537 8007
rect 4571 8004 4583 8007
rect 9858 8004 9864 8016
rect 4571 7976 9864 8004
rect 4571 7973 4583 7976
rect 4525 7967 4583 7973
rect 9858 7964 9864 7976
rect 9916 7964 9922 8016
rect 12986 8013 12992 8016
rect 12980 8004 12992 8013
rect 12947 7976 12992 8004
rect 12980 7967 12992 7976
rect 12986 7964 12992 7967
rect 13044 7964 13050 8016
rect 17972 8004 18000 8035
rect 18138 8032 18144 8044
rect 18196 8032 18202 8084
rect 18233 8075 18291 8081
rect 18233 8041 18245 8075
rect 18279 8072 18291 8075
rect 18414 8072 18420 8084
rect 18279 8044 18420 8072
rect 18279 8041 18291 8044
rect 18233 8035 18291 8041
rect 18414 8032 18420 8044
rect 18472 8032 18478 8084
rect 16500 7976 18000 8004
rect 19052 8007 19110 8013
rect 1670 7936 1676 7948
rect 1583 7908 1676 7936
rect 1670 7896 1676 7908
rect 1728 7936 1734 7948
rect 2777 7939 2835 7945
rect 2777 7936 2789 7939
rect 1728 7908 2789 7936
rect 1728 7896 1734 7908
rect 2777 7905 2789 7908
rect 2823 7905 2835 7939
rect 2777 7899 2835 7905
rect 4246 7896 4252 7948
rect 4304 7936 4310 7948
rect 5445 7939 5503 7945
rect 5445 7936 5457 7939
rect 4304 7908 5457 7936
rect 4304 7896 4310 7908
rect 5445 7905 5457 7908
rect 5491 7905 5503 7939
rect 8202 7936 8208 7948
rect 8163 7908 8208 7936
rect 5445 7899 5503 7905
rect 8202 7896 8208 7908
rect 8260 7896 8266 7948
rect 12069 7939 12127 7945
rect 12069 7936 12081 7939
rect 11164 7908 12081 7936
rect 11164 7880 11192 7908
rect 12069 7905 12081 7908
rect 12115 7905 12127 7939
rect 12069 7899 12127 7905
rect 12713 7939 12771 7945
rect 12713 7905 12725 7939
rect 12759 7936 12771 7939
rect 12802 7936 12808 7948
rect 12759 7908 12808 7936
rect 12759 7905 12771 7908
rect 12713 7899 12771 7905
rect 12802 7896 12808 7908
rect 12860 7896 12866 7948
rect 15933 7939 15991 7945
rect 15933 7905 15945 7939
rect 15979 7905 15991 7939
rect 15933 7899 15991 7905
rect 2869 7871 2927 7877
rect 2869 7837 2881 7871
rect 2915 7837 2927 7871
rect 3050 7868 3056 7880
rect 3011 7840 3056 7868
rect 2869 7831 2927 7837
rect 2884 7800 2912 7831
rect 3050 7828 3056 7840
rect 3108 7828 3114 7880
rect 3418 7868 3424 7880
rect 3379 7840 3424 7868
rect 3418 7828 3424 7840
rect 3476 7828 3482 7880
rect 4614 7828 4620 7880
rect 4672 7868 4678 7880
rect 4672 7840 4717 7868
rect 4672 7828 4678 7840
rect 5258 7828 5264 7880
rect 5316 7868 5322 7880
rect 5537 7871 5595 7877
rect 5537 7868 5549 7871
rect 5316 7840 5549 7868
rect 5316 7828 5322 7840
rect 5537 7837 5549 7840
rect 5583 7837 5595 7871
rect 5718 7868 5724 7880
rect 5679 7840 5724 7868
rect 5537 7831 5595 7837
rect 5718 7828 5724 7840
rect 5776 7828 5782 7880
rect 10873 7871 10931 7877
rect 10873 7868 10885 7871
rect 7576 7840 10885 7868
rect 3326 7800 3332 7812
rect 2884 7772 3332 7800
rect 1302 7692 1308 7744
rect 1360 7732 1366 7744
rect 2041 7735 2099 7741
rect 2041 7732 2053 7735
rect 1360 7704 2053 7732
rect 1360 7692 1366 7704
rect 2041 7701 2053 7704
rect 2087 7732 2099 7735
rect 2884 7732 2912 7772
rect 3326 7760 3332 7772
rect 3384 7760 3390 7812
rect 4062 7760 4068 7812
rect 4120 7800 4126 7812
rect 7576 7800 7604 7840
rect 10873 7837 10885 7840
rect 10919 7868 10931 7871
rect 11146 7868 11152 7880
rect 10919 7840 11152 7868
rect 10919 7837 10931 7840
rect 10873 7831 10931 7837
rect 11146 7828 11152 7840
rect 11204 7828 11210 7880
rect 11238 7828 11244 7880
rect 11296 7868 11302 7880
rect 12253 7871 12311 7877
rect 12253 7868 12265 7871
rect 11296 7840 12265 7868
rect 11296 7828 11302 7840
rect 12253 7837 12265 7840
rect 12299 7837 12311 7871
rect 15948 7868 15976 7899
rect 16206 7868 16212 7880
rect 12253 7831 12311 7837
rect 14844 7840 15976 7868
rect 16119 7840 16212 7868
rect 7742 7800 7748 7812
rect 4120 7772 7604 7800
rect 7655 7772 7748 7800
rect 4120 7760 4126 7772
rect 2087 7704 2912 7732
rect 5077 7735 5135 7741
rect 2087 7701 2099 7704
rect 2041 7695 2099 7701
rect 5077 7701 5089 7735
rect 5123 7732 5135 7735
rect 6822 7732 6828 7744
rect 5123 7704 6828 7732
rect 5123 7701 5135 7704
rect 5077 7695 5135 7701
rect 6822 7692 6828 7704
rect 6880 7692 6886 7744
rect 6914 7692 6920 7744
rect 6972 7732 6978 7744
rect 7668 7741 7696 7772
rect 7742 7760 7748 7772
rect 7800 7800 7806 7812
rect 8481 7803 8539 7809
rect 8481 7800 8493 7803
rect 7800 7772 8493 7800
rect 7800 7760 7806 7772
rect 8481 7769 8493 7772
rect 8527 7769 8539 7803
rect 8481 7763 8539 7769
rect 7653 7735 7711 7741
rect 7653 7732 7665 7735
rect 6972 7704 7665 7732
rect 6972 7692 6978 7704
rect 7653 7701 7665 7704
rect 7699 7701 7711 7735
rect 7653 7695 7711 7701
rect 9214 7692 9220 7744
rect 9272 7732 9278 7744
rect 9490 7732 9496 7744
rect 9272 7704 9496 7732
rect 9272 7692 9278 7704
rect 9490 7692 9496 7704
rect 9548 7692 9554 7744
rect 10042 7692 10048 7744
rect 10100 7732 10106 7744
rect 10413 7735 10471 7741
rect 10413 7732 10425 7735
rect 10100 7704 10425 7732
rect 10100 7692 10106 7704
rect 10413 7701 10425 7704
rect 10459 7732 10471 7735
rect 10962 7732 10968 7744
rect 10459 7704 10968 7732
rect 10459 7701 10471 7704
rect 10413 7695 10471 7701
rect 10962 7692 10968 7704
rect 11020 7692 11026 7744
rect 11698 7732 11704 7744
rect 11659 7704 11704 7732
rect 11698 7692 11704 7704
rect 11756 7692 11762 7744
rect 12268 7732 12296 7831
rect 14844 7744 14872 7840
rect 16206 7828 16212 7840
rect 16264 7868 16270 7880
rect 16500 7868 16528 7976
rect 19052 7973 19064 8007
rect 19098 8004 19110 8007
rect 19978 8004 19984 8016
rect 19098 7976 19984 8004
rect 19098 7973 19110 7976
rect 19052 7967 19110 7973
rect 19978 7964 19984 7976
rect 20036 7964 20042 8016
rect 16850 7945 16856 7948
rect 16844 7899 16856 7945
rect 16908 7936 16914 7948
rect 16908 7908 16944 7936
rect 16850 7896 16856 7899
rect 16908 7896 16914 7908
rect 17862 7896 17868 7948
rect 17920 7936 17926 7948
rect 18785 7939 18843 7945
rect 18785 7936 18797 7939
rect 17920 7908 18797 7936
rect 17920 7896 17926 7908
rect 18785 7905 18797 7908
rect 18831 7936 18843 7939
rect 19426 7936 19432 7948
rect 18831 7908 19432 7936
rect 18831 7905 18843 7908
rect 18785 7899 18843 7905
rect 19426 7896 19432 7908
rect 19484 7896 19490 7948
rect 16264 7840 16528 7868
rect 16264 7828 16270 7840
rect 16574 7828 16580 7880
rect 16632 7868 16638 7880
rect 16632 7840 16677 7868
rect 16632 7828 16638 7840
rect 14093 7735 14151 7741
rect 14093 7732 14105 7735
rect 12268 7704 14105 7732
rect 14093 7701 14105 7704
rect 14139 7701 14151 7735
rect 14826 7732 14832 7744
rect 14787 7704 14832 7732
rect 14093 7695 14151 7701
rect 14826 7692 14832 7704
rect 14884 7692 14890 7744
rect 15562 7732 15568 7744
rect 15523 7704 15568 7732
rect 15562 7692 15568 7704
rect 15620 7692 15626 7744
rect 20162 7732 20168 7744
rect 20123 7704 20168 7732
rect 20162 7692 20168 7704
rect 20220 7692 20226 7744
rect 1104 7642 21896 7664
rect 1104 7590 4447 7642
rect 4499 7590 4511 7642
rect 4563 7590 4575 7642
rect 4627 7590 4639 7642
rect 4691 7590 11378 7642
rect 11430 7590 11442 7642
rect 11494 7590 11506 7642
rect 11558 7590 11570 7642
rect 11622 7590 18308 7642
rect 18360 7590 18372 7642
rect 18424 7590 18436 7642
rect 18488 7590 18500 7642
rect 18552 7590 21896 7642
rect 1104 7568 21896 7590
rect 2409 7531 2467 7537
rect 2409 7497 2421 7531
rect 2455 7528 2467 7531
rect 2590 7528 2596 7540
rect 2455 7500 2596 7528
rect 2455 7497 2467 7500
rect 2409 7491 2467 7497
rect 2590 7488 2596 7500
rect 2648 7488 2654 7540
rect 4246 7528 4252 7540
rect 4207 7500 4252 7528
rect 4246 7488 4252 7500
rect 4304 7488 4310 7540
rect 5258 7528 5264 7540
rect 5219 7500 5264 7528
rect 5258 7488 5264 7500
rect 5316 7488 5322 7540
rect 8202 7528 8208 7540
rect 7852 7500 8208 7528
rect 2961 7395 3019 7401
rect 2961 7361 2973 7395
rect 3007 7392 3019 7395
rect 3050 7392 3056 7404
rect 3007 7364 3056 7392
rect 3007 7361 3019 7364
rect 2961 7355 3019 7361
rect 3050 7352 3056 7364
rect 3108 7352 3114 7404
rect 4154 7352 4160 7404
rect 4212 7392 4218 7404
rect 4709 7395 4767 7401
rect 4709 7392 4721 7395
rect 4212 7364 4721 7392
rect 4212 7352 4218 7364
rect 4709 7361 4721 7364
rect 4755 7361 4767 7395
rect 4709 7355 4767 7361
rect 4893 7395 4951 7401
rect 4893 7361 4905 7395
rect 4939 7392 4951 7395
rect 5442 7392 5448 7404
rect 4939 7364 5448 7392
rect 4939 7361 4951 7364
rect 4893 7355 4951 7361
rect 5442 7352 5448 7364
rect 5500 7392 5506 7404
rect 7852 7401 7880 7500
rect 8202 7488 8208 7500
rect 8260 7488 8266 7540
rect 9217 7531 9275 7537
rect 9217 7497 9229 7531
rect 9263 7528 9275 7531
rect 9306 7528 9312 7540
rect 9263 7500 9312 7528
rect 9263 7497 9275 7500
rect 9217 7491 9275 7497
rect 9306 7488 9312 7500
rect 9364 7488 9370 7540
rect 9490 7488 9496 7540
rect 9548 7528 9554 7540
rect 9677 7531 9735 7537
rect 9677 7528 9689 7531
rect 9548 7500 9689 7528
rect 9548 7488 9554 7500
rect 9677 7497 9689 7500
rect 9723 7497 9735 7531
rect 9677 7491 9735 7497
rect 9766 7488 9772 7540
rect 9824 7528 9830 7540
rect 16390 7528 16396 7540
rect 9824 7500 16396 7528
rect 9824 7488 9830 7500
rect 16390 7488 16396 7500
rect 16448 7488 16454 7540
rect 20438 7488 20444 7540
rect 20496 7528 20502 7540
rect 21085 7531 21143 7537
rect 21085 7528 21097 7531
rect 20496 7500 21097 7528
rect 20496 7488 20502 7500
rect 21085 7497 21097 7500
rect 21131 7497 21143 7531
rect 21085 7491 21143 7497
rect 16758 7420 16764 7472
rect 16816 7460 16822 7472
rect 16816 7432 17172 7460
rect 16816 7420 16822 7432
rect 5813 7395 5871 7401
rect 5813 7392 5825 7395
rect 5500 7364 5825 7392
rect 5500 7352 5506 7364
rect 5813 7361 5825 7364
rect 5859 7361 5871 7395
rect 5813 7355 5871 7361
rect 7837 7395 7895 7401
rect 7837 7361 7849 7395
rect 7883 7361 7895 7395
rect 7837 7355 7895 7361
rect 15562 7352 15568 7404
rect 15620 7392 15626 7404
rect 17144 7401 17172 7432
rect 17037 7395 17095 7401
rect 17037 7392 17049 7395
rect 15620 7364 17049 7392
rect 15620 7352 15626 7364
rect 17037 7361 17049 7364
rect 17083 7361 17095 7395
rect 17037 7355 17095 7361
rect 17129 7395 17187 7401
rect 17129 7361 17141 7395
rect 17175 7361 17187 7395
rect 19426 7392 19432 7404
rect 19387 7364 19432 7392
rect 17129 7355 17187 7361
rect 19426 7352 19432 7364
rect 19484 7352 19490 7404
rect 2777 7327 2835 7333
rect 2777 7293 2789 7327
rect 2823 7324 2835 7327
rect 3418 7324 3424 7336
rect 2823 7296 3424 7324
rect 2823 7293 2835 7296
rect 2777 7287 2835 7293
rect 3418 7284 3424 7296
rect 3476 7284 3482 7336
rect 5626 7324 5632 7336
rect 5539 7296 5632 7324
rect 5626 7284 5632 7296
rect 5684 7324 5690 7336
rect 10502 7324 10508 7336
rect 5684 7296 10508 7324
rect 5684 7284 5690 7296
rect 10502 7284 10508 7296
rect 10560 7284 10566 7336
rect 10689 7327 10747 7333
rect 10689 7293 10701 7327
rect 10735 7293 10747 7327
rect 10689 7287 10747 7293
rect 10956 7327 11014 7333
rect 10956 7293 10968 7327
rect 11002 7324 11014 7327
rect 11238 7324 11244 7336
rect 11002 7296 11244 7324
rect 11002 7293 11014 7296
rect 10956 7287 11014 7293
rect 3789 7259 3847 7265
rect 3789 7225 3801 7259
rect 3835 7256 3847 7259
rect 4617 7259 4675 7265
rect 4617 7256 4629 7259
rect 3835 7228 4629 7256
rect 3835 7225 3847 7228
rect 3789 7219 3847 7225
rect 4617 7225 4629 7228
rect 4663 7225 4675 7259
rect 4617 7219 4675 7225
rect 7742 7216 7748 7268
rect 7800 7256 7806 7268
rect 8082 7259 8140 7265
rect 8082 7256 8094 7259
rect 7800 7228 8094 7256
rect 7800 7216 7806 7228
rect 8082 7225 8094 7228
rect 8128 7225 8140 7259
rect 10594 7256 10600 7268
rect 8082 7219 8140 7225
rect 8220 7228 10600 7256
rect 1394 7188 1400 7200
rect 1355 7160 1400 7188
rect 1394 7148 1400 7160
rect 1452 7148 1458 7200
rect 2038 7188 2044 7200
rect 1999 7160 2044 7188
rect 2038 7148 2044 7160
rect 2096 7188 2102 7200
rect 2869 7191 2927 7197
rect 2869 7188 2881 7191
rect 2096 7160 2881 7188
rect 2096 7148 2102 7160
rect 2869 7157 2881 7160
rect 2915 7188 2927 7191
rect 3142 7188 3148 7200
rect 2915 7160 3148 7188
rect 2915 7157 2927 7160
rect 2869 7151 2927 7157
rect 3142 7148 3148 7160
rect 3200 7148 3206 7200
rect 5721 7191 5779 7197
rect 5721 7157 5733 7191
rect 5767 7188 5779 7191
rect 5810 7188 5816 7200
rect 5767 7160 5816 7188
rect 5767 7157 5779 7160
rect 5721 7151 5779 7157
rect 5810 7148 5816 7160
rect 5868 7188 5874 7200
rect 6273 7191 6331 7197
rect 6273 7188 6285 7191
rect 5868 7160 6285 7188
rect 5868 7148 5874 7160
rect 6273 7157 6285 7160
rect 6319 7188 6331 7191
rect 8220 7188 8248 7228
rect 10594 7216 10600 7228
rect 10652 7216 10658 7268
rect 10704 7256 10732 7287
rect 11238 7284 11244 7296
rect 11296 7284 11302 7336
rect 12894 7324 12900 7336
rect 11348 7296 12900 7324
rect 11348 7256 11376 7296
rect 12894 7284 12900 7296
rect 12952 7324 12958 7336
rect 13722 7324 13728 7336
rect 12952 7296 13728 7324
rect 12952 7284 12958 7296
rect 13722 7284 13728 7296
rect 13780 7324 13786 7336
rect 14001 7327 14059 7333
rect 14001 7324 14013 7327
rect 13780 7296 14013 7324
rect 13780 7284 13786 7296
rect 14001 7293 14013 7296
rect 14047 7293 14059 7327
rect 14001 7287 14059 7293
rect 14268 7327 14326 7333
rect 14268 7293 14280 7327
rect 14314 7324 14326 7327
rect 14550 7324 14556 7336
rect 14314 7296 14556 7324
rect 14314 7293 14326 7296
rect 14268 7287 14326 7293
rect 14550 7284 14556 7296
rect 14608 7284 14614 7336
rect 16945 7327 17003 7333
rect 16945 7293 16957 7327
rect 16991 7324 17003 7327
rect 18046 7324 18052 7336
rect 16991 7296 18052 7324
rect 16991 7293 17003 7296
rect 16945 7287 17003 7293
rect 18046 7284 18052 7296
rect 18104 7284 18110 7336
rect 19696 7327 19754 7333
rect 19696 7293 19708 7327
rect 19742 7324 19754 7327
rect 20162 7324 20168 7336
rect 19742 7296 20168 7324
rect 19742 7293 19754 7296
rect 19696 7287 19754 7293
rect 20162 7284 20168 7296
rect 20220 7284 20226 7336
rect 10704 7228 11376 7256
rect 12710 7216 12716 7268
rect 12768 7256 12774 7268
rect 13078 7256 13084 7268
rect 12768 7228 13084 7256
rect 12768 7216 12774 7228
rect 13078 7216 13084 7228
rect 13136 7256 13142 7268
rect 13136 7228 19196 7256
rect 13136 7216 13142 7228
rect 19168 7200 19196 7228
rect 12066 7188 12072 7200
rect 6319 7160 8248 7188
rect 12027 7160 12072 7188
rect 6319 7157 6331 7160
rect 6273 7151 6331 7157
rect 12066 7148 12072 7160
rect 12124 7148 12130 7200
rect 15378 7188 15384 7200
rect 15339 7160 15384 7188
rect 15378 7148 15384 7160
rect 15436 7148 15442 7200
rect 16574 7188 16580 7200
rect 16535 7160 16580 7188
rect 16574 7148 16580 7160
rect 16632 7148 16638 7200
rect 19150 7188 19156 7200
rect 19111 7160 19156 7188
rect 19150 7148 19156 7160
rect 19208 7148 19214 7200
rect 20254 7148 20260 7200
rect 20312 7188 20318 7200
rect 20809 7191 20867 7197
rect 20809 7188 20821 7191
rect 20312 7160 20821 7188
rect 20312 7148 20318 7160
rect 20809 7157 20821 7160
rect 20855 7157 20867 7191
rect 20809 7151 20867 7157
rect 1104 7098 21896 7120
rect 1104 7046 7912 7098
rect 7964 7046 7976 7098
rect 8028 7046 8040 7098
rect 8092 7046 8104 7098
rect 8156 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 15035 7098
rect 15087 7046 21896 7098
rect 1104 7024 21896 7046
rect 1394 6944 1400 6996
rect 1452 6984 1458 6996
rect 2041 6987 2099 6993
rect 2041 6984 2053 6987
rect 1452 6956 2053 6984
rect 1452 6944 1458 6956
rect 2041 6953 2053 6956
rect 2087 6953 2099 6987
rect 4154 6984 4160 6996
rect 4115 6956 4160 6984
rect 2041 6947 2099 6953
rect 4154 6944 4160 6956
rect 4212 6944 4218 6996
rect 5718 6944 5724 6996
rect 5776 6984 5782 6996
rect 5813 6987 5871 6993
rect 5813 6984 5825 6987
rect 5776 6956 5825 6984
rect 5776 6944 5782 6956
rect 5813 6953 5825 6956
rect 5859 6953 5871 6987
rect 7742 6984 7748 6996
rect 7703 6956 7748 6984
rect 5813 6947 5871 6953
rect 4890 6916 4896 6928
rect 4632 6888 4896 6916
rect 1946 6848 1952 6860
rect 1907 6820 1952 6848
rect 1946 6808 1952 6820
rect 2004 6808 2010 6860
rect 2774 6808 2780 6860
rect 2832 6848 2838 6860
rect 4062 6848 4068 6860
rect 2832 6820 4068 6848
rect 2832 6808 2838 6820
rect 4062 6808 4068 6820
rect 4120 6848 4126 6860
rect 4433 6851 4491 6857
rect 4433 6848 4445 6851
rect 4120 6820 4445 6848
rect 4120 6808 4126 6820
rect 4433 6817 4445 6820
rect 4479 6848 4491 6851
rect 4632 6848 4660 6888
rect 4890 6876 4896 6888
rect 4948 6876 4954 6928
rect 4479 6820 4660 6848
rect 4700 6851 4758 6857
rect 4479 6817 4491 6820
rect 4433 6811 4491 6817
rect 4700 6817 4712 6851
rect 4746 6848 4758 6851
rect 5442 6848 5448 6860
rect 4746 6820 5448 6848
rect 4746 6817 4758 6820
rect 4700 6811 4758 6817
rect 5442 6808 5448 6820
rect 5500 6808 5506 6860
rect 5828 6848 5856 6947
rect 7742 6944 7748 6956
rect 7800 6944 7806 6996
rect 8941 6987 8999 6993
rect 8941 6953 8953 6987
rect 8987 6984 8999 6987
rect 9030 6984 9036 6996
rect 8987 6956 9036 6984
rect 8987 6953 8999 6956
rect 8941 6947 8999 6953
rect 9030 6944 9036 6956
rect 9088 6984 9094 6996
rect 9677 6987 9735 6993
rect 9677 6984 9689 6987
rect 9088 6956 9689 6984
rect 9088 6944 9094 6956
rect 9677 6953 9689 6956
rect 9723 6984 9735 6987
rect 10502 6984 10508 6996
rect 9723 6956 10508 6984
rect 9723 6953 9735 6956
rect 9677 6947 9735 6953
rect 10502 6944 10508 6956
rect 10560 6944 10566 6996
rect 11698 6944 11704 6996
rect 11756 6984 11762 6996
rect 12345 6987 12403 6993
rect 12345 6984 12357 6987
rect 11756 6956 12357 6984
rect 11756 6944 11762 6956
rect 12345 6953 12357 6956
rect 12391 6953 12403 6987
rect 12345 6947 12403 6953
rect 12802 6944 12808 6996
rect 12860 6984 12866 6996
rect 16761 6987 16819 6993
rect 12860 6956 16712 6984
rect 12860 6944 12866 6956
rect 12250 6916 12256 6928
rect 8956 6888 9628 6916
rect 12211 6888 12256 6916
rect 6270 6848 6276 6860
rect 5828 6820 6276 6848
rect 6270 6808 6276 6820
rect 6328 6848 6334 6860
rect 6621 6851 6679 6857
rect 6621 6848 6633 6851
rect 6328 6820 6633 6848
rect 6328 6808 6334 6820
rect 6621 6817 6633 6820
rect 6667 6817 6679 6851
rect 6621 6811 6679 6817
rect 7098 6808 7104 6860
rect 7156 6848 7162 6860
rect 8021 6851 8079 6857
rect 8021 6848 8033 6851
rect 7156 6820 8033 6848
rect 7156 6808 7162 6820
rect 8021 6817 8033 6820
rect 8067 6848 8079 6851
rect 8956 6848 8984 6888
rect 8067 6820 8984 6848
rect 9033 6851 9091 6857
rect 8067 6817 8079 6820
rect 8021 6811 8079 6817
rect 9033 6817 9045 6851
rect 9079 6848 9091 6851
rect 9490 6848 9496 6860
rect 9079 6820 9496 6848
rect 9079 6817 9091 6820
rect 9033 6811 9091 6817
rect 9490 6808 9496 6820
rect 9548 6808 9554 6860
rect 9600 6848 9628 6888
rect 12250 6876 12256 6888
rect 12308 6876 12314 6928
rect 12526 6876 12532 6928
rect 12584 6916 12590 6928
rect 14001 6919 14059 6925
rect 14001 6916 14013 6919
rect 12584 6888 14013 6916
rect 12584 6876 12590 6888
rect 14001 6885 14013 6888
rect 14047 6916 14059 6919
rect 14274 6916 14280 6928
rect 14047 6888 14280 6916
rect 14047 6885 14059 6888
rect 14001 6879 14059 6885
rect 14274 6876 14280 6888
rect 14332 6916 14338 6928
rect 14642 6916 14648 6928
rect 14332 6888 14648 6916
rect 14332 6876 14338 6888
rect 14642 6876 14648 6888
rect 14700 6876 14706 6928
rect 16684 6916 16712 6956
rect 16761 6953 16773 6987
rect 16807 6984 16819 6987
rect 16850 6984 16856 6996
rect 16807 6956 16856 6984
rect 16807 6953 16819 6956
rect 16761 6947 16819 6953
rect 16850 6944 16856 6956
rect 16908 6944 16914 6996
rect 19150 6944 19156 6996
rect 19208 6984 19214 6996
rect 19981 6987 20039 6993
rect 19981 6984 19993 6987
rect 19208 6956 19993 6984
rect 19208 6944 19214 6956
rect 19981 6953 19993 6956
rect 20027 6953 20039 6987
rect 19981 6947 20039 6953
rect 18969 6919 19027 6925
rect 15580 6888 16436 6916
rect 16684 6888 18736 6916
rect 10318 6848 10324 6860
rect 9600 6820 10324 6848
rect 10318 6808 10324 6820
rect 10376 6808 10382 6860
rect 10496 6851 10554 6857
rect 10496 6817 10508 6851
rect 10542 6848 10554 6851
rect 12066 6848 12072 6860
rect 10542 6820 12072 6848
rect 10542 6817 10554 6820
rect 10496 6811 10554 6817
rect 12066 6808 12072 6820
rect 12124 6848 12130 6860
rect 15580 6848 15608 6888
rect 12124 6820 12480 6848
rect 12124 6808 12130 6820
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6780 2283 6783
rect 3050 6780 3056 6792
rect 2271 6752 3056 6780
rect 2271 6749 2283 6752
rect 2225 6743 2283 6749
rect 3050 6740 3056 6752
rect 3108 6740 3114 6792
rect 6365 6783 6423 6789
rect 6365 6749 6377 6783
rect 6411 6749 6423 6783
rect 6365 6743 6423 6749
rect 9217 6783 9275 6789
rect 9217 6749 9229 6783
rect 9263 6780 9275 6783
rect 9306 6780 9312 6792
rect 9263 6752 9312 6780
rect 9263 6749 9275 6752
rect 9217 6743 9275 6749
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6644 1639 6647
rect 1854 6644 1860 6656
rect 1627 6616 1860 6644
rect 1627 6613 1639 6616
rect 1581 6607 1639 6613
rect 1854 6604 1860 6616
rect 1912 6604 1918 6656
rect 2685 6647 2743 6653
rect 2685 6613 2697 6647
rect 2731 6644 2743 6647
rect 3142 6644 3148 6656
rect 2731 6616 3148 6644
rect 2731 6613 2743 6616
rect 2685 6607 2743 6613
rect 3142 6604 3148 6616
rect 3200 6604 3206 6656
rect 6380 6644 6408 6743
rect 9306 6740 9312 6752
rect 9364 6740 9370 6792
rect 12452 6789 12480 6820
rect 15212 6820 15608 6848
rect 15648 6851 15706 6857
rect 10229 6783 10287 6789
rect 10229 6749 10241 6783
rect 10275 6749 10287 6783
rect 10229 6743 10287 6749
rect 12437 6783 12495 6789
rect 12437 6749 12449 6783
rect 12483 6749 12495 6783
rect 12437 6743 12495 6749
rect 8202 6672 8208 6724
rect 8260 6712 8266 6724
rect 10134 6712 10140 6724
rect 8260 6684 10140 6712
rect 8260 6672 8266 6684
rect 10134 6672 10140 6684
rect 10192 6712 10198 6724
rect 10244 6712 10272 6743
rect 13630 6740 13636 6792
rect 13688 6780 13694 6792
rect 14461 6783 14519 6789
rect 14461 6780 14473 6783
rect 13688 6752 14473 6780
rect 13688 6740 13694 6752
rect 14461 6749 14473 6752
rect 14507 6780 14519 6783
rect 15212 6780 15240 6820
rect 15648 6817 15660 6851
rect 15694 6848 15706 6851
rect 16206 6848 16212 6860
rect 15694 6820 16212 6848
rect 15694 6817 15706 6820
rect 15648 6811 15706 6817
rect 16206 6808 16212 6820
rect 16264 6808 16270 6860
rect 14507 6752 15240 6780
rect 14507 6749 14519 6752
rect 14461 6743 14519 6749
rect 15286 6740 15292 6792
rect 15344 6780 15350 6792
rect 15381 6783 15439 6789
rect 15381 6780 15393 6783
rect 15344 6752 15393 6780
rect 15344 6740 15350 6752
rect 15381 6749 15393 6752
rect 15427 6749 15439 6783
rect 16408 6780 16436 6888
rect 18598 6848 18604 6860
rect 16776 6820 18604 6848
rect 16776 6780 16804 6820
rect 18598 6808 18604 6820
rect 18656 6808 18662 6860
rect 18708 6848 18736 6888
rect 18969 6885 18981 6919
rect 19015 6916 19027 6919
rect 19015 6888 20944 6916
rect 19015 6885 19027 6888
rect 18969 6879 19027 6885
rect 19702 6848 19708 6860
rect 18708 6820 19708 6848
rect 19702 6808 19708 6820
rect 19760 6808 19766 6860
rect 20073 6851 20131 6857
rect 20073 6817 20085 6851
rect 20119 6848 20131 6851
rect 20438 6848 20444 6860
rect 20119 6820 20444 6848
rect 20119 6817 20131 6820
rect 20073 6811 20131 6817
rect 20438 6808 20444 6820
rect 20496 6808 20502 6860
rect 20916 6857 20944 6888
rect 20901 6851 20959 6857
rect 20901 6817 20913 6851
rect 20947 6817 20959 6851
rect 20901 6811 20959 6817
rect 16408 6752 16804 6780
rect 17037 6783 17095 6789
rect 15381 6743 15439 6749
rect 17037 6749 17049 6783
rect 17083 6780 17095 6783
rect 17126 6780 17132 6792
rect 17083 6752 17132 6780
rect 17083 6749 17095 6752
rect 17037 6743 17095 6749
rect 10192 6684 10272 6712
rect 10192 6672 10198 6684
rect 8220 6644 8248 6672
rect 6380 6616 8248 6644
rect 8573 6647 8631 6653
rect 8573 6613 8585 6647
rect 8619 6644 8631 6647
rect 9582 6644 9588 6656
rect 8619 6616 9588 6644
rect 8619 6613 8631 6616
rect 8573 6607 8631 6613
rect 9582 6604 9588 6616
rect 9640 6604 9646 6656
rect 10962 6604 10968 6656
rect 11020 6644 11026 6656
rect 11609 6647 11667 6653
rect 11609 6644 11621 6647
rect 11020 6616 11621 6644
rect 11020 6604 11026 6616
rect 11609 6613 11621 6616
rect 11655 6613 11667 6647
rect 11882 6644 11888 6656
rect 11843 6616 11888 6644
rect 11609 6607 11667 6613
rect 11882 6604 11888 6616
rect 11940 6604 11946 6656
rect 15396 6644 15424 6743
rect 17126 6740 17132 6752
rect 17184 6740 17190 6792
rect 18138 6740 18144 6792
rect 18196 6780 18202 6792
rect 18874 6780 18880 6792
rect 18196 6752 18880 6780
rect 18196 6740 18202 6752
rect 18874 6740 18880 6752
rect 18932 6740 18938 6792
rect 19061 6783 19119 6789
rect 19061 6749 19073 6783
rect 19107 6749 19119 6783
rect 19061 6743 19119 6749
rect 19245 6783 19303 6789
rect 19245 6749 19257 6783
rect 19291 6780 19303 6783
rect 19291 6752 20024 6780
rect 19291 6749 19303 6752
rect 19245 6743 19303 6749
rect 19076 6712 19104 6743
rect 19613 6715 19671 6721
rect 19613 6712 19625 6715
rect 19076 6684 19625 6712
rect 19613 6681 19625 6684
rect 19659 6681 19671 6715
rect 19996 6712 20024 6752
rect 20162 6740 20168 6792
rect 20220 6780 20226 6792
rect 20220 6752 20265 6780
rect 20220 6740 20226 6752
rect 20254 6712 20260 6724
rect 19996 6684 20260 6712
rect 19613 6675 19671 6681
rect 20254 6672 20260 6684
rect 20312 6672 20318 6724
rect 16482 6644 16488 6656
rect 15396 6616 16488 6644
rect 16482 6604 16488 6616
rect 16540 6604 16546 6656
rect 18601 6647 18659 6653
rect 18601 6613 18613 6647
rect 18647 6644 18659 6647
rect 18874 6644 18880 6656
rect 18647 6616 18880 6644
rect 18647 6613 18659 6616
rect 18601 6607 18659 6613
rect 18874 6604 18880 6616
rect 18932 6604 18938 6656
rect 1104 6554 21896 6576
rect 1104 6502 4447 6554
rect 4499 6502 4511 6554
rect 4563 6502 4575 6554
rect 4627 6502 4639 6554
rect 4691 6502 11378 6554
rect 11430 6502 11442 6554
rect 11494 6502 11506 6554
rect 11558 6502 11570 6554
rect 11622 6502 18308 6554
rect 18360 6502 18372 6554
rect 18424 6502 18436 6554
rect 18488 6502 18500 6554
rect 18552 6502 21896 6554
rect 1104 6480 21896 6502
rect 5534 6400 5540 6452
rect 5592 6440 5598 6452
rect 9585 6443 9643 6449
rect 9585 6440 9597 6443
rect 5592 6412 9597 6440
rect 5592 6400 5598 6412
rect 9585 6409 9597 6412
rect 9631 6409 9643 6443
rect 9858 6440 9864 6452
rect 9819 6412 9864 6440
rect 9585 6403 9643 6409
rect 3970 6332 3976 6384
rect 4028 6372 4034 6384
rect 4985 6375 5043 6381
rect 4985 6372 4997 6375
rect 4028 6344 4997 6372
rect 4028 6332 4034 6344
rect 4985 6341 4997 6344
rect 5031 6372 5043 6375
rect 5626 6372 5632 6384
rect 5031 6344 5632 6372
rect 5031 6341 5043 6344
rect 4985 6335 5043 6341
rect 5626 6332 5632 6344
rect 5684 6332 5690 6384
rect 6454 6332 6460 6384
rect 6512 6372 6518 6384
rect 8110 6372 8116 6384
rect 6512 6344 8116 6372
rect 6512 6332 6518 6344
rect 8110 6332 8116 6344
rect 8168 6332 8174 6384
rect 9600 6372 9628 6403
rect 9858 6400 9864 6412
rect 9916 6400 9922 6452
rect 11885 6443 11943 6449
rect 11885 6409 11897 6443
rect 11931 6440 11943 6443
rect 11974 6440 11980 6452
rect 11931 6412 11980 6440
rect 11931 6409 11943 6412
rect 11885 6403 11943 6409
rect 11974 6400 11980 6412
rect 12032 6400 12038 6452
rect 18138 6440 18144 6452
rect 18099 6412 18144 6440
rect 18138 6400 18144 6412
rect 18196 6400 18202 6452
rect 18969 6443 19027 6449
rect 18969 6409 18981 6443
rect 19015 6440 19027 6443
rect 20346 6440 20352 6452
rect 19015 6412 20352 6440
rect 19015 6409 19027 6412
rect 18969 6403 19027 6409
rect 20346 6400 20352 6412
rect 20404 6400 20410 6452
rect 9600 6344 10456 6372
rect 2133 6307 2191 6313
rect 2133 6273 2145 6307
rect 2179 6304 2191 6307
rect 2866 6304 2872 6316
rect 2179 6276 2872 6304
rect 2179 6273 2191 6276
rect 2133 6267 2191 6273
rect 2866 6264 2872 6276
rect 2924 6264 2930 6316
rect 3050 6304 3056 6316
rect 3011 6276 3056 6304
rect 3050 6264 3056 6276
rect 3108 6264 3114 6316
rect 6270 6304 6276 6316
rect 6231 6276 6276 6304
rect 6270 6264 6276 6276
rect 6328 6264 6334 6316
rect 7374 6304 7380 6316
rect 7335 6276 7380 6304
rect 7374 6264 7380 6276
rect 7432 6264 7438 6316
rect 8202 6304 8208 6316
rect 8163 6276 8208 6304
rect 8202 6264 8208 6276
rect 8260 6264 8266 6316
rect 9582 6264 9588 6316
rect 9640 6304 9646 6316
rect 10428 6313 10456 6344
rect 10594 6332 10600 6384
rect 10652 6372 10658 6384
rect 11609 6375 11667 6381
rect 11609 6372 11621 6375
rect 10652 6344 11621 6372
rect 10652 6332 10658 6344
rect 11609 6341 11621 6344
rect 11655 6341 11667 6375
rect 11609 6335 11667 6341
rect 13173 6375 13231 6381
rect 13173 6341 13185 6375
rect 13219 6372 13231 6375
rect 14366 6372 14372 6384
rect 13219 6344 14372 6372
rect 13219 6341 13231 6344
rect 13173 6335 13231 6341
rect 14366 6332 14372 6344
rect 14424 6332 14430 6384
rect 18156 6372 18184 6400
rect 16224 6344 18184 6372
rect 10321 6307 10379 6313
rect 10321 6304 10333 6307
rect 9640 6276 10333 6304
rect 9640 6264 9646 6276
rect 10321 6273 10333 6276
rect 10367 6273 10379 6307
rect 10321 6267 10379 6273
rect 10413 6307 10471 6313
rect 10413 6273 10425 6307
rect 10459 6273 10471 6307
rect 10413 6267 10471 6273
rect 10502 6264 10508 6316
rect 10560 6304 10566 6316
rect 13630 6304 13636 6316
rect 10560 6276 13636 6304
rect 10560 6264 10566 6276
rect 13630 6264 13636 6276
rect 13688 6264 13694 6316
rect 13814 6304 13820 6316
rect 13727 6276 13820 6304
rect 13814 6264 13820 6276
rect 13872 6304 13878 6316
rect 16224 6313 16252 6344
rect 14737 6307 14795 6313
rect 14737 6304 14749 6307
rect 13872 6276 14749 6304
rect 13872 6264 13878 6276
rect 14737 6273 14749 6276
rect 14783 6273 14795 6307
rect 14737 6267 14795 6273
rect 16209 6307 16267 6313
rect 16209 6273 16221 6307
rect 16255 6273 16267 6307
rect 16209 6267 16267 6273
rect 16298 6264 16304 6316
rect 16356 6304 16362 6316
rect 16393 6307 16451 6313
rect 16393 6304 16405 6307
rect 16356 6276 16405 6304
rect 16356 6264 16362 6276
rect 16393 6273 16405 6276
rect 16439 6304 16451 6307
rect 17310 6304 17316 6316
rect 16439 6276 17316 6304
rect 16439 6273 16451 6276
rect 16393 6267 16451 6273
rect 17310 6264 17316 6276
rect 17368 6264 17374 6316
rect 19613 6307 19671 6313
rect 19613 6273 19625 6307
rect 19659 6304 19671 6307
rect 19886 6304 19892 6316
rect 19659 6276 19892 6304
rect 19659 6273 19671 6276
rect 19613 6267 19671 6273
rect 19886 6264 19892 6276
rect 19944 6264 19950 6316
rect 1854 6236 1860 6248
rect 1815 6208 1860 6236
rect 1854 6196 1860 6208
rect 1912 6196 1918 6248
rect 7190 6236 7196 6248
rect 7103 6208 7196 6236
rect 7190 6196 7196 6208
rect 7248 6236 7254 6248
rect 7929 6239 7987 6245
rect 7929 6236 7941 6239
rect 7248 6208 7941 6236
rect 7248 6196 7254 6208
rect 7929 6205 7941 6208
rect 7975 6236 7987 6239
rect 12710 6236 12716 6248
rect 7975 6208 12716 6236
rect 7975 6205 7987 6208
rect 7929 6199 7987 6205
rect 12710 6196 12716 6208
rect 12768 6196 12774 6248
rect 15381 6239 15439 6245
rect 15381 6236 15393 6239
rect 12820 6208 15393 6236
rect 2869 6171 2927 6177
rect 2869 6137 2881 6171
rect 2915 6168 2927 6171
rect 3142 6168 3148 6180
rect 2915 6140 3148 6168
rect 2915 6137 2927 6140
rect 2869 6131 2927 6137
rect 3142 6128 3148 6140
rect 3200 6128 3206 6180
rect 6270 6128 6276 6180
rect 6328 6168 6334 6180
rect 8472 6171 8530 6177
rect 6328 6140 8432 6168
rect 6328 6128 6334 6140
rect 1486 6100 1492 6112
rect 1447 6072 1492 6100
rect 1486 6060 1492 6072
rect 1544 6060 1550 6112
rect 1949 6103 2007 6109
rect 1949 6069 1961 6103
rect 1995 6100 2007 6103
rect 2501 6103 2559 6109
rect 2501 6100 2513 6103
rect 1995 6072 2513 6100
rect 1995 6069 2007 6072
rect 1949 6063 2007 6069
rect 2501 6069 2513 6072
rect 2547 6069 2559 6103
rect 2501 6063 2559 6069
rect 2961 6103 3019 6109
rect 2961 6069 2973 6103
rect 3007 6100 3019 6103
rect 3602 6100 3608 6112
rect 3007 6072 3608 6100
rect 3007 6069 3019 6072
rect 2961 6063 3019 6069
rect 3602 6060 3608 6072
rect 3660 6060 3666 6112
rect 5445 6103 5503 6109
rect 5445 6069 5457 6103
rect 5491 6100 5503 6103
rect 5534 6100 5540 6112
rect 5491 6072 5540 6100
rect 5491 6069 5503 6072
rect 5445 6063 5503 6069
rect 5534 6060 5540 6072
rect 5592 6060 5598 6112
rect 5718 6100 5724 6112
rect 5679 6072 5724 6100
rect 5718 6060 5724 6072
rect 5776 6060 5782 6112
rect 6086 6100 6092 6112
rect 6047 6072 6092 6100
rect 6086 6060 6092 6072
rect 6144 6060 6150 6112
rect 6181 6103 6239 6109
rect 6181 6069 6193 6103
rect 6227 6100 6239 6103
rect 6825 6103 6883 6109
rect 6825 6100 6837 6103
rect 6227 6072 6837 6100
rect 6227 6069 6239 6072
rect 6181 6063 6239 6069
rect 6825 6069 6837 6072
rect 6871 6069 6883 6103
rect 6825 6063 6883 6069
rect 7098 6060 7104 6112
rect 7156 6100 7162 6112
rect 7285 6103 7343 6109
rect 7285 6100 7297 6103
rect 7156 6072 7297 6100
rect 7156 6060 7162 6072
rect 7285 6069 7297 6072
rect 7331 6069 7343 6103
rect 8404 6100 8432 6140
rect 8472 6137 8484 6171
rect 8518 6168 8530 6171
rect 9306 6168 9312 6180
rect 8518 6140 9312 6168
rect 8518 6137 8530 6140
rect 8472 6131 8530 6137
rect 9306 6128 9312 6140
rect 9364 6128 9370 6180
rect 11609 6171 11667 6177
rect 9416 6140 11560 6168
rect 9416 6100 9444 6140
rect 10226 6100 10232 6112
rect 8404 6072 9444 6100
rect 10187 6072 10232 6100
rect 7285 6063 7343 6069
rect 10226 6060 10232 6072
rect 10284 6060 10290 6112
rect 10686 6060 10692 6112
rect 10744 6100 10750 6112
rect 11422 6100 11428 6112
rect 10744 6072 11428 6100
rect 10744 6060 10750 6072
rect 11422 6060 11428 6072
rect 11480 6060 11486 6112
rect 11532 6100 11560 6140
rect 11609 6137 11621 6171
rect 11655 6168 11667 6171
rect 12820 6168 12848 6208
rect 15381 6205 15393 6208
rect 15427 6236 15439 6239
rect 16117 6239 16175 6245
rect 16117 6236 16129 6239
rect 15427 6208 16129 6236
rect 15427 6205 15439 6208
rect 15381 6199 15439 6205
rect 16117 6205 16129 6208
rect 16163 6205 16175 6239
rect 17126 6236 17132 6248
rect 17087 6208 17132 6236
rect 16117 6199 16175 6205
rect 17126 6196 17132 6208
rect 17184 6196 17190 6248
rect 17218 6196 17224 6248
rect 17276 6236 17282 6248
rect 17678 6236 17684 6248
rect 17276 6208 17684 6236
rect 17276 6196 17282 6208
rect 17678 6196 17684 6208
rect 17736 6196 17742 6248
rect 19334 6196 19340 6248
rect 19392 6196 19398 6248
rect 19426 6196 19432 6248
rect 19484 6236 19490 6248
rect 20254 6245 20260 6248
rect 19981 6239 20039 6245
rect 19981 6236 19993 6239
rect 19484 6208 19993 6236
rect 19484 6196 19490 6208
rect 19981 6205 19993 6208
rect 20027 6205 20039 6239
rect 20248 6236 20260 6245
rect 20215 6208 20260 6236
rect 19981 6199 20039 6205
rect 20248 6199 20260 6208
rect 20254 6196 20260 6199
rect 20312 6196 20318 6248
rect 11655 6140 12848 6168
rect 12897 6171 12955 6177
rect 11655 6137 11667 6140
rect 11609 6131 11667 6137
rect 12897 6137 12909 6171
rect 12943 6168 12955 6171
rect 13541 6171 13599 6177
rect 13541 6168 13553 6171
rect 12943 6140 13553 6168
rect 12943 6137 12955 6140
rect 12897 6131 12955 6137
rect 13541 6137 13553 6140
rect 13587 6137 13599 6171
rect 19352 6168 19380 6196
rect 19794 6168 19800 6180
rect 19352 6140 19800 6168
rect 13541 6131 13599 6137
rect 12912 6100 12940 6131
rect 19794 6128 19800 6140
rect 19852 6128 19858 6180
rect 14182 6100 14188 6112
rect 11532 6072 12940 6100
rect 14143 6072 14188 6100
rect 14182 6060 14188 6072
rect 14240 6060 14246 6112
rect 14550 6100 14556 6112
rect 14511 6072 14556 6100
rect 14550 6060 14556 6072
rect 14608 6060 14614 6112
rect 14642 6060 14648 6112
rect 14700 6100 14706 6112
rect 15746 6100 15752 6112
rect 14700 6072 14745 6100
rect 15707 6072 15752 6100
rect 14700 6060 14706 6072
rect 15746 6060 15752 6072
rect 15804 6060 15810 6112
rect 16482 6060 16488 6112
rect 16540 6100 16546 6112
rect 16761 6103 16819 6109
rect 16761 6100 16773 6103
rect 16540 6072 16773 6100
rect 16540 6060 16546 6072
rect 16761 6069 16773 6072
rect 16807 6069 16819 6103
rect 18690 6100 18696 6112
rect 18651 6072 18696 6100
rect 16761 6063 16819 6069
rect 18690 6060 18696 6072
rect 18748 6060 18754 6112
rect 19334 6100 19340 6112
rect 19295 6072 19340 6100
rect 19334 6060 19340 6072
rect 19392 6060 19398 6112
rect 19426 6060 19432 6112
rect 19484 6100 19490 6112
rect 21358 6100 21364 6112
rect 19484 6072 19529 6100
rect 21319 6072 21364 6100
rect 19484 6060 19490 6072
rect 21358 6060 21364 6072
rect 21416 6060 21422 6112
rect 1104 6010 21896 6032
rect 1104 5958 7912 6010
rect 7964 5958 7976 6010
rect 8028 5958 8040 6010
rect 8092 5958 8104 6010
rect 8156 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 15035 6010
rect 15087 5958 21896 6010
rect 1104 5936 21896 5958
rect 1857 5899 1915 5905
rect 1857 5865 1869 5899
rect 1903 5896 1915 5899
rect 1946 5896 1952 5908
rect 1903 5868 1952 5896
rect 1903 5865 1915 5868
rect 1857 5859 1915 5865
rect 1946 5856 1952 5868
rect 2004 5856 2010 5908
rect 6086 5856 6092 5908
rect 6144 5896 6150 5908
rect 6181 5899 6239 5905
rect 6181 5896 6193 5899
rect 6144 5868 6193 5896
rect 6144 5856 6150 5868
rect 6181 5865 6193 5868
rect 6227 5865 6239 5899
rect 6181 5859 6239 5865
rect 6822 5856 6828 5908
rect 6880 5896 6886 5908
rect 7561 5899 7619 5905
rect 7561 5896 7573 5899
rect 6880 5868 7573 5896
rect 6880 5856 6886 5868
rect 7561 5865 7573 5868
rect 7607 5865 7619 5899
rect 7561 5859 7619 5865
rect 8573 5899 8631 5905
rect 8573 5865 8585 5899
rect 8619 5896 8631 5899
rect 10226 5896 10232 5908
rect 8619 5868 10232 5896
rect 8619 5865 8631 5868
rect 8573 5859 8631 5865
rect 10226 5856 10232 5868
rect 10284 5856 10290 5908
rect 11790 5896 11796 5908
rect 10888 5868 11796 5896
rect 2584 5831 2642 5837
rect 2584 5797 2596 5831
rect 2630 5828 2642 5831
rect 2866 5828 2872 5840
rect 2630 5800 2872 5828
rect 2630 5797 2642 5800
rect 2584 5791 2642 5797
rect 2866 5788 2872 5800
rect 2924 5788 2930 5840
rect 4062 5828 4068 5840
rect 3620 5800 4068 5828
rect 3620 5760 3648 5800
rect 4062 5788 4068 5800
rect 4120 5788 4126 5840
rect 5718 5788 5724 5840
rect 5776 5828 5782 5840
rect 7653 5831 7711 5837
rect 7653 5828 7665 5831
rect 5776 5800 7665 5828
rect 5776 5788 5782 5800
rect 7653 5797 7665 5800
rect 7699 5797 7711 5831
rect 9401 5831 9459 5837
rect 9401 5828 9413 5831
rect 7653 5791 7711 5797
rect 7760 5800 9413 5828
rect 4321 5763 4379 5769
rect 4321 5760 4333 5763
rect 2332 5732 3648 5760
rect 3712 5732 4333 5760
rect 1578 5652 1584 5704
rect 1636 5692 1642 5704
rect 2332 5701 2360 5732
rect 2317 5695 2375 5701
rect 2317 5692 2329 5695
rect 1636 5664 2329 5692
rect 1636 5652 1642 5664
rect 2317 5661 2329 5664
rect 2363 5661 2375 5695
rect 2317 5655 2375 5661
rect 2958 5516 2964 5568
rect 3016 5556 3022 5568
rect 3712 5565 3740 5732
rect 4321 5729 4333 5732
rect 4367 5729 4379 5763
rect 4321 5723 4379 5729
rect 5534 5720 5540 5772
rect 5592 5760 5598 5772
rect 6546 5760 6552 5772
rect 5592 5732 6552 5760
rect 5592 5720 5598 5732
rect 6546 5720 6552 5732
rect 6604 5760 6610 5772
rect 7760 5760 7788 5800
rect 9401 5797 9413 5800
rect 9447 5797 9459 5831
rect 9401 5791 9459 5797
rect 9582 5788 9588 5840
rect 9640 5828 9646 5840
rect 10888 5828 10916 5868
rect 11790 5856 11796 5868
rect 11848 5856 11854 5908
rect 11974 5856 11980 5908
rect 12032 5856 12038 5908
rect 14550 5896 14556 5908
rect 14511 5868 14556 5896
rect 14550 5856 14556 5868
rect 14608 5856 14614 5908
rect 16482 5896 16488 5908
rect 16443 5868 16488 5896
rect 16482 5856 16488 5868
rect 16540 5856 16546 5908
rect 17218 5896 17224 5908
rect 17179 5868 17224 5896
rect 17218 5856 17224 5868
rect 17276 5856 17282 5908
rect 18233 5899 18291 5905
rect 18233 5865 18245 5899
rect 18279 5896 18291 5899
rect 18690 5896 18696 5908
rect 18279 5868 18696 5896
rect 18279 5865 18291 5868
rect 18233 5859 18291 5865
rect 18690 5856 18696 5868
rect 18748 5856 18754 5908
rect 19334 5856 19340 5908
rect 19392 5896 19398 5908
rect 19613 5899 19671 5905
rect 19613 5896 19625 5899
rect 19392 5868 19625 5896
rect 19392 5856 19398 5868
rect 19613 5865 19625 5868
rect 19659 5865 19671 5899
rect 19613 5859 19671 5865
rect 20073 5899 20131 5905
rect 20073 5865 20085 5899
rect 20119 5896 20131 5899
rect 20622 5896 20628 5908
rect 20119 5868 20628 5896
rect 20119 5865 20131 5868
rect 20073 5859 20131 5865
rect 9640 5800 10916 5828
rect 11057 5831 11115 5837
rect 9640 5788 9646 5800
rect 11057 5797 11069 5831
rect 11103 5828 11115 5831
rect 11992 5828 12020 5856
rect 11103 5800 12020 5828
rect 11103 5797 11115 5800
rect 11057 5791 11115 5797
rect 12526 5788 12532 5840
rect 12584 5828 12590 5840
rect 17954 5828 17960 5840
rect 12584 5800 17960 5828
rect 12584 5788 12590 5800
rect 17954 5788 17960 5800
rect 18012 5788 18018 5840
rect 19702 5828 19708 5840
rect 19352 5800 19708 5828
rect 6604 5732 7788 5760
rect 8941 5763 8999 5769
rect 6604 5720 6610 5732
rect 8941 5729 8953 5763
rect 8987 5760 8999 5763
rect 9600 5760 9628 5788
rect 8987 5732 9628 5760
rect 10321 5763 10379 5769
rect 8987 5729 8999 5732
rect 8941 5723 8999 5729
rect 10321 5729 10333 5763
rect 10367 5760 10379 5763
rect 10686 5760 10692 5772
rect 10367 5732 10692 5760
rect 10367 5729 10379 5732
rect 10321 5723 10379 5729
rect 10686 5720 10692 5732
rect 10744 5760 10750 5772
rect 10965 5763 11023 5769
rect 10965 5760 10977 5763
rect 10744 5732 10977 5760
rect 10744 5720 10750 5732
rect 10965 5729 10977 5732
rect 11011 5729 11023 5763
rect 11974 5760 11980 5772
rect 11935 5732 11980 5760
rect 10965 5723 11023 5729
rect 11974 5720 11980 5732
rect 12032 5720 12038 5772
rect 12084 5732 12296 5760
rect 4062 5692 4068 5704
rect 4023 5664 4068 5692
rect 4062 5652 4068 5664
rect 4120 5652 4126 5704
rect 6270 5652 6276 5704
rect 6328 5692 6334 5704
rect 6641 5695 6699 5701
rect 6641 5692 6653 5695
rect 6328 5664 6653 5692
rect 6328 5652 6334 5664
rect 6641 5661 6653 5664
rect 6687 5661 6699 5695
rect 6641 5655 6699 5661
rect 6825 5695 6883 5701
rect 6825 5661 6837 5695
rect 6871 5692 6883 5695
rect 7374 5692 7380 5704
rect 6871 5664 7380 5692
rect 6871 5661 6883 5664
rect 6825 5655 6883 5661
rect 5442 5624 5448 5636
rect 5355 5596 5448 5624
rect 5442 5584 5448 5596
rect 5500 5624 5506 5636
rect 6840 5624 6868 5655
rect 7374 5652 7380 5664
rect 7432 5652 7438 5704
rect 7742 5692 7748 5704
rect 7703 5664 7748 5692
rect 7742 5652 7748 5664
rect 7800 5652 7806 5704
rect 8570 5652 8576 5704
rect 8628 5692 8634 5704
rect 9033 5695 9091 5701
rect 9033 5692 9045 5695
rect 8628 5664 9045 5692
rect 8628 5652 8634 5664
rect 9033 5661 9045 5664
rect 9079 5661 9091 5695
rect 9033 5655 9091 5661
rect 9217 5695 9275 5701
rect 9217 5661 9229 5695
rect 9263 5692 9275 5695
rect 9306 5692 9312 5704
rect 9263 5664 9312 5692
rect 9263 5661 9275 5664
rect 9217 5655 9275 5661
rect 9306 5652 9312 5664
rect 9364 5652 9370 5704
rect 9401 5695 9459 5701
rect 9401 5661 9413 5695
rect 9447 5692 9459 5695
rect 10594 5692 10600 5704
rect 9447 5664 10600 5692
rect 9447 5661 9459 5664
rect 9401 5655 9459 5661
rect 10594 5652 10600 5664
rect 10652 5652 10658 5704
rect 11241 5695 11299 5701
rect 11241 5661 11253 5695
rect 11287 5661 11299 5695
rect 11241 5655 11299 5661
rect 5500 5596 6868 5624
rect 7193 5627 7251 5633
rect 5500 5584 5506 5596
rect 7193 5593 7205 5627
rect 7239 5624 7251 5627
rect 10318 5624 10324 5636
rect 7239 5596 10324 5624
rect 7239 5593 7251 5596
rect 7193 5587 7251 5593
rect 10318 5584 10324 5596
rect 10376 5584 10382 5636
rect 10962 5584 10968 5636
rect 11020 5624 11026 5636
rect 11256 5624 11284 5655
rect 11422 5652 11428 5704
rect 11480 5692 11486 5704
rect 12084 5701 12112 5732
rect 12069 5695 12127 5701
rect 12069 5692 12081 5695
rect 11480 5664 12081 5692
rect 11480 5652 11486 5664
rect 12069 5661 12081 5664
rect 12115 5661 12127 5695
rect 12069 5655 12127 5661
rect 12161 5695 12219 5701
rect 12161 5661 12173 5695
rect 12207 5661 12219 5695
rect 12268 5692 12296 5732
rect 12434 5720 12440 5772
rect 12492 5760 12498 5772
rect 12894 5760 12900 5772
rect 12492 5732 12900 5760
rect 12492 5720 12498 5732
rect 12894 5720 12900 5732
rect 12952 5720 12958 5772
rect 13164 5763 13222 5769
rect 13164 5729 13176 5763
rect 13210 5760 13222 5763
rect 13722 5760 13728 5772
rect 13210 5732 13728 5760
rect 13210 5729 13222 5732
rect 13164 5723 13222 5729
rect 13722 5720 13728 5732
rect 13780 5720 13786 5772
rect 15746 5720 15752 5772
rect 15804 5760 15810 5772
rect 16577 5763 16635 5769
rect 16577 5760 16589 5763
rect 15804 5732 16589 5760
rect 15804 5720 15810 5732
rect 16577 5729 16589 5732
rect 16623 5729 16635 5763
rect 18325 5763 18383 5769
rect 16577 5723 16635 5729
rect 16684 5732 18276 5760
rect 12802 5692 12808 5704
rect 12268 5664 12808 5692
rect 12161 5655 12219 5661
rect 12176 5624 12204 5655
rect 12802 5652 12808 5664
rect 12860 5652 12866 5704
rect 15378 5652 15384 5704
rect 15436 5692 15442 5704
rect 16684 5692 16712 5732
rect 15436 5664 16712 5692
rect 16761 5695 16819 5701
rect 15436 5652 15442 5664
rect 16761 5661 16773 5695
rect 16807 5692 16819 5695
rect 16850 5692 16856 5704
rect 16807 5664 16856 5692
rect 16807 5661 16819 5664
rect 16761 5655 16819 5661
rect 16850 5652 16856 5664
rect 16908 5652 16914 5704
rect 18248 5692 18276 5732
rect 18325 5729 18337 5763
rect 18371 5760 18383 5763
rect 19058 5760 19064 5772
rect 18371 5732 19064 5760
rect 18371 5729 18383 5732
rect 18325 5723 18383 5729
rect 19058 5720 19064 5732
rect 19116 5720 19122 5772
rect 19352 5769 19380 5800
rect 19702 5788 19708 5800
rect 19760 5828 19766 5840
rect 20088 5828 20116 5859
rect 20622 5856 20628 5868
rect 20680 5856 20686 5908
rect 19760 5800 20116 5828
rect 19760 5788 19766 5800
rect 19337 5763 19395 5769
rect 19337 5729 19349 5763
rect 19383 5729 19395 5763
rect 19978 5760 19984 5772
rect 19939 5732 19984 5760
rect 19337 5723 19395 5729
rect 19978 5720 19984 5732
rect 20036 5720 20042 5772
rect 18417 5695 18475 5701
rect 18417 5692 18429 5695
rect 18248 5664 18429 5692
rect 18417 5661 18429 5664
rect 18463 5692 18475 5695
rect 18598 5692 18604 5704
rect 18463 5664 18604 5692
rect 18463 5661 18475 5664
rect 18417 5655 18475 5661
rect 18598 5652 18604 5664
rect 18656 5652 18662 5704
rect 20254 5692 20260 5704
rect 20215 5664 20260 5692
rect 20254 5652 20260 5664
rect 20312 5652 20318 5704
rect 15289 5627 15347 5633
rect 15289 5624 15301 5627
rect 11020 5596 12204 5624
rect 14108 5596 15301 5624
rect 11020 5584 11026 5596
rect 3697 5559 3755 5565
rect 3697 5556 3709 5559
rect 3016 5528 3709 5556
rect 3016 5516 3022 5528
rect 3697 5525 3709 5528
rect 3743 5525 3755 5559
rect 3697 5519 3755 5525
rect 5905 5559 5963 5565
rect 5905 5525 5917 5559
rect 5951 5556 5963 5559
rect 6270 5556 6276 5568
rect 5951 5528 6276 5556
rect 5951 5525 5963 5528
rect 5905 5519 5963 5525
rect 6270 5516 6276 5528
rect 6328 5516 6334 5568
rect 8297 5559 8355 5565
rect 8297 5525 8309 5559
rect 8343 5556 8355 5559
rect 8570 5556 8576 5568
rect 8343 5528 8576 5556
rect 8343 5525 8355 5528
rect 8297 5519 8355 5525
rect 8570 5516 8576 5528
rect 8628 5516 8634 5568
rect 9582 5516 9588 5568
rect 9640 5556 9646 5568
rect 9677 5559 9735 5565
rect 9677 5556 9689 5559
rect 9640 5528 9689 5556
rect 9640 5516 9646 5528
rect 9677 5525 9689 5528
rect 9723 5525 9735 5559
rect 9677 5519 9735 5525
rect 10597 5559 10655 5565
rect 10597 5525 10609 5559
rect 10643 5556 10655 5559
rect 11238 5556 11244 5568
rect 10643 5528 11244 5556
rect 10643 5525 10655 5528
rect 10597 5519 10655 5525
rect 11238 5516 11244 5528
rect 11296 5516 11302 5568
rect 11609 5559 11667 5565
rect 11609 5525 11621 5559
rect 11655 5556 11667 5559
rect 11698 5556 11704 5568
rect 11655 5528 11704 5556
rect 11655 5525 11667 5528
rect 11609 5519 11667 5525
rect 11698 5516 11704 5528
rect 11756 5516 11762 5568
rect 11790 5516 11796 5568
rect 11848 5556 11854 5568
rect 14108 5556 14136 5596
rect 15289 5593 15301 5596
rect 15335 5624 15347 5627
rect 15470 5624 15476 5636
rect 15335 5596 15476 5624
rect 15335 5593 15347 5596
rect 15289 5587 15347 5593
rect 15470 5584 15476 5596
rect 15528 5584 15534 5636
rect 17865 5627 17923 5633
rect 17865 5593 17877 5627
rect 17911 5624 17923 5627
rect 19150 5624 19156 5636
rect 17911 5596 19156 5624
rect 17911 5593 17923 5596
rect 17865 5587 17923 5593
rect 19150 5584 19156 5596
rect 19208 5584 19214 5636
rect 14274 5556 14280 5568
rect 11848 5528 14136 5556
rect 14235 5528 14280 5556
rect 11848 5516 11854 5528
rect 14274 5516 14280 5528
rect 14332 5516 14338 5568
rect 16117 5559 16175 5565
rect 16117 5525 16129 5559
rect 16163 5556 16175 5559
rect 17034 5556 17040 5568
rect 16163 5528 17040 5556
rect 16163 5525 16175 5528
rect 16117 5519 16175 5525
rect 17034 5516 17040 5528
rect 17092 5516 17098 5568
rect 18969 5559 19027 5565
rect 18969 5525 18981 5559
rect 19015 5556 19027 5559
rect 19058 5556 19064 5568
rect 19015 5528 19064 5556
rect 19015 5525 19027 5528
rect 18969 5519 19027 5525
rect 19058 5516 19064 5528
rect 19116 5516 19122 5568
rect 21266 5556 21272 5568
rect 21227 5528 21272 5556
rect 21266 5516 21272 5528
rect 21324 5516 21330 5568
rect 1104 5466 21896 5488
rect 1104 5414 4447 5466
rect 4499 5414 4511 5466
rect 4563 5414 4575 5466
rect 4627 5414 4639 5466
rect 4691 5414 11378 5466
rect 11430 5414 11442 5466
rect 11494 5414 11506 5466
rect 11558 5414 11570 5466
rect 11622 5414 18308 5466
rect 18360 5414 18372 5466
rect 18424 5414 18436 5466
rect 18488 5414 18500 5466
rect 18552 5414 21896 5466
rect 1104 5392 21896 5414
rect 3789 5355 3847 5361
rect 3789 5321 3801 5355
rect 3835 5352 3847 5355
rect 9950 5352 9956 5364
rect 3835 5324 9956 5352
rect 3835 5321 3847 5324
rect 3789 5315 3847 5321
rect 9950 5312 9956 5324
rect 10008 5312 10014 5364
rect 11146 5312 11152 5364
rect 11204 5352 11210 5364
rect 12342 5352 12348 5364
rect 11204 5324 12348 5352
rect 11204 5312 11210 5324
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 13814 5352 13820 5364
rect 13775 5324 13820 5352
rect 13814 5312 13820 5324
rect 13872 5312 13878 5364
rect 16022 5312 16028 5364
rect 16080 5352 16086 5364
rect 16117 5355 16175 5361
rect 16117 5352 16129 5355
rect 16080 5324 16129 5352
rect 16080 5312 16086 5324
rect 16117 5321 16129 5324
rect 16163 5321 16175 5355
rect 16117 5315 16175 5321
rect 16390 5312 16396 5364
rect 16448 5352 16454 5364
rect 16485 5355 16543 5361
rect 16485 5352 16497 5355
rect 16448 5324 16497 5352
rect 16448 5312 16454 5324
rect 16485 5321 16497 5324
rect 16531 5321 16543 5355
rect 16485 5315 16543 5321
rect 19426 5312 19432 5364
rect 19484 5352 19490 5364
rect 19705 5355 19763 5361
rect 19705 5352 19717 5355
rect 19484 5324 19717 5352
rect 19484 5312 19490 5324
rect 19705 5321 19717 5324
rect 19751 5321 19763 5355
rect 19705 5315 19763 5321
rect 1489 5287 1547 5293
rect 1489 5253 1501 5287
rect 1535 5284 1547 5287
rect 2774 5284 2780 5296
rect 1535 5256 2780 5284
rect 1535 5253 1547 5256
rect 1489 5247 1547 5253
rect 2774 5244 2780 5256
rect 2832 5244 2838 5296
rect 3878 5244 3884 5296
rect 3936 5284 3942 5296
rect 5261 5287 5319 5293
rect 5261 5284 5273 5287
rect 3936 5256 5273 5284
rect 3936 5244 3942 5256
rect 5261 5253 5273 5256
rect 5307 5284 5319 5287
rect 6454 5284 6460 5296
rect 5307 5256 6460 5284
rect 5307 5253 5319 5256
rect 5261 5247 5319 5253
rect 6454 5244 6460 5256
rect 6512 5244 6518 5296
rect 9398 5244 9404 5296
rect 9456 5284 9462 5296
rect 9582 5284 9588 5296
rect 9456 5256 9588 5284
rect 9456 5244 9462 5256
rect 9582 5244 9588 5256
rect 9640 5244 9646 5296
rect 15286 5244 15292 5296
rect 15344 5284 15350 5296
rect 17862 5284 17868 5296
rect 15344 5256 17868 5284
rect 15344 5244 15350 5256
rect 17862 5244 17868 5256
rect 17920 5284 17926 5296
rect 17920 5256 18092 5284
rect 17920 5244 17926 5256
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5216 2191 5219
rect 2958 5216 2964 5228
rect 2179 5188 2964 5216
rect 2179 5185 2191 5188
rect 2133 5179 2191 5185
rect 2958 5176 2964 5188
rect 3016 5176 3022 5228
rect 3050 5176 3056 5228
rect 3108 5216 3114 5228
rect 3973 5219 4031 5225
rect 3108 5188 3153 5216
rect 3108 5176 3114 5188
rect 3973 5185 3985 5219
rect 4019 5216 4031 5219
rect 4154 5216 4160 5228
rect 4019 5188 4160 5216
rect 4019 5185 4031 5188
rect 3973 5179 4031 5185
rect 1486 5108 1492 5160
rect 1544 5148 1550 5160
rect 1857 5151 1915 5157
rect 1857 5148 1869 5151
rect 1544 5120 1869 5148
rect 1544 5108 1550 5120
rect 1857 5117 1869 5120
rect 1903 5117 1915 5151
rect 1857 5111 1915 5117
rect 198 5040 204 5092
rect 256 5080 262 5092
rect 2869 5083 2927 5089
rect 2869 5080 2881 5083
rect 256 5052 2881 5080
rect 256 5040 262 5052
rect 2869 5049 2881 5052
rect 2915 5049 2927 5083
rect 2869 5043 2927 5049
rect 2961 5083 3019 5089
rect 2961 5049 2973 5083
rect 3007 5080 3019 5083
rect 3988 5080 4016 5179
rect 4154 5176 4160 5188
rect 4212 5176 4218 5228
rect 5718 5176 5724 5228
rect 5776 5216 5782 5228
rect 6089 5219 6147 5225
rect 6089 5216 6101 5219
rect 5776 5188 6101 5216
rect 5776 5176 5782 5188
rect 6089 5185 6101 5188
rect 6135 5185 6147 5219
rect 6089 5179 6147 5185
rect 10134 5176 10140 5228
rect 10192 5216 10198 5228
rect 10413 5219 10471 5225
rect 10413 5216 10425 5219
rect 10192 5188 10425 5216
rect 10192 5176 10198 5188
rect 10413 5185 10425 5188
rect 10459 5185 10471 5219
rect 10413 5179 10471 5185
rect 14274 5176 14280 5228
rect 14332 5216 14338 5228
rect 14645 5219 14703 5225
rect 14645 5216 14657 5219
rect 14332 5188 14657 5216
rect 14332 5176 14338 5188
rect 14645 5185 14657 5188
rect 14691 5185 14703 5219
rect 14645 5179 14703 5185
rect 15378 5176 15384 5228
rect 15436 5216 15442 5228
rect 18064 5225 18092 5256
rect 15657 5219 15715 5225
rect 15657 5216 15669 5219
rect 15436 5188 15669 5216
rect 15436 5176 15442 5188
rect 15657 5185 15669 5188
rect 15703 5185 15715 5219
rect 15657 5179 15715 5185
rect 18049 5219 18107 5225
rect 18049 5185 18061 5219
rect 18095 5185 18107 5219
rect 18049 5179 18107 5185
rect 19150 5176 19156 5228
rect 19208 5216 19214 5228
rect 20165 5219 20223 5225
rect 20165 5216 20177 5219
rect 19208 5188 20177 5216
rect 19208 5176 19214 5188
rect 20165 5185 20177 5188
rect 20211 5185 20223 5219
rect 20165 5179 20223 5185
rect 20254 5176 20260 5228
rect 20312 5216 20318 5228
rect 20312 5188 20405 5216
rect 20312 5176 20318 5188
rect 5905 5151 5963 5157
rect 5905 5117 5917 5151
rect 5951 5148 5963 5151
rect 5994 5148 6000 5160
rect 5951 5120 6000 5148
rect 5951 5117 5963 5120
rect 5905 5111 5963 5117
rect 5994 5108 6000 5120
rect 6052 5108 6058 5160
rect 10680 5151 10738 5157
rect 10680 5117 10692 5151
rect 10726 5148 10738 5151
rect 10962 5148 10968 5160
rect 10726 5120 10968 5148
rect 10726 5117 10738 5120
rect 10680 5111 10738 5117
rect 10962 5108 10968 5120
rect 11020 5108 11026 5160
rect 12434 5148 12440 5160
rect 12395 5120 12440 5148
rect 12434 5108 12440 5120
rect 12492 5108 12498 5160
rect 14182 5108 14188 5160
rect 14240 5148 14246 5160
rect 14461 5151 14519 5157
rect 14461 5148 14473 5151
rect 14240 5120 14473 5148
rect 14240 5108 14246 5120
rect 14461 5117 14473 5120
rect 14507 5117 14519 5151
rect 15470 5148 15476 5160
rect 15431 5120 15476 5148
rect 14461 5111 14519 5117
rect 15470 5108 15476 5120
rect 15528 5108 15534 5160
rect 20073 5151 20131 5157
rect 20073 5148 20085 5151
rect 18156 5120 20085 5148
rect 3007 5052 4016 5080
rect 3007 5049 3019 5052
rect 2961 5043 3019 5049
rect 1949 5015 2007 5021
rect 1949 4981 1961 5015
rect 1995 5012 2007 5015
rect 2222 5012 2228 5024
rect 1995 4984 2228 5012
rect 1995 4981 2007 4984
rect 1949 4975 2007 4981
rect 2222 4972 2228 4984
rect 2280 4972 2286 5024
rect 2501 5015 2559 5021
rect 2501 4981 2513 5015
rect 2547 5012 2559 5015
rect 2682 5012 2688 5024
rect 2547 4984 2688 5012
rect 2547 4981 2559 4984
rect 2501 4975 2559 4981
rect 2682 4972 2688 4984
rect 2740 4972 2746 5024
rect 2884 5012 2912 5043
rect 4062 5040 4068 5092
rect 4120 5080 4126 5092
rect 7561 5083 7619 5089
rect 7561 5080 7573 5083
rect 4120 5052 7573 5080
rect 4120 5040 4126 5052
rect 7561 5049 7573 5052
rect 7607 5080 7619 5083
rect 8202 5080 8208 5092
rect 7607 5052 8208 5080
rect 7607 5049 7619 5052
rect 7561 5043 7619 5049
rect 8202 5040 8208 5052
rect 8260 5040 8266 5092
rect 12682 5083 12740 5089
rect 12682 5080 12694 5083
rect 11808 5052 12694 5080
rect 3513 5015 3571 5021
rect 3513 5012 3525 5015
rect 2884 4984 3525 5012
rect 3513 4981 3525 4984
rect 3559 5012 3571 5015
rect 3789 5015 3847 5021
rect 3789 5012 3801 5015
rect 3559 4984 3801 5012
rect 3559 4981 3571 4984
rect 3513 4975 3571 4981
rect 3789 4981 3801 4984
rect 3835 4981 3847 5015
rect 5534 5012 5540 5024
rect 5495 4984 5540 5012
rect 3789 4975 3847 4981
rect 5534 4972 5540 4984
rect 5592 4972 5598 5024
rect 5997 5015 6055 5021
rect 5997 4981 6009 5015
rect 6043 5012 6055 5015
rect 6454 5012 6460 5024
rect 6043 4984 6460 5012
rect 6043 4981 6055 4984
rect 5997 4975 6055 4981
rect 6454 4972 6460 4984
rect 6512 4972 6518 5024
rect 11606 4972 11612 5024
rect 11664 5012 11670 5024
rect 11808 5021 11836 5052
rect 12682 5049 12694 5052
rect 12728 5049 12740 5083
rect 12682 5043 12740 5049
rect 14366 5040 14372 5092
rect 14424 5080 14430 5092
rect 14553 5083 14611 5089
rect 14553 5080 14565 5083
rect 14424 5052 14565 5080
rect 14424 5040 14430 5052
rect 14553 5049 14565 5052
rect 14599 5049 14611 5083
rect 18156 5080 18184 5120
rect 20073 5117 20085 5120
rect 20119 5117 20131 5151
rect 20272 5148 20300 5176
rect 20073 5111 20131 5117
rect 20180 5120 20300 5148
rect 20809 5151 20867 5157
rect 14553 5043 14611 5049
rect 15120 5052 18184 5080
rect 18316 5083 18374 5089
rect 11793 5015 11851 5021
rect 11793 5012 11805 5015
rect 11664 4984 11805 5012
rect 11664 4972 11670 4984
rect 11793 4981 11805 4984
rect 11839 4981 11851 5015
rect 11793 4975 11851 4981
rect 13906 4972 13912 5024
rect 13964 5012 13970 5024
rect 15120 5021 15148 5052
rect 18316 5049 18328 5083
rect 18362 5080 18374 5083
rect 18598 5080 18604 5092
rect 18362 5052 18604 5080
rect 18362 5049 18374 5052
rect 18316 5043 18374 5049
rect 18598 5040 18604 5052
rect 18656 5040 18662 5092
rect 20180 5080 20208 5120
rect 20809 5117 20821 5151
rect 20855 5148 20867 5151
rect 21266 5148 21272 5160
rect 20855 5120 21272 5148
rect 20855 5117 20867 5120
rect 20809 5111 20867 5117
rect 21266 5108 21272 5120
rect 21324 5108 21330 5160
rect 19444 5052 20208 5080
rect 19444 5024 19472 5052
rect 14093 5015 14151 5021
rect 14093 5012 14105 5015
rect 13964 4984 14105 5012
rect 13964 4972 13970 4984
rect 14093 4981 14105 4984
rect 14139 4981 14151 5015
rect 14093 4975 14151 4981
rect 15105 5015 15163 5021
rect 15105 4981 15117 5015
rect 15151 4981 15163 5015
rect 15105 4975 15163 4981
rect 15562 4972 15568 5024
rect 15620 5012 15626 5024
rect 19426 5012 19432 5024
rect 15620 4984 15665 5012
rect 19387 4984 19432 5012
rect 15620 4972 15626 4984
rect 19426 4972 19432 4984
rect 19484 4972 19490 5024
rect 20438 4972 20444 5024
rect 20496 5012 20502 5024
rect 20993 5015 21051 5021
rect 20993 5012 21005 5015
rect 20496 4984 21005 5012
rect 20496 4972 20502 4984
rect 20993 4981 21005 4984
rect 21039 4981 21051 5015
rect 20993 4975 21051 4981
rect 1104 4922 21896 4944
rect 1104 4870 7912 4922
rect 7964 4870 7976 4922
rect 8028 4870 8040 4922
rect 8092 4870 8104 4922
rect 8156 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 15035 4922
rect 15087 4870 21896 4922
rect 1104 4848 21896 4870
rect 2222 4808 2228 4820
rect 2183 4780 2228 4808
rect 2222 4768 2228 4780
rect 2280 4768 2286 4820
rect 2682 4808 2688 4820
rect 2643 4780 2688 4808
rect 2682 4768 2688 4780
rect 2740 4768 2746 4820
rect 3970 4768 3976 4820
rect 4028 4808 4034 4820
rect 4157 4811 4215 4817
rect 4157 4808 4169 4811
rect 4028 4780 4169 4808
rect 4028 4768 4034 4780
rect 4157 4777 4169 4780
rect 4203 4808 4215 4811
rect 5169 4811 5227 4817
rect 5169 4808 5181 4811
rect 4203 4780 5181 4808
rect 4203 4777 4215 4780
rect 4157 4771 4215 4777
rect 5169 4777 5181 4780
rect 5215 4777 5227 4811
rect 5169 4771 5227 4777
rect 5626 4768 5632 4820
rect 5684 4808 5690 4820
rect 6273 4811 6331 4817
rect 6273 4808 6285 4811
rect 5684 4780 6285 4808
rect 5684 4768 5690 4780
rect 6273 4777 6285 4780
rect 6319 4808 6331 4811
rect 7009 4811 7067 4817
rect 7009 4808 7021 4811
rect 6319 4780 7021 4808
rect 6319 4777 6331 4780
rect 6273 4771 6331 4777
rect 7009 4777 7021 4780
rect 7055 4808 7067 4811
rect 7190 4808 7196 4820
rect 7055 4780 7196 4808
rect 7055 4777 7067 4780
rect 7009 4771 7067 4777
rect 7190 4768 7196 4780
rect 7248 4768 7254 4820
rect 8202 4768 8208 4820
rect 8260 4808 8266 4820
rect 8297 4811 8355 4817
rect 8297 4808 8309 4811
rect 8260 4780 8309 4808
rect 8260 4768 8266 4780
rect 8297 4777 8309 4780
rect 8343 4777 8355 4811
rect 8297 4771 8355 4777
rect 8389 4811 8447 4817
rect 8389 4777 8401 4811
rect 8435 4808 8447 4811
rect 10778 4808 10784 4820
rect 8435 4780 10784 4808
rect 8435 4777 8447 4780
rect 8389 4771 8447 4777
rect 6365 4743 6423 4749
rect 6365 4709 6377 4743
rect 6411 4740 6423 4743
rect 7466 4740 7472 4752
rect 6411 4712 7472 4740
rect 6411 4709 6423 4712
rect 6365 4703 6423 4709
rect 7466 4700 7472 4712
rect 7524 4700 7530 4752
rect 7653 4743 7711 4749
rect 7653 4709 7665 4743
rect 7699 4740 7711 4743
rect 8404 4740 8432 4771
rect 10778 4768 10784 4780
rect 10836 4768 10842 4820
rect 11333 4811 11391 4817
rect 11333 4777 11345 4811
rect 11379 4808 11391 4811
rect 11698 4808 11704 4820
rect 11379 4780 11704 4808
rect 11379 4777 11391 4780
rect 11333 4771 11391 4777
rect 11698 4768 11704 4780
rect 11756 4768 11762 4820
rect 11974 4808 11980 4820
rect 11935 4780 11980 4808
rect 11974 4768 11980 4780
rect 12032 4768 12038 4820
rect 12342 4768 12348 4820
rect 12400 4808 12406 4820
rect 13538 4808 13544 4820
rect 12400 4780 13544 4808
rect 12400 4768 12406 4780
rect 13538 4768 13544 4780
rect 13596 4768 13602 4820
rect 17129 4811 17187 4817
rect 17129 4777 17141 4811
rect 17175 4808 17187 4811
rect 17310 4808 17316 4820
rect 17175 4780 17316 4808
rect 17175 4777 17187 4780
rect 17129 4771 17187 4777
rect 17310 4768 17316 4780
rect 17368 4768 17374 4820
rect 19978 4768 19984 4820
rect 20036 4808 20042 4820
rect 20349 4811 20407 4817
rect 20349 4808 20361 4811
rect 20036 4780 20361 4808
rect 20036 4768 20042 4780
rect 20349 4777 20361 4780
rect 20395 4777 20407 4811
rect 20349 4771 20407 4777
rect 7699 4712 8432 4740
rect 7699 4709 7711 4712
rect 7653 4703 7711 4709
rect 2593 4675 2651 4681
rect 2593 4641 2605 4675
rect 2639 4672 2651 4675
rect 3142 4672 3148 4684
rect 2639 4644 3148 4672
rect 2639 4641 2651 4644
rect 2593 4635 2651 4641
rect 3142 4632 3148 4644
rect 3200 4632 3206 4684
rect 3602 4632 3608 4684
rect 3660 4672 3666 4684
rect 7668 4672 7696 4703
rect 8570 4700 8576 4752
rect 8628 4700 8634 4752
rect 11238 4700 11244 4752
rect 11296 4740 11302 4752
rect 11425 4743 11483 4749
rect 11425 4740 11437 4743
rect 11296 4712 11437 4740
rect 11296 4700 11302 4712
rect 11425 4709 11437 4712
rect 11471 4709 11483 4743
rect 11425 4703 11483 4709
rect 18960 4743 19018 4749
rect 18960 4709 18972 4743
rect 19006 4740 19018 4743
rect 19426 4740 19432 4752
rect 19006 4712 19432 4740
rect 19006 4709 19018 4712
rect 18960 4703 19018 4709
rect 19426 4700 19432 4712
rect 19484 4700 19490 4752
rect 3660 4644 7696 4672
rect 8588 4672 8616 4700
rect 14737 4675 14795 4681
rect 14737 4672 14749 4675
rect 8588 4644 14749 4672
rect 3660 4632 3666 4644
rect 14737 4641 14749 4644
rect 14783 4672 14795 4675
rect 15562 4672 15568 4684
rect 14783 4644 15568 4672
rect 14783 4641 14795 4644
rect 14737 4635 14795 4641
rect 15562 4632 15568 4644
rect 15620 4632 15626 4684
rect 16016 4675 16074 4681
rect 16016 4641 16028 4675
rect 16062 4672 16074 4675
rect 16482 4672 16488 4684
rect 16062 4644 16488 4672
rect 16062 4641 16074 4644
rect 16016 4635 16074 4641
rect 16482 4632 16488 4644
rect 16540 4632 16546 4684
rect 17862 4632 17868 4684
rect 17920 4672 17926 4684
rect 18693 4675 18751 4681
rect 18693 4672 18705 4675
rect 17920 4644 18705 4672
rect 17920 4632 17926 4644
rect 18693 4641 18705 4644
rect 18739 4672 18751 4675
rect 19334 4672 19340 4684
rect 18739 4644 19340 4672
rect 18739 4641 18751 4644
rect 18693 4635 18751 4641
rect 19334 4632 19340 4644
rect 19392 4632 19398 4684
rect 20622 4632 20628 4684
rect 20680 4672 20686 4684
rect 20901 4675 20959 4681
rect 20901 4672 20913 4675
rect 20680 4644 20913 4672
rect 20680 4632 20686 4644
rect 20901 4641 20913 4644
rect 20947 4641 20959 4675
rect 20901 4635 20959 4641
rect 2866 4604 2872 4616
rect 2827 4576 2872 4604
rect 2866 4564 2872 4576
rect 2924 4564 2930 4616
rect 2958 4564 2964 4616
rect 3016 4604 3022 4616
rect 3620 4604 3648 4632
rect 3016 4576 3648 4604
rect 5261 4607 5319 4613
rect 3016 4564 3022 4576
rect 5261 4573 5273 4607
rect 5307 4573 5319 4607
rect 5261 4567 5319 4573
rect 5445 4607 5503 4613
rect 5445 4573 5457 4607
rect 5491 4604 5503 4607
rect 5718 4604 5724 4616
rect 5491 4576 5724 4604
rect 5491 4573 5503 4576
rect 5445 4567 5503 4573
rect 3418 4496 3424 4548
rect 3476 4536 3482 4548
rect 4433 4539 4491 4545
rect 4433 4536 4445 4539
rect 3476 4508 4445 4536
rect 3476 4496 3482 4508
rect 4433 4505 4445 4508
rect 4479 4536 4491 4539
rect 5276 4536 5304 4567
rect 5718 4564 5724 4576
rect 5776 4604 5782 4616
rect 6457 4607 6515 4613
rect 6457 4604 6469 4607
rect 5776 4576 6469 4604
rect 5776 4564 5782 4576
rect 6457 4573 6469 4576
rect 6503 4573 6515 4607
rect 6457 4567 6515 4573
rect 8573 4607 8631 4613
rect 8573 4573 8585 4607
rect 8619 4573 8631 4607
rect 8938 4604 8944 4616
rect 8899 4576 8944 4604
rect 8573 4567 8631 4573
rect 5810 4536 5816 4548
rect 4479 4508 5816 4536
rect 4479 4505 4491 4508
rect 4433 4499 4491 4505
rect 5810 4496 5816 4508
rect 5868 4496 5874 4548
rect 8588 4536 8616 4567
rect 8938 4564 8944 4576
rect 8996 4564 9002 4616
rect 11606 4604 11612 4616
rect 11567 4576 11612 4604
rect 11606 4564 11612 4576
rect 11664 4564 11670 4616
rect 15286 4564 15292 4616
rect 15344 4604 15350 4616
rect 15749 4607 15807 4613
rect 15749 4604 15761 4607
rect 15344 4576 15761 4604
rect 15344 4564 15350 4576
rect 15749 4573 15761 4576
rect 15795 4573 15807 4607
rect 15749 4567 15807 4573
rect 8846 4536 8852 4548
rect 8588 4508 8852 4536
rect 8846 4496 8852 4508
rect 8904 4496 8910 4548
rect 19886 4496 19892 4548
rect 19944 4536 19950 4548
rect 20073 4539 20131 4545
rect 20073 4536 20085 4539
rect 19944 4508 20085 4536
rect 19944 4496 19950 4508
rect 20073 4505 20085 4508
rect 20119 4505 20131 4539
rect 20073 4499 20131 4505
rect 3329 4471 3387 4477
rect 3329 4437 3341 4471
rect 3375 4468 3387 4471
rect 3602 4468 3608 4480
rect 3375 4440 3608 4468
rect 3375 4437 3387 4440
rect 3329 4431 3387 4437
rect 3602 4428 3608 4440
rect 3660 4428 3666 4480
rect 4798 4468 4804 4480
rect 4759 4440 4804 4468
rect 4798 4428 4804 4440
rect 4856 4428 4862 4480
rect 5902 4468 5908 4480
rect 5863 4440 5908 4468
rect 5902 4428 5908 4440
rect 5960 4428 5966 4480
rect 7834 4428 7840 4480
rect 7892 4468 7898 4480
rect 7929 4471 7987 4477
rect 7929 4468 7941 4471
rect 7892 4440 7941 4468
rect 7892 4428 7898 4440
rect 7929 4437 7941 4440
rect 7975 4437 7987 4471
rect 7929 4431 7987 4437
rect 10965 4471 11023 4477
rect 10965 4437 10977 4471
rect 11011 4468 11023 4471
rect 11698 4468 11704 4480
rect 11011 4440 11704 4468
rect 11011 4437 11023 4440
rect 10965 4431 11023 4437
rect 11698 4428 11704 4440
rect 11756 4428 11762 4480
rect 15381 4471 15439 4477
rect 15381 4437 15393 4471
rect 15427 4468 15439 4471
rect 15470 4468 15476 4480
rect 15427 4440 15476 4468
rect 15427 4437 15439 4440
rect 15381 4431 15439 4437
rect 15470 4428 15476 4440
rect 15528 4428 15534 4480
rect 19978 4428 19984 4480
rect 20036 4468 20042 4480
rect 21085 4471 21143 4477
rect 21085 4468 21097 4471
rect 20036 4440 21097 4468
rect 20036 4428 20042 4440
rect 21085 4437 21097 4440
rect 21131 4437 21143 4471
rect 21085 4431 21143 4437
rect 1104 4378 21896 4400
rect 1104 4326 4447 4378
rect 4499 4326 4511 4378
rect 4563 4326 4575 4378
rect 4627 4326 4639 4378
rect 4691 4326 11378 4378
rect 11430 4326 11442 4378
rect 11494 4326 11506 4378
rect 11558 4326 11570 4378
rect 11622 4326 18308 4378
rect 18360 4326 18372 4378
rect 18424 4326 18436 4378
rect 18488 4326 18500 4378
rect 18552 4326 21896 4378
rect 1104 4304 21896 4326
rect 2866 4264 2872 4276
rect 2827 4236 2872 4264
rect 2866 4224 2872 4236
rect 2924 4224 2930 4276
rect 3142 4264 3148 4276
rect 3103 4236 3148 4264
rect 3142 4224 3148 4236
rect 3200 4224 3206 4276
rect 6825 4267 6883 4273
rect 6825 4233 6837 4267
rect 6871 4264 6883 4267
rect 7466 4264 7472 4276
rect 6871 4236 7472 4264
rect 6871 4233 6883 4236
rect 6825 4227 6883 4233
rect 7466 4224 7472 4236
rect 7524 4224 7530 4276
rect 8570 4264 8576 4276
rect 7944 4236 8576 4264
rect 3878 4156 3884 4208
rect 3936 4196 3942 4208
rect 7742 4196 7748 4208
rect 3936 4168 7748 4196
rect 3936 4156 3942 4168
rect 7742 4156 7748 4168
rect 7800 4156 7806 4208
rect 2961 4131 3019 4137
rect 2961 4097 2973 4131
rect 3007 4128 3019 4131
rect 3602 4128 3608 4140
rect 3007 4100 3608 4128
rect 3007 4097 3019 4100
rect 2961 4091 3019 4097
rect 3602 4088 3608 4100
rect 3660 4088 3666 4140
rect 3697 4131 3755 4137
rect 3697 4097 3709 4131
rect 3743 4097 3755 4131
rect 3697 4091 3755 4097
rect 1486 4060 1492 4072
rect 1447 4032 1492 4060
rect 1486 4020 1492 4032
rect 1544 4020 1550 4072
rect 1756 4063 1814 4069
rect 1756 4029 1768 4063
rect 1802 4060 1814 4063
rect 3050 4060 3056 4072
rect 1802 4032 3056 4060
rect 1802 4029 1814 4032
rect 1756 4023 1814 4029
rect 3050 4020 3056 4032
rect 3108 4060 3114 4072
rect 3712 4060 3740 4091
rect 4798 4088 4804 4140
rect 4856 4128 4862 4140
rect 5353 4131 5411 4137
rect 5353 4128 5365 4131
rect 4856 4100 5365 4128
rect 4856 4088 4862 4100
rect 5353 4097 5365 4100
rect 5399 4097 5411 4131
rect 5353 4091 5411 4097
rect 5442 4088 5448 4140
rect 5500 4128 5506 4140
rect 5994 4128 6000 4140
rect 5500 4100 5545 4128
rect 5955 4100 6000 4128
rect 5500 4088 5506 4100
rect 5994 4088 6000 4100
rect 6052 4088 6058 4140
rect 7650 4128 7656 4140
rect 6104 4100 7656 4128
rect 3108 4032 3740 4060
rect 5261 4063 5319 4069
rect 3108 4020 3114 4032
rect 5261 4029 5273 4063
rect 5307 4060 5319 4063
rect 5534 4060 5540 4072
rect 5307 4032 5540 4060
rect 5307 4029 5319 4032
rect 5261 4023 5319 4029
rect 5534 4020 5540 4032
rect 5592 4020 5598 4072
rect 1026 3952 1032 4004
rect 1084 3992 1090 4004
rect 2961 3995 3019 4001
rect 2961 3992 2973 3995
rect 1084 3964 2973 3992
rect 1084 3952 1090 3964
rect 2961 3961 2973 3964
rect 3007 3961 3019 3995
rect 3513 3995 3571 4001
rect 3513 3992 3525 3995
rect 2961 3955 3019 3961
rect 3160 3964 3525 3992
rect 2682 3884 2688 3936
rect 2740 3924 2746 3936
rect 3160 3924 3188 3964
rect 3513 3961 3525 3964
rect 3559 3961 3571 3995
rect 3513 3955 3571 3961
rect 3602 3952 3608 4004
rect 3660 3992 3666 4004
rect 3660 3964 5304 3992
rect 3660 3952 3666 3964
rect 4890 3924 4896 3936
rect 2740 3896 3188 3924
rect 4851 3896 4896 3924
rect 2740 3884 2746 3896
rect 4890 3884 4896 3896
rect 4948 3884 4954 3936
rect 5276 3924 5304 3964
rect 5350 3952 5356 4004
rect 5408 3992 5414 4004
rect 6104 3992 6132 4100
rect 7650 4088 7656 4100
rect 7708 4088 7714 4140
rect 7834 4128 7840 4140
rect 7795 4100 7840 4128
rect 7834 4088 7840 4100
rect 7892 4088 7898 4140
rect 6454 4020 6460 4072
rect 6512 4060 6518 4072
rect 7944 4060 7972 4236
rect 8570 4224 8576 4236
rect 8628 4224 8634 4276
rect 10134 4264 10140 4276
rect 9416 4236 10140 4264
rect 8386 4196 8392 4208
rect 8036 4168 8392 4196
rect 8036 4137 8064 4168
rect 8386 4156 8392 4168
rect 8444 4156 8450 4208
rect 8021 4131 8079 4137
rect 8021 4097 8033 4131
rect 8067 4097 8079 4131
rect 8021 4091 8079 4097
rect 6512 4032 7972 4060
rect 8389 4063 8447 4069
rect 6512 4020 6518 4032
rect 8389 4029 8401 4063
rect 8435 4060 8447 4063
rect 8478 4060 8484 4072
rect 8435 4032 8484 4060
rect 8435 4029 8447 4032
rect 8389 4023 8447 4029
rect 8478 4020 8484 4032
rect 8536 4060 8542 4072
rect 9416 4060 9444 4236
rect 10134 4224 10140 4236
rect 10192 4224 10198 4276
rect 11238 4224 11244 4276
rect 11296 4264 11302 4276
rect 17954 4264 17960 4276
rect 11296 4236 17960 4264
rect 11296 4224 11302 4236
rect 17954 4224 17960 4236
rect 18012 4224 18018 4276
rect 19337 4267 19395 4273
rect 19337 4233 19349 4267
rect 19383 4264 19395 4267
rect 20622 4264 20628 4276
rect 19383 4236 20628 4264
rect 19383 4233 19395 4236
rect 19337 4227 19395 4233
rect 20622 4224 20628 4236
rect 20680 4224 20686 4276
rect 13262 4196 13268 4208
rect 8536 4032 9444 4060
rect 9508 4168 13268 4196
rect 8536 4020 8542 4032
rect 5408 3964 6132 3992
rect 8656 3995 8714 4001
rect 5408 3952 5414 3964
rect 8656 3961 8668 3995
rect 8702 3992 8714 3995
rect 8846 3992 8852 4004
rect 8702 3964 8852 3992
rect 8702 3961 8714 3964
rect 8656 3955 8714 3961
rect 8846 3952 8852 3964
rect 8904 3952 8910 4004
rect 7282 3924 7288 3936
rect 5276 3896 7288 3924
rect 7282 3884 7288 3896
rect 7340 3884 7346 3936
rect 7377 3927 7435 3933
rect 7377 3893 7389 3927
rect 7423 3924 7435 3927
rect 7650 3924 7656 3936
rect 7423 3896 7656 3924
rect 7423 3893 7435 3896
rect 7377 3887 7435 3893
rect 7650 3884 7656 3896
rect 7708 3884 7714 3936
rect 7745 3927 7803 3933
rect 7745 3893 7757 3927
rect 7791 3924 7803 3927
rect 8202 3924 8208 3936
rect 7791 3896 8208 3924
rect 7791 3893 7803 3896
rect 7745 3887 7803 3893
rect 8202 3884 8208 3896
rect 8260 3884 8266 3936
rect 8754 3884 8760 3936
rect 8812 3924 8818 3936
rect 9508 3924 9536 4168
rect 13262 4156 13268 4168
rect 13320 4156 13326 4208
rect 14921 4199 14979 4205
rect 14921 4165 14933 4199
rect 14967 4165 14979 4199
rect 14921 4159 14979 4165
rect 12434 4088 12440 4140
rect 12492 4128 12498 4140
rect 13541 4131 13599 4137
rect 13541 4128 13553 4131
rect 12492 4100 13553 4128
rect 12492 4088 12498 4100
rect 13541 4097 13553 4100
rect 13587 4097 13599 4131
rect 14936 4128 14964 4159
rect 15562 4128 15568 4140
rect 14936 4100 15568 4128
rect 13541 4091 13599 4097
rect 15562 4088 15568 4100
rect 15620 4128 15626 4140
rect 15841 4131 15899 4137
rect 15841 4128 15853 4131
rect 15620 4100 15853 4128
rect 15620 4088 15626 4100
rect 15841 4097 15853 4100
rect 15887 4128 15899 4131
rect 16761 4131 16819 4137
rect 16761 4128 16773 4131
rect 15887 4100 16773 4128
rect 15887 4097 15899 4100
rect 15841 4091 15899 4097
rect 16761 4097 16773 4100
rect 16807 4097 16819 4131
rect 16761 4091 16819 4097
rect 18969 4131 19027 4137
rect 18969 4097 18981 4131
rect 19015 4128 19027 4131
rect 19242 4128 19248 4140
rect 19015 4100 19248 4128
rect 19015 4097 19027 4100
rect 18969 4091 19027 4097
rect 19242 4088 19248 4100
rect 19300 4088 19306 4140
rect 19334 4088 19340 4140
rect 19392 4128 19398 4140
rect 19613 4131 19671 4137
rect 19613 4128 19625 4131
rect 19392 4100 19625 4128
rect 19392 4088 19398 4100
rect 19613 4097 19625 4100
rect 19659 4097 19671 4131
rect 19613 4091 19671 4097
rect 13808 4063 13866 4069
rect 13808 4029 13820 4063
rect 13854 4060 13866 4063
rect 14274 4060 14280 4072
rect 13854 4032 14280 4060
rect 13854 4029 13866 4032
rect 13808 4023 13866 4029
rect 14274 4020 14280 4032
rect 14332 4020 14338 4072
rect 15657 4063 15715 4069
rect 15657 4029 15669 4063
rect 15703 4060 15715 4063
rect 16390 4060 16396 4072
rect 15703 4032 16396 4060
rect 15703 4029 15715 4032
rect 15657 4023 15715 4029
rect 16390 4020 16396 4032
rect 16448 4020 16454 4072
rect 19886 4069 19892 4072
rect 16669 4063 16727 4069
rect 16669 4060 16681 4063
rect 16500 4032 16681 4060
rect 16022 3952 16028 4004
rect 16080 3992 16086 4004
rect 16500 3992 16528 4032
rect 16669 4029 16681 4032
rect 16715 4029 16727 4063
rect 19880 4060 19892 4069
rect 19847 4032 19892 4060
rect 16669 4023 16727 4029
rect 19880 4023 19892 4032
rect 19886 4020 19892 4023
rect 19944 4020 19950 4072
rect 16080 3964 16528 3992
rect 16577 3995 16635 4001
rect 16080 3952 16086 3964
rect 16577 3961 16589 3995
rect 16623 3992 16635 3995
rect 17221 3995 17279 4001
rect 17221 3992 17233 3995
rect 16623 3964 17233 3992
rect 16623 3961 16635 3964
rect 16577 3955 16635 3961
rect 17221 3961 17233 3964
rect 17267 3961 17279 3995
rect 17221 3955 17279 3961
rect 18601 3995 18659 4001
rect 18601 3961 18613 3995
rect 18647 3992 18659 3995
rect 20714 3992 20720 4004
rect 18647 3964 20720 3992
rect 18647 3961 18659 3964
rect 18601 3955 18659 3961
rect 20714 3952 20720 3964
rect 20772 3952 20778 4004
rect 9766 3924 9772 3936
rect 8812 3896 9536 3924
rect 9727 3896 9772 3924
rect 8812 3884 8818 3896
rect 9766 3884 9772 3896
rect 9824 3884 9830 3936
rect 15194 3924 15200 3936
rect 15155 3896 15200 3924
rect 15194 3884 15200 3896
rect 15252 3884 15258 3936
rect 15470 3884 15476 3936
rect 15528 3924 15534 3936
rect 15565 3927 15623 3933
rect 15565 3924 15577 3927
rect 15528 3896 15577 3924
rect 15528 3884 15534 3896
rect 15565 3893 15577 3896
rect 15611 3893 15623 3927
rect 15565 3887 15623 3893
rect 15838 3884 15844 3936
rect 15896 3924 15902 3936
rect 16209 3927 16267 3933
rect 16209 3924 16221 3927
rect 15896 3896 16221 3924
rect 15896 3884 15902 3896
rect 16209 3893 16221 3896
rect 16255 3893 16267 3927
rect 16209 3887 16267 3893
rect 16298 3884 16304 3936
rect 16356 3924 16362 3936
rect 20993 3927 21051 3933
rect 20993 3924 21005 3927
rect 16356 3896 21005 3924
rect 16356 3884 16362 3896
rect 20993 3893 21005 3896
rect 21039 3893 21051 3927
rect 20993 3887 21051 3893
rect 21361 3927 21419 3933
rect 21361 3893 21373 3927
rect 21407 3924 21419 3927
rect 21818 3924 21824 3936
rect 21407 3896 21824 3924
rect 21407 3893 21419 3896
rect 21361 3887 21419 3893
rect 21818 3884 21824 3896
rect 21876 3884 21882 3936
rect 1104 3834 21896 3856
rect 1104 3782 7912 3834
rect 7964 3782 7976 3834
rect 8028 3782 8040 3834
rect 8092 3782 8104 3834
rect 8156 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 15035 3834
rect 15087 3782 21896 3834
rect 1104 3760 21896 3782
rect 3050 3720 3056 3732
rect 3011 3692 3056 3720
rect 3050 3680 3056 3692
rect 3108 3680 3114 3732
rect 5258 3720 5264 3732
rect 5219 3692 5264 3720
rect 5258 3680 5264 3692
rect 5316 3680 5322 3732
rect 5721 3723 5779 3729
rect 5721 3689 5733 3723
rect 5767 3720 5779 3723
rect 5902 3720 5908 3732
rect 5767 3692 5908 3720
rect 5767 3689 5779 3692
rect 5721 3683 5779 3689
rect 5902 3680 5908 3692
rect 5960 3680 5966 3732
rect 8202 3720 8208 3732
rect 8163 3692 8208 3720
rect 8202 3680 8208 3692
rect 8260 3680 8266 3732
rect 8573 3723 8631 3729
rect 8573 3689 8585 3723
rect 8619 3720 8631 3723
rect 8938 3720 8944 3732
rect 8619 3692 8944 3720
rect 8619 3689 8631 3692
rect 8573 3683 8631 3689
rect 8938 3680 8944 3692
rect 8996 3680 9002 3732
rect 9490 3680 9496 3732
rect 9548 3720 9554 3732
rect 10689 3723 10747 3729
rect 10689 3720 10701 3723
rect 9548 3692 10701 3720
rect 9548 3680 9554 3692
rect 10689 3689 10701 3692
rect 10735 3720 10747 3723
rect 11238 3720 11244 3732
rect 10735 3692 11244 3720
rect 10735 3689 10747 3692
rect 10689 3683 10747 3689
rect 11238 3680 11244 3692
rect 11296 3680 11302 3732
rect 16298 3720 16304 3732
rect 11532 3692 16304 3720
rect 566 3612 572 3664
rect 624 3652 630 3664
rect 5534 3652 5540 3664
rect 624 3624 5540 3652
rect 624 3612 630 3624
rect 5534 3612 5540 3624
rect 5592 3612 5598 3664
rect 5629 3655 5687 3661
rect 5629 3621 5641 3655
rect 5675 3652 5687 3655
rect 5810 3652 5816 3664
rect 5675 3624 5816 3652
rect 5675 3621 5687 3624
rect 5629 3615 5687 3621
rect 5810 3612 5816 3624
rect 5868 3612 5874 3664
rect 9217 3655 9275 3661
rect 9217 3652 9229 3655
rect 6472 3624 9229 3652
rect 1486 3544 1492 3596
rect 1544 3584 1550 3596
rect 1673 3587 1731 3593
rect 1673 3584 1685 3587
rect 1544 3556 1685 3584
rect 1544 3544 1550 3556
rect 1673 3553 1685 3556
rect 1719 3584 1731 3587
rect 1762 3584 1768 3596
rect 1719 3556 1768 3584
rect 1719 3553 1731 3556
rect 1673 3547 1731 3553
rect 1762 3544 1768 3556
rect 1820 3544 1826 3596
rect 1946 3593 1952 3596
rect 1929 3587 1952 3593
rect 1929 3553 1941 3587
rect 1929 3547 1952 3553
rect 1946 3544 1952 3547
rect 2004 3544 2010 3596
rect 4062 3544 4068 3596
rect 4120 3584 4126 3596
rect 6365 3587 6423 3593
rect 6365 3584 6377 3587
rect 4120 3556 6377 3584
rect 4120 3544 4126 3556
rect 6365 3553 6377 3556
rect 6411 3553 6423 3587
rect 6365 3547 6423 3553
rect 5442 3476 5448 3528
rect 5500 3516 5506 3528
rect 5813 3519 5871 3525
rect 5813 3516 5825 3519
rect 5500 3488 5825 3516
rect 5500 3476 5506 3488
rect 5813 3485 5825 3488
rect 5859 3485 5871 3519
rect 6472 3516 6500 3624
rect 9217 3621 9229 3624
rect 9263 3652 9275 3655
rect 10502 3652 10508 3664
rect 9263 3624 10508 3652
rect 9263 3621 9275 3624
rect 9217 3615 9275 3621
rect 10502 3612 10508 3624
rect 10560 3612 10566 3664
rect 6632 3587 6690 3593
rect 6632 3553 6644 3587
rect 6678 3584 6690 3587
rect 9490 3584 9496 3596
rect 6678 3556 9496 3584
rect 6678 3553 6690 3556
rect 6632 3547 6690 3553
rect 9490 3544 9496 3556
rect 9548 3544 9554 3596
rect 9950 3584 9956 3596
rect 9911 3556 9956 3584
rect 9950 3544 9956 3556
rect 10008 3584 10014 3596
rect 10597 3587 10655 3593
rect 10597 3584 10609 3587
rect 10008 3556 10609 3584
rect 10008 3544 10014 3556
rect 10597 3553 10609 3556
rect 10643 3553 10655 3587
rect 10597 3547 10655 3553
rect 5813 3479 5871 3485
rect 6380 3488 6500 3516
rect 2774 3408 2780 3460
rect 2832 3448 2838 3460
rect 2958 3448 2964 3460
rect 2832 3420 2964 3448
rect 2832 3408 2838 3420
rect 2958 3408 2964 3420
rect 3016 3408 3022 3460
rect 6380 3448 6408 3488
rect 7742 3476 7748 3528
rect 7800 3516 7806 3528
rect 8665 3519 8723 3525
rect 8665 3516 8677 3519
rect 7800 3488 8677 3516
rect 7800 3476 7806 3488
rect 8665 3485 8677 3488
rect 8711 3516 8723 3519
rect 8754 3516 8760 3528
rect 8711 3488 8760 3516
rect 8711 3485 8723 3488
rect 8665 3479 8723 3485
rect 8754 3476 8760 3488
rect 8812 3476 8818 3528
rect 8846 3476 8852 3528
rect 8904 3516 8910 3528
rect 10778 3516 10784 3528
rect 8904 3488 10784 3516
rect 8904 3476 8910 3488
rect 10778 3476 10784 3488
rect 10836 3516 10842 3528
rect 10873 3519 10931 3525
rect 10873 3516 10885 3519
rect 10836 3488 10885 3516
rect 10836 3476 10842 3488
rect 10873 3485 10885 3488
rect 10919 3516 10931 3519
rect 11532 3516 11560 3692
rect 16298 3680 16304 3692
rect 16356 3680 16362 3732
rect 16482 3680 16488 3732
rect 16540 3720 16546 3732
rect 16669 3723 16727 3729
rect 16669 3720 16681 3723
rect 16540 3692 16681 3720
rect 16540 3680 16546 3692
rect 16669 3689 16681 3692
rect 16715 3689 16727 3723
rect 16669 3683 16727 3689
rect 19794 3680 19800 3732
rect 19852 3720 19858 3732
rect 20530 3720 20536 3732
rect 19852 3692 20536 3720
rect 19852 3680 19858 3692
rect 20530 3680 20536 3692
rect 20588 3680 20594 3732
rect 15562 3661 15568 3664
rect 15556 3652 15568 3661
rect 15523 3624 15568 3652
rect 15556 3615 15568 3624
rect 15562 3612 15568 3615
rect 15620 3612 15626 3664
rect 11698 3584 11704 3596
rect 11659 3556 11704 3584
rect 11698 3544 11704 3556
rect 11756 3544 11762 3596
rect 12437 3587 12495 3593
rect 12437 3584 12449 3587
rect 11808 3556 12449 3584
rect 10919 3488 11560 3516
rect 10919 3485 10931 3488
rect 10873 3479 10931 3485
rect 3344 3420 6408 3448
rect 1946 3340 1952 3392
rect 2004 3380 2010 3392
rect 2682 3380 2688 3392
rect 2004 3352 2688 3380
rect 2004 3340 2010 3352
rect 2682 3340 2688 3352
rect 2740 3380 2746 3392
rect 3344 3389 3372 3420
rect 7374 3408 7380 3460
rect 7432 3448 7438 3460
rect 7432 3420 7880 3448
rect 7432 3408 7438 3420
rect 3329 3383 3387 3389
rect 3329 3380 3341 3383
rect 2740 3352 3341 3380
rect 2740 3340 2746 3352
rect 3329 3349 3341 3352
rect 3375 3349 3387 3383
rect 3329 3343 3387 3349
rect 3786 3340 3792 3392
rect 3844 3380 3850 3392
rect 6086 3380 6092 3392
rect 3844 3352 6092 3380
rect 3844 3340 3850 3352
rect 6086 3340 6092 3352
rect 6144 3340 6150 3392
rect 6730 3340 6736 3392
rect 6788 3380 6794 3392
rect 7745 3383 7803 3389
rect 7745 3380 7757 3383
rect 6788 3352 7757 3380
rect 6788 3340 6794 3352
rect 7745 3349 7757 3352
rect 7791 3349 7803 3383
rect 7852 3380 7880 3420
rect 8110 3408 8116 3460
rect 8168 3448 8174 3460
rect 8478 3448 8484 3460
rect 8168 3420 8484 3448
rect 8168 3408 8174 3420
rect 8478 3408 8484 3420
rect 8536 3408 8542 3460
rect 10318 3408 10324 3460
rect 10376 3448 10382 3460
rect 11808 3448 11836 3556
rect 12437 3553 12449 3556
rect 12483 3553 12495 3587
rect 12437 3547 12495 3553
rect 12802 3544 12808 3596
rect 12860 3584 12866 3596
rect 13173 3587 13231 3593
rect 13173 3584 13185 3587
rect 12860 3556 13185 3584
rect 12860 3544 12866 3556
rect 13173 3553 13185 3556
rect 13219 3553 13231 3587
rect 13173 3547 13231 3553
rect 13446 3544 13452 3596
rect 13504 3584 13510 3596
rect 13725 3587 13783 3593
rect 13725 3584 13737 3587
rect 13504 3556 13737 3584
rect 13504 3544 13510 3556
rect 13725 3553 13737 3556
rect 13771 3553 13783 3587
rect 15286 3584 15292 3596
rect 15247 3556 15292 3584
rect 13725 3547 13783 3553
rect 15286 3544 15292 3556
rect 15344 3544 15350 3596
rect 16574 3544 16580 3596
rect 16632 3584 16638 3596
rect 17129 3587 17187 3593
rect 17129 3584 17141 3587
rect 16632 3556 17141 3584
rect 16632 3544 16638 3556
rect 17129 3553 17141 3556
rect 17175 3553 17187 3587
rect 17129 3547 17187 3553
rect 18049 3587 18107 3593
rect 18049 3553 18061 3587
rect 18095 3584 18107 3587
rect 18138 3584 18144 3596
rect 18095 3556 18144 3584
rect 18095 3553 18107 3556
rect 18049 3547 18107 3553
rect 18138 3544 18144 3556
rect 18196 3544 18202 3596
rect 18874 3584 18880 3596
rect 18835 3556 18880 3584
rect 18874 3544 18880 3556
rect 18932 3544 18938 3596
rect 19242 3544 19248 3596
rect 19300 3584 19306 3596
rect 19889 3587 19947 3593
rect 19889 3584 19901 3587
rect 19300 3556 19901 3584
rect 19300 3544 19306 3556
rect 19889 3553 19901 3556
rect 19935 3553 19947 3587
rect 19889 3547 19947 3553
rect 20901 3587 20959 3593
rect 20901 3553 20913 3587
rect 20947 3584 20959 3587
rect 21818 3584 21824 3596
rect 20947 3556 21824 3584
rect 20947 3553 20959 3556
rect 20901 3547 20959 3553
rect 21818 3544 21824 3556
rect 21876 3544 21882 3596
rect 11977 3519 12035 3525
rect 11977 3485 11989 3519
rect 12023 3485 12035 3519
rect 11977 3479 12035 3485
rect 12713 3519 12771 3525
rect 12713 3485 12725 3519
rect 12759 3516 12771 3519
rect 13354 3516 13360 3528
rect 12759 3488 13360 3516
rect 12759 3485 12771 3488
rect 12713 3479 12771 3485
rect 10376 3420 11836 3448
rect 10376 3408 10382 3420
rect 9674 3380 9680 3392
rect 7852 3352 9680 3380
rect 7745 3343 7803 3349
rect 9674 3340 9680 3352
rect 9732 3340 9738 3392
rect 10134 3340 10140 3392
rect 10192 3380 10198 3392
rect 10229 3383 10287 3389
rect 10229 3380 10241 3383
rect 10192 3352 10241 3380
rect 10192 3340 10198 3352
rect 10229 3349 10241 3352
rect 10275 3349 10287 3383
rect 11992 3380 12020 3479
rect 13354 3476 13360 3488
rect 13412 3476 13418 3528
rect 17218 3476 17224 3528
rect 17276 3516 17282 3528
rect 17313 3519 17371 3525
rect 17313 3516 17325 3519
rect 17276 3488 17325 3516
rect 17276 3476 17282 3488
rect 17313 3485 17325 3488
rect 17359 3485 17371 3519
rect 17313 3479 17371 3485
rect 19153 3519 19211 3525
rect 19153 3485 19165 3519
rect 19199 3516 19211 3519
rect 19518 3516 19524 3528
rect 19199 3488 19524 3516
rect 19199 3485 19211 3488
rect 19153 3479 19211 3485
rect 19518 3476 19524 3488
rect 19576 3476 19582 3528
rect 13262 3380 13268 3392
rect 11992 3352 13268 3380
rect 10229 3343 10287 3349
rect 13262 3340 13268 3352
rect 13320 3340 13326 3392
rect 13357 3383 13415 3389
rect 13357 3349 13369 3383
rect 13403 3380 13415 3383
rect 13722 3380 13728 3392
rect 13403 3352 13728 3380
rect 13403 3349 13415 3352
rect 13357 3343 13415 3349
rect 13722 3340 13728 3352
rect 13780 3340 13786 3392
rect 13909 3383 13967 3389
rect 13909 3349 13921 3383
rect 13955 3380 13967 3383
rect 14550 3380 14556 3392
rect 13955 3352 14556 3380
rect 13955 3349 13967 3352
rect 13909 3343 13967 3349
rect 14550 3340 14556 3352
rect 14608 3340 14614 3392
rect 17770 3340 17776 3392
rect 17828 3380 17834 3392
rect 18233 3383 18291 3389
rect 18233 3380 18245 3383
rect 17828 3352 18245 3380
rect 17828 3340 17834 3352
rect 18233 3349 18245 3352
rect 18279 3349 18291 3383
rect 18233 3343 18291 3349
rect 19610 3340 19616 3392
rect 19668 3380 19674 3392
rect 20073 3383 20131 3389
rect 20073 3380 20085 3383
rect 19668 3352 20085 3380
rect 19668 3340 19674 3352
rect 20073 3349 20085 3352
rect 20119 3349 20131 3383
rect 20073 3343 20131 3349
rect 21085 3383 21143 3389
rect 21085 3349 21097 3383
rect 21131 3380 21143 3383
rect 22278 3380 22284 3392
rect 21131 3352 22284 3380
rect 21131 3349 21143 3352
rect 21085 3343 21143 3349
rect 22278 3340 22284 3352
rect 22336 3340 22342 3392
rect 1104 3290 21896 3312
rect 1104 3238 4447 3290
rect 4499 3238 4511 3290
rect 4563 3238 4575 3290
rect 4627 3238 4639 3290
rect 4691 3238 11378 3290
rect 11430 3238 11442 3290
rect 11494 3238 11506 3290
rect 11558 3238 11570 3290
rect 11622 3238 18308 3290
rect 18360 3238 18372 3290
rect 18424 3238 18436 3290
rect 18488 3238 18500 3290
rect 18552 3238 21896 3290
rect 1104 3216 21896 3238
rect 3510 3136 3516 3188
rect 3568 3176 3574 3188
rect 5442 3176 5448 3188
rect 3568 3148 5448 3176
rect 3568 3136 3574 3148
rect 5442 3136 5448 3148
rect 5500 3176 5506 3188
rect 5813 3179 5871 3185
rect 5813 3176 5825 3179
rect 5500 3148 5825 3176
rect 5500 3136 5506 3148
rect 5813 3145 5825 3148
rect 5859 3145 5871 3179
rect 9490 3176 9496 3188
rect 5813 3139 5871 3145
rect 6932 3148 9076 3176
rect 9451 3148 9496 3176
rect 4154 3108 4160 3120
rect 4115 3080 4160 3108
rect 4154 3068 4160 3080
rect 4212 3068 4218 3120
rect 5534 3068 5540 3120
rect 5592 3108 5598 3120
rect 6638 3108 6644 3120
rect 5592 3080 6644 3108
rect 5592 3068 5598 3080
rect 6638 3068 6644 3080
rect 6696 3068 6702 3120
rect 4062 3000 4068 3052
rect 4120 3040 4126 3052
rect 4433 3043 4491 3049
rect 4433 3040 4445 3043
rect 4120 3012 4445 3040
rect 4120 3000 4126 3012
rect 4433 3009 4445 3012
rect 4479 3009 4491 3043
rect 4433 3003 4491 3009
rect 1762 2932 1768 2984
rect 1820 2972 1826 2984
rect 2777 2975 2835 2981
rect 2777 2972 2789 2975
rect 1820 2944 2789 2972
rect 1820 2932 1826 2944
rect 2777 2941 2789 2944
rect 2823 2972 2835 2975
rect 4080 2972 4108 3000
rect 2823 2944 4108 2972
rect 4700 2975 4758 2981
rect 2823 2941 2835 2944
rect 2777 2935 2835 2941
rect 4700 2941 4712 2975
rect 4746 2972 4758 2975
rect 5718 2972 5724 2984
rect 4746 2944 5724 2972
rect 4746 2941 4758 2944
rect 4700 2935 4758 2941
rect 5718 2932 5724 2944
rect 5776 2972 5782 2984
rect 5902 2972 5908 2984
rect 5776 2944 5908 2972
rect 5776 2932 5782 2944
rect 5902 2932 5908 2944
rect 5960 2932 5966 2984
rect 6181 2975 6239 2981
rect 6181 2941 6193 2975
rect 6227 2972 6239 2975
rect 6270 2972 6276 2984
rect 6227 2944 6276 2972
rect 6227 2941 6239 2944
rect 6181 2935 6239 2941
rect 6270 2932 6276 2944
rect 6328 2932 6334 2984
rect 6822 2972 6828 2984
rect 6783 2944 6828 2972
rect 6822 2932 6828 2944
rect 6880 2932 6886 2984
rect 3044 2907 3102 2913
rect 3044 2873 3056 2907
rect 3090 2904 3102 2907
rect 3510 2904 3516 2916
rect 3090 2876 3516 2904
rect 3090 2873 3102 2876
rect 3044 2867 3102 2873
rect 3510 2864 3516 2876
rect 3568 2864 3574 2916
rect 6932 2904 6960 3148
rect 7742 3108 7748 3120
rect 7703 3080 7748 3108
rect 7742 3068 7748 3080
rect 7800 3068 7806 3120
rect 9048 3108 9076 3148
rect 9490 3136 9496 3148
rect 9548 3136 9554 3188
rect 19058 3176 19064 3188
rect 9600 3148 19064 3176
rect 9600 3108 9628 3148
rect 19058 3136 19064 3148
rect 19116 3136 19122 3188
rect 9048 3080 9628 3108
rect 13081 3111 13139 3117
rect 13081 3077 13093 3111
rect 13127 3108 13139 3111
rect 15470 3108 15476 3120
rect 13127 3080 15476 3108
rect 13127 3077 13139 3080
rect 13081 3071 13139 3077
rect 15470 3068 15476 3080
rect 15528 3068 15534 3120
rect 16482 3108 16488 3120
rect 16132 3080 16488 3108
rect 8110 3040 8116 3052
rect 8071 3012 8116 3040
rect 8110 3000 8116 3012
rect 8168 3000 8174 3052
rect 9674 3000 9680 3052
rect 9732 3040 9738 3052
rect 9953 3043 10011 3049
rect 9953 3040 9965 3043
rect 9732 3012 9965 3040
rect 9732 3000 9738 3012
rect 9953 3009 9965 3012
rect 9999 3040 10011 3043
rect 10686 3040 10692 3052
rect 9999 3012 10692 3040
rect 9999 3009 10011 3012
rect 9953 3003 10011 3009
rect 10686 3000 10692 3012
rect 10744 3000 10750 3052
rect 10778 3000 10784 3052
rect 10836 3040 10842 3052
rect 10836 3012 10881 3040
rect 10980 3012 13216 3040
rect 10836 3000 10842 3012
rect 7101 2975 7159 2981
rect 7101 2941 7113 2975
rect 7147 2972 7159 2975
rect 10980 2972 11008 3012
rect 7147 2944 11008 2972
rect 11241 2975 11299 2981
rect 7147 2941 7159 2944
rect 7101 2935 7159 2941
rect 11241 2941 11253 2975
rect 11287 2941 11299 2975
rect 11241 2935 11299 2941
rect 8386 2913 8392 2916
rect 5828 2876 6960 2904
rect 3878 2796 3884 2848
rect 3936 2836 3942 2848
rect 5828 2836 5856 2876
rect 8380 2867 8392 2913
rect 8444 2904 8450 2916
rect 8444 2876 9628 2904
rect 8386 2864 8392 2867
rect 8444 2864 8450 2876
rect 3936 2808 5856 2836
rect 9600 2836 9628 2876
rect 9674 2864 9680 2916
rect 9732 2904 9738 2916
rect 11256 2904 11284 2935
rect 11882 2932 11888 2984
rect 11940 2972 11946 2984
rect 13188 2981 13216 3012
rect 13262 3000 13268 3052
rect 13320 3040 13326 3052
rect 13320 3012 14688 3040
rect 13320 3000 13326 3012
rect 12437 2975 12495 2981
rect 12437 2972 12449 2975
rect 11940 2944 12449 2972
rect 11940 2932 11946 2944
rect 12437 2941 12449 2944
rect 12483 2941 12495 2975
rect 12437 2935 12495 2941
rect 13173 2975 13231 2981
rect 13173 2941 13185 2975
rect 13219 2941 13231 2975
rect 13906 2972 13912 2984
rect 13867 2944 13912 2972
rect 13173 2935 13231 2941
rect 13906 2932 13912 2944
rect 13964 2932 13970 2984
rect 14660 2981 14688 3012
rect 15194 3000 15200 3052
rect 15252 3040 15258 3052
rect 16132 3049 16160 3080
rect 16482 3068 16488 3080
rect 16540 3068 16546 3120
rect 15933 3043 15991 3049
rect 15933 3040 15945 3043
rect 15252 3012 15945 3040
rect 15252 3000 15258 3012
rect 15933 3009 15945 3012
rect 15979 3009 15991 3043
rect 15933 3003 15991 3009
rect 16117 3043 16175 3049
rect 16117 3009 16129 3043
rect 16163 3009 16175 3043
rect 16117 3003 16175 3009
rect 18138 3000 18144 3052
rect 18196 3040 18202 3052
rect 18233 3043 18291 3049
rect 18233 3040 18245 3043
rect 18196 3012 18245 3040
rect 18196 3000 18202 3012
rect 18233 3009 18245 3012
rect 18279 3009 18291 3043
rect 19426 3040 19432 3052
rect 18233 3003 18291 3009
rect 18800 3012 19432 3040
rect 14645 2975 14703 2981
rect 14645 2941 14657 2975
rect 14691 2941 14703 2975
rect 16485 2975 16543 2981
rect 16485 2972 16497 2975
rect 14645 2935 14703 2941
rect 15488 2944 16497 2972
rect 9732 2876 11284 2904
rect 11517 2907 11575 2913
rect 9732 2864 9738 2876
rect 11517 2873 11529 2907
rect 11563 2904 11575 2907
rect 11790 2904 11796 2916
rect 11563 2876 11796 2904
rect 11563 2873 11575 2876
rect 11517 2867 11575 2873
rect 11790 2864 11796 2876
rect 11848 2864 11854 2916
rect 12713 2907 12771 2913
rect 12713 2873 12725 2907
rect 12759 2904 12771 2907
rect 13814 2904 13820 2916
rect 12759 2876 13820 2904
rect 12759 2873 12771 2876
rect 12713 2867 12771 2873
rect 13814 2864 13820 2876
rect 13872 2864 13878 2916
rect 14185 2907 14243 2913
rect 14185 2873 14197 2907
rect 14231 2904 14243 2907
rect 14734 2904 14740 2916
rect 14231 2876 14740 2904
rect 14231 2873 14243 2876
rect 14185 2867 14243 2873
rect 14734 2864 14740 2876
rect 14792 2864 14798 2916
rect 9766 2836 9772 2848
rect 9600 2808 9772 2836
rect 3936 2796 3942 2808
rect 9766 2796 9772 2808
rect 9824 2796 9830 2848
rect 10226 2836 10232 2848
rect 10187 2808 10232 2836
rect 10226 2796 10232 2808
rect 10284 2796 10290 2848
rect 10502 2796 10508 2848
rect 10560 2836 10566 2848
rect 10597 2839 10655 2845
rect 10597 2836 10609 2839
rect 10560 2808 10609 2836
rect 10560 2796 10566 2808
rect 10597 2805 10609 2808
rect 10643 2836 10655 2839
rect 13081 2839 13139 2845
rect 13081 2836 13093 2839
rect 10643 2808 13093 2836
rect 10643 2805 10655 2808
rect 10597 2799 10655 2805
rect 13081 2805 13093 2808
rect 13127 2805 13139 2839
rect 13081 2799 13139 2805
rect 13262 2796 13268 2848
rect 13320 2836 13326 2848
rect 13357 2839 13415 2845
rect 13357 2836 13369 2839
rect 13320 2808 13369 2836
rect 13320 2796 13326 2808
rect 13357 2805 13369 2808
rect 13403 2805 13415 2839
rect 13357 2799 13415 2805
rect 14829 2839 14887 2845
rect 14829 2805 14841 2839
rect 14875 2836 14887 2839
rect 15378 2836 15384 2848
rect 14875 2808 15384 2836
rect 14875 2805 14887 2808
rect 14829 2799 14887 2805
rect 15378 2796 15384 2808
rect 15436 2796 15442 2848
rect 15488 2845 15516 2944
rect 16485 2941 16497 2944
rect 16531 2941 16543 2975
rect 16485 2935 16543 2941
rect 17034 2932 17040 2984
rect 17092 2972 17098 2984
rect 17221 2975 17279 2981
rect 17221 2972 17233 2975
rect 17092 2944 17233 2972
rect 17092 2932 17098 2944
rect 17221 2941 17233 2944
rect 17267 2941 17279 2975
rect 18046 2972 18052 2984
rect 18007 2944 18052 2972
rect 17221 2935 17279 2941
rect 18046 2932 18052 2944
rect 18104 2932 18110 2984
rect 18800 2981 18828 3012
rect 19426 3000 19432 3012
rect 19484 3000 19490 3052
rect 20806 3040 20812 3052
rect 20767 3012 20812 3040
rect 20806 3000 20812 3012
rect 20864 3000 20870 3052
rect 18785 2975 18843 2981
rect 18785 2941 18797 2975
rect 18831 2941 18843 2975
rect 19518 2972 19524 2984
rect 19479 2944 19524 2972
rect 18785 2935 18843 2941
rect 19518 2932 19524 2944
rect 19576 2932 19582 2984
rect 20349 2975 20407 2981
rect 20349 2941 20361 2975
rect 20395 2972 20407 2975
rect 20714 2972 20720 2984
rect 20395 2944 20720 2972
rect 20395 2941 20407 2944
rect 20349 2935 20407 2941
rect 20714 2932 20720 2944
rect 20772 2972 20778 2984
rect 22738 2972 22744 2984
rect 20772 2944 22744 2972
rect 20772 2932 20778 2944
rect 22738 2932 22744 2944
rect 22796 2932 22802 2984
rect 15838 2904 15844 2916
rect 15799 2876 15844 2904
rect 15838 2864 15844 2876
rect 15896 2864 15902 2916
rect 16574 2864 16580 2916
rect 16632 2904 16638 2916
rect 16761 2907 16819 2913
rect 16761 2904 16773 2907
rect 16632 2876 16773 2904
rect 16632 2864 16638 2876
rect 16761 2873 16773 2876
rect 16807 2873 16819 2907
rect 16761 2867 16819 2873
rect 16850 2864 16856 2916
rect 16908 2904 16914 2916
rect 17497 2907 17555 2913
rect 17497 2904 17509 2907
rect 16908 2876 17509 2904
rect 16908 2864 16914 2876
rect 17497 2873 17509 2876
rect 17543 2873 17555 2907
rect 17497 2867 17555 2873
rect 18506 2864 18512 2916
rect 18564 2904 18570 2916
rect 19061 2907 19119 2913
rect 19061 2904 19073 2907
rect 18564 2876 19073 2904
rect 18564 2864 18570 2876
rect 19061 2873 19073 2876
rect 19107 2873 19119 2907
rect 19061 2867 19119 2873
rect 15473 2839 15531 2845
rect 15473 2805 15485 2839
rect 15519 2805 15531 2839
rect 15473 2799 15531 2805
rect 18598 2796 18604 2848
rect 18656 2836 18662 2848
rect 19705 2839 19763 2845
rect 19705 2836 19717 2839
rect 18656 2808 19717 2836
rect 18656 2796 18662 2808
rect 19705 2805 19717 2808
rect 19751 2805 19763 2839
rect 19705 2799 19763 2805
rect 1104 2746 21896 2768
rect 1104 2694 7912 2746
rect 7964 2694 7976 2746
rect 8028 2694 8040 2746
rect 8092 2694 8104 2746
rect 8156 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 15035 2746
rect 15087 2694 21896 2746
rect 1104 2672 21896 2694
rect 4890 2592 4896 2644
rect 4948 2632 4954 2644
rect 5077 2635 5135 2641
rect 5077 2632 5089 2635
rect 4948 2604 5089 2632
rect 4948 2592 4954 2604
rect 5077 2601 5089 2604
rect 5123 2601 5135 2635
rect 5077 2595 5135 2601
rect 5169 2635 5227 2641
rect 5169 2601 5181 2635
rect 5215 2632 5227 2635
rect 5258 2632 5264 2644
rect 5215 2604 5264 2632
rect 5215 2601 5227 2604
rect 5169 2595 5227 2601
rect 5258 2592 5264 2604
rect 5316 2592 5322 2644
rect 5810 2592 5816 2644
rect 5868 2632 5874 2644
rect 5868 2604 5913 2632
rect 5868 2592 5874 2604
rect 7650 2592 7656 2644
rect 7708 2632 7714 2644
rect 9033 2635 9091 2641
rect 9033 2632 9045 2635
rect 7708 2604 9045 2632
rect 7708 2592 7714 2604
rect 9033 2601 9045 2604
rect 9079 2601 9091 2635
rect 9033 2595 9091 2601
rect 9125 2635 9183 2641
rect 9125 2601 9137 2635
rect 9171 2632 9183 2635
rect 9769 2635 9827 2641
rect 9769 2632 9781 2635
rect 9171 2604 9781 2632
rect 9171 2601 9183 2604
rect 9125 2595 9183 2601
rect 9769 2601 9781 2604
rect 9815 2601 9827 2635
rect 9769 2595 9827 2601
rect 10137 2635 10195 2641
rect 10137 2601 10149 2635
rect 10183 2632 10195 2635
rect 10226 2632 10232 2644
rect 10183 2604 10232 2632
rect 10183 2601 10195 2604
rect 10137 2595 10195 2601
rect 10226 2592 10232 2604
rect 10284 2592 10290 2644
rect 19058 2632 19064 2644
rect 19019 2604 19064 2632
rect 19058 2592 19064 2604
rect 19116 2592 19122 2644
rect 6181 2567 6239 2573
rect 6181 2564 6193 2567
rect 2976 2536 6193 2564
rect 2777 2499 2835 2505
rect 2777 2465 2789 2499
rect 2823 2496 2835 2499
rect 2866 2496 2872 2508
rect 2823 2468 2872 2496
rect 2823 2465 2835 2468
rect 2777 2459 2835 2465
rect 2866 2456 2872 2468
rect 2924 2456 2930 2508
rect 2406 2252 2412 2304
rect 2464 2292 2470 2304
rect 2976 2292 3004 2536
rect 6181 2533 6193 2536
rect 6227 2564 6239 2567
rect 6546 2564 6552 2576
rect 6227 2536 6552 2564
rect 6227 2533 6239 2536
rect 6181 2527 6239 2533
rect 6546 2524 6552 2536
rect 6604 2564 6610 2576
rect 6917 2567 6975 2573
rect 6917 2564 6929 2567
rect 6604 2536 6929 2564
rect 6604 2524 6610 2536
rect 6917 2533 6929 2536
rect 6963 2533 6975 2567
rect 12802 2564 12808 2576
rect 6917 2527 6975 2533
rect 7668 2536 12808 2564
rect 3053 2431 3111 2437
rect 3053 2397 3065 2431
rect 3099 2397 3111 2431
rect 3053 2391 3111 2397
rect 3068 2360 3096 2391
rect 4154 2388 4160 2440
rect 4212 2428 4218 2440
rect 5261 2431 5319 2437
rect 5261 2428 5273 2431
rect 4212 2400 5273 2428
rect 4212 2388 4218 2400
rect 5261 2397 5273 2400
rect 5307 2397 5319 2431
rect 6270 2428 6276 2440
rect 6231 2400 6276 2428
rect 5261 2391 5319 2397
rect 6270 2388 6276 2400
rect 6328 2388 6334 2440
rect 6457 2431 6515 2437
rect 6457 2397 6469 2431
rect 6503 2428 6515 2431
rect 6730 2428 6736 2440
rect 6503 2400 6736 2428
rect 6503 2397 6515 2400
rect 6457 2391 6515 2397
rect 6730 2388 6736 2400
rect 6788 2388 6794 2440
rect 7668 2360 7696 2536
rect 12802 2524 12808 2536
rect 12860 2524 12866 2576
rect 12897 2567 12955 2573
rect 12897 2533 12909 2567
rect 12943 2564 12955 2567
rect 13446 2564 13452 2576
rect 12943 2536 13452 2564
rect 12943 2533 12955 2536
rect 12897 2527 12955 2533
rect 13446 2524 13452 2536
rect 13504 2524 13510 2576
rect 19076 2564 19104 2592
rect 19076 2536 20024 2564
rect 10134 2456 10140 2508
rect 10192 2496 10198 2508
rect 10229 2499 10287 2505
rect 10229 2496 10241 2499
rect 10192 2468 10241 2496
rect 10192 2456 10198 2468
rect 10229 2465 10241 2468
rect 10275 2465 10287 2499
rect 11790 2496 11796 2508
rect 11751 2468 11796 2496
rect 10229 2459 10287 2465
rect 11790 2456 11796 2468
rect 11848 2456 11854 2508
rect 12618 2496 12624 2508
rect 12579 2468 12624 2496
rect 12618 2456 12624 2468
rect 12676 2456 12682 2508
rect 13354 2496 13360 2508
rect 13315 2468 13360 2496
rect 13354 2456 13360 2468
rect 13412 2456 13418 2508
rect 13814 2456 13820 2508
rect 13872 2496 13878 2508
rect 13909 2499 13967 2505
rect 13909 2496 13921 2499
rect 13872 2468 13921 2496
rect 13872 2456 13878 2468
rect 13909 2465 13921 2468
rect 13955 2465 13967 2499
rect 14734 2496 14740 2508
rect 14695 2468 14740 2496
rect 13909 2459 13967 2465
rect 14734 2456 14740 2468
rect 14792 2456 14798 2508
rect 16117 2499 16175 2505
rect 16117 2465 16129 2499
rect 16163 2496 16175 2499
rect 16574 2496 16580 2508
rect 16163 2468 16580 2496
rect 16163 2465 16175 2468
rect 16117 2459 16175 2465
rect 16574 2456 16580 2468
rect 16632 2456 16638 2508
rect 16669 2499 16727 2505
rect 16669 2465 16681 2499
rect 16715 2496 16727 2499
rect 16850 2496 16856 2508
rect 16715 2468 16856 2496
rect 16715 2465 16727 2468
rect 16669 2459 16727 2465
rect 16850 2456 16856 2468
rect 16908 2456 16914 2508
rect 17218 2496 17224 2508
rect 17179 2468 17224 2496
rect 17218 2456 17224 2468
rect 17276 2456 17282 2508
rect 18506 2496 18512 2508
rect 18467 2468 18512 2496
rect 18506 2456 18512 2468
rect 18564 2456 18570 2508
rect 19429 2499 19487 2505
rect 19429 2465 19441 2499
rect 19475 2496 19487 2499
rect 19794 2496 19800 2508
rect 19475 2468 19800 2496
rect 19475 2465 19487 2468
rect 19429 2459 19487 2465
rect 19794 2456 19800 2468
rect 19852 2456 19858 2508
rect 19996 2505 20024 2536
rect 19981 2499 20039 2505
rect 19981 2465 19993 2499
rect 20027 2465 20039 2499
rect 19981 2459 20039 2465
rect 20533 2499 20591 2505
rect 20533 2465 20545 2499
rect 20579 2496 20591 2499
rect 20622 2496 20628 2508
rect 20579 2468 20628 2496
rect 20579 2465 20591 2468
rect 20533 2459 20591 2465
rect 20622 2456 20628 2468
rect 20680 2496 20686 2508
rect 21177 2499 21235 2505
rect 21177 2496 21189 2499
rect 20680 2468 21189 2496
rect 20680 2456 20686 2468
rect 21177 2465 21189 2468
rect 21223 2465 21235 2499
rect 21177 2459 21235 2465
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2428 9367 2431
rect 9582 2428 9588 2440
rect 9355 2400 9588 2428
rect 9355 2397 9367 2400
rect 9309 2391 9367 2397
rect 9582 2388 9588 2400
rect 9640 2388 9646 2440
rect 9766 2388 9772 2440
rect 9824 2428 9830 2440
rect 10321 2431 10379 2437
rect 10321 2428 10333 2431
rect 9824 2400 10333 2428
rect 9824 2388 9830 2400
rect 10321 2397 10333 2400
rect 10367 2397 10379 2431
rect 10321 2391 10379 2397
rect 3068 2332 7696 2360
rect 8665 2363 8723 2369
rect 8665 2329 8677 2363
rect 8711 2360 8723 2363
rect 9674 2360 9680 2372
rect 8711 2332 9680 2360
rect 8711 2329 8723 2332
rect 8665 2323 8723 2329
rect 9674 2320 9680 2332
rect 9732 2320 9738 2372
rect 14093 2363 14151 2369
rect 14093 2329 14105 2363
rect 14139 2360 14151 2363
rect 15010 2360 15016 2372
rect 14139 2332 15016 2360
rect 14139 2329 14151 2332
rect 14093 2323 14151 2329
rect 15010 2320 15016 2332
rect 15068 2320 15074 2372
rect 20165 2363 20223 2369
rect 20165 2329 20177 2363
rect 20211 2360 20223 2363
rect 21358 2360 21364 2372
rect 20211 2332 21364 2360
rect 20211 2329 20223 2332
rect 20165 2323 20223 2329
rect 21358 2320 21364 2332
rect 21416 2320 21422 2372
rect 2464 2264 3004 2292
rect 4709 2295 4767 2301
rect 2464 2252 2470 2264
rect 4709 2261 4721 2295
rect 4755 2292 4767 2295
rect 6822 2292 6828 2304
rect 4755 2264 6828 2292
rect 4755 2261 4767 2264
rect 4709 2255 4767 2261
rect 6822 2252 6828 2264
rect 6880 2252 6886 2304
rect 11977 2295 12035 2301
rect 11977 2261 11989 2295
rect 12023 2292 12035 2295
rect 12802 2292 12808 2304
rect 12023 2264 12808 2292
rect 12023 2261 12035 2264
rect 11977 2255 12035 2261
rect 12802 2252 12808 2264
rect 12860 2252 12866 2304
rect 13541 2295 13599 2301
rect 13541 2261 13553 2295
rect 13587 2292 13599 2295
rect 13998 2292 14004 2304
rect 13587 2264 14004 2292
rect 13587 2261 13599 2264
rect 13541 2255 13599 2261
rect 13998 2252 14004 2264
rect 14056 2252 14062 2304
rect 14921 2295 14979 2301
rect 14921 2261 14933 2295
rect 14967 2292 14979 2295
rect 15930 2292 15936 2304
rect 14967 2264 15936 2292
rect 14967 2261 14979 2264
rect 14921 2255 14979 2261
rect 15930 2252 15936 2264
rect 15988 2252 15994 2304
rect 16301 2295 16359 2301
rect 16301 2261 16313 2295
rect 16347 2292 16359 2295
rect 16390 2292 16396 2304
rect 16347 2264 16396 2292
rect 16347 2261 16359 2264
rect 16301 2255 16359 2261
rect 16390 2252 16396 2264
rect 16448 2252 16454 2304
rect 16850 2292 16856 2304
rect 16811 2264 16856 2292
rect 16850 2252 16856 2264
rect 16908 2252 16914 2304
rect 17310 2252 17316 2304
rect 17368 2292 17374 2304
rect 17405 2295 17463 2301
rect 17405 2292 17417 2295
rect 17368 2264 17417 2292
rect 17368 2252 17374 2264
rect 17405 2261 17417 2264
rect 17451 2261 17463 2295
rect 17405 2255 17463 2261
rect 18138 2252 18144 2304
rect 18196 2292 18202 2304
rect 18693 2295 18751 2301
rect 18693 2292 18705 2295
rect 18196 2264 18705 2292
rect 18196 2252 18202 2264
rect 18693 2261 18705 2264
rect 18739 2261 18751 2295
rect 18693 2255 18751 2261
rect 19150 2252 19156 2304
rect 19208 2292 19214 2304
rect 19613 2295 19671 2301
rect 19613 2292 19625 2295
rect 19208 2264 19625 2292
rect 19208 2252 19214 2264
rect 19613 2261 19625 2264
rect 19659 2261 19671 2295
rect 19613 2255 19671 2261
rect 20717 2295 20775 2301
rect 20717 2261 20729 2295
rect 20763 2292 20775 2295
rect 20898 2292 20904 2304
rect 20763 2264 20904 2292
rect 20763 2261 20775 2264
rect 20717 2255 20775 2261
rect 20898 2252 20904 2264
rect 20956 2252 20962 2304
rect 1104 2202 21896 2224
rect 1104 2150 4447 2202
rect 4499 2150 4511 2202
rect 4563 2150 4575 2202
rect 4627 2150 4639 2202
rect 4691 2150 11378 2202
rect 11430 2150 11442 2202
rect 11494 2150 11506 2202
rect 11558 2150 11570 2202
rect 11622 2150 18308 2202
rect 18360 2150 18372 2202
rect 18424 2150 18436 2202
rect 18488 2150 18500 2202
rect 18552 2150 21896 2202
rect 1104 2128 21896 2150
rect 5902 2048 5908 2100
rect 5960 2088 5966 2100
rect 6730 2088 6736 2100
rect 5960 2060 6736 2088
rect 5960 2048 5966 2060
rect 6730 2048 6736 2060
rect 6788 2048 6794 2100
rect 1486 1980 1492 2032
rect 1544 2020 1550 2032
rect 6270 2020 6276 2032
rect 1544 1992 6276 2020
rect 1544 1980 1550 1992
rect 6270 1980 6276 1992
rect 6328 1980 6334 2032
rect 5994 1504 6000 1556
rect 6052 1544 6058 1556
rect 8662 1544 8668 1556
rect 6052 1516 8668 1544
rect 6052 1504 6058 1516
rect 8662 1504 8668 1516
rect 8720 1504 8726 1556
<< via1 >>
rect 4447 20646 4499 20698
rect 4511 20646 4563 20698
rect 4575 20646 4627 20698
rect 4639 20646 4691 20698
rect 11378 20646 11430 20698
rect 11442 20646 11494 20698
rect 11506 20646 11558 20698
rect 11570 20646 11622 20698
rect 18308 20646 18360 20698
rect 18372 20646 18424 20698
rect 18436 20646 18488 20698
rect 18500 20646 18552 20698
rect 2780 20544 2832 20596
rect 20628 20544 20680 20596
rect 2872 20476 2924 20528
rect 7656 20408 7708 20460
rect 10048 20340 10100 20392
rect 19984 20340 20036 20392
rect 20260 20204 20312 20256
rect 20812 20204 20864 20256
rect 7912 20102 7964 20154
rect 7976 20102 8028 20154
rect 8040 20102 8092 20154
rect 8104 20102 8156 20154
rect 14843 20102 14895 20154
rect 14907 20102 14959 20154
rect 14971 20102 15023 20154
rect 15035 20102 15087 20154
rect 1952 20043 2004 20052
rect 1952 20009 1961 20043
rect 1961 20009 1995 20043
rect 1995 20009 2004 20043
rect 1952 20000 2004 20009
rect 20444 20043 20496 20052
rect 20444 20009 20453 20043
rect 20453 20009 20487 20043
rect 20487 20009 20496 20043
rect 20444 20000 20496 20009
rect 21088 20043 21140 20052
rect 21088 20009 21097 20043
rect 21097 20009 21131 20043
rect 21131 20009 21140 20043
rect 21088 20000 21140 20009
rect 6828 19864 6880 19916
rect 20168 19864 20220 19916
rect 20812 19864 20864 19916
rect 2872 19796 2924 19848
rect 7104 19796 7156 19848
rect 8392 19796 8444 19848
rect 5908 19728 5960 19780
rect 2044 19660 2096 19712
rect 3608 19703 3660 19712
rect 3608 19669 3617 19703
rect 3617 19669 3651 19703
rect 3651 19669 3660 19703
rect 3608 19660 3660 19669
rect 7564 19703 7616 19712
rect 7564 19669 7573 19703
rect 7573 19669 7607 19703
rect 7607 19669 7616 19703
rect 7564 19660 7616 19669
rect 19892 19703 19944 19712
rect 19892 19669 19901 19703
rect 19901 19669 19935 19703
rect 19935 19669 19944 19703
rect 19892 19660 19944 19669
rect 4447 19558 4499 19610
rect 4511 19558 4563 19610
rect 4575 19558 4627 19610
rect 4639 19558 4691 19610
rect 11378 19558 11430 19610
rect 11442 19558 11494 19610
rect 11506 19558 11558 19610
rect 11570 19558 11622 19610
rect 18308 19558 18360 19610
rect 18372 19558 18424 19610
rect 18436 19558 18488 19610
rect 18500 19558 18552 19610
rect 1952 19499 2004 19508
rect 1952 19465 1961 19499
rect 1961 19465 1995 19499
rect 1995 19465 2004 19499
rect 1952 19456 2004 19465
rect 9496 19456 9548 19508
rect 20444 19499 20496 19508
rect 20444 19465 20453 19499
rect 20453 19465 20487 19499
rect 20487 19465 20496 19499
rect 20444 19456 20496 19465
rect 19892 19320 19944 19372
rect 2044 19252 2096 19304
rect 3148 19295 3200 19304
rect 3148 19261 3157 19295
rect 3157 19261 3191 19295
rect 3191 19261 3200 19295
rect 3148 19252 3200 19261
rect 7564 19252 7616 19304
rect 8116 19295 8168 19304
rect 8116 19261 8125 19295
rect 8125 19261 8159 19295
rect 8159 19261 8168 19295
rect 8116 19252 8168 19261
rect 8392 19295 8444 19304
rect 8392 19261 8426 19295
rect 8426 19261 8444 19295
rect 8392 19252 8444 19261
rect 2964 19116 3016 19168
rect 3516 19184 3568 19236
rect 5724 19184 5776 19236
rect 3608 19116 3660 19168
rect 5080 19116 5132 19168
rect 6828 19116 6880 19168
rect 7564 19159 7616 19168
rect 7564 19125 7573 19159
rect 7573 19125 7607 19159
rect 7607 19125 7616 19159
rect 7564 19116 7616 19125
rect 10416 19295 10468 19304
rect 10416 19261 10425 19295
rect 10425 19261 10459 19295
rect 10459 19261 10468 19295
rect 10416 19252 10468 19261
rect 11980 19252 12032 19304
rect 18880 19295 18932 19304
rect 18880 19261 18889 19295
rect 18889 19261 18923 19295
rect 18923 19261 18932 19295
rect 18880 19252 18932 19261
rect 19340 19252 19392 19304
rect 20260 19295 20312 19304
rect 20260 19261 20269 19295
rect 20269 19261 20303 19295
rect 20303 19261 20312 19295
rect 20260 19252 20312 19261
rect 13360 19184 13412 19236
rect 19248 19184 19300 19236
rect 9496 19159 9548 19168
rect 9496 19125 9505 19159
rect 9505 19125 9539 19159
rect 9539 19125 9548 19159
rect 9496 19116 9548 19125
rect 11796 19159 11848 19168
rect 11796 19125 11805 19159
rect 11805 19125 11839 19159
rect 11839 19125 11848 19159
rect 11796 19116 11848 19125
rect 14740 19116 14792 19168
rect 15568 19116 15620 19168
rect 19156 19116 19208 19168
rect 20996 19159 21048 19168
rect 20996 19125 21005 19159
rect 21005 19125 21039 19159
rect 21039 19125 21048 19159
rect 20996 19116 21048 19125
rect 7912 19014 7964 19066
rect 7976 19014 8028 19066
rect 8040 19014 8092 19066
rect 8104 19014 8156 19066
rect 14843 19014 14895 19066
rect 14907 19014 14959 19066
rect 14971 19014 15023 19066
rect 15035 19014 15087 19066
rect 1952 18955 2004 18964
rect 1952 18921 1961 18955
rect 1961 18921 1995 18955
rect 1995 18921 2004 18955
rect 1952 18912 2004 18921
rect 2780 18912 2832 18964
rect 3056 18955 3108 18964
rect 3056 18921 3065 18955
rect 3065 18921 3099 18955
rect 3099 18921 3108 18955
rect 3056 18912 3108 18921
rect 3608 18912 3660 18964
rect 5448 18912 5500 18964
rect 8392 18912 8444 18964
rect 9496 18912 9548 18964
rect 17224 18912 17276 18964
rect 21088 18955 21140 18964
rect 21088 18921 21097 18955
rect 21097 18921 21131 18955
rect 21131 18921 21140 18955
rect 21088 18912 21140 18921
rect 6184 18844 6236 18896
rect 2872 18819 2924 18828
rect 2872 18785 2881 18819
rect 2881 18785 2915 18819
rect 2915 18785 2924 18819
rect 2872 18776 2924 18785
rect 3608 18776 3660 18828
rect 3148 18708 3200 18760
rect 3240 18640 3292 18692
rect 4344 18708 4396 18760
rect 4988 18776 5040 18828
rect 8208 18844 8260 18896
rect 10416 18844 10468 18896
rect 15292 18844 15344 18896
rect 8944 18776 8996 18828
rect 11796 18776 11848 18828
rect 14648 18819 14700 18828
rect 11980 18751 12032 18760
rect 11980 18717 11989 18751
rect 11989 18717 12023 18751
rect 12023 18717 12032 18751
rect 11980 18708 12032 18717
rect 13360 18683 13412 18692
rect 3700 18572 3752 18624
rect 13360 18649 13369 18683
rect 13369 18649 13403 18683
rect 13403 18649 13412 18683
rect 13360 18640 13412 18649
rect 14648 18785 14657 18819
rect 14657 18785 14691 18819
rect 14691 18785 14700 18819
rect 14648 18776 14700 18785
rect 14740 18751 14792 18760
rect 14740 18717 14749 18751
rect 14749 18717 14783 18751
rect 14783 18717 14792 18751
rect 14740 18708 14792 18717
rect 17408 18844 17460 18896
rect 20168 18887 20220 18896
rect 20168 18853 20177 18887
rect 20177 18853 20211 18887
rect 20211 18853 20220 18887
rect 20168 18844 20220 18853
rect 15568 18819 15620 18828
rect 15568 18785 15602 18819
rect 15602 18785 15620 18819
rect 15568 18776 15620 18785
rect 20076 18776 20128 18828
rect 20352 18708 20404 18760
rect 15200 18640 15252 18692
rect 5540 18572 5592 18624
rect 6920 18572 6972 18624
rect 14188 18615 14240 18624
rect 14188 18581 14197 18615
rect 14197 18581 14231 18615
rect 14231 18581 14240 18615
rect 14188 18572 14240 18581
rect 16028 18572 16080 18624
rect 19340 18572 19392 18624
rect 4447 18470 4499 18522
rect 4511 18470 4563 18522
rect 4575 18470 4627 18522
rect 4639 18470 4691 18522
rect 11378 18470 11430 18522
rect 11442 18470 11494 18522
rect 11506 18470 11558 18522
rect 11570 18470 11622 18522
rect 18308 18470 18360 18522
rect 18372 18470 18424 18522
rect 18436 18470 18488 18522
rect 18500 18470 18552 18522
rect 1952 18411 2004 18420
rect 1952 18377 1961 18411
rect 1961 18377 1995 18411
rect 1995 18377 2004 18411
rect 1952 18368 2004 18377
rect 3608 18368 3660 18420
rect 4988 18411 5040 18420
rect 4988 18377 4997 18411
rect 4997 18377 5031 18411
rect 5031 18377 5040 18411
rect 4988 18368 5040 18377
rect 7564 18368 7616 18420
rect 20444 18411 20496 18420
rect 20444 18377 20453 18411
rect 20453 18377 20487 18411
rect 20487 18377 20496 18411
rect 20444 18368 20496 18377
rect 3148 18164 3200 18216
rect 8392 18232 8444 18284
rect 10416 18275 10468 18284
rect 10416 18241 10425 18275
rect 10425 18241 10459 18275
rect 10459 18241 10468 18275
rect 10416 18232 10468 18241
rect 14740 18232 14792 18284
rect 16028 18275 16080 18284
rect 16028 18241 16037 18275
rect 16037 18241 16071 18275
rect 16071 18241 16080 18275
rect 16028 18232 16080 18241
rect 14188 18164 14240 18216
rect 20536 18164 20588 18216
rect 2964 18071 3016 18080
rect 2964 18037 2973 18071
rect 2973 18037 3007 18071
rect 3007 18037 3016 18071
rect 2964 18028 3016 18037
rect 3056 18071 3108 18080
rect 3056 18037 3065 18071
rect 3065 18037 3099 18071
rect 3099 18037 3108 18071
rect 5080 18096 5132 18148
rect 5908 18096 5960 18148
rect 9588 18096 9640 18148
rect 10968 18096 11020 18148
rect 14740 18096 14792 18148
rect 17040 18096 17092 18148
rect 3056 18028 3108 18037
rect 8208 18028 8260 18080
rect 8484 18071 8536 18080
rect 8484 18037 8493 18071
rect 8493 18037 8527 18071
rect 8527 18037 8536 18071
rect 8484 18028 8536 18037
rect 8576 18071 8628 18080
rect 8576 18037 8585 18071
rect 8585 18037 8619 18071
rect 8619 18037 8628 18071
rect 9220 18071 9272 18080
rect 8576 18028 8628 18037
rect 9220 18037 9229 18071
rect 9229 18037 9263 18071
rect 9263 18037 9272 18071
rect 9220 18028 9272 18037
rect 10508 18028 10560 18080
rect 12164 18028 12216 18080
rect 13544 18028 13596 18080
rect 13820 18028 13872 18080
rect 17132 18028 17184 18080
rect 19800 18028 19852 18080
rect 20996 18071 21048 18080
rect 20996 18037 21005 18071
rect 21005 18037 21039 18071
rect 21039 18037 21048 18071
rect 20996 18028 21048 18037
rect 7912 17926 7964 17978
rect 7976 17926 8028 17978
rect 8040 17926 8092 17978
rect 8104 17926 8156 17978
rect 14843 17926 14895 17978
rect 14907 17926 14959 17978
rect 14971 17926 15023 17978
rect 15035 17926 15087 17978
rect 1676 17867 1728 17876
rect 1676 17833 1685 17867
rect 1685 17833 1719 17867
rect 1719 17833 1728 17867
rect 1676 17824 1728 17833
rect 2964 17867 3016 17876
rect 2964 17833 2973 17867
rect 2973 17833 3007 17867
rect 3007 17833 3016 17867
rect 2964 17824 3016 17833
rect 4344 17824 4396 17876
rect 8576 17824 8628 17876
rect 12440 17824 12492 17876
rect 14648 17824 14700 17876
rect 15292 17867 15344 17876
rect 15292 17833 15301 17867
rect 15301 17833 15335 17867
rect 15335 17833 15344 17867
rect 15292 17824 15344 17833
rect 17040 17824 17092 17876
rect 17500 17824 17552 17876
rect 19892 17824 19944 17876
rect 3424 17799 3476 17808
rect 3424 17765 3433 17799
rect 3433 17765 3467 17799
rect 3467 17765 3476 17799
rect 3424 17756 3476 17765
rect 6092 17756 6144 17808
rect 6184 17756 6236 17808
rect 8208 17756 8260 17808
rect 9220 17756 9272 17808
rect 10416 17756 10468 17808
rect 10508 17756 10560 17808
rect 11888 17756 11940 17808
rect 1492 17731 1544 17740
rect 1492 17697 1501 17731
rect 1501 17697 1535 17731
rect 1535 17697 1544 17731
rect 1492 17688 1544 17697
rect 3240 17688 3292 17740
rect 4160 17688 4212 17740
rect 7012 17688 7064 17740
rect 8300 17688 8352 17740
rect 8760 17731 8812 17740
rect 8760 17697 8769 17731
rect 8769 17697 8803 17731
rect 8803 17697 8812 17731
rect 8760 17688 8812 17697
rect 9680 17731 9732 17740
rect 9680 17697 9689 17731
rect 9689 17697 9723 17731
rect 9723 17697 9732 17731
rect 9680 17688 9732 17697
rect 9772 17688 9824 17740
rect 11704 17688 11756 17740
rect 1768 17620 1820 17672
rect 3516 17663 3568 17672
rect 3516 17629 3525 17663
rect 3525 17629 3559 17663
rect 3559 17629 3568 17663
rect 3516 17620 3568 17629
rect 4988 17663 5040 17672
rect 4988 17629 4997 17663
rect 4997 17629 5031 17663
rect 5031 17629 5040 17663
rect 4988 17620 5040 17629
rect 5080 17663 5132 17672
rect 5080 17629 5089 17663
rect 5089 17629 5123 17663
rect 5123 17629 5132 17663
rect 5080 17620 5132 17629
rect 5540 17620 5592 17672
rect 8944 17663 8996 17672
rect 8944 17629 8953 17663
rect 8953 17629 8987 17663
rect 8987 17629 8996 17663
rect 8944 17620 8996 17629
rect 10692 17620 10744 17672
rect 12256 17663 12308 17672
rect 12256 17629 12265 17663
rect 12265 17629 12299 17663
rect 12299 17629 12308 17663
rect 12256 17620 12308 17629
rect 13452 17756 13504 17808
rect 13268 17688 13320 17740
rect 13728 17731 13780 17740
rect 13728 17697 13737 17731
rect 13737 17697 13771 17731
rect 13771 17697 13780 17731
rect 13728 17688 13780 17697
rect 3608 17484 3660 17536
rect 9496 17552 9548 17604
rect 7196 17484 7248 17536
rect 10968 17484 11020 17536
rect 11152 17484 11204 17536
rect 13636 17620 13688 17672
rect 14004 17756 14056 17808
rect 20076 17799 20128 17808
rect 17408 17731 17460 17740
rect 14280 17620 14332 17672
rect 15844 17663 15896 17672
rect 15844 17629 15853 17663
rect 15853 17629 15887 17663
rect 15887 17629 15896 17663
rect 16856 17663 16908 17672
rect 15844 17620 15896 17629
rect 16856 17629 16865 17663
rect 16865 17629 16899 17663
rect 16899 17629 16908 17663
rect 16856 17620 16908 17629
rect 17408 17697 17417 17731
rect 17417 17697 17451 17731
rect 17451 17697 17460 17731
rect 17408 17688 17460 17697
rect 17500 17688 17552 17740
rect 17684 17731 17736 17740
rect 17684 17697 17718 17731
rect 17718 17697 17736 17731
rect 17684 17688 17736 17697
rect 17960 17688 18012 17740
rect 19340 17688 19392 17740
rect 14280 17484 14332 17536
rect 16396 17527 16448 17536
rect 16396 17493 16405 17527
rect 16405 17493 16439 17527
rect 16439 17493 16448 17527
rect 16396 17484 16448 17493
rect 20076 17765 20085 17799
rect 20085 17765 20119 17799
rect 20119 17765 20128 17799
rect 20076 17756 20128 17765
rect 19616 17688 19668 17740
rect 20260 17688 20312 17740
rect 19892 17484 19944 17536
rect 21088 17527 21140 17536
rect 21088 17493 21097 17527
rect 21097 17493 21131 17527
rect 21131 17493 21140 17527
rect 21088 17484 21140 17493
rect 4447 17382 4499 17434
rect 4511 17382 4563 17434
rect 4575 17382 4627 17434
rect 4639 17382 4691 17434
rect 11378 17382 11430 17434
rect 11442 17382 11494 17434
rect 11506 17382 11558 17434
rect 11570 17382 11622 17434
rect 18308 17382 18360 17434
rect 18372 17382 18424 17434
rect 18436 17382 18488 17434
rect 18500 17382 18552 17434
rect 2780 17280 2832 17332
rect 3056 17280 3108 17332
rect 4988 17280 5040 17332
rect 7012 17323 7064 17332
rect 7012 17289 7021 17323
rect 7021 17289 7055 17323
rect 7055 17289 7064 17323
rect 7012 17280 7064 17289
rect 8484 17280 8536 17332
rect 9496 17280 9548 17332
rect 10140 17280 10192 17332
rect 13820 17280 13872 17332
rect 14740 17280 14792 17332
rect 1492 17255 1544 17264
rect 1492 17221 1501 17255
rect 1501 17221 1535 17255
rect 1535 17221 1544 17255
rect 1492 17212 1544 17221
rect 3608 17212 3660 17264
rect 3516 17144 3568 17196
rect 4160 17187 4212 17196
rect 4160 17153 4169 17187
rect 4169 17153 4203 17187
rect 4203 17153 4212 17187
rect 4160 17144 4212 17153
rect 7196 17144 7248 17196
rect 2228 17076 2280 17128
rect 2320 17119 2372 17128
rect 2320 17085 2329 17119
rect 2329 17085 2363 17119
rect 2363 17085 2372 17119
rect 2320 17076 2372 17085
rect 3332 17076 3384 17128
rect 10784 17212 10836 17264
rect 19708 17280 19760 17332
rect 8392 17144 8444 17196
rect 8944 17144 8996 17196
rect 10968 17144 11020 17196
rect 12440 17187 12492 17196
rect 12440 17153 12449 17187
rect 12449 17153 12483 17187
rect 12483 17153 12492 17187
rect 12440 17144 12492 17153
rect 10324 17076 10376 17128
rect 11152 17076 11204 17128
rect 12072 17076 12124 17128
rect 17500 17212 17552 17264
rect 17960 17212 18012 17264
rect 13452 17144 13504 17196
rect 15844 17144 15896 17196
rect 16488 17144 16540 17196
rect 17132 17144 17184 17196
rect 5356 17008 5408 17060
rect 6828 17008 6880 17060
rect 7288 17008 7340 17060
rect 8208 17008 8260 17060
rect 16396 17076 16448 17128
rect 17408 17076 17460 17128
rect 17776 17076 17828 17128
rect 19892 17076 19944 17128
rect 1952 16983 2004 16992
rect 1952 16949 1961 16983
rect 1961 16949 1995 16983
rect 1995 16949 2004 16983
rect 1952 16940 2004 16949
rect 3516 16983 3568 16992
rect 3516 16949 3525 16983
rect 3525 16949 3559 16983
rect 3559 16949 3568 16983
rect 3516 16940 3568 16949
rect 5540 16983 5592 16992
rect 5540 16949 5549 16983
rect 5549 16949 5583 16983
rect 5583 16949 5592 16983
rect 5540 16940 5592 16949
rect 8760 16940 8812 16992
rect 9312 16940 9364 16992
rect 9956 16940 10008 16992
rect 10232 16983 10284 16992
rect 10232 16949 10241 16983
rect 10241 16949 10275 16983
rect 10275 16949 10284 16983
rect 10232 16940 10284 16949
rect 10968 16940 11020 16992
rect 11244 16983 11296 16992
rect 11244 16949 11253 16983
rect 11253 16949 11287 16983
rect 11287 16949 11296 16983
rect 11244 16940 11296 16949
rect 12992 16940 13044 16992
rect 13452 16940 13504 16992
rect 15568 16983 15620 16992
rect 15568 16949 15577 16983
rect 15577 16949 15611 16983
rect 15611 16949 15620 16983
rect 15568 16940 15620 16949
rect 18052 17008 18104 17060
rect 19064 17008 19116 17060
rect 20904 17008 20956 17060
rect 17224 16983 17276 16992
rect 17224 16949 17233 16983
rect 17233 16949 17267 16983
rect 17267 16949 17276 16983
rect 17224 16940 17276 16949
rect 17684 16940 17736 16992
rect 20628 16940 20680 16992
rect 7912 16838 7964 16890
rect 7976 16838 8028 16890
rect 8040 16838 8092 16890
rect 8104 16838 8156 16890
rect 14843 16838 14895 16890
rect 14907 16838 14959 16890
rect 14971 16838 15023 16890
rect 15035 16838 15087 16890
rect 5540 16779 5592 16788
rect 5540 16745 5549 16779
rect 5549 16745 5583 16779
rect 5583 16745 5592 16779
rect 5540 16736 5592 16745
rect 7564 16736 7616 16788
rect 8208 16736 8260 16788
rect 10968 16779 11020 16788
rect 10968 16745 10977 16779
rect 10977 16745 11011 16779
rect 11011 16745 11020 16779
rect 10968 16736 11020 16745
rect 11244 16736 11296 16788
rect 13452 16779 13504 16788
rect 13452 16745 13461 16779
rect 13461 16745 13495 16779
rect 13495 16745 13504 16779
rect 13452 16736 13504 16745
rect 15568 16736 15620 16788
rect 16856 16736 16908 16788
rect 19248 16736 19300 16788
rect 21272 16736 21324 16788
rect 5908 16711 5960 16720
rect 1768 16643 1820 16652
rect 1768 16609 1777 16643
rect 1777 16609 1811 16643
rect 1811 16609 1820 16643
rect 1768 16600 1820 16609
rect 5908 16677 5917 16711
rect 5917 16677 5951 16711
rect 5951 16677 5960 16711
rect 5908 16668 5960 16677
rect 6828 16668 6880 16720
rect 10232 16668 10284 16720
rect 7288 16600 7340 16652
rect 10508 16600 10560 16652
rect 6092 16575 6144 16584
rect 6092 16541 6101 16575
rect 6101 16541 6135 16575
rect 6135 16541 6144 16575
rect 6092 16532 6144 16541
rect 9772 16532 9824 16584
rect 10876 16532 10928 16584
rect 11704 16532 11756 16584
rect 2504 16507 2556 16516
rect 2504 16473 2513 16507
rect 2513 16473 2547 16507
rect 2547 16473 2556 16507
rect 2504 16464 2556 16473
rect 3516 16464 3568 16516
rect 3700 16464 3752 16516
rect 9036 16464 9088 16516
rect 1860 16396 1912 16448
rect 2320 16396 2372 16448
rect 6000 16396 6052 16448
rect 7288 16439 7340 16448
rect 7288 16405 7297 16439
rect 7297 16405 7331 16439
rect 7331 16405 7340 16439
rect 7288 16396 7340 16405
rect 9956 16439 10008 16448
rect 9956 16405 9965 16439
rect 9965 16405 9999 16439
rect 9999 16405 10008 16439
rect 9956 16396 10008 16405
rect 10324 16439 10376 16448
rect 10324 16405 10333 16439
rect 10333 16405 10367 16439
rect 10367 16405 10376 16439
rect 10324 16396 10376 16405
rect 12072 16600 12124 16652
rect 13820 16643 13872 16652
rect 13820 16609 13829 16643
rect 13829 16609 13863 16643
rect 13863 16609 13872 16643
rect 13820 16600 13872 16609
rect 16856 16600 16908 16652
rect 17224 16600 17276 16652
rect 12164 16532 12216 16584
rect 12992 16507 13044 16516
rect 12992 16473 13001 16507
rect 13001 16473 13035 16507
rect 13035 16473 13044 16507
rect 12992 16464 13044 16473
rect 15200 16532 15252 16584
rect 16672 16575 16724 16584
rect 16672 16541 16681 16575
rect 16681 16541 16715 16575
rect 16715 16541 16724 16575
rect 16672 16532 16724 16541
rect 17868 16575 17920 16584
rect 14004 16396 14056 16448
rect 16488 16464 16540 16516
rect 17868 16541 17877 16575
rect 17877 16541 17911 16575
rect 17911 16541 17920 16575
rect 17868 16532 17920 16541
rect 18972 16600 19024 16652
rect 19524 16600 19576 16652
rect 19708 16600 19760 16652
rect 20720 16600 20772 16652
rect 20904 16643 20956 16652
rect 20904 16609 20913 16643
rect 20913 16609 20947 16643
rect 20947 16609 20956 16643
rect 20904 16600 20956 16609
rect 17684 16464 17736 16516
rect 17040 16396 17092 16448
rect 18972 16439 19024 16448
rect 18972 16405 18981 16439
rect 18981 16405 19015 16439
rect 19015 16405 19024 16439
rect 18972 16396 19024 16405
rect 4447 16294 4499 16346
rect 4511 16294 4563 16346
rect 4575 16294 4627 16346
rect 4639 16294 4691 16346
rect 11378 16294 11430 16346
rect 11442 16294 11494 16346
rect 11506 16294 11558 16346
rect 11570 16294 11622 16346
rect 18308 16294 18360 16346
rect 18372 16294 18424 16346
rect 18436 16294 18488 16346
rect 18500 16294 18552 16346
rect 3332 16192 3384 16244
rect 4252 16192 4304 16244
rect 6092 16192 6144 16244
rect 7104 16235 7156 16244
rect 7104 16201 7113 16235
rect 7113 16201 7147 16235
rect 7147 16201 7156 16235
rect 7104 16192 7156 16201
rect 8392 16192 8444 16244
rect 10324 16192 10376 16244
rect 13544 16192 13596 16244
rect 16672 16192 16724 16244
rect 17960 16192 18012 16244
rect 18144 16192 18196 16244
rect 18696 16192 18748 16244
rect 1676 16167 1728 16176
rect 1676 16133 1685 16167
rect 1685 16133 1719 16167
rect 1719 16133 1728 16167
rect 1676 16124 1728 16133
rect 2228 16099 2280 16108
rect 2228 16065 2237 16099
rect 2237 16065 2271 16099
rect 2271 16065 2280 16099
rect 2228 16056 2280 16065
rect 9496 16124 9548 16176
rect 13820 16124 13872 16176
rect 8392 16056 8444 16108
rect 11704 16056 11756 16108
rect 18972 16056 19024 16108
rect 20260 16099 20312 16108
rect 20260 16065 20269 16099
rect 20269 16065 20303 16099
rect 20303 16065 20312 16099
rect 20260 16056 20312 16065
rect 4344 15988 4396 16040
rect 4436 16031 4488 16040
rect 4436 15997 4445 16031
rect 4445 15997 4479 16031
rect 4479 15997 4488 16031
rect 4436 15988 4488 15997
rect 5632 15988 5684 16040
rect 7288 15988 7340 16040
rect 8484 16031 8536 16040
rect 8484 15997 8493 16031
rect 8493 15997 8527 16031
rect 8527 15997 8536 16031
rect 8484 15988 8536 15997
rect 9680 15988 9732 16040
rect 13820 15988 13872 16040
rect 20720 15988 20772 16040
rect 4712 15963 4764 15972
rect 4712 15929 4746 15963
rect 4746 15929 4764 15963
rect 4712 15920 4764 15929
rect 7380 15920 7432 15972
rect 8852 15920 8904 15972
rect 9864 15920 9916 15972
rect 16396 15920 16448 15972
rect 5816 15852 5868 15904
rect 6644 15852 6696 15904
rect 10876 15852 10928 15904
rect 16856 15852 16908 15904
rect 19708 15895 19760 15904
rect 19708 15861 19717 15895
rect 19717 15861 19751 15895
rect 19751 15861 19760 15895
rect 19708 15852 19760 15861
rect 20628 15852 20680 15904
rect 7912 15750 7964 15802
rect 7976 15750 8028 15802
rect 8040 15750 8092 15802
rect 8104 15750 8156 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 15035 15750 15087 15802
rect 1952 15691 2004 15700
rect 1952 15657 1961 15691
rect 1961 15657 1995 15691
rect 1995 15657 2004 15691
rect 1952 15648 2004 15657
rect 2412 15512 2464 15564
rect 3056 15555 3108 15564
rect 3056 15521 3065 15555
rect 3065 15521 3099 15555
rect 3099 15521 3108 15555
rect 3056 15512 3108 15521
rect 2320 15444 2372 15496
rect 3148 15487 3200 15496
rect 1584 15376 1636 15428
rect 3148 15453 3157 15487
rect 3157 15453 3191 15487
rect 3191 15453 3200 15487
rect 3148 15444 3200 15453
rect 4712 15648 4764 15700
rect 6920 15648 6972 15700
rect 8484 15648 8536 15700
rect 13820 15691 13872 15700
rect 13820 15657 13829 15691
rect 13829 15657 13863 15691
rect 13863 15657 13872 15691
rect 13820 15648 13872 15657
rect 15384 15648 15436 15700
rect 18880 15648 18932 15700
rect 19064 15691 19116 15700
rect 19064 15657 19073 15691
rect 19073 15657 19107 15691
rect 19107 15657 19116 15691
rect 19064 15648 19116 15657
rect 20444 15691 20496 15700
rect 20444 15657 20453 15691
rect 20453 15657 20487 15691
rect 20487 15657 20496 15691
rect 20444 15648 20496 15657
rect 21088 15691 21140 15700
rect 21088 15657 21097 15691
rect 21097 15657 21131 15691
rect 21131 15657 21140 15691
rect 21088 15648 21140 15657
rect 4436 15580 4488 15632
rect 12164 15580 12216 15632
rect 16028 15580 16080 15632
rect 4160 15512 4212 15564
rect 5632 15512 5684 15564
rect 6920 15512 6972 15564
rect 11980 15512 12032 15564
rect 14188 15555 14240 15564
rect 14188 15521 14197 15555
rect 14197 15521 14231 15555
rect 14231 15521 14240 15555
rect 14188 15512 14240 15521
rect 15660 15512 15712 15564
rect 17776 15512 17828 15564
rect 17960 15555 18012 15564
rect 17960 15521 17994 15555
rect 17994 15521 18012 15555
rect 17960 15512 18012 15521
rect 19708 15512 19760 15564
rect 20444 15512 20496 15564
rect 13820 15444 13872 15496
rect 14556 15444 14608 15496
rect 19340 15487 19392 15496
rect 19340 15453 19349 15487
rect 19349 15453 19383 15487
rect 19383 15453 19392 15487
rect 19340 15444 19392 15453
rect 7380 15376 7432 15428
rect 12348 15376 12400 15428
rect 15200 15376 15252 15428
rect 2412 15351 2464 15360
rect 2412 15317 2421 15351
rect 2421 15317 2455 15351
rect 2455 15317 2464 15351
rect 2412 15308 2464 15317
rect 6828 15308 6880 15360
rect 7472 15308 7524 15360
rect 16948 15351 17000 15360
rect 16948 15317 16957 15351
rect 16957 15317 16991 15351
rect 16991 15317 17000 15351
rect 16948 15308 17000 15317
rect 19892 15351 19944 15360
rect 19892 15317 19901 15351
rect 19901 15317 19935 15351
rect 19935 15317 19944 15351
rect 19892 15308 19944 15317
rect 4447 15206 4499 15258
rect 4511 15206 4563 15258
rect 4575 15206 4627 15258
rect 4639 15206 4691 15258
rect 11378 15206 11430 15258
rect 11442 15206 11494 15258
rect 11506 15206 11558 15258
rect 11570 15206 11622 15258
rect 18308 15206 18360 15258
rect 18372 15206 18424 15258
rect 18436 15206 18488 15258
rect 18500 15206 18552 15258
rect 5632 15104 5684 15156
rect 8852 15104 8904 15156
rect 11980 15104 12032 15156
rect 8484 15011 8536 15020
rect 8484 14977 8493 15011
rect 8493 14977 8527 15011
rect 8527 14977 8536 15011
rect 8484 14968 8536 14977
rect 9680 14968 9732 15020
rect 12716 14968 12768 15020
rect 15200 14968 15252 15020
rect 15936 14968 15988 15020
rect 1768 14943 1820 14952
rect 1768 14909 1777 14943
rect 1777 14909 1811 14943
rect 1811 14909 1820 14943
rect 1768 14900 1820 14909
rect 2320 14900 2372 14952
rect 2780 14875 2832 14884
rect 2780 14841 2814 14875
rect 2814 14841 2832 14875
rect 9864 14900 9916 14952
rect 2780 14832 2832 14841
rect 6920 14832 6972 14884
rect 7472 14832 7524 14884
rect 1952 14807 2004 14816
rect 1952 14773 1961 14807
rect 1961 14773 1995 14807
rect 1995 14773 2004 14807
rect 1952 14764 2004 14773
rect 3884 14807 3936 14816
rect 3884 14773 3893 14807
rect 3893 14773 3927 14807
rect 3927 14773 3936 14807
rect 3884 14764 3936 14773
rect 4160 14764 4212 14816
rect 6460 14764 6512 14816
rect 10232 14764 10284 14816
rect 15384 14900 15436 14952
rect 19064 15036 19116 15088
rect 17960 14968 18012 15020
rect 18788 14968 18840 15020
rect 19248 14968 19300 15020
rect 20812 14943 20864 14952
rect 20812 14909 20821 14943
rect 20821 14909 20855 14943
rect 20855 14909 20864 14943
rect 20812 14900 20864 14909
rect 13452 14875 13504 14884
rect 13452 14841 13486 14875
rect 13486 14841 13504 14875
rect 13452 14832 13504 14841
rect 13912 14764 13964 14816
rect 14556 14807 14608 14816
rect 14556 14773 14565 14807
rect 14565 14773 14599 14807
rect 14599 14773 14608 14807
rect 14556 14764 14608 14773
rect 14740 14764 14792 14816
rect 15200 14807 15252 14816
rect 15200 14773 15209 14807
rect 15209 14773 15243 14807
rect 15243 14773 15252 14807
rect 15200 14764 15252 14773
rect 15844 14764 15896 14816
rect 19340 14832 19392 14884
rect 19432 14764 19484 14816
rect 20076 14764 20128 14816
rect 20260 14807 20312 14816
rect 20260 14773 20269 14807
rect 20269 14773 20303 14807
rect 20303 14773 20312 14807
rect 20260 14764 20312 14773
rect 20996 14807 21048 14816
rect 20996 14773 21005 14807
rect 21005 14773 21039 14807
rect 21039 14773 21048 14807
rect 20996 14764 21048 14773
rect 7912 14662 7964 14714
rect 7976 14662 8028 14714
rect 8040 14662 8092 14714
rect 8104 14662 8156 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 15035 14662 15087 14714
rect 3056 14560 3108 14612
rect 3148 14560 3200 14612
rect 5816 14603 5868 14612
rect 5816 14569 5825 14603
rect 5825 14569 5859 14603
rect 5859 14569 5868 14603
rect 5816 14560 5868 14569
rect 7656 14560 7708 14612
rect 14188 14560 14240 14612
rect 15200 14560 15252 14612
rect 19432 14603 19484 14612
rect 19432 14569 19441 14603
rect 19441 14569 19475 14603
rect 19475 14569 19484 14603
rect 19432 14560 19484 14569
rect 1768 14492 1820 14544
rect 7380 14492 7432 14544
rect 12348 14492 12400 14544
rect 14740 14492 14792 14544
rect 17960 14492 18012 14544
rect 20720 14492 20772 14544
rect 20812 14492 20864 14544
rect 1584 14467 1636 14476
rect 1584 14433 1593 14467
rect 1593 14433 1627 14467
rect 1627 14433 1636 14467
rect 1584 14424 1636 14433
rect 2228 14424 2280 14476
rect 4160 14424 4212 14476
rect 6184 14467 6236 14476
rect 6184 14433 6193 14467
rect 6193 14433 6227 14467
rect 6227 14433 6236 14467
rect 6184 14424 6236 14433
rect 9680 14467 9732 14476
rect 9680 14433 9689 14467
rect 9689 14433 9723 14467
rect 9723 14433 9732 14467
rect 9680 14424 9732 14433
rect 10232 14424 10284 14476
rect 11980 14467 12032 14476
rect 11980 14433 11989 14467
rect 11989 14433 12023 14467
rect 12023 14433 12032 14467
rect 11980 14424 12032 14433
rect 15200 14424 15252 14476
rect 15384 14424 15436 14476
rect 15660 14424 15712 14476
rect 2504 14356 2556 14408
rect 3884 14356 3936 14408
rect 4068 14356 4120 14408
rect 6460 14399 6512 14408
rect 6460 14365 6469 14399
rect 6469 14365 6503 14399
rect 6503 14365 6512 14399
rect 6460 14356 6512 14365
rect 7104 14356 7156 14408
rect 7472 14399 7524 14408
rect 7472 14365 7481 14399
rect 7481 14365 7515 14399
rect 7515 14365 7524 14399
rect 7472 14356 7524 14365
rect 14096 14399 14148 14408
rect 14096 14365 14105 14399
rect 14105 14365 14139 14399
rect 14139 14365 14148 14399
rect 14096 14356 14148 14365
rect 13452 14288 13504 14340
rect 14372 14356 14424 14408
rect 15752 14399 15804 14408
rect 15752 14365 15761 14399
rect 15761 14365 15795 14399
rect 15795 14365 15804 14399
rect 15752 14356 15804 14365
rect 16764 14288 16816 14340
rect 19248 14424 19300 14476
rect 19708 14424 19760 14476
rect 20076 14424 20128 14476
rect 5264 14220 5316 14272
rect 9864 14220 9916 14272
rect 15752 14220 15804 14272
rect 18788 14263 18840 14272
rect 18788 14229 18797 14263
rect 18797 14229 18831 14263
rect 18831 14229 18840 14263
rect 18788 14220 18840 14229
rect 20168 14220 20220 14272
rect 20444 14263 20496 14272
rect 20444 14229 20453 14263
rect 20453 14229 20487 14263
rect 20487 14229 20496 14263
rect 20444 14220 20496 14229
rect 4447 14118 4499 14170
rect 4511 14118 4563 14170
rect 4575 14118 4627 14170
rect 4639 14118 4691 14170
rect 11378 14118 11430 14170
rect 11442 14118 11494 14170
rect 11506 14118 11558 14170
rect 11570 14118 11622 14170
rect 18308 14118 18360 14170
rect 18372 14118 18424 14170
rect 18436 14118 18488 14170
rect 18500 14118 18552 14170
rect 1860 14059 1912 14068
rect 1860 14025 1869 14059
rect 1869 14025 1903 14059
rect 1903 14025 1912 14059
rect 1860 14016 1912 14025
rect 2228 14059 2280 14068
rect 2228 14025 2237 14059
rect 2237 14025 2271 14059
rect 2271 14025 2280 14059
rect 2228 14016 2280 14025
rect 4068 14059 4120 14068
rect 4068 14025 4077 14059
rect 4077 14025 4111 14059
rect 4111 14025 4120 14059
rect 4068 14016 4120 14025
rect 7104 14059 7156 14068
rect 7104 14025 7113 14059
rect 7113 14025 7147 14059
rect 7147 14025 7156 14059
rect 7104 14016 7156 14025
rect 8300 14059 8352 14068
rect 8300 14025 8309 14059
rect 8309 14025 8343 14059
rect 8343 14025 8352 14059
rect 8300 14016 8352 14025
rect 14096 14016 14148 14068
rect 15844 14059 15896 14068
rect 15844 14025 15853 14059
rect 15853 14025 15887 14059
rect 15887 14025 15896 14059
rect 15844 14016 15896 14025
rect 18052 14016 18104 14068
rect 20260 14016 20312 14068
rect 21088 14059 21140 14068
rect 21088 14025 21097 14059
rect 21097 14025 21131 14059
rect 21131 14025 21140 14059
rect 21088 14016 21140 14025
rect 13820 13991 13872 14000
rect 13820 13957 13829 13991
rect 13829 13957 13863 13991
rect 13863 13957 13872 13991
rect 13820 13948 13872 13957
rect 13912 13948 13964 14000
rect 18144 13991 18196 14000
rect 2780 13923 2832 13932
rect 2780 13889 2789 13923
rect 2789 13889 2823 13923
rect 2823 13889 2832 13923
rect 2780 13880 2832 13889
rect 2964 13880 3016 13932
rect 5172 13880 5224 13932
rect 6000 13880 6052 13932
rect 2136 13812 2188 13864
rect 7012 13880 7064 13932
rect 8208 13880 8260 13932
rect 8852 13923 8904 13932
rect 8852 13889 8861 13923
rect 8861 13889 8895 13923
rect 8895 13889 8904 13923
rect 8852 13880 8904 13889
rect 9864 13923 9916 13932
rect 9864 13889 9873 13923
rect 9873 13889 9907 13923
rect 9907 13889 9916 13923
rect 9864 13880 9916 13889
rect 10324 13880 10376 13932
rect 8300 13812 8352 13864
rect 10416 13812 10468 13864
rect 11796 13880 11848 13932
rect 12348 13880 12400 13932
rect 14372 13923 14424 13932
rect 14372 13889 14381 13923
rect 14381 13889 14415 13923
rect 14415 13889 14424 13923
rect 14372 13880 14424 13889
rect 11704 13855 11756 13864
rect 2688 13719 2740 13728
rect 2688 13685 2697 13719
rect 2697 13685 2731 13719
rect 2731 13685 2740 13719
rect 2688 13676 2740 13685
rect 4528 13719 4580 13728
rect 4528 13685 4537 13719
rect 4537 13685 4571 13719
rect 4571 13685 4580 13719
rect 6368 13744 6420 13796
rect 11704 13821 11713 13855
rect 11713 13821 11747 13855
rect 11747 13821 11756 13855
rect 11704 13812 11756 13821
rect 15292 13812 15344 13864
rect 18144 13957 18153 13991
rect 18153 13957 18187 13991
rect 18187 13957 18196 13991
rect 18144 13948 18196 13957
rect 16764 13880 16816 13932
rect 18972 13880 19024 13932
rect 19248 13880 19300 13932
rect 18788 13812 18840 13864
rect 20812 13812 20864 13864
rect 4528 13676 4580 13685
rect 5264 13676 5316 13728
rect 7656 13676 7708 13728
rect 8668 13719 8720 13728
rect 8668 13685 8677 13719
rect 8677 13685 8711 13719
rect 8711 13685 8720 13719
rect 8668 13676 8720 13685
rect 9680 13719 9732 13728
rect 9680 13685 9689 13719
rect 9689 13685 9723 13719
rect 9723 13685 9732 13719
rect 9680 13676 9732 13685
rect 9772 13719 9824 13728
rect 9772 13685 9781 13719
rect 9781 13685 9815 13719
rect 9815 13685 9824 13719
rect 11888 13744 11940 13796
rect 15476 13744 15528 13796
rect 19432 13744 19484 13796
rect 19984 13744 20036 13796
rect 20444 13744 20496 13796
rect 9772 13676 9824 13685
rect 11152 13676 11204 13728
rect 14188 13719 14240 13728
rect 14188 13685 14197 13719
rect 14197 13685 14231 13719
rect 14231 13685 14240 13719
rect 14188 13676 14240 13685
rect 15844 13676 15896 13728
rect 16212 13719 16264 13728
rect 16212 13685 16221 13719
rect 16221 13685 16255 13719
rect 16255 13685 16264 13719
rect 16212 13676 16264 13685
rect 16304 13719 16356 13728
rect 16304 13685 16313 13719
rect 16313 13685 16347 13719
rect 16347 13685 16356 13719
rect 17224 13719 17276 13728
rect 16304 13676 16356 13685
rect 17224 13685 17233 13719
rect 17233 13685 17267 13719
rect 17267 13685 17276 13719
rect 17224 13676 17276 13685
rect 19340 13719 19392 13728
rect 19340 13685 19349 13719
rect 19349 13685 19383 13719
rect 19383 13685 19392 13719
rect 19340 13676 19392 13685
rect 20260 13719 20312 13728
rect 20260 13685 20269 13719
rect 20269 13685 20303 13719
rect 20303 13685 20312 13719
rect 20260 13676 20312 13685
rect 7912 13574 7964 13626
rect 7976 13574 8028 13626
rect 8040 13574 8092 13626
rect 8104 13574 8156 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 15035 13574 15087 13626
rect 2688 13472 2740 13524
rect 4252 13472 4304 13524
rect 4528 13472 4580 13524
rect 6184 13472 6236 13524
rect 6920 13472 6972 13524
rect 9772 13472 9824 13524
rect 14188 13472 14240 13524
rect 15292 13515 15344 13524
rect 15292 13481 15301 13515
rect 15301 13481 15335 13515
rect 15335 13481 15344 13515
rect 15292 13472 15344 13481
rect 16304 13515 16356 13524
rect 16304 13481 16313 13515
rect 16313 13481 16347 13515
rect 16347 13481 16356 13515
rect 16304 13472 16356 13481
rect 17224 13472 17276 13524
rect 3148 13404 3200 13456
rect 3700 13336 3752 13388
rect 4344 13404 4396 13456
rect 5080 13404 5132 13456
rect 6368 13404 6420 13456
rect 7012 13404 7064 13456
rect 12624 13447 12676 13456
rect 12624 13413 12633 13447
rect 12633 13413 12667 13447
rect 12667 13413 12676 13447
rect 12624 13404 12676 13413
rect 13268 13404 13320 13456
rect 4988 13336 5040 13388
rect 5448 13336 5500 13388
rect 7104 13379 7156 13388
rect 4804 13268 4856 13320
rect 5264 13268 5316 13320
rect 5172 13200 5224 13252
rect 7104 13345 7113 13379
rect 7113 13345 7147 13379
rect 7147 13345 7156 13379
rect 7104 13336 7156 13345
rect 8208 13336 8260 13388
rect 8300 13379 8352 13388
rect 8300 13345 8309 13379
rect 8309 13345 8343 13379
rect 8343 13345 8352 13379
rect 8300 13336 8352 13345
rect 8760 13336 8812 13388
rect 10048 13379 10100 13388
rect 10048 13345 10057 13379
rect 10057 13345 10091 13379
rect 10091 13345 10100 13379
rect 10048 13336 10100 13345
rect 11244 13336 11296 13388
rect 12808 13336 12860 13388
rect 14096 13379 14148 13388
rect 14096 13345 14105 13379
rect 14105 13345 14139 13379
rect 14139 13345 14148 13379
rect 14096 13336 14148 13345
rect 17408 13404 17460 13456
rect 16672 13379 16724 13388
rect 7196 13311 7248 13320
rect 7196 13277 7205 13311
rect 7205 13277 7239 13311
rect 7239 13277 7248 13311
rect 7196 13268 7248 13277
rect 7472 13268 7524 13320
rect 10140 13311 10192 13320
rect 10140 13277 10149 13311
rect 10149 13277 10183 13311
rect 10183 13277 10192 13311
rect 10140 13268 10192 13277
rect 10232 13311 10284 13320
rect 10232 13277 10241 13311
rect 10241 13277 10275 13311
rect 10275 13277 10284 13311
rect 10232 13268 10284 13277
rect 11152 13268 11204 13320
rect 11796 13311 11848 13320
rect 11796 13277 11805 13311
rect 11805 13277 11839 13311
rect 11839 13277 11848 13311
rect 11796 13268 11848 13277
rect 12900 13268 12952 13320
rect 15752 13311 15804 13320
rect 15752 13277 15761 13311
rect 15761 13277 15795 13311
rect 15795 13277 15804 13311
rect 15752 13268 15804 13277
rect 15936 13311 15988 13320
rect 15936 13277 15945 13311
rect 15945 13277 15979 13311
rect 15979 13277 15988 13311
rect 15936 13268 15988 13277
rect 16672 13345 16681 13379
rect 16681 13345 16715 13379
rect 16715 13345 16724 13379
rect 16672 13336 16724 13345
rect 19340 13472 19392 13524
rect 18788 13379 18840 13388
rect 18788 13345 18797 13379
rect 18797 13345 18831 13379
rect 18831 13345 18840 13379
rect 18788 13336 18840 13345
rect 20812 13404 20864 13456
rect 20720 13336 20772 13388
rect 11888 13200 11940 13252
rect 13912 13243 13964 13252
rect 2136 13175 2188 13184
rect 2136 13141 2145 13175
rect 2145 13141 2179 13175
rect 2179 13141 2188 13175
rect 2136 13132 2188 13141
rect 3148 13132 3200 13184
rect 3424 13175 3476 13184
rect 3424 13141 3433 13175
rect 3433 13141 3467 13175
rect 3467 13141 3476 13175
rect 3424 13132 3476 13141
rect 7656 13132 7708 13184
rect 8300 13132 8352 13184
rect 13636 13132 13688 13184
rect 13912 13209 13921 13243
rect 13921 13209 13955 13243
rect 13955 13209 13964 13243
rect 13912 13200 13964 13209
rect 15568 13200 15620 13252
rect 16488 13200 16540 13252
rect 18604 13268 18656 13320
rect 18880 13311 18932 13320
rect 18880 13277 18889 13311
rect 18889 13277 18923 13311
rect 18923 13277 18932 13311
rect 18880 13268 18932 13277
rect 19156 13268 19208 13320
rect 18696 13200 18748 13252
rect 18972 13200 19024 13252
rect 19984 13311 20036 13320
rect 19984 13277 19993 13311
rect 19993 13277 20027 13311
rect 20027 13277 20036 13311
rect 21088 13311 21140 13320
rect 19984 13268 20036 13277
rect 21088 13277 21097 13311
rect 21097 13277 21131 13311
rect 21131 13277 21140 13311
rect 21088 13268 21140 13277
rect 18144 13132 18196 13184
rect 20260 13132 20312 13184
rect 4447 13030 4499 13082
rect 4511 13030 4563 13082
rect 4575 13030 4627 13082
rect 4639 13030 4691 13082
rect 11378 13030 11430 13082
rect 11442 13030 11494 13082
rect 11506 13030 11558 13082
rect 11570 13030 11622 13082
rect 18308 13030 18360 13082
rect 18372 13030 18424 13082
rect 18436 13030 18488 13082
rect 18500 13030 18552 13082
rect 2504 12928 2556 12980
rect 4160 12928 4212 12980
rect 7380 12971 7432 12980
rect 7380 12937 7389 12971
rect 7389 12937 7423 12971
rect 7423 12937 7432 12971
rect 7380 12928 7432 12937
rect 8668 12928 8720 12980
rect 15660 12971 15712 12980
rect 2964 12792 3016 12844
rect 3608 12792 3660 12844
rect 5172 12835 5224 12844
rect 5172 12801 5181 12835
rect 5181 12801 5215 12835
rect 5215 12801 5224 12835
rect 5172 12792 5224 12801
rect 5448 12792 5500 12844
rect 7472 12792 7524 12844
rect 8116 12792 8168 12844
rect 10416 12860 10468 12912
rect 11152 12903 11204 12912
rect 11152 12869 11161 12903
rect 11161 12869 11195 12903
rect 11195 12869 11204 12903
rect 11152 12860 11204 12869
rect 11244 12860 11296 12912
rect 12900 12860 12952 12912
rect 15660 12937 15669 12971
rect 15669 12937 15703 12971
rect 15703 12937 15712 12971
rect 15660 12928 15712 12937
rect 18788 12928 18840 12980
rect 18880 12928 18932 12980
rect 9864 12792 9916 12844
rect 10140 12792 10192 12844
rect 13084 12792 13136 12844
rect 15752 12860 15804 12912
rect 18604 12860 18656 12912
rect 4068 12724 4120 12776
rect 4712 12656 4764 12708
rect 4988 12699 5040 12708
rect 4988 12665 4997 12699
rect 4997 12665 5031 12699
rect 5031 12665 5040 12699
rect 4988 12656 5040 12665
rect 2596 12631 2648 12640
rect 2596 12597 2605 12631
rect 2605 12597 2639 12631
rect 2639 12597 2648 12631
rect 2596 12588 2648 12597
rect 2688 12631 2740 12640
rect 2688 12597 2697 12631
rect 2697 12597 2731 12631
rect 2731 12597 2740 12631
rect 2688 12588 2740 12597
rect 8576 12724 8628 12776
rect 13360 12724 13412 12776
rect 13820 12724 13872 12776
rect 16488 12792 16540 12844
rect 16672 12724 16724 12776
rect 17132 12792 17184 12844
rect 18052 12792 18104 12844
rect 19156 12860 19208 12912
rect 18696 12767 18748 12776
rect 7656 12656 7708 12708
rect 8116 12656 8168 12708
rect 10600 12656 10652 12708
rect 11888 12656 11940 12708
rect 8484 12588 8536 12640
rect 9680 12588 9732 12640
rect 9956 12588 10008 12640
rect 12440 12631 12492 12640
rect 12440 12597 12449 12631
rect 12449 12597 12483 12631
rect 12483 12597 12492 12631
rect 12440 12588 12492 12597
rect 13912 12588 13964 12640
rect 14188 12656 14240 12708
rect 17684 12656 17736 12708
rect 18696 12733 18705 12767
rect 18705 12733 18739 12767
rect 18739 12733 18748 12767
rect 18696 12724 18748 12733
rect 19708 12792 19760 12844
rect 19984 12792 20036 12844
rect 20260 12792 20312 12844
rect 20996 12767 21048 12776
rect 20996 12733 21005 12767
rect 21005 12733 21039 12767
rect 21039 12733 21048 12767
rect 20996 12724 21048 12733
rect 19524 12656 19576 12708
rect 18052 12588 18104 12640
rect 18144 12588 18196 12640
rect 19248 12588 19300 12640
rect 19340 12588 19392 12640
rect 20536 12631 20588 12640
rect 20536 12597 20545 12631
rect 20545 12597 20579 12631
rect 20579 12597 20588 12631
rect 20536 12588 20588 12597
rect 20904 12631 20956 12640
rect 20904 12597 20913 12631
rect 20913 12597 20947 12631
rect 20947 12597 20956 12631
rect 20904 12588 20956 12597
rect 7912 12486 7964 12538
rect 7976 12486 8028 12538
rect 8040 12486 8092 12538
rect 8104 12486 8156 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 15035 12486 15087 12538
rect 2688 12384 2740 12436
rect 4712 12427 4764 12436
rect 4712 12393 4721 12427
rect 4721 12393 4755 12427
rect 4755 12393 4764 12427
rect 4712 12384 4764 12393
rect 3332 12248 3384 12300
rect 4344 12248 4396 12300
rect 7196 12427 7248 12436
rect 7196 12393 7205 12427
rect 7205 12393 7239 12427
rect 7239 12393 7248 12427
rect 7196 12384 7248 12393
rect 9680 12427 9732 12436
rect 9680 12393 9689 12427
rect 9689 12393 9723 12427
rect 9723 12393 9732 12427
rect 9680 12384 9732 12393
rect 5540 12316 5592 12368
rect 10692 12384 10744 12436
rect 12900 12384 12952 12436
rect 13360 12384 13412 12436
rect 14188 12427 14240 12436
rect 6460 12248 6512 12300
rect 10968 12316 11020 12368
rect 12716 12316 12768 12368
rect 13820 12316 13872 12368
rect 14188 12393 14197 12427
rect 14197 12393 14231 12427
rect 14231 12393 14240 12427
rect 14188 12384 14240 12393
rect 16212 12384 16264 12436
rect 16764 12384 16816 12436
rect 17132 12384 17184 12436
rect 18052 12427 18104 12436
rect 18052 12393 18061 12427
rect 18061 12393 18095 12427
rect 18095 12393 18104 12427
rect 18052 12384 18104 12393
rect 18604 12384 18656 12436
rect 18972 12384 19024 12436
rect 19432 12384 19484 12436
rect 21180 12384 21232 12436
rect 16948 12316 17000 12368
rect 5448 12180 5500 12232
rect 7196 12180 7248 12232
rect 7748 12223 7800 12232
rect 7748 12189 7757 12223
rect 7757 12189 7791 12223
rect 7791 12189 7800 12223
rect 7748 12180 7800 12189
rect 3792 12044 3844 12096
rect 6644 12112 6696 12164
rect 9956 12112 10008 12164
rect 6460 12087 6512 12096
rect 6460 12053 6469 12087
rect 6469 12053 6503 12087
rect 6503 12053 6512 12087
rect 6460 12044 6512 12053
rect 6736 12044 6788 12096
rect 11152 12248 11204 12300
rect 11612 12248 11664 12300
rect 10232 12223 10284 12232
rect 10232 12189 10241 12223
rect 10241 12189 10275 12223
rect 10275 12189 10284 12223
rect 10232 12180 10284 12189
rect 12900 12248 12952 12300
rect 12164 12112 12216 12164
rect 12256 12044 12308 12096
rect 12716 12112 12768 12164
rect 15936 12248 15988 12300
rect 18144 12248 18196 12300
rect 15660 12112 15712 12164
rect 19248 12316 19300 12368
rect 18604 12223 18656 12232
rect 18604 12189 18613 12223
rect 18613 12189 18647 12223
rect 18647 12189 18656 12223
rect 18604 12180 18656 12189
rect 21088 12248 21140 12300
rect 19984 12223 20036 12232
rect 19248 12112 19300 12164
rect 19708 12112 19760 12164
rect 19984 12189 19993 12223
rect 19993 12189 20027 12223
rect 20027 12189 20036 12223
rect 19984 12180 20036 12189
rect 14648 12044 14700 12096
rect 19892 12044 19944 12096
rect 20720 12044 20772 12096
rect 20996 12044 21048 12096
rect 4447 11942 4499 11994
rect 4511 11942 4563 11994
rect 4575 11942 4627 11994
rect 4639 11942 4691 11994
rect 11378 11942 11430 11994
rect 11442 11942 11494 11994
rect 11506 11942 11558 11994
rect 11570 11942 11622 11994
rect 18308 11942 18360 11994
rect 18372 11942 18424 11994
rect 18436 11942 18488 11994
rect 18500 11942 18552 11994
rect 2872 11840 2924 11892
rect 3608 11883 3660 11892
rect 3608 11849 3617 11883
rect 3617 11849 3651 11883
rect 3651 11849 3660 11883
rect 3608 11840 3660 11849
rect 7104 11840 7156 11892
rect 8484 11883 8536 11892
rect 8484 11849 8493 11883
rect 8493 11849 8527 11883
rect 8527 11849 8536 11883
rect 8484 11840 8536 11849
rect 9772 11840 9824 11892
rect 11888 11840 11940 11892
rect 12624 11840 12676 11892
rect 14648 11840 14700 11892
rect 14740 11840 14792 11892
rect 20720 11840 20772 11892
rect 4068 11772 4120 11824
rect 12532 11772 12584 11824
rect 19064 11772 19116 11824
rect 3516 11704 3568 11756
rect 6920 11704 6972 11756
rect 7748 11704 7800 11756
rect 10232 11704 10284 11756
rect 11152 11747 11204 11756
rect 11152 11713 11161 11747
rect 11161 11713 11195 11747
rect 11195 11713 11204 11747
rect 11152 11704 11204 11713
rect 13912 11747 13964 11756
rect 1952 11636 2004 11688
rect 2320 11636 2372 11688
rect 3240 11636 3292 11688
rect 3884 11636 3936 11688
rect 5080 11636 5132 11688
rect 7196 11679 7248 11688
rect 7196 11645 7205 11679
rect 7205 11645 7239 11679
rect 7239 11645 7248 11679
rect 7196 11636 7248 11645
rect 8300 11636 8352 11688
rect 11980 11636 12032 11688
rect 2872 11568 2924 11620
rect 3608 11500 3660 11552
rect 4344 11543 4396 11552
rect 4344 11509 4353 11543
rect 4353 11509 4387 11543
rect 4387 11509 4396 11543
rect 4344 11500 4396 11509
rect 7104 11500 7156 11552
rect 7564 11500 7616 11552
rect 8852 11543 8904 11552
rect 8852 11509 8861 11543
rect 8861 11509 8895 11543
rect 8895 11509 8904 11543
rect 8852 11500 8904 11509
rect 9128 11500 9180 11552
rect 11796 11568 11848 11620
rect 12164 11568 12216 11620
rect 12348 11568 12400 11620
rect 13912 11713 13921 11747
rect 13921 11713 13955 11747
rect 13955 11713 13964 11747
rect 13912 11704 13964 11713
rect 14188 11704 14240 11756
rect 17408 11704 17460 11756
rect 17960 11704 18012 11756
rect 13728 11636 13780 11688
rect 17776 11636 17828 11688
rect 18236 11704 18288 11756
rect 18604 11747 18656 11756
rect 18604 11713 18613 11747
rect 18613 11713 18647 11747
rect 18647 11713 18656 11747
rect 18604 11704 18656 11713
rect 19340 11704 19392 11756
rect 19892 11704 19944 11756
rect 18420 11679 18472 11688
rect 13636 11568 13688 11620
rect 16764 11568 16816 11620
rect 18420 11645 18429 11679
rect 18429 11645 18463 11679
rect 18463 11645 18472 11679
rect 18420 11636 18472 11645
rect 18512 11636 18564 11688
rect 9956 11543 10008 11552
rect 9956 11509 9965 11543
rect 9965 11509 9999 11543
rect 9999 11509 10008 11543
rect 9956 11500 10008 11509
rect 11888 11543 11940 11552
rect 11888 11509 11897 11543
rect 11897 11509 11931 11543
rect 11931 11509 11940 11543
rect 11888 11500 11940 11509
rect 11980 11500 12032 11552
rect 18236 11568 18288 11620
rect 20996 11636 21048 11688
rect 20260 11611 20312 11620
rect 20260 11577 20294 11611
rect 20294 11577 20312 11611
rect 20260 11568 20312 11577
rect 20628 11568 20680 11620
rect 17684 11500 17736 11552
rect 18144 11500 18196 11552
rect 18972 11500 19024 11552
rect 19248 11500 19300 11552
rect 21364 11543 21416 11552
rect 21364 11509 21373 11543
rect 21373 11509 21407 11543
rect 21407 11509 21416 11543
rect 21364 11500 21416 11509
rect 7912 11398 7964 11450
rect 7976 11398 8028 11450
rect 8040 11398 8092 11450
rect 8104 11398 8156 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 15035 11398 15087 11450
rect 2596 11296 2648 11348
rect 2872 11296 2924 11348
rect 3240 11339 3292 11348
rect 3240 11305 3249 11339
rect 3249 11305 3283 11339
rect 3283 11305 3292 11339
rect 3240 11296 3292 11305
rect 5448 11296 5500 11348
rect 6920 11339 6972 11348
rect 6920 11305 6929 11339
rect 6929 11305 6963 11339
rect 6963 11305 6972 11339
rect 6920 11296 6972 11305
rect 8852 11296 8904 11348
rect 1952 11271 2004 11280
rect 1952 11237 1961 11271
rect 1961 11237 1995 11271
rect 1995 11237 2004 11271
rect 1952 11228 2004 11237
rect 4896 11228 4948 11280
rect 5080 11228 5132 11280
rect 14740 11296 14792 11348
rect 15200 11296 15252 11348
rect 17592 11296 17644 11348
rect 1584 11092 1636 11144
rect 2964 11160 3016 11212
rect 5172 11160 5224 11212
rect 6644 11160 6696 11212
rect 4160 11092 4212 11144
rect 3516 11067 3568 11076
rect 3516 11033 3525 11067
rect 3525 11033 3559 11067
rect 3559 11033 3568 11067
rect 3516 11024 3568 11033
rect 3700 10956 3752 11008
rect 6828 11092 6880 11144
rect 7748 11160 7800 11212
rect 8024 11135 8076 11144
rect 8024 11101 8033 11135
rect 8033 11101 8067 11135
rect 8067 11101 8076 11135
rect 8024 11092 8076 11101
rect 13084 11228 13136 11280
rect 14556 11228 14608 11280
rect 12440 11160 12492 11212
rect 12532 11160 12584 11212
rect 15200 11160 15252 11212
rect 15936 11160 15988 11212
rect 7288 11024 7340 11076
rect 8208 11024 8260 11076
rect 9128 11024 9180 11076
rect 13360 11092 13412 11144
rect 13636 11092 13688 11144
rect 19064 11296 19116 11348
rect 20904 11296 20956 11348
rect 18788 11228 18840 11280
rect 19156 11228 19208 11280
rect 18052 11203 18104 11212
rect 18052 11169 18061 11203
rect 18061 11169 18095 11203
rect 18095 11169 18104 11203
rect 18052 11160 18104 11169
rect 17960 11092 18012 11144
rect 18144 11135 18196 11144
rect 18144 11101 18153 11135
rect 18153 11101 18187 11135
rect 18187 11101 18196 11135
rect 18144 11092 18196 11101
rect 14648 11024 14700 11076
rect 16672 11067 16724 11076
rect 16672 11033 16681 11067
rect 16681 11033 16715 11067
rect 16715 11033 16724 11067
rect 16672 11024 16724 11033
rect 16856 11024 16908 11076
rect 19708 11160 19760 11212
rect 19156 11092 19208 11144
rect 19892 11135 19944 11144
rect 19892 11101 19901 11135
rect 19901 11101 19935 11135
rect 19935 11101 19944 11135
rect 19892 11092 19944 11101
rect 20260 11092 20312 11144
rect 20444 11092 20496 11144
rect 19248 11067 19300 11076
rect 19248 11033 19257 11067
rect 19257 11033 19291 11067
rect 19291 11033 19300 11067
rect 19248 11024 19300 11033
rect 19524 11024 19576 11076
rect 20076 11024 20128 11076
rect 6552 10999 6604 11008
rect 6552 10965 6561 10999
rect 6561 10965 6595 10999
rect 6595 10965 6604 10999
rect 6552 10956 6604 10965
rect 6920 10956 6972 11008
rect 12808 10999 12860 11008
rect 12808 10965 12817 10999
rect 12817 10965 12851 10999
rect 12851 10965 12860 10999
rect 12808 10956 12860 10965
rect 15476 10956 15528 11008
rect 18880 10956 18932 11008
rect 4447 10854 4499 10906
rect 4511 10854 4563 10906
rect 4575 10854 4627 10906
rect 4639 10854 4691 10906
rect 11378 10854 11430 10906
rect 11442 10854 11494 10906
rect 11506 10854 11558 10906
rect 11570 10854 11622 10906
rect 18308 10854 18360 10906
rect 18372 10854 18424 10906
rect 18436 10854 18488 10906
rect 18500 10854 18552 10906
rect 1584 10795 1636 10804
rect 1584 10761 1593 10795
rect 1593 10761 1627 10795
rect 1627 10761 1636 10795
rect 1584 10752 1636 10761
rect 2780 10795 2832 10804
rect 2780 10761 2789 10795
rect 2789 10761 2823 10795
rect 2823 10761 2832 10795
rect 2780 10752 2832 10761
rect 4068 10752 4120 10804
rect 5172 10752 5224 10804
rect 12532 10795 12584 10804
rect 8024 10684 8076 10736
rect 1860 10591 1912 10600
rect 1860 10557 1869 10591
rect 1869 10557 1903 10591
rect 1903 10557 1912 10591
rect 1860 10548 1912 10557
rect 6644 10616 6696 10668
rect 12532 10761 12541 10795
rect 12541 10761 12575 10795
rect 12575 10761 12584 10795
rect 12532 10752 12584 10761
rect 13360 10752 13412 10804
rect 16028 10752 16080 10804
rect 19984 10752 20036 10804
rect 20628 10795 20680 10804
rect 20628 10761 20637 10795
rect 20637 10761 20671 10795
rect 20671 10761 20680 10795
rect 20628 10752 20680 10761
rect 10784 10684 10836 10736
rect 14096 10684 14148 10736
rect 6552 10548 6604 10600
rect 6920 10480 6972 10532
rect 4160 10412 4212 10464
rect 5724 10455 5776 10464
rect 5724 10421 5733 10455
rect 5733 10421 5767 10455
rect 5767 10421 5776 10455
rect 5724 10412 5776 10421
rect 10140 10659 10192 10668
rect 10140 10625 10149 10659
rect 10149 10625 10183 10659
rect 10183 10625 10192 10659
rect 10140 10616 10192 10625
rect 14740 10616 14792 10668
rect 18144 10616 18196 10668
rect 7288 10591 7340 10600
rect 7288 10557 7322 10591
rect 7322 10557 7340 10591
rect 7288 10548 7340 10557
rect 12440 10548 12492 10600
rect 14556 10548 14608 10600
rect 17684 10548 17736 10600
rect 17868 10548 17920 10600
rect 18604 10659 18656 10668
rect 18604 10625 18613 10659
rect 18613 10625 18647 10659
rect 18647 10625 18656 10659
rect 18604 10616 18656 10625
rect 19064 10548 19116 10600
rect 8300 10412 8352 10464
rect 13820 10480 13872 10532
rect 19156 10480 19208 10532
rect 14004 10455 14056 10464
rect 14004 10421 14013 10455
rect 14013 10421 14047 10455
rect 14047 10421 14056 10455
rect 14004 10412 14056 10421
rect 14372 10455 14424 10464
rect 14372 10421 14381 10455
rect 14381 10421 14415 10455
rect 14415 10421 14424 10455
rect 14372 10412 14424 10421
rect 17132 10455 17184 10464
rect 17132 10421 17141 10455
rect 17141 10421 17175 10455
rect 17175 10421 17184 10455
rect 17132 10412 17184 10421
rect 18144 10412 18196 10464
rect 7912 10310 7964 10362
rect 7976 10310 8028 10362
rect 8040 10310 8092 10362
rect 8104 10310 8156 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 15035 10310 15087 10362
rect 1860 10208 1912 10260
rect 4896 10251 4948 10260
rect 4896 10217 4905 10251
rect 4905 10217 4939 10251
rect 4939 10217 4948 10251
rect 4896 10208 4948 10217
rect 7748 10208 7800 10260
rect 14372 10208 14424 10260
rect 4068 10140 4120 10192
rect 14556 10140 14608 10192
rect 14648 10140 14700 10192
rect 17868 10140 17920 10192
rect 2688 10115 2740 10124
rect 2688 10081 2697 10115
rect 2697 10081 2731 10115
rect 2731 10081 2740 10115
rect 2688 10072 2740 10081
rect 5724 10072 5776 10124
rect 6460 10072 6512 10124
rect 2780 10047 2832 10056
rect 2780 10013 2789 10047
rect 2789 10013 2823 10047
rect 2823 10013 2832 10047
rect 2780 10004 2832 10013
rect 3424 10004 3476 10056
rect 5172 10004 5224 10056
rect 6368 10047 6420 10056
rect 6368 10013 6377 10047
rect 6377 10013 6411 10047
rect 6411 10013 6420 10047
rect 6368 10004 6420 10013
rect 6644 10004 6696 10056
rect 2412 9936 2464 9988
rect 6920 9936 6972 9988
rect 7288 9936 7340 9988
rect 8300 10072 8352 10124
rect 10232 10072 10284 10124
rect 11244 10072 11296 10124
rect 13084 10072 13136 10124
rect 15660 10115 15712 10124
rect 12992 10047 13044 10056
rect 10968 9868 11020 9920
rect 12992 10013 13001 10047
rect 13001 10013 13035 10047
rect 13035 10013 13044 10047
rect 12992 10004 13044 10013
rect 15660 10081 15669 10115
rect 15669 10081 15703 10115
rect 15703 10081 15712 10115
rect 15660 10072 15712 10081
rect 16580 10072 16632 10124
rect 16764 10115 16816 10124
rect 16764 10081 16798 10115
rect 16798 10081 16816 10115
rect 16764 10072 16816 10081
rect 18604 10140 18656 10192
rect 19156 10208 19208 10260
rect 20260 10183 20312 10192
rect 20260 10149 20269 10183
rect 20269 10149 20303 10183
rect 20303 10149 20312 10183
rect 20260 10140 20312 10149
rect 20904 10072 20956 10124
rect 16212 9936 16264 9988
rect 20720 10004 20772 10056
rect 21364 10004 21416 10056
rect 12716 9911 12768 9920
rect 12716 9877 12725 9911
rect 12725 9877 12759 9911
rect 12759 9877 12768 9911
rect 12716 9868 12768 9877
rect 14740 9868 14792 9920
rect 16672 9868 16724 9920
rect 19708 9868 19760 9920
rect 4447 9766 4499 9818
rect 4511 9766 4563 9818
rect 4575 9766 4627 9818
rect 4639 9766 4691 9818
rect 11378 9766 11430 9818
rect 11442 9766 11494 9818
rect 11506 9766 11558 9818
rect 11570 9766 11622 9818
rect 18308 9766 18360 9818
rect 18372 9766 18424 9818
rect 18436 9766 18488 9818
rect 18500 9766 18552 9818
rect 4068 9664 4120 9716
rect 6368 9664 6420 9716
rect 12532 9664 12584 9716
rect 17868 9664 17920 9716
rect 9496 9596 9548 9648
rect 16856 9596 16908 9648
rect 18052 9639 18104 9648
rect 18052 9605 18061 9639
rect 18061 9605 18095 9639
rect 18095 9605 18104 9639
rect 18052 9596 18104 9605
rect 7288 9528 7340 9580
rect 9956 9528 10008 9580
rect 10140 9571 10192 9580
rect 10140 9537 10149 9571
rect 10149 9537 10183 9571
rect 10183 9537 10192 9571
rect 10140 9528 10192 9537
rect 11244 9528 11296 9580
rect 14096 9528 14148 9580
rect 8208 9460 8260 9512
rect 2872 9392 2924 9444
rect 3976 9392 4028 9444
rect 9588 9460 9640 9512
rect 2504 9324 2556 9376
rect 3424 9367 3476 9376
rect 3424 9333 3433 9367
rect 3433 9333 3467 9367
rect 3467 9333 3476 9367
rect 3424 9324 3476 9333
rect 6460 9367 6512 9376
rect 6460 9333 6469 9367
rect 6469 9333 6503 9367
rect 6503 9333 6512 9367
rect 6460 9324 6512 9333
rect 6828 9324 6880 9376
rect 7380 9324 7432 9376
rect 8208 9324 8260 9376
rect 8392 9367 8444 9376
rect 8392 9333 8401 9367
rect 8401 9333 8435 9367
rect 8435 9333 8444 9367
rect 8392 9324 8444 9333
rect 9404 9367 9456 9376
rect 9404 9333 9413 9367
rect 9413 9333 9447 9367
rect 9447 9333 9456 9367
rect 9404 9324 9456 9333
rect 12992 9460 13044 9512
rect 9772 9392 9824 9444
rect 10324 9392 10376 9444
rect 9956 9367 10008 9376
rect 9956 9333 9965 9367
rect 9965 9333 9999 9367
rect 9999 9333 10008 9367
rect 9956 9324 10008 9333
rect 10784 9324 10836 9376
rect 11796 9392 11848 9444
rect 14740 9460 14792 9512
rect 15660 9528 15712 9580
rect 16212 9571 16264 9580
rect 16212 9537 16221 9571
rect 16221 9537 16255 9571
rect 16255 9537 16264 9571
rect 16212 9528 16264 9537
rect 18328 9528 18380 9580
rect 18604 9571 18656 9580
rect 18604 9537 18613 9571
rect 18613 9537 18647 9571
rect 18647 9537 18656 9571
rect 18604 9528 18656 9537
rect 17592 9503 17644 9512
rect 12624 9324 12676 9376
rect 13728 9392 13780 9444
rect 17592 9469 17601 9503
rect 17601 9469 17635 9503
rect 17635 9469 17644 9503
rect 17592 9460 17644 9469
rect 18144 9460 18196 9512
rect 20720 9460 20772 9512
rect 14556 9324 14608 9376
rect 15200 9324 15252 9376
rect 15660 9367 15712 9376
rect 15660 9333 15669 9367
rect 15669 9333 15703 9367
rect 15703 9333 15712 9367
rect 15660 9324 15712 9333
rect 16856 9324 16908 9376
rect 18788 9324 18840 9376
rect 19984 9324 20036 9376
rect 7912 9222 7964 9274
rect 7976 9222 8028 9274
rect 8040 9222 8092 9274
rect 8104 9222 8156 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 15035 9222 15087 9274
rect 2688 9120 2740 9172
rect 4988 9120 5040 9172
rect 2504 9052 2556 9104
rect 2596 9027 2648 9036
rect 2596 8993 2605 9027
rect 2605 8993 2639 9027
rect 2639 8993 2648 9027
rect 2596 8984 2648 8993
rect 2688 8959 2740 8968
rect 2688 8925 2697 8959
rect 2697 8925 2731 8959
rect 2731 8925 2740 8959
rect 2688 8916 2740 8925
rect 2872 8959 2924 8968
rect 2872 8925 2881 8959
rect 2881 8925 2915 8959
rect 2915 8925 2924 8959
rect 2872 8916 2924 8925
rect 3424 9052 3476 9104
rect 7196 9120 7248 9172
rect 7380 9163 7432 9172
rect 7380 9129 7389 9163
rect 7389 9129 7423 9163
rect 7423 9129 7432 9163
rect 7380 9120 7432 9129
rect 7748 9120 7800 9172
rect 8852 9120 8904 9172
rect 9312 9120 9364 9172
rect 9956 9120 10008 9172
rect 10324 9120 10376 9172
rect 7472 9052 7524 9104
rect 15660 9120 15712 9172
rect 20536 9120 20588 9172
rect 20904 9163 20956 9172
rect 20904 9129 20913 9163
rect 20913 9129 20947 9163
rect 20947 9129 20956 9163
rect 20904 9120 20956 9129
rect 4160 8984 4212 9036
rect 6552 8984 6604 9036
rect 7288 8984 7340 9036
rect 5448 8916 5500 8968
rect 6920 8916 6972 8968
rect 7380 8916 7432 8968
rect 8392 8916 8444 8968
rect 8668 8916 8720 8968
rect 9496 8984 9548 9036
rect 9864 8984 9916 9036
rect 10048 9027 10100 9036
rect 10048 8993 10057 9027
rect 10057 8993 10091 9027
rect 10091 8993 10100 9027
rect 10048 8984 10100 8993
rect 10324 8984 10376 9036
rect 11152 9027 11204 9036
rect 11152 8993 11161 9027
rect 11161 8993 11195 9027
rect 11195 8993 11204 9027
rect 11152 8984 11204 8993
rect 8760 8848 8812 8900
rect 9312 8848 9364 8900
rect 10968 8916 11020 8968
rect 19156 9052 19208 9104
rect 20076 9052 20128 9104
rect 21180 9052 21232 9104
rect 11428 8984 11480 9036
rect 11796 9027 11848 9036
rect 11796 8993 11805 9027
rect 11805 8993 11839 9027
rect 11839 8993 11848 9027
rect 11796 8984 11848 8993
rect 15200 8984 15252 9036
rect 13084 8916 13136 8968
rect 14740 8959 14792 8968
rect 14740 8925 14749 8959
rect 14749 8925 14783 8959
rect 14783 8925 14792 8959
rect 14740 8916 14792 8925
rect 13820 8848 13872 8900
rect 16396 8848 16448 8900
rect 19064 8848 19116 8900
rect 13084 8780 13136 8832
rect 13728 8823 13780 8832
rect 13728 8789 13737 8823
rect 13737 8789 13771 8823
rect 13771 8789 13780 8823
rect 13728 8780 13780 8789
rect 14464 8780 14516 8832
rect 16580 8780 16632 8832
rect 16672 8780 16724 8832
rect 20720 8916 20772 8968
rect 19800 8823 19852 8832
rect 19800 8789 19809 8823
rect 19809 8789 19843 8823
rect 19843 8789 19852 8823
rect 19800 8780 19852 8789
rect 4447 8678 4499 8730
rect 4511 8678 4563 8730
rect 4575 8678 4627 8730
rect 4639 8678 4691 8730
rect 11378 8678 11430 8730
rect 11442 8678 11494 8730
rect 11506 8678 11558 8730
rect 11570 8678 11622 8730
rect 18308 8678 18360 8730
rect 18372 8678 18424 8730
rect 18436 8678 18488 8730
rect 18500 8678 18552 8730
rect 2872 8576 2924 8628
rect 4896 8576 4948 8628
rect 5448 8576 5500 8628
rect 6828 8619 6880 8628
rect 6828 8585 6837 8619
rect 6837 8585 6871 8619
rect 6871 8585 6880 8619
rect 6828 8576 6880 8585
rect 7288 8576 7340 8628
rect 9772 8576 9824 8628
rect 10140 8619 10192 8628
rect 10140 8585 10149 8619
rect 10149 8585 10183 8619
rect 10183 8585 10192 8619
rect 10140 8576 10192 8585
rect 10600 8619 10652 8628
rect 10600 8585 10609 8619
rect 10609 8585 10643 8619
rect 10643 8585 10652 8619
rect 10600 8576 10652 8585
rect 11704 8576 11756 8628
rect 16672 8576 16724 8628
rect 16764 8576 16816 8628
rect 17500 8576 17552 8628
rect 4344 8508 4396 8560
rect 4620 8508 4672 8560
rect 5540 8440 5592 8492
rect 6184 8440 6236 8492
rect 8668 8508 8720 8560
rect 11428 8508 11480 8560
rect 16488 8508 16540 8560
rect 7472 8483 7524 8492
rect 7472 8449 7481 8483
rect 7481 8449 7515 8483
rect 7515 8449 7524 8483
rect 7472 8440 7524 8449
rect 8300 8440 8352 8492
rect 11244 8440 11296 8492
rect 12716 8440 12768 8492
rect 12992 8440 13044 8492
rect 14464 8483 14516 8492
rect 14464 8449 14473 8483
rect 14473 8449 14507 8483
rect 14507 8449 14516 8483
rect 14464 8440 14516 8449
rect 14832 8440 14884 8492
rect 2504 8372 2556 8424
rect 4988 8372 5040 8424
rect 8208 8372 8260 8424
rect 9312 8372 9364 8424
rect 10600 8372 10652 8424
rect 13176 8415 13228 8424
rect 13176 8381 13185 8415
rect 13185 8381 13219 8415
rect 13219 8381 13228 8415
rect 13176 8372 13228 8381
rect 14004 8372 14056 8424
rect 19524 8508 19576 8560
rect 18144 8440 18196 8492
rect 19800 8483 19852 8492
rect 19800 8449 19809 8483
rect 19809 8449 19843 8483
rect 19843 8449 19852 8483
rect 19800 8440 19852 8449
rect 19984 8483 20036 8492
rect 19984 8449 19993 8483
rect 19993 8449 20027 8483
rect 20027 8449 20036 8483
rect 19984 8440 20036 8449
rect 19708 8415 19760 8424
rect 3056 8304 3108 8356
rect 5080 8304 5132 8356
rect 12532 8304 12584 8356
rect 13084 8347 13136 8356
rect 13084 8313 13093 8347
rect 13093 8313 13127 8347
rect 13127 8313 13136 8347
rect 13084 8304 13136 8313
rect 13728 8304 13780 8356
rect 19708 8381 19717 8415
rect 19717 8381 19751 8415
rect 19751 8381 19760 8415
rect 19708 8372 19760 8381
rect 16212 8304 16264 8356
rect 16672 8304 16724 8356
rect 19616 8304 19668 8356
rect 2320 8236 2372 8288
rect 3608 8236 3660 8288
rect 6920 8236 6972 8288
rect 11336 8279 11388 8288
rect 11336 8245 11345 8279
rect 11345 8245 11379 8279
rect 11379 8245 11388 8279
rect 11336 8236 11388 8245
rect 11428 8236 11480 8288
rect 12256 8236 12308 8288
rect 12716 8279 12768 8288
rect 12716 8245 12725 8279
rect 12725 8245 12759 8279
rect 12759 8245 12768 8279
rect 12716 8236 12768 8245
rect 14188 8236 14240 8288
rect 14648 8236 14700 8288
rect 17776 8236 17828 8288
rect 18052 8279 18104 8288
rect 18052 8245 18061 8279
rect 18061 8245 18095 8279
rect 18095 8245 18104 8279
rect 18052 8236 18104 8245
rect 18420 8279 18472 8288
rect 18420 8245 18429 8279
rect 18429 8245 18463 8279
rect 18463 8245 18472 8279
rect 18420 8236 18472 8245
rect 7912 8134 7964 8186
rect 7976 8134 8028 8186
rect 8040 8134 8092 8186
rect 8104 8134 8156 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 15035 8134 15087 8186
rect 1584 8032 1636 8084
rect 2688 8032 2740 8084
rect 2780 8032 2832 8084
rect 4344 8032 4396 8084
rect 8300 8032 8352 8084
rect 11336 8032 11388 8084
rect 12716 8032 12768 8084
rect 13176 8032 13228 8084
rect 14648 8032 14700 8084
rect 16488 8032 16540 8084
rect 16580 8032 16632 8084
rect 17868 8032 17920 8084
rect 9864 7964 9916 8016
rect 12992 8007 13044 8016
rect 12992 7973 13026 8007
rect 13026 7973 13044 8007
rect 12992 7964 13044 7973
rect 18144 8032 18196 8084
rect 18420 8032 18472 8084
rect 1676 7896 1728 7948
rect 4252 7896 4304 7948
rect 8208 7939 8260 7948
rect 8208 7905 8217 7939
rect 8217 7905 8251 7939
rect 8251 7905 8260 7939
rect 8208 7896 8260 7905
rect 12808 7896 12860 7948
rect 3056 7871 3108 7880
rect 3056 7837 3065 7871
rect 3065 7837 3099 7871
rect 3099 7837 3108 7871
rect 3056 7828 3108 7837
rect 3424 7871 3476 7880
rect 3424 7837 3433 7871
rect 3433 7837 3467 7871
rect 3467 7837 3476 7871
rect 3424 7828 3476 7837
rect 4620 7871 4672 7880
rect 4620 7837 4629 7871
rect 4629 7837 4663 7871
rect 4663 7837 4672 7871
rect 4620 7828 4672 7837
rect 5264 7828 5316 7880
rect 5724 7871 5776 7880
rect 5724 7837 5733 7871
rect 5733 7837 5767 7871
rect 5767 7837 5776 7871
rect 5724 7828 5776 7837
rect 1308 7692 1360 7744
rect 3332 7760 3384 7812
rect 4068 7760 4120 7812
rect 11152 7828 11204 7880
rect 11244 7828 11296 7880
rect 16212 7871 16264 7880
rect 6828 7692 6880 7744
rect 6920 7692 6972 7744
rect 7748 7760 7800 7812
rect 9220 7692 9272 7744
rect 9496 7692 9548 7744
rect 10048 7692 10100 7744
rect 10968 7692 11020 7744
rect 11704 7735 11756 7744
rect 11704 7701 11713 7735
rect 11713 7701 11747 7735
rect 11747 7701 11756 7735
rect 11704 7692 11756 7701
rect 16212 7837 16221 7871
rect 16221 7837 16255 7871
rect 16255 7837 16264 7871
rect 19984 7964 20036 8016
rect 16856 7939 16908 7948
rect 16856 7905 16890 7939
rect 16890 7905 16908 7939
rect 16856 7896 16908 7905
rect 17868 7896 17920 7948
rect 19432 7896 19484 7948
rect 16212 7828 16264 7837
rect 16580 7871 16632 7880
rect 16580 7837 16589 7871
rect 16589 7837 16623 7871
rect 16623 7837 16632 7871
rect 16580 7828 16632 7837
rect 14832 7735 14884 7744
rect 14832 7701 14841 7735
rect 14841 7701 14875 7735
rect 14875 7701 14884 7735
rect 14832 7692 14884 7701
rect 15568 7735 15620 7744
rect 15568 7701 15577 7735
rect 15577 7701 15611 7735
rect 15611 7701 15620 7735
rect 15568 7692 15620 7701
rect 20168 7735 20220 7744
rect 20168 7701 20177 7735
rect 20177 7701 20211 7735
rect 20211 7701 20220 7735
rect 20168 7692 20220 7701
rect 4447 7590 4499 7642
rect 4511 7590 4563 7642
rect 4575 7590 4627 7642
rect 4639 7590 4691 7642
rect 11378 7590 11430 7642
rect 11442 7590 11494 7642
rect 11506 7590 11558 7642
rect 11570 7590 11622 7642
rect 18308 7590 18360 7642
rect 18372 7590 18424 7642
rect 18436 7590 18488 7642
rect 18500 7590 18552 7642
rect 2596 7488 2648 7540
rect 4252 7531 4304 7540
rect 4252 7497 4261 7531
rect 4261 7497 4295 7531
rect 4295 7497 4304 7531
rect 4252 7488 4304 7497
rect 5264 7531 5316 7540
rect 5264 7497 5273 7531
rect 5273 7497 5307 7531
rect 5307 7497 5316 7531
rect 5264 7488 5316 7497
rect 3056 7352 3108 7404
rect 4160 7352 4212 7404
rect 5448 7352 5500 7404
rect 8208 7488 8260 7540
rect 9312 7488 9364 7540
rect 9496 7488 9548 7540
rect 9772 7488 9824 7540
rect 16396 7488 16448 7540
rect 20444 7488 20496 7540
rect 16764 7420 16816 7472
rect 15568 7352 15620 7404
rect 19432 7395 19484 7404
rect 19432 7361 19441 7395
rect 19441 7361 19475 7395
rect 19475 7361 19484 7395
rect 19432 7352 19484 7361
rect 3424 7284 3476 7336
rect 5632 7327 5684 7336
rect 5632 7293 5641 7327
rect 5641 7293 5675 7327
rect 5675 7293 5684 7327
rect 5632 7284 5684 7293
rect 10508 7284 10560 7336
rect 7748 7216 7800 7268
rect 1400 7191 1452 7200
rect 1400 7157 1409 7191
rect 1409 7157 1443 7191
rect 1443 7157 1452 7191
rect 1400 7148 1452 7157
rect 2044 7191 2096 7200
rect 2044 7157 2053 7191
rect 2053 7157 2087 7191
rect 2087 7157 2096 7191
rect 2044 7148 2096 7157
rect 3148 7148 3200 7200
rect 5816 7148 5868 7200
rect 10600 7216 10652 7268
rect 11244 7284 11296 7336
rect 12900 7284 12952 7336
rect 13728 7284 13780 7336
rect 14556 7284 14608 7336
rect 18052 7284 18104 7336
rect 20168 7284 20220 7336
rect 12716 7216 12768 7268
rect 13084 7216 13136 7268
rect 12072 7191 12124 7200
rect 12072 7157 12081 7191
rect 12081 7157 12115 7191
rect 12115 7157 12124 7191
rect 12072 7148 12124 7157
rect 15384 7191 15436 7200
rect 15384 7157 15393 7191
rect 15393 7157 15427 7191
rect 15427 7157 15436 7191
rect 15384 7148 15436 7157
rect 16580 7191 16632 7200
rect 16580 7157 16589 7191
rect 16589 7157 16623 7191
rect 16623 7157 16632 7191
rect 16580 7148 16632 7157
rect 19156 7191 19208 7200
rect 19156 7157 19165 7191
rect 19165 7157 19199 7191
rect 19199 7157 19208 7191
rect 19156 7148 19208 7157
rect 20260 7148 20312 7200
rect 7912 7046 7964 7098
rect 7976 7046 8028 7098
rect 8040 7046 8092 7098
rect 8104 7046 8156 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 15035 7046 15087 7098
rect 1400 6944 1452 6996
rect 4160 6987 4212 6996
rect 4160 6953 4169 6987
rect 4169 6953 4203 6987
rect 4203 6953 4212 6987
rect 4160 6944 4212 6953
rect 5724 6944 5776 6996
rect 7748 6987 7800 6996
rect 1952 6851 2004 6860
rect 1952 6817 1961 6851
rect 1961 6817 1995 6851
rect 1995 6817 2004 6851
rect 1952 6808 2004 6817
rect 2780 6808 2832 6860
rect 4068 6808 4120 6860
rect 4896 6876 4948 6928
rect 5448 6808 5500 6860
rect 7748 6953 7757 6987
rect 7757 6953 7791 6987
rect 7791 6953 7800 6987
rect 7748 6944 7800 6953
rect 9036 6944 9088 6996
rect 10508 6944 10560 6996
rect 11704 6944 11756 6996
rect 12808 6944 12860 6996
rect 12256 6919 12308 6928
rect 6276 6808 6328 6860
rect 7104 6808 7156 6860
rect 9496 6808 9548 6860
rect 12256 6885 12265 6919
rect 12265 6885 12299 6919
rect 12299 6885 12308 6919
rect 12256 6876 12308 6885
rect 12532 6876 12584 6928
rect 14280 6876 14332 6928
rect 14648 6876 14700 6928
rect 16856 6944 16908 6996
rect 19156 6944 19208 6996
rect 10324 6808 10376 6860
rect 12072 6808 12124 6860
rect 3056 6740 3108 6792
rect 1860 6604 1912 6656
rect 3148 6604 3200 6656
rect 9312 6740 9364 6792
rect 8208 6672 8260 6724
rect 10140 6672 10192 6724
rect 13636 6740 13688 6792
rect 16212 6808 16264 6860
rect 15292 6740 15344 6792
rect 18604 6808 18656 6860
rect 19708 6808 19760 6860
rect 20444 6808 20496 6860
rect 9588 6604 9640 6656
rect 10968 6604 11020 6656
rect 11888 6647 11940 6656
rect 11888 6613 11897 6647
rect 11897 6613 11931 6647
rect 11931 6613 11940 6647
rect 11888 6604 11940 6613
rect 17132 6740 17184 6792
rect 18144 6740 18196 6792
rect 18880 6740 18932 6792
rect 20168 6783 20220 6792
rect 20168 6749 20177 6783
rect 20177 6749 20211 6783
rect 20211 6749 20220 6783
rect 20168 6740 20220 6749
rect 20260 6672 20312 6724
rect 16488 6604 16540 6656
rect 18880 6604 18932 6656
rect 4447 6502 4499 6554
rect 4511 6502 4563 6554
rect 4575 6502 4627 6554
rect 4639 6502 4691 6554
rect 11378 6502 11430 6554
rect 11442 6502 11494 6554
rect 11506 6502 11558 6554
rect 11570 6502 11622 6554
rect 18308 6502 18360 6554
rect 18372 6502 18424 6554
rect 18436 6502 18488 6554
rect 18500 6502 18552 6554
rect 5540 6400 5592 6452
rect 9864 6443 9916 6452
rect 3976 6332 4028 6384
rect 5632 6332 5684 6384
rect 6460 6332 6512 6384
rect 8116 6332 8168 6384
rect 9864 6409 9873 6443
rect 9873 6409 9907 6443
rect 9907 6409 9916 6443
rect 9864 6400 9916 6409
rect 11980 6400 12032 6452
rect 18144 6443 18196 6452
rect 18144 6409 18153 6443
rect 18153 6409 18187 6443
rect 18187 6409 18196 6443
rect 18144 6400 18196 6409
rect 20352 6400 20404 6452
rect 2872 6264 2924 6316
rect 3056 6307 3108 6316
rect 3056 6273 3065 6307
rect 3065 6273 3099 6307
rect 3099 6273 3108 6307
rect 3056 6264 3108 6273
rect 6276 6307 6328 6316
rect 6276 6273 6285 6307
rect 6285 6273 6319 6307
rect 6319 6273 6328 6307
rect 6276 6264 6328 6273
rect 7380 6307 7432 6316
rect 7380 6273 7389 6307
rect 7389 6273 7423 6307
rect 7423 6273 7432 6307
rect 7380 6264 7432 6273
rect 8208 6307 8260 6316
rect 8208 6273 8217 6307
rect 8217 6273 8251 6307
rect 8251 6273 8260 6307
rect 8208 6264 8260 6273
rect 9588 6264 9640 6316
rect 10600 6332 10652 6384
rect 14372 6332 14424 6384
rect 10508 6264 10560 6316
rect 13636 6307 13688 6316
rect 13636 6273 13645 6307
rect 13645 6273 13679 6307
rect 13679 6273 13688 6307
rect 13636 6264 13688 6273
rect 13820 6307 13872 6316
rect 13820 6273 13829 6307
rect 13829 6273 13863 6307
rect 13863 6273 13872 6307
rect 13820 6264 13872 6273
rect 16304 6264 16356 6316
rect 17316 6307 17368 6316
rect 17316 6273 17325 6307
rect 17325 6273 17359 6307
rect 17359 6273 17368 6307
rect 17316 6264 17368 6273
rect 19892 6264 19944 6316
rect 1860 6239 1912 6248
rect 1860 6205 1869 6239
rect 1869 6205 1903 6239
rect 1903 6205 1912 6239
rect 1860 6196 1912 6205
rect 7196 6239 7248 6248
rect 7196 6205 7205 6239
rect 7205 6205 7239 6239
rect 7239 6205 7248 6239
rect 7196 6196 7248 6205
rect 12716 6196 12768 6248
rect 3148 6128 3200 6180
rect 6276 6128 6328 6180
rect 1492 6103 1544 6112
rect 1492 6069 1501 6103
rect 1501 6069 1535 6103
rect 1535 6069 1544 6103
rect 1492 6060 1544 6069
rect 3608 6103 3660 6112
rect 3608 6069 3617 6103
rect 3617 6069 3651 6103
rect 3651 6069 3660 6103
rect 3608 6060 3660 6069
rect 5540 6060 5592 6112
rect 5724 6103 5776 6112
rect 5724 6069 5733 6103
rect 5733 6069 5767 6103
rect 5767 6069 5776 6103
rect 5724 6060 5776 6069
rect 6092 6103 6144 6112
rect 6092 6069 6101 6103
rect 6101 6069 6135 6103
rect 6135 6069 6144 6103
rect 6092 6060 6144 6069
rect 7104 6060 7156 6112
rect 9312 6128 9364 6180
rect 10232 6103 10284 6112
rect 10232 6069 10241 6103
rect 10241 6069 10275 6103
rect 10275 6069 10284 6103
rect 10232 6060 10284 6069
rect 10692 6060 10744 6112
rect 11428 6103 11480 6112
rect 11428 6069 11437 6103
rect 11437 6069 11471 6103
rect 11471 6069 11480 6103
rect 11428 6060 11480 6069
rect 17132 6239 17184 6248
rect 17132 6205 17141 6239
rect 17141 6205 17175 6239
rect 17175 6205 17184 6239
rect 17132 6196 17184 6205
rect 17224 6239 17276 6248
rect 17224 6205 17233 6239
rect 17233 6205 17267 6239
rect 17267 6205 17276 6239
rect 17224 6196 17276 6205
rect 17684 6196 17736 6248
rect 19340 6196 19392 6248
rect 19432 6196 19484 6248
rect 20260 6239 20312 6248
rect 20260 6205 20294 6239
rect 20294 6205 20312 6239
rect 20260 6196 20312 6205
rect 19800 6128 19852 6180
rect 14188 6103 14240 6112
rect 14188 6069 14197 6103
rect 14197 6069 14231 6103
rect 14231 6069 14240 6103
rect 14188 6060 14240 6069
rect 14556 6103 14608 6112
rect 14556 6069 14565 6103
rect 14565 6069 14599 6103
rect 14599 6069 14608 6103
rect 14556 6060 14608 6069
rect 14648 6103 14700 6112
rect 14648 6069 14657 6103
rect 14657 6069 14691 6103
rect 14691 6069 14700 6103
rect 15752 6103 15804 6112
rect 14648 6060 14700 6069
rect 15752 6069 15761 6103
rect 15761 6069 15795 6103
rect 15795 6069 15804 6103
rect 15752 6060 15804 6069
rect 16488 6060 16540 6112
rect 18696 6103 18748 6112
rect 18696 6069 18705 6103
rect 18705 6069 18739 6103
rect 18739 6069 18748 6103
rect 18696 6060 18748 6069
rect 19340 6103 19392 6112
rect 19340 6069 19349 6103
rect 19349 6069 19383 6103
rect 19383 6069 19392 6103
rect 19340 6060 19392 6069
rect 19432 6103 19484 6112
rect 19432 6069 19441 6103
rect 19441 6069 19475 6103
rect 19475 6069 19484 6103
rect 21364 6103 21416 6112
rect 19432 6060 19484 6069
rect 21364 6069 21373 6103
rect 21373 6069 21407 6103
rect 21407 6069 21416 6103
rect 21364 6060 21416 6069
rect 7912 5958 7964 6010
rect 7976 5958 8028 6010
rect 8040 5958 8092 6010
rect 8104 5958 8156 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 15035 5958 15087 6010
rect 1952 5856 2004 5908
rect 6092 5856 6144 5908
rect 6828 5856 6880 5908
rect 10232 5856 10284 5908
rect 2872 5788 2924 5840
rect 4068 5788 4120 5840
rect 5724 5788 5776 5840
rect 1584 5652 1636 5704
rect 2964 5516 3016 5568
rect 5540 5720 5592 5772
rect 6552 5763 6604 5772
rect 6552 5729 6561 5763
rect 6561 5729 6595 5763
rect 6595 5729 6604 5763
rect 9588 5788 9640 5840
rect 11796 5856 11848 5908
rect 11980 5856 12032 5908
rect 14556 5899 14608 5908
rect 14556 5865 14565 5899
rect 14565 5865 14599 5899
rect 14599 5865 14608 5899
rect 14556 5856 14608 5865
rect 16488 5899 16540 5908
rect 16488 5865 16497 5899
rect 16497 5865 16531 5899
rect 16531 5865 16540 5899
rect 16488 5856 16540 5865
rect 17224 5899 17276 5908
rect 17224 5865 17233 5899
rect 17233 5865 17267 5899
rect 17267 5865 17276 5899
rect 17224 5856 17276 5865
rect 18696 5856 18748 5908
rect 19340 5856 19392 5908
rect 12532 5788 12584 5840
rect 17960 5788 18012 5840
rect 6552 5720 6604 5729
rect 10692 5720 10744 5772
rect 11980 5763 12032 5772
rect 11980 5729 11989 5763
rect 11989 5729 12023 5763
rect 12023 5729 12032 5763
rect 11980 5720 12032 5729
rect 4068 5695 4120 5704
rect 4068 5661 4077 5695
rect 4077 5661 4111 5695
rect 4111 5661 4120 5695
rect 4068 5652 4120 5661
rect 6276 5652 6328 5704
rect 5448 5627 5500 5636
rect 5448 5593 5457 5627
rect 5457 5593 5491 5627
rect 5491 5593 5500 5627
rect 7380 5652 7432 5704
rect 7748 5695 7800 5704
rect 7748 5661 7757 5695
rect 7757 5661 7791 5695
rect 7791 5661 7800 5695
rect 7748 5652 7800 5661
rect 8576 5652 8628 5704
rect 9312 5652 9364 5704
rect 10600 5652 10652 5704
rect 5448 5584 5500 5593
rect 10324 5584 10376 5636
rect 10968 5584 11020 5636
rect 11428 5652 11480 5704
rect 12440 5720 12492 5772
rect 12900 5763 12952 5772
rect 12900 5729 12909 5763
rect 12909 5729 12943 5763
rect 12943 5729 12952 5763
rect 12900 5720 12952 5729
rect 13728 5720 13780 5772
rect 15752 5720 15804 5772
rect 12808 5652 12860 5704
rect 15384 5652 15436 5704
rect 16856 5652 16908 5704
rect 19064 5720 19116 5772
rect 19708 5788 19760 5840
rect 20628 5856 20680 5908
rect 19984 5763 20036 5772
rect 19984 5729 19993 5763
rect 19993 5729 20027 5763
rect 20027 5729 20036 5763
rect 19984 5720 20036 5729
rect 18604 5652 18656 5704
rect 20260 5695 20312 5704
rect 20260 5661 20269 5695
rect 20269 5661 20303 5695
rect 20303 5661 20312 5695
rect 20260 5652 20312 5661
rect 6276 5516 6328 5568
rect 8576 5516 8628 5568
rect 9588 5516 9640 5568
rect 11244 5516 11296 5568
rect 11704 5516 11756 5568
rect 11796 5516 11848 5568
rect 15476 5584 15528 5636
rect 19156 5584 19208 5636
rect 14280 5559 14332 5568
rect 14280 5525 14289 5559
rect 14289 5525 14323 5559
rect 14323 5525 14332 5559
rect 14280 5516 14332 5525
rect 17040 5516 17092 5568
rect 19064 5516 19116 5568
rect 21272 5559 21324 5568
rect 21272 5525 21281 5559
rect 21281 5525 21315 5559
rect 21315 5525 21324 5559
rect 21272 5516 21324 5525
rect 4447 5414 4499 5466
rect 4511 5414 4563 5466
rect 4575 5414 4627 5466
rect 4639 5414 4691 5466
rect 11378 5414 11430 5466
rect 11442 5414 11494 5466
rect 11506 5414 11558 5466
rect 11570 5414 11622 5466
rect 18308 5414 18360 5466
rect 18372 5414 18424 5466
rect 18436 5414 18488 5466
rect 18500 5414 18552 5466
rect 9956 5312 10008 5364
rect 11152 5312 11204 5364
rect 12348 5312 12400 5364
rect 13820 5355 13872 5364
rect 13820 5321 13829 5355
rect 13829 5321 13863 5355
rect 13863 5321 13872 5355
rect 13820 5312 13872 5321
rect 16028 5312 16080 5364
rect 16396 5312 16448 5364
rect 19432 5312 19484 5364
rect 2780 5244 2832 5296
rect 3884 5244 3936 5296
rect 6460 5244 6512 5296
rect 9404 5244 9456 5296
rect 9588 5244 9640 5296
rect 15292 5244 15344 5296
rect 17868 5244 17920 5296
rect 2964 5176 3016 5228
rect 3056 5219 3108 5228
rect 3056 5185 3065 5219
rect 3065 5185 3099 5219
rect 3099 5185 3108 5219
rect 3056 5176 3108 5185
rect 1492 5108 1544 5160
rect 204 5040 256 5092
rect 4160 5176 4212 5228
rect 5724 5176 5776 5228
rect 10140 5176 10192 5228
rect 14280 5176 14332 5228
rect 15384 5176 15436 5228
rect 19156 5176 19208 5228
rect 20260 5219 20312 5228
rect 20260 5185 20269 5219
rect 20269 5185 20303 5219
rect 20303 5185 20312 5219
rect 20260 5176 20312 5185
rect 6000 5108 6052 5160
rect 10968 5108 11020 5160
rect 12440 5151 12492 5160
rect 12440 5117 12449 5151
rect 12449 5117 12483 5151
rect 12483 5117 12492 5151
rect 12440 5108 12492 5117
rect 14188 5108 14240 5160
rect 15476 5151 15528 5160
rect 15476 5117 15485 5151
rect 15485 5117 15519 5151
rect 15519 5117 15528 5151
rect 15476 5108 15528 5117
rect 2228 4972 2280 5024
rect 2688 4972 2740 5024
rect 4068 5040 4120 5092
rect 8208 5040 8260 5092
rect 5540 5015 5592 5024
rect 5540 4981 5549 5015
rect 5549 4981 5583 5015
rect 5583 4981 5592 5015
rect 5540 4972 5592 4981
rect 6460 4972 6512 5024
rect 11612 4972 11664 5024
rect 14372 5040 14424 5092
rect 13912 4972 13964 5024
rect 18604 5040 18656 5092
rect 21272 5108 21324 5160
rect 15568 5015 15620 5024
rect 15568 4981 15577 5015
rect 15577 4981 15611 5015
rect 15611 4981 15620 5015
rect 19432 5015 19484 5024
rect 15568 4972 15620 4981
rect 19432 4981 19441 5015
rect 19441 4981 19475 5015
rect 19475 4981 19484 5015
rect 19432 4972 19484 4981
rect 20444 4972 20496 5024
rect 7912 4870 7964 4922
rect 7976 4870 8028 4922
rect 8040 4870 8092 4922
rect 8104 4870 8156 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 15035 4870 15087 4922
rect 2228 4811 2280 4820
rect 2228 4777 2237 4811
rect 2237 4777 2271 4811
rect 2271 4777 2280 4811
rect 2228 4768 2280 4777
rect 2688 4811 2740 4820
rect 2688 4777 2697 4811
rect 2697 4777 2731 4811
rect 2731 4777 2740 4811
rect 2688 4768 2740 4777
rect 3976 4768 4028 4820
rect 5632 4768 5684 4820
rect 7196 4768 7248 4820
rect 8208 4768 8260 4820
rect 7472 4700 7524 4752
rect 10784 4768 10836 4820
rect 11704 4768 11756 4820
rect 11980 4811 12032 4820
rect 11980 4777 11989 4811
rect 11989 4777 12023 4811
rect 12023 4777 12032 4811
rect 11980 4768 12032 4777
rect 12348 4768 12400 4820
rect 13544 4768 13596 4820
rect 17316 4768 17368 4820
rect 19984 4768 20036 4820
rect 3148 4632 3200 4684
rect 3608 4632 3660 4684
rect 8576 4700 8628 4752
rect 11244 4700 11296 4752
rect 19432 4700 19484 4752
rect 15568 4632 15620 4684
rect 16488 4632 16540 4684
rect 17868 4632 17920 4684
rect 19340 4632 19392 4684
rect 20628 4632 20680 4684
rect 2872 4607 2924 4616
rect 2872 4573 2881 4607
rect 2881 4573 2915 4607
rect 2915 4573 2924 4607
rect 2872 4564 2924 4573
rect 2964 4564 3016 4616
rect 3424 4496 3476 4548
rect 5724 4564 5776 4616
rect 8944 4607 8996 4616
rect 5816 4496 5868 4548
rect 8944 4573 8953 4607
rect 8953 4573 8987 4607
rect 8987 4573 8996 4607
rect 8944 4564 8996 4573
rect 11612 4607 11664 4616
rect 11612 4573 11621 4607
rect 11621 4573 11655 4607
rect 11655 4573 11664 4607
rect 11612 4564 11664 4573
rect 15292 4564 15344 4616
rect 8852 4496 8904 4548
rect 19892 4496 19944 4548
rect 3608 4428 3660 4480
rect 4804 4471 4856 4480
rect 4804 4437 4813 4471
rect 4813 4437 4847 4471
rect 4847 4437 4856 4471
rect 4804 4428 4856 4437
rect 5908 4471 5960 4480
rect 5908 4437 5917 4471
rect 5917 4437 5951 4471
rect 5951 4437 5960 4471
rect 5908 4428 5960 4437
rect 7840 4428 7892 4480
rect 11704 4428 11756 4480
rect 15476 4428 15528 4480
rect 19984 4428 20036 4480
rect 4447 4326 4499 4378
rect 4511 4326 4563 4378
rect 4575 4326 4627 4378
rect 4639 4326 4691 4378
rect 11378 4326 11430 4378
rect 11442 4326 11494 4378
rect 11506 4326 11558 4378
rect 11570 4326 11622 4378
rect 18308 4326 18360 4378
rect 18372 4326 18424 4378
rect 18436 4326 18488 4378
rect 18500 4326 18552 4378
rect 2872 4267 2924 4276
rect 2872 4233 2881 4267
rect 2881 4233 2915 4267
rect 2915 4233 2924 4267
rect 2872 4224 2924 4233
rect 3148 4267 3200 4276
rect 3148 4233 3157 4267
rect 3157 4233 3191 4267
rect 3191 4233 3200 4267
rect 3148 4224 3200 4233
rect 7472 4224 7524 4276
rect 3884 4156 3936 4208
rect 7748 4156 7800 4208
rect 3608 4088 3660 4140
rect 1492 4063 1544 4072
rect 1492 4029 1501 4063
rect 1501 4029 1535 4063
rect 1535 4029 1544 4063
rect 1492 4020 1544 4029
rect 3056 4020 3108 4072
rect 4804 4088 4856 4140
rect 5448 4131 5500 4140
rect 5448 4097 5457 4131
rect 5457 4097 5491 4131
rect 5491 4097 5500 4131
rect 6000 4131 6052 4140
rect 5448 4088 5500 4097
rect 6000 4097 6009 4131
rect 6009 4097 6043 4131
rect 6043 4097 6052 4131
rect 6000 4088 6052 4097
rect 5540 4020 5592 4072
rect 1032 3952 1084 4004
rect 2688 3884 2740 3936
rect 3608 3995 3660 4004
rect 3608 3961 3617 3995
rect 3617 3961 3651 3995
rect 3651 3961 3660 3995
rect 3608 3952 3660 3961
rect 4896 3927 4948 3936
rect 4896 3893 4905 3927
rect 4905 3893 4939 3927
rect 4939 3893 4948 3927
rect 4896 3884 4948 3893
rect 5356 3952 5408 4004
rect 7656 4088 7708 4140
rect 7840 4131 7892 4140
rect 7840 4097 7849 4131
rect 7849 4097 7883 4131
rect 7883 4097 7892 4131
rect 7840 4088 7892 4097
rect 6460 4020 6512 4072
rect 8576 4224 8628 4276
rect 8392 4156 8444 4208
rect 8484 4020 8536 4072
rect 10140 4224 10192 4276
rect 11244 4224 11296 4276
rect 17960 4224 18012 4276
rect 20628 4224 20680 4276
rect 8852 3952 8904 4004
rect 7288 3884 7340 3936
rect 7656 3884 7708 3936
rect 8208 3884 8260 3936
rect 8760 3884 8812 3936
rect 13268 4156 13320 4208
rect 12440 4088 12492 4140
rect 15568 4088 15620 4140
rect 19248 4088 19300 4140
rect 19340 4088 19392 4140
rect 14280 4020 14332 4072
rect 16396 4020 16448 4072
rect 16028 3952 16080 4004
rect 19892 4063 19944 4072
rect 19892 4029 19926 4063
rect 19926 4029 19944 4063
rect 19892 4020 19944 4029
rect 20720 3952 20772 4004
rect 9772 3927 9824 3936
rect 9772 3893 9781 3927
rect 9781 3893 9815 3927
rect 9815 3893 9824 3927
rect 9772 3884 9824 3893
rect 15200 3927 15252 3936
rect 15200 3893 15209 3927
rect 15209 3893 15243 3927
rect 15243 3893 15252 3927
rect 15200 3884 15252 3893
rect 15476 3884 15528 3936
rect 15844 3884 15896 3936
rect 16304 3884 16356 3936
rect 21824 3884 21876 3936
rect 7912 3782 7964 3834
rect 7976 3782 8028 3834
rect 8040 3782 8092 3834
rect 8104 3782 8156 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 15035 3782 15087 3834
rect 3056 3723 3108 3732
rect 3056 3689 3065 3723
rect 3065 3689 3099 3723
rect 3099 3689 3108 3723
rect 3056 3680 3108 3689
rect 5264 3723 5316 3732
rect 5264 3689 5273 3723
rect 5273 3689 5307 3723
rect 5307 3689 5316 3723
rect 5264 3680 5316 3689
rect 5908 3680 5960 3732
rect 8208 3723 8260 3732
rect 8208 3689 8217 3723
rect 8217 3689 8251 3723
rect 8251 3689 8260 3723
rect 8208 3680 8260 3689
rect 8944 3680 8996 3732
rect 9496 3680 9548 3732
rect 11244 3723 11296 3732
rect 11244 3689 11253 3723
rect 11253 3689 11287 3723
rect 11287 3689 11296 3723
rect 11244 3680 11296 3689
rect 572 3612 624 3664
rect 5540 3612 5592 3664
rect 5816 3612 5868 3664
rect 1492 3544 1544 3596
rect 1768 3544 1820 3596
rect 1952 3587 2004 3596
rect 1952 3553 1975 3587
rect 1975 3553 2004 3587
rect 1952 3544 2004 3553
rect 4068 3544 4120 3596
rect 5448 3476 5500 3528
rect 10508 3612 10560 3664
rect 9496 3544 9548 3596
rect 9956 3587 10008 3596
rect 9956 3553 9965 3587
rect 9965 3553 9999 3587
rect 9999 3553 10008 3587
rect 9956 3544 10008 3553
rect 2780 3408 2832 3460
rect 2964 3408 3016 3460
rect 7748 3476 7800 3528
rect 8760 3476 8812 3528
rect 8852 3519 8904 3528
rect 8852 3485 8861 3519
rect 8861 3485 8895 3519
rect 8895 3485 8904 3519
rect 8852 3476 8904 3485
rect 10784 3476 10836 3528
rect 16304 3680 16356 3732
rect 16488 3680 16540 3732
rect 19800 3680 19852 3732
rect 20536 3723 20588 3732
rect 20536 3689 20545 3723
rect 20545 3689 20579 3723
rect 20579 3689 20588 3723
rect 20536 3680 20588 3689
rect 15568 3655 15620 3664
rect 15568 3621 15602 3655
rect 15602 3621 15620 3655
rect 15568 3612 15620 3621
rect 11704 3587 11756 3596
rect 11704 3553 11713 3587
rect 11713 3553 11747 3587
rect 11747 3553 11756 3587
rect 11704 3544 11756 3553
rect 1952 3340 2004 3392
rect 2688 3340 2740 3392
rect 7380 3408 7432 3460
rect 3792 3340 3844 3392
rect 6092 3340 6144 3392
rect 6736 3340 6788 3392
rect 8116 3408 8168 3460
rect 8484 3408 8536 3460
rect 10324 3408 10376 3460
rect 12808 3544 12860 3596
rect 13452 3544 13504 3596
rect 15292 3587 15344 3596
rect 15292 3553 15301 3587
rect 15301 3553 15335 3587
rect 15335 3553 15344 3587
rect 15292 3544 15344 3553
rect 16580 3544 16632 3596
rect 18144 3544 18196 3596
rect 18880 3587 18932 3596
rect 18880 3553 18889 3587
rect 18889 3553 18923 3587
rect 18923 3553 18932 3587
rect 18880 3544 18932 3553
rect 19248 3544 19300 3596
rect 21824 3544 21876 3596
rect 9680 3340 9732 3392
rect 10140 3340 10192 3392
rect 13360 3476 13412 3528
rect 17224 3476 17276 3528
rect 19524 3476 19576 3528
rect 13268 3340 13320 3392
rect 13728 3340 13780 3392
rect 14556 3340 14608 3392
rect 17776 3340 17828 3392
rect 19616 3340 19668 3392
rect 22284 3340 22336 3392
rect 4447 3238 4499 3290
rect 4511 3238 4563 3290
rect 4575 3238 4627 3290
rect 4639 3238 4691 3290
rect 11378 3238 11430 3290
rect 11442 3238 11494 3290
rect 11506 3238 11558 3290
rect 11570 3238 11622 3290
rect 18308 3238 18360 3290
rect 18372 3238 18424 3290
rect 18436 3238 18488 3290
rect 18500 3238 18552 3290
rect 3516 3136 3568 3188
rect 5448 3136 5500 3188
rect 9496 3179 9548 3188
rect 4160 3111 4212 3120
rect 4160 3077 4169 3111
rect 4169 3077 4203 3111
rect 4203 3077 4212 3111
rect 4160 3068 4212 3077
rect 5540 3068 5592 3120
rect 6644 3068 6696 3120
rect 4068 3000 4120 3052
rect 1768 2932 1820 2984
rect 5724 2932 5776 2984
rect 5908 2932 5960 2984
rect 6276 2932 6328 2984
rect 6828 2975 6880 2984
rect 6828 2941 6837 2975
rect 6837 2941 6871 2975
rect 6871 2941 6880 2975
rect 6828 2932 6880 2941
rect 3516 2864 3568 2916
rect 7748 3111 7800 3120
rect 7748 3077 7757 3111
rect 7757 3077 7791 3111
rect 7791 3077 7800 3111
rect 7748 3068 7800 3077
rect 9496 3145 9505 3179
rect 9505 3145 9539 3179
rect 9539 3145 9548 3179
rect 9496 3136 9548 3145
rect 19064 3136 19116 3188
rect 15476 3068 15528 3120
rect 8116 3043 8168 3052
rect 8116 3009 8125 3043
rect 8125 3009 8159 3043
rect 8159 3009 8168 3043
rect 8116 3000 8168 3009
rect 9680 3000 9732 3052
rect 10692 3043 10744 3052
rect 10692 3009 10701 3043
rect 10701 3009 10735 3043
rect 10735 3009 10744 3043
rect 10692 3000 10744 3009
rect 10784 3043 10836 3052
rect 10784 3009 10793 3043
rect 10793 3009 10827 3043
rect 10827 3009 10836 3043
rect 10784 3000 10836 3009
rect 3884 2796 3936 2848
rect 8392 2907 8444 2916
rect 8392 2873 8426 2907
rect 8426 2873 8444 2907
rect 8392 2864 8444 2873
rect 9680 2864 9732 2916
rect 11888 2932 11940 2984
rect 13268 3000 13320 3052
rect 13912 2975 13964 2984
rect 13912 2941 13921 2975
rect 13921 2941 13955 2975
rect 13955 2941 13964 2975
rect 13912 2932 13964 2941
rect 15200 3000 15252 3052
rect 16488 3068 16540 3120
rect 18144 3000 18196 3052
rect 11796 2864 11848 2916
rect 13820 2864 13872 2916
rect 14740 2864 14792 2916
rect 9772 2796 9824 2848
rect 10232 2839 10284 2848
rect 10232 2805 10241 2839
rect 10241 2805 10275 2839
rect 10275 2805 10284 2839
rect 10232 2796 10284 2805
rect 10508 2796 10560 2848
rect 13268 2796 13320 2848
rect 15384 2796 15436 2848
rect 17040 2932 17092 2984
rect 18052 2975 18104 2984
rect 18052 2941 18061 2975
rect 18061 2941 18095 2975
rect 18095 2941 18104 2975
rect 18052 2932 18104 2941
rect 19432 3000 19484 3052
rect 20812 3043 20864 3052
rect 20812 3009 20821 3043
rect 20821 3009 20855 3043
rect 20855 3009 20864 3043
rect 20812 3000 20864 3009
rect 19524 2975 19576 2984
rect 19524 2941 19533 2975
rect 19533 2941 19567 2975
rect 19567 2941 19576 2975
rect 19524 2932 19576 2941
rect 20720 2932 20772 2984
rect 22744 2932 22796 2984
rect 15844 2907 15896 2916
rect 15844 2873 15853 2907
rect 15853 2873 15887 2907
rect 15887 2873 15896 2907
rect 15844 2864 15896 2873
rect 16580 2864 16632 2916
rect 16856 2864 16908 2916
rect 18512 2864 18564 2916
rect 18604 2796 18656 2848
rect 7912 2694 7964 2746
rect 7976 2694 8028 2746
rect 8040 2694 8092 2746
rect 8104 2694 8156 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 15035 2694 15087 2746
rect 4896 2592 4948 2644
rect 5264 2592 5316 2644
rect 5816 2635 5868 2644
rect 5816 2601 5825 2635
rect 5825 2601 5859 2635
rect 5859 2601 5868 2635
rect 5816 2592 5868 2601
rect 7656 2592 7708 2644
rect 10232 2592 10284 2644
rect 19064 2635 19116 2644
rect 19064 2601 19073 2635
rect 19073 2601 19107 2635
rect 19107 2601 19116 2635
rect 19064 2592 19116 2601
rect 2872 2456 2924 2508
rect 2412 2252 2464 2304
rect 6552 2524 6604 2576
rect 4160 2388 4212 2440
rect 6276 2431 6328 2440
rect 6276 2397 6285 2431
rect 6285 2397 6319 2431
rect 6319 2397 6328 2431
rect 6276 2388 6328 2397
rect 6736 2388 6788 2440
rect 12808 2524 12860 2576
rect 13452 2524 13504 2576
rect 10140 2456 10192 2508
rect 11796 2499 11848 2508
rect 11796 2465 11805 2499
rect 11805 2465 11839 2499
rect 11839 2465 11848 2499
rect 11796 2456 11848 2465
rect 12624 2499 12676 2508
rect 12624 2465 12633 2499
rect 12633 2465 12667 2499
rect 12667 2465 12676 2499
rect 12624 2456 12676 2465
rect 13360 2499 13412 2508
rect 13360 2465 13369 2499
rect 13369 2465 13403 2499
rect 13403 2465 13412 2499
rect 13360 2456 13412 2465
rect 13820 2456 13872 2508
rect 14740 2499 14792 2508
rect 14740 2465 14749 2499
rect 14749 2465 14783 2499
rect 14783 2465 14792 2499
rect 14740 2456 14792 2465
rect 16580 2456 16632 2508
rect 16856 2456 16908 2508
rect 17224 2499 17276 2508
rect 17224 2465 17233 2499
rect 17233 2465 17267 2499
rect 17267 2465 17276 2499
rect 17224 2456 17276 2465
rect 18512 2499 18564 2508
rect 18512 2465 18521 2499
rect 18521 2465 18555 2499
rect 18555 2465 18564 2499
rect 18512 2456 18564 2465
rect 19800 2456 19852 2508
rect 20628 2456 20680 2508
rect 9588 2388 9640 2440
rect 9772 2388 9824 2440
rect 9680 2320 9732 2372
rect 15016 2320 15068 2372
rect 21364 2320 21416 2372
rect 6828 2252 6880 2304
rect 12808 2252 12860 2304
rect 14004 2252 14056 2304
rect 15936 2252 15988 2304
rect 16396 2252 16448 2304
rect 16856 2295 16908 2304
rect 16856 2261 16865 2295
rect 16865 2261 16899 2295
rect 16899 2261 16908 2295
rect 16856 2252 16908 2261
rect 17316 2252 17368 2304
rect 18144 2252 18196 2304
rect 19156 2252 19208 2304
rect 20904 2252 20956 2304
rect 4447 2150 4499 2202
rect 4511 2150 4563 2202
rect 4575 2150 4627 2202
rect 4639 2150 4691 2202
rect 11378 2150 11430 2202
rect 11442 2150 11494 2202
rect 11506 2150 11558 2202
rect 11570 2150 11622 2202
rect 18308 2150 18360 2202
rect 18372 2150 18424 2202
rect 18436 2150 18488 2202
rect 18500 2150 18552 2202
rect 5908 2048 5960 2100
rect 6736 2048 6788 2100
rect 1492 1980 1544 2032
rect 6276 1980 6328 2032
rect 6000 1504 6052 1556
rect 8668 1504 8720 1556
<< metal2 >>
rect 3330 22672 3386 22681
rect 3330 22607 3386 22616
rect 2870 22264 2926 22273
rect 2870 22199 2926 22208
rect 2778 21720 2834 21729
rect 2778 21655 2834 21664
rect 1950 21312 2006 21321
rect 1950 21247 2006 21256
rect 1964 20058 1992 21247
rect 2792 20602 2820 21655
rect 2780 20596 2832 20602
rect 2780 20538 2832 20544
rect 2884 20534 2912 22199
rect 3054 20768 3110 20777
rect 3054 20703 3110 20712
rect 2872 20528 2924 20534
rect 2872 20470 2924 20476
rect 2962 20360 3018 20369
rect 2962 20295 3018 20304
rect 1952 20052 2004 20058
rect 1952 19994 2004 20000
rect 2872 19848 2924 19854
rect 1950 19816 2006 19825
rect 2872 19790 2924 19796
rect 1950 19751 2006 19760
rect 1964 19514 1992 19751
rect 2044 19712 2096 19718
rect 2044 19654 2096 19660
rect 1952 19508 2004 19514
rect 1952 19450 2004 19456
rect 2056 19310 2084 19654
rect 2778 19408 2834 19417
rect 2778 19343 2834 19352
rect 2044 19304 2096 19310
rect 2044 19246 2096 19252
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 1964 18873 1992 18906
rect 1950 18864 2006 18873
rect 1950 18799 2006 18808
rect 1950 18456 2006 18465
rect 1950 18391 1952 18400
rect 2004 18391 2006 18400
rect 1952 18362 2004 18368
rect 1674 18048 1730 18057
rect 1674 17983 1730 17992
rect 1688 17882 1716 17983
rect 1676 17876 1728 17882
rect 1676 17818 1728 17824
rect 1492 17740 1544 17746
rect 1492 17682 1544 17688
rect 1504 17270 1532 17682
rect 1768 17672 1820 17678
rect 1768 17614 1820 17620
rect 1492 17264 1544 17270
rect 1492 17206 1544 17212
rect 1780 16658 1808 17614
rect 1950 17096 2006 17105
rect 1950 17031 2006 17040
rect 1964 16998 1992 17031
rect 1952 16992 2004 16998
rect 1952 16934 2004 16940
rect 1768 16652 1820 16658
rect 1768 16594 1820 16600
rect 1860 16448 1912 16454
rect 1860 16390 1912 16396
rect 1676 16176 1728 16182
rect 1674 16144 1676 16153
rect 1728 16144 1730 16153
rect 1674 16079 1730 16088
rect 1584 15428 1636 15434
rect 1584 15370 1636 15376
rect 1596 14482 1624 15370
rect 1872 15201 1900 16390
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 1964 15609 1992 15642
rect 1950 15600 2006 15609
rect 1950 15535 2006 15544
rect 1858 15192 1914 15201
rect 1858 15127 1914 15136
rect 1768 14952 1820 14958
rect 1768 14894 1820 14900
rect 1780 14550 1808 14894
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 1858 14648 1914 14657
rect 1858 14583 1914 14592
rect 1768 14544 1820 14550
rect 1768 14486 1820 14492
rect 1584 14476 1636 14482
rect 1584 14418 1636 14424
rect 1872 14074 1900 14583
rect 1964 14249 1992 14758
rect 1950 14240 2006 14249
rect 1950 14175 2006 14184
rect 1860 14068 1912 14074
rect 1860 14010 1912 14016
rect 1952 11688 2004 11694
rect 1952 11630 2004 11636
rect 1964 11286 1992 11630
rect 1952 11280 2004 11286
rect 1952 11222 2004 11228
rect 1584 11144 1636 11150
rect 1584 11086 1636 11092
rect 1596 10810 1624 11086
rect 1584 10804 1636 10810
rect 1584 10746 1636 10752
rect 1596 8090 1624 10746
rect 1860 10600 1912 10606
rect 1860 10542 1912 10548
rect 1872 10266 1900 10542
rect 1860 10260 1912 10266
rect 1860 10202 1912 10208
rect 2056 9217 2084 19246
rect 2792 18970 2820 19343
rect 2780 18964 2832 18970
rect 2780 18906 2832 18912
rect 2884 18834 2912 19790
rect 2976 19174 3004 20295
rect 2964 19168 3016 19174
rect 2964 19110 3016 19116
rect 3068 18970 3096 20703
rect 3148 19304 3200 19310
rect 3148 19246 3200 19252
rect 3056 18964 3108 18970
rect 3056 18906 3108 18912
rect 2872 18828 2924 18834
rect 2872 18770 2924 18776
rect 3160 18766 3188 19246
rect 3148 18760 3200 18766
rect 3148 18702 3200 18708
rect 3160 18222 3188 18702
rect 3240 18692 3292 18698
rect 3240 18634 3292 18640
rect 3148 18216 3200 18222
rect 3148 18158 3200 18164
rect 2964 18080 3016 18086
rect 2964 18022 3016 18028
rect 3056 18080 3108 18086
rect 3056 18022 3108 18028
rect 2976 17882 3004 18022
rect 2964 17876 3016 17882
rect 2964 17818 3016 17824
rect 2778 17504 2834 17513
rect 2778 17439 2834 17448
rect 2792 17338 2820 17439
rect 3068 17338 3096 18022
rect 3252 17746 3280 18634
rect 3240 17740 3292 17746
rect 3240 17682 3292 17688
rect 2780 17332 2832 17338
rect 2780 17274 2832 17280
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 3344 17134 3372 22607
rect 5722 22200 5778 23000
rect 17222 22200 17278 23000
rect 18694 22672 18750 22681
rect 18694 22607 18750 22616
rect 4421 20700 4717 20720
rect 4477 20698 4501 20700
rect 4557 20698 4581 20700
rect 4637 20698 4661 20700
rect 4499 20646 4501 20698
rect 4563 20646 4575 20698
rect 4637 20646 4639 20698
rect 4477 20644 4501 20646
rect 4557 20644 4581 20646
rect 4637 20644 4661 20646
rect 4421 20624 4717 20644
rect 3608 19712 3660 19718
rect 3608 19654 3660 19660
rect 3516 19236 3568 19242
rect 3516 19178 3568 19184
rect 3424 17808 3476 17814
rect 3424 17750 3476 17756
rect 2228 17128 2280 17134
rect 2228 17070 2280 17076
rect 2320 17128 2372 17134
rect 2320 17070 2372 17076
rect 3332 17128 3384 17134
rect 3332 17070 3384 17076
rect 2240 16114 2268 17070
rect 2332 16454 2360 17070
rect 2502 16552 2558 16561
rect 2502 16487 2504 16496
rect 2556 16487 2558 16496
rect 2504 16458 2556 16464
rect 2320 16448 2372 16454
rect 2320 16390 2372 16396
rect 3344 16250 3372 17070
rect 3332 16244 3384 16250
rect 3332 16186 3384 16192
rect 2228 16108 2280 16114
rect 2228 16050 2280 16056
rect 2412 15564 2464 15570
rect 2412 15506 2464 15512
rect 3056 15564 3108 15570
rect 3056 15506 3108 15512
rect 2320 15496 2372 15502
rect 2320 15438 2372 15444
rect 2332 14958 2360 15438
rect 2424 15366 2452 15506
rect 2412 15360 2464 15366
rect 2412 15302 2464 15308
rect 2320 14952 2372 14958
rect 2320 14894 2372 14900
rect 2228 14476 2280 14482
rect 2228 14418 2280 14424
rect 2240 14074 2268 14418
rect 2228 14068 2280 14074
rect 2228 14010 2280 14016
rect 2136 13864 2188 13870
rect 2136 13806 2188 13812
rect 2148 13190 2176 13806
rect 2136 13184 2188 13190
rect 2136 13126 2188 13132
rect 2148 12209 2176 13126
rect 2134 12200 2190 12209
rect 2134 12135 2190 12144
rect 2332 11694 2360 14894
rect 2320 11688 2372 11694
rect 2320 11630 2372 11636
rect 2424 9994 2452 15302
rect 2780 14884 2832 14890
rect 2780 14826 2832 14832
rect 2504 14408 2556 14414
rect 2504 14350 2556 14356
rect 2516 12986 2544 14350
rect 2792 13938 2820 14826
rect 3068 14618 3096 15506
rect 3148 15496 3200 15502
rect 3148 15438 3200 15444
rect 3160 14618 3188 15438
rect 3056 14612 3108 14618
rect 3056 14554 3108 14560
rect 3148 14612 3200 14618
rect 3148 14554 3200 14560
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 2964 13932 3016 13938
rect 2964 13874 3016 13880
rect 2870 13832 2926 13841
rect 2870 13767 2926 13776
rect 2688 13728 2740 13734
rect 2688 13670 2740 13676
rect 2700 13530 2728 13670
rect 2688 13524 2740 13530
rect 2688 13466 2740 13472
rect 2778 13288 2834 13297
rect 2778 13223 2834 13232
rect 2504 12980 2556 12986
rect 2504 12922 2556 12928
rect 2596 12640 2648 12646
rect 2596 12582 2648 12588
rect 2688 12640 2740 12646
rect 2688 12582 2740 12588
rect 2608 11354 2636 12582
rect 2700 12442 2728 12582
rect 2688 12436 2740 12442
rect 2688 12378 2740 12384
rect 2596 11348 2648 11354
rect 2596 11290 2648 11296
rect 2792 10810 2820 13223
rect 2884 11898 2912 13767
rect 2976 12850 3004 13874
rect 3148 13456 3200 13462
rect 3148 13398 3200 13404
rect 3160 13190 3188 13398
rect 3436 13190 3464 17750
rect 3528 17678 3556 19178
rect 3620 19174 3648 19654
rect 4421 19612 4717 19632
rect 4477 19610 4501 19612
rect 4557 19610 4581 19612
rect 4637 19610 4661 19612
rect 4499 19558 4501 19610
rect 4563 19558 4575 19610
rect 4637 19558 4639 19610
rect 4477 19556 4501 19558
rect 4557 19556 4581 19558
rect 4637 19556 4661 19558
rect 4421 19536 4717 19556
rect 5736 19242 5764 22200
rect 11352 20700 11648 20720
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11430 20646 11432 20698
rect 11494 20646 11506 20698
rect 11568 20646 11570 20698
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11352 20624 11648 20644
rect 7656 20460 7708 20466
rect 7656 20402 7708 20408
rect 6828 19916 6880 19922
rect 6828 19858 6880 19864
rect 5908 19780 5960 19786
rect 5908 19722 5960 19728
rect 5724 19236 5776 19242
rect 5724 19178 5776 19184
rect 3608 19168 3660 19174
rect 3608 19110 3660 19116
rect 5080 19168 5132 19174
rect 5080 19110 5132 19116
rect 3620 18970 3648 19110
rect 3608 18964 3660 18970
rect 3608 18906 3660 18912
rect 3608 18828 3660 18834
rect 3608 18770 3660 18776
rect 4988 18828 5040 18834
rect 4988 18770 5040 18776
rect 3620 18426 3648 18770
rect 4344 18760 4396 18766
rect 4344 18702 4396 18708
rect 3700 18624 3752 18630
rect 3700 18566 3752 18572
rect 3608 18420 3660 18426
rect 3608 18362 3660 18368
rect 3516 17672 3568 17678
rect 3516 17614 3568 17620
rect 3528 17202 3556 17614
rect 3608 17536 3660 17542
rect 3608 17478 3660 17484
rect 3620 17270 3648 17478
rect 3608 17264 3660 17270
rect 3608 17206 3660 17212
rect 3516 17196 3568 17202
rect 3516 17138 3568 17144
rect 3516 16992 3568 16998
rect 3516 16934 3568 16940
rect 3528 16522 3556 16934
rect 3712 16522 3740 18566
rect 4356 17882 4384 18702
rect 4421 18524 4717 18544
rect 4477 18522 4501 18524
rect 4557 18522 4581 18524
rect 4637 18522 4661 18524
rect 4499 18470 4501 18522
rect 4563 18470 4575 18522
rect 4637 18470 4639 18522
rect 4477 18468 4501 18470
rect 4557 18468 4581 18470
rect 4637 18468 4661 18470
rect 4421 18448 4717 18468
rect 5000 18426 5028 18770
rect 4988 18420 5040 18426
rect 4988 18362 5040 18368
rect 5092 18154 5120 19110
rect 5448 18964 5500 18970
rect 5448 18906 5500 18912
rect 5080 18148 5132 18154
rect 5080 18090 5132 18096
rect 4344 17876 4396 17882
rect 4344 17818 4396 17824
rect 4160 17740 4212 17746
rect 4160 17682 4212 17688
rect 4172 17202 4200 17682
rect 5092 17678 5120 18090
rect 4988 17672 5040 17678
rect 4988 17614 5040 17620
rect 5080 17672 5132 17678
rect 5080 17614 5132 17620
rect 4421 17436 4717 17456
rect 4477 17434 4501 17436
rect 4557 17434 4581 17436
rect 4637 17434 4661 17436
rect 4499 17382 4501 17434
rect 4563 17382 4575 17434
rect 4637 17382 4639 17434
rect 4477 17380 4501 17382
rect 4557 17380 4581 17382
rect 4637 17380 4661 17382
rect 4421 17360 4717 17380
rect 5000 17338 5028 17614
rect 4988 17332 5040 17338
rect 4988 17274 5040 17280
rect 4160 17196 4212 17202
rect 4160 17138 4212 17144
rect 5356 17060 5408 17066
rect 5356 17002 5408 17008
rect 3516 16516 3568 16522
rect 3516 16458 3568 16464
rect 3700 16516 3752 16522
rect 3700 16458 3752 16464
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 3424 13184 3476 13190
rect 3424 13126 3476 13132
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 2872 11620 2924 11626
rect 2872 11562 2924 11568
rect 2884 11354 2912 11562
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 2884 11200 2912 11290
rect 2964 11212 3016 11218
rect 2884 11172 2964 11200
rect 2964 11154 3016 11160
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 2412 9988 2464 9994
rect 2412 9930 2464 9936
rect 2504 9376 2556 9382
rect 2504 9318 2556 9324
rect 2042 9208 2098 9217
rect 2042 9143 2098 9152
rect 2516 9110 2544 9318
rect 2700 9178 2728 10066
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 2504 9104 2556 9110
rect 2504 9046 2556 9052
rect 2516 8430 2544 9046
rect 2596 9036 2648 9042
rect 2596 8978 2648 8984
rect 2504 8424 2556 8430
rect 2504 8366 2556 8372
rect 2320 8288 2372 8294
rect 2320 8230 2372 8236
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 1676 7948 1728 7954
rect 1676 7890 1728 7896
rect 1308 7744 1360 7750
rect 1308 7686 1360 7692
rect 204 5092 256 5098
rect 204 5034 256 5040
rect 216 800 244 5034
rect 1032 4004 1084 4010
rect 1032 3946 1084 3952
rect 572 3664 624 3670
rect 572 3606 624 3612
rect 584 800 612 3606
rect 1044 800 1072 3946
rect 1320 1601 1348 7686
rect 1400 7200 1452 7206
rect 1398 7168 1400 7177
rect 1452 7168 1454 7177
rect 1398 7103 1454 7112
rect 1412 7002 1440 7103
rect 1400 6996 1452 7002
rect 1400 6938 1452 6944
rect 1492 6112 1544 6118
rect 1492 6054 1544 6060
rect 1504 5166 1532 6054
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 1492 5160 1544 5166
rect 1492 5102 1544 5108
rect 1596 4978 1624 5646
rect 1504 4950 1624 4978
rect 1504 4078 1532 4950
rect 1492 4072 1544 4078
rect 1492 4014 1544 4020
rect 1504 3602 1532 4014
rect 1492 3596 1544 3602
rect 1492 3538 1544 3544
rect 1688 2553 1716 7890
rect 2044 7200 2096 7206
rect 2044 7142 2096 7148
rect 1952 6860 2004 6866
rect 1952 6802 2004 6808
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1872 6254 1900 6598
rect 1860 6248 1912 6254
rect 1860 6190 1912 6196
rect 1964 5914 1992 6802
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 1950 3632 2006 3641
rect 1768 3596 1820 3602
rect 1950 3567 1952 3576
rect 1768 3538 1820 3544
rect 2004 3567 2006 3576
rect 1952 3538 2004 3544
rect 1780 2990 1808 3538
rect 2056 3505 2084 7142
rect 2228 5024 2280 5030
rect 2228 4966 2280 4972
rect 2240 4826 2268 4966
rect 2228 4820 2280 4826
rect 2228 4762 2280 4768
rect 2042 3496 2098 3505
rect 2042 3431 2098 3440
rect 1952 3392 2004 3398
rect 1952 3334 2004 3340
rect 1768 2984 1820 2990
rect 1768 2926 1820 2932
rect 1674 2544 1730 2553
rect 1674 2479 1730 2488
rect 1492 2032 1544 2038
rect 1492 1974 1544 1980
rect 1306 1592 1362 1601
rect 1306 1527 1362 1536
rect 1504 800 1532 1974
rect 1964 800 1992 3334
rect 202 0 258 800
rect 570 0 626 800
rect 1030 0 1086 800
rect 1490 0 1546 800
rect 1950 0 2006 800
rect 2332 649 2360 8230
rect 2516 7426 2544 8366
rect 2608 7546 2636 8978
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2700 8090 2728 8910
rect 2792 8090 2820 9998
rect 2872 9444 2924 9450
rect 2872 9386 2924 9392
rect 2884 8974 2912 9386
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2884 8634 2912 8910
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 3056 8356 3108 8362
rect 3056 8298 3108 8304
rect 3068 8265 3096 8298
rect 3054 8256 3110 8265
rect 3054 8191 3110 8200
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 3068 7886 3096 8191
rect 3056 7880 3108 7886
rect 3056 7822 3108 7828
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 2516 7398 2820 7426
rect 3068 7410 3096 7822
rect 2792 6866 2820 7398
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 3160 7206 3188 13126
rect 3332 12300 3384 12306
rect 3528 12288 3556 16458
rect 4421 16348 4717 16368
rect 4477 16346 4501 16348
rect 4557 16346 4581 16348
rect 4637 16346 4661 16348
rect 4499 16294 4501 16346
rect 4563 16294 4575 16346
rect 4637 16294 4639 16346
rect 4477 16292 4501 16294
rect 4557 16292 4581 16294
rect 4637 16292 4661 16294
rect 4421 16272 4717 16292
rect 4252 16244 4304 16250
rect 4252 16186 4304 16192
rect 4160 15564 4212 15570
rect 4160 15506 4212 15512
rect 4172 14822 4200 15506
rect 3884 14816 3936 14822
rect 3884 14758 3936 14764
rect 4160 14816 4212 14822
rect 4160 14758 4212 14764
rect 3896 14414 3924 14758
rect 4160 14476 4212 14482
rect 4160 14418 4212 14424
rect 3884 14408 3936 14414
rect 3884 14350 3936 14356
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 4080 14074 4108 14350
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 3700 13388 3752 13394
rect 3700 13330 3752 13336
rect 3608 12844 3660 12850
rect 3608 12786 3660 12792
rect 3384 12260 3556 12288
rect 3332 12242 3384 12248
rect 3240 11688 3292 11694
rect 3240 11630 3292 11636
rect 3252 11354 3280 11630
rect 3240 11348 3292 11354
rect 3240 11290 3292 11296
rect 3344 7818 3372 12242
rect 3620 11898 3648 12786
rect 3608 11892 3660 11898
rect 3608 11834 3660 11840
rect 3516 11756 3568 11762
rect 3516 11698 3568 11704
rect 3528 11082 3556 11698
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3516 11076 3568 11082
rect 3516 11018 3568 11024
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 3436 9382 3464 9998
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3436 9110 3464 9318
rect 3424 9104 3476 9110
rect 3424 9046 3476 9052
rect 3424 7880 3476 7886
rect 3424 7822 3476 7828
rect 3332 7812 3384 7818
rect 3332 7754 3384 7760
rect 3436 7342 3464 7822
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 3148 7200 3200 7206
rect 3148 7142 3200 7148
rect 2780 6860 2832 6866
rect 2780 6802 2832 6808
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 3068 6322 3096 6734
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 3160 6361 3188 6598
rect 3146 6352 3202 6361
rect 2872 6316 2924 6322
rect 2872 6258 2924 6264
rect 3056 6316 3108 6322
rect 3146 6287 3202 6296
rect 3056 6258 3108 6264
rect 2884 5846 2912 6258
rect 2872 5840 2924 5846
rect 2872 5782 2924 5788
rect 2780 5296 2832 5302
rect 2780 5238 2832 5244
rect 2688 5024 2740 5030
rect 2688 4966 2740 4972
rect 2700 4826 2728 4966
rect 2688 4820 2740 4826
rect 2688 4762 2740 4768
rect 2792 4162 2820 5238
rect 2884 4622 2912 5782
rect 2964 5568 3016 5574
rect 2964 5510 3016 5516
rect 2976 5234 3004 5510
rect 3068 5234 3096 6258
rect 3160 6186 3188 6287
rect 3148 6180 3200 6186
rect 3148 6122 3200 6128
rect 2964 5228 3016 5234
rect 2964 5170 3016 5176
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 2872 4616 2924 4622
rect 2872 4558 2924 4564
rect 2964 4616 3016 4622
rect 2964 4558 3016 4564
rect 2884 4282 2912 4558
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 2792 4134 2912 4162
rect 2688 3936 2740 3942
rect 2688 3878 2740 3884
rect 2700 3398 2728 3878
rect 2780 3460 2832 3466
rect 2780 3402 2832 3408
rect 2688 3392 2740 3398
rect 2688 3334 2740 3340
rect 2412 2304 2464 2310
rect 2412 2246 2464 2252
rect 2424 800 2452 2246
rect 2792 1442 2820 3402
rect 2884 2514 2912 4134
rect 2976 3466 3004 4558
rect 3068 4078 3096 5170
rect 3148 4684 3200 4690
rect 3148 4626 3200 4632
rect 3160 4282 3188 4626
rect 3424 4548 3476 4554
rect 3344 4508 3424 4536
rect 3148 4276 3200 4282
rect 3148 4218 3200 4224
rect 3056 4072 3108 4078
rect 3056 4014 3108 4020
rect 3068 3738 3096 4014
rect 3056 3732 3108 3738
rect 3056 3674 3108 3680
rect 2964 3460 3016 3466
rect 2964 3402 3016 3408
rect 2872 2508 2924 2514
rect 2872 2450 2924 2456
rect 2792 1414 2912 1442
rect 2884 800 2912 1414
rect 3344 800 3372 4508
rect 3424 4490 3476 4496
rect 3528 3890 3556 11018
rect 3620 8294 3648 11494
rect 3712 11014 3740 13330
rect 4172 12986 4200 14418
rect 4264 13530 4292 16186
rect 4344 16040 4396 16046
rect 4344 15982 4396 15988
rect 4436 16040 4488 16046
rect 4436 15982 4488 15988
rect 4252 13524 4304 13530
rect 4252 13466 4304 13472
rect 4356 13462 4384 15982
rect 4448 15638 4476 15982
rect 4712 15972 4764 15978
rect 4712 15914 4764 15920
rect 4724 15706 4752 15914
rect 4712 15700 4764 15706
rect 4712 15642 4764 15648
rect 4436 15632 4488 15638
rect 4436 15574 4488 15580
rect 4421 15260 4717 15280
rect 4477 15258 4501 15260
rect 4557 15258 4581 15260
rect 4637 15258 4661 15260
rect 4499 15206 4501 15258
rect 4563 15206 4575 15258
rect 4637 15206 4639 15258
rect 4477 15204 4501 15206
rect 4557 15204 4581 15206
rect 4637 15204 4661 15206
rect 4421 15184 4717 15204
rect 5264 14272 5316 14278
rect 5264 14214 5316 14220
rect 4421 14172 4717 14192
rect 4477 14170 4501 14172
rect 4557 14170 4581 14172
rect 4637 14170 4661 14172
rect 4499 14118 4501 14170
rect 4563 14118 4575 14170
rect 4637 14118 4639 14170
rect 4477 14116 4501 14118
rect 4557 14116 4581 14118
rect 4637 14116 4661 14118
rect 4421 14096 4717 14116
rect 5172 13932 5224 13938
rect 5172 13874 5224 13880
rect 4528 13728 4580 13734
rect 4528 13670 4580 13676
rect 4540 13530 4568 13670
rect 4528 13524 4580 13530
rect 4528 13466 4580 13472
rect 4344 13456 4396 13462
rect 4344 13398 4396 13404
rect 5080 13456 5132 13462
rect 5080 13398 5132 13404
rect 4988 13388 5040 13394
rect 4988 13330 5040 13336
rect 4804 13320 4856 13326
rect 4804 13262 4856 13268
rect 4421 13084 4717 13104
rect 4477 13082 4501 13084
rect 4557 13082 4581 13084
rect 4637 13082 4661 13084
rect 4499 13030 4501 13082
rect 4563 13030 4575 13082
rect 4637 13030 4639 13082
rect 4477 13028 4501 13030
rect 4557 13028 4581 13030
rect 4637 13028 4661 13030
rect 4421 13008 4717 13028
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 4066 12880 4122 12889
rect 4066 12815 4122 12824
rect 4080 12782 4108 12815
rect 4068 12776 4120 12782
rect 4068 12718 4120 12724
rect 4712 12708 4764 12714
rect 4712 12650 4764 12656
rect 4724 12442 4752 12650
rect 4712 12436 4764 12442
rect 4712 12378 4764 12384
rect 3882 12336 3938 12345
rect 3882 12271 3938 12280
rect 4344 12300 4396 12306
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3700 11008 3752 11014
rect 3700 10950 3752 10956
rect 3608 8288 3660 8294
rect 3608 8230 3660 8236
rect 3608 6112 3660 6118
rect 3608 6054 3660 6060
rect 3620 4690 3648 6054
rect 3608 4684 3660 4690
rect 3608 4626 3660 4632
rect 3608 4480 3660 4486
rect 3608 4422 3660 4428
rect 3620 4146 3648 4422
rect 3608 4140 3660 4146
rect 3608 4082 3660 4088
rect 3620 4010 3648 4082
rect 3608 4004 3660 4010
rect 3608 3946 3660 3952
rect 3528 3862 3648 3890
rect 3516 3188 3568 3194
rect 3516 3130 3568 3136
rect 3528 2922 3556 3130
rect 3516 2916 3568 2922
rect 3516 2858 3568 2864
rect 3620 2009 3648 3862
rect 3712 2961 3740 10950
rect 3804 4026 3832 12038
rect 3896 11694 3924 12271
rect 4344 12242 4396 12248
rect 4066 11928 4122 11937
rect 4066 11863 4122 11872
rect 4080 11830 4108 11863
rect 4068 11824 4120 11830
rect 4068 11766 4120 11772
rect 3884 11688 3936 11694
rect 3884 11630 3936 11636
rect 4356 11558 4384 12242
rect 4421 11996 4717 12016
rect 4477 11994 4501 11996
rect 4557 11994 4581 11996
rect 4637 11994 4661 11996
rect 4499 11942 4501 11994
rect 4563 11942 4575 11994
rect 4637 11942 4639 11994
rect 4477 11940 4501 11942
rect 4557 11940 4581 11942
rect 4637 11940 4661 11942
rect 4421 11920 4717 11940
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 4066 10976 4122 10985
rect 4066 10911 4122 10920
rect 4080 10810 4108 10911
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 4172 10470 4200 11086
rect 4421 10908 4717 10928
rect 4477 10906 4501 10908
rect 4557 10906 4581 10908
rect 4637 10906 4661 10908
rect 4499 10854 4501 10906
rect 4563 10854 4575 10906
rect 4637 10854 4639 10906
rect 4477 10852 4501 10854
rect 4557 10852 4581 10854
rect 4637 10852 4661 10854
rect 4421 10832 4717 10852
rect 4160 10464 4212 10470
rect 4066 10432 4122 10441
rect 4160 10406 4212 10412
rect 4066 10367 4122 10376
rect 4080 10198 4108 10367
rect 4068 10192 4120 10198
rect 4068 10134 4120 10140
rect 4066 10024 4122 10033
rect 4066 9959 4122 9968
rect 4080 9722 4108 9959
rect 4068 9716 4120 9722
rect 4068 9658 4120 9664
rect 3976 9444 4028 9450
rect 3976 9386 4028 9392
rect 3988 7721 4016 9386
rect 4066 9072 4122 9081
rect 4172 9042 4200 10406
rect 4421 9820 4717 9840
rect 4477 9818 4501 9820
rect 4557 9818 4581 9820
rect 4637 9818 4661 9820
rect 4499 9766 4501 9818
rect 4563 9766 4575 9818
rect 4637 9766 4639 9818
rect 4477 9764 4501 9766
rect 4557 9764 4581 9766
rect 4637 9764 4661 9766
rect 4421 9744 4717 9764
rect 4250 9616 4306 9625
rect 4250 9551 4306 9560
rect 4066 9007 4122 9016
rect 4160 9036 4212 9042
rect 4080 8378 4108 9007
rect 4160 8978 4212 8984
rect 4264 8673 4292 9551
rect 4421 8732 4717 8752
rect 4477 8730 4501 8732
rect 4557 8730 4581 8732
rect 4637 8730 4661 8732
rect 4499 8678 4501 8730
rect 4563 8678 4575 8730
rect 4637 8678 4639 8730
rect 4477 8676 4501 8678
rect 4557 8676 4581 8678
rect 4637 8676 4661 8678
rect 4250 8664 4306 8673
rect 4421 8656 4717 8676
rect 4250 8599 4306 8608
rect 4344 8560 4396 8566
rect 4344 8502 4396 8508
rect 4620 8560 4672 8566
rect 4620 8502 4672 8508
rect 4080 8350 4200 8378
rect 4066 8120 4122 8129
rect 4066 8055 4122 8064
rect 4080 7818 4108 8055
rect 4068 7812 4120 7818
rect 4068 7754 4120 7760
rect 3974 7712 4030 7721
rect 3974 7647 4030 7656
rect 4172 7410 4200 8350
rect 4356 8090 4384 8502
rect 4344 8084 4396 8090
rect 4344 8026 4396 8032
rect 4252 7948 4304 7954
rect 4252 7890 4304 7896
rect 4264 7546 4292 7890
rect 4632 7886 4660 8502
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4421 7644 4717 7664
rect 4477 7642 4501 7644
rect 4557 7642 4581 7644
rect 4637 7642 4661 7644
rect 4499 7590 4501 7642
rect 4563 7590 4575 7642
rect 4637 7590 4639 7642
rect 4477 7588 4501 7590
rect 4557 7588 4581 7590
rect 4637 7588 4661 7590
rect 4421 7568 4717 7588
rect 4252 7540 4304 7546
rect 4816 7528 4844 13262
rect 5000 12714 5028 13330
rect 4988 12708 5040 12714
rect 5092 12696 5120 13398
rect 5184 13258 5212 13874
rect 5276 13734 5304 14214
rect 5264 13728 5316 13734
rect 5264 13670 5316 13676
rect 5276 13326 5304 13670
rect 5264 13320 5316 13326
rect 5264 13262 5316 13268
rect 5172 13252 5224 13258
rect 5172 13194 5224 13200
rect 5184 12850 5212 13194
rect 5172 12844 5224 12850
rect 5172 12786 5224 12792
rect 5092 12668 5304 12696
rect 4988 12650 5040 12656
rect 4896 11280 4948 11286
rect 4896 11222 4948 11228
rect 4908 10266 4936 11222
rect 4896 10260 4948 10266
rect 4896 10202 4948 10208
rect 5000 9178 5028 12650
rect 5080 11688 5132 11694
rect 5080 11630 5132 11636
rect 5092 11286 5120 11630
rect 5080 11280 5132 11286
rect 5080 11222 5132 11228
rect 5172 11212 5224 11218
rect 5172 11154 5224 11160
rect 5184 10810 5212 11154
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 5184 10062 5212 10746
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 5276 9908 5304 12668
rect 5184 9880 5304 9908
rect 5078 9480 5134 9489
rect 5078 9415 5134 9424
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 4252 7482 4304 7488
rect 4356 7500 4844 7528
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4172 7002 4200 7346
rect 4160 6996 4212 7002
rect 4160 6938 4212 6944
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 3974 6760 4030 6769
rect 3974 6695 4030 6704
rect 3988 6390 4016 6695
rect 3976 6384 4028 6390
rect 3976 6326 4028 6332
rect 4080 5846 4108 6802
rect 4158 6216 4214 6225
rect 4158 6151 4214 6160
rect 4068 5840 4120 5846
rect 3882 5808 3938 5817
rect 4068 5782 4120 5788
rect 3882 5743 3938 5752
rect 3896 5302 3924 5743
rect 4080 5710 4108 5782
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 3974 5264 4030 5273
rect 4172 5234 4200 6151
rect 3974 5199 4030 5208
rect 4160 5228 4212 5234
rect 3882 4856 3938 4865
rect 3988 4826 4016 5199
rect 4160 5170 4212 5176
rect 4068 5092 4120 5098
rect 4068 5034 4120 5040
rect 3882 4791 3938 4800
rect 3976 4820 4028 4826
rect 3896 4214 3924 4791
rect 3976 4762 4028 4768
rect 4080 4457 4108 5034
rect 4066 4448 4122 4457
rect 4066 4383 4122 4392
rect 3884 4208 3936 4214
rect 3884 4150 3936 4156
rect 3804 3998 4016 4026
rect 3882 3904 3938 3913
rect 3882 3839 3938 3848
rect 3792 3392 3844 3398
rect 3792 3334 3844 3340
rect 3698 2952 3754 2961
rect 3698 2887 3754 2896
rect 3606 2000 3662 2009
rect 3606 1935 3662 1944
rect 3804 800 3832 3334
rect 3896 2854 3924 3839
rect 3884 2848 3936 2854
rect 3884 2790 3936 2796
rect 3988 1057 4016 3998
rect 4158 3632 4214 3641
rect 4068 3596 4120 3602
rect 4158 3567 4214 3576
rect 4068 3538 4120 3544
rect 4080 3058 4108 3538
rect 4172 3126 4200 3567
rect 4160 3120 4212 3126
rect 4160 3062 4212 3068
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 4172 2446 4200 3062
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 3974 1048 4030 1057
rect 3974 983 4030 992
rect 4356 898 4384 7500
rect 4908 6934 4936 8570
rect 5000 8430 5028 9114
rect 4988 8424 5040 8430
rect 4988 8366 5040 8372
rect 5092 8362 5120 9415
rect 5080 8356 5132 8362
rect 5080 8298 5132 8304
rect 4896 6928 4948 6934
rect 4896 6870 4948 6876
rect 4421 6556 4717 6576
rect 4477 6554 4501 6556
rect 4557 6554 4581 6556
rect 4637 6554 4661 6556
rect 4499 6502 4501 6554
rect 4563 6502 4575 6554
rect 4637 6502 4639 6554
rect 4477 6500 4501 6502
rect 4557 6500 4581 6502
rect 4637 6500 4661 6502
rect 4421 6480 4717 6500
rect 5184 6089 5212 9880
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 5276 7546 5304 7822
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5170 6080 5226 6089
rect 5170 6015 5226 6024
rect 4421 5468 4717 5488
rect 4477 5466 4501 5468
rect 4557 5466 4581 5468
rect 4637 5466 4661 5468
rect 4499 5414 4501 5466
rect 4563 5414 4575 5466
rect 4637 5414 4639 5466
rect 4477 5412 4501 5414
rect 4557 5412 4581 5414
rect 4637 5412 4661 5414
rect 4421 5392 4717 5412
rect 5368 5386 5396 17002
rect 5460 13394 5488 18906
rect 5540 18624 5592 18630
rect 5540 18566 5592 18572
rect 5552 17678 5580 18566
rect 5920 18154 5948 19722
rect 6840 19174 6868 19858
rect 7104 19848 7156 19854
rect 7104 19790 7156 19796
rect 6828 19168 6880 19174
rect 6828 19110 6880 19116
rect 6184 18896 6236 18902
rect 6184 18838 6236 18844
rect 5908 18148 5960 18154
rect 5908 18090 5960 18096
rect 5540 17672 5592 17678
rect 5540 17614 5592 17620
rect 5552 17082 5580 17614
rect 5552 17054 5672 17082
rect 5540 16992 5592 16998
rect 5540 16934 5592 16940
rect 5552 16794 5580 16934
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 5644 16046 5672 17054
rect 5920 16726 5948 18090
rect 6196 17814 6224 18838
rect 6920 18624 6972 18630
rect 6920 18566 6972 18572
rect 6092 17808 6144 17814
rect 6092 17750 6144 17756
rect 6184 17808 6236 17814
rect 6184 17750 6236 17756
rect 5908 16720 5960 16726
rect 5908 16662 5960 16668
rect 6104 16590 6132 17750
rect 6828 17060 6880 17066
rect 6828 17002 6880 17008
rect 6840 16726 6868 17002
rect 6828 16720 6880 16726
rect 6828 16662 6880 16668
rect 6092 16584 6144 16590
rect 6092 16526 6144 16532
rect 6000 16448 6052 16454
rect 6000 16390 6052 16396
rect 5632 16040 5684 16046
rect 5632 15982 5684 15988
rect 5644 15570 5672 15982
rect 5816 15904 5868 15910
rect 5816 15846 5868 15852
rect 5632 15564 5684 15570
rect 5632 15506 5684 15512
rect 5644 15162 5672 15506
rect 5632 15156 5684 15162
rect 5632 15098 5684 15104
rect 5828 14618 5856 15846
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 6012 13938 6040 16390
rect 6104 16250 6132 16526
rect 6092 16244 6144 16250
rect 6092 16186 6144 16192
rect 6644 15904 6696 15910
rect 6644 15846 6696 15852
rect 6460 14816 6512 14822
rect 6460 14758 6512 14764
rect 6184 14476 6236 14482
rect 6184 14418 6236 14424
rect 6000 13932 6052 13938
rect 6000 13874 6052 13880
rect 6196 13530 6224 14418
rect 6472 14414 6500 14758
rect 6460 14408 6512 14414
rect 6460 14350 6512 14356
rect 6368 13796 6420 13802
rect 6368 13738 6420 13744
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 6380 13462 6408 13738
rect 6368 13456 6420 13462
rect 6368 13398 6420 13404
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 5448 12844 5500 12850
rect 5448 12786 5500 12792
rect 5460 12238 5488 12786
rect 5540 12368 5592 12374
rect 5540 12310 5592 12316
rect 5448 12232 5500 12238
rect 5448 12174 5500 12180
rect 5460 11354 5488 12174
rect 5552 11393 5580 12310
rect 6460 12300 6512 12306
rect 6460 12242 6512 12248
rect 6472 12102 6500 12242
rect 6656 12170 6684 15846
rect 6932 15722 6960 18566
rect 7012 17740 7064 17746
rect 7012 17682 7064 17688
rect 7024 17338 7052 17682
rect 7012 17332 7064 17338
rect 7012 17274 7064 17280
rect 7116 16250 7144 19790
rect 7564 19712 7616 19718
rect 7564 19654 7616 19660
rect 7576 19310 7604 19654
rect 7564 19304 7616 19310
rect 7564 19246 7616 19252
rect 7564 19168 7616 19174
rect 7564 19110 7616 19116
rect 7576 18426 7604 19110
rect 7564 18420 7616 18426
rect 7564 18362 7616 18368
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7208 17202 7236 17478
rect 7196 17196 7248 17202
rect 7196 17138 7248 17144
rect 7288 17060 7340 17066
rect 7288 17002 7340 17008
rect 7300 16658 7328 17002
rect 7564 16788 7616 16794
rect 7564 16730 7616 16736
rect 7288 16652 7340 16658
rect 7288 16594 7340 16600
rect 7300 16454 7328 16594
rect 7288 16448 7340 16454
rect 7288 16390 7340 16396
rect 7104 16244 7156 16250
rect 7104 16186 7156 16192
rect 7300 16046 7328 16390
rect 7288 16040 7340 16046
rect 7288 15982 7340 15988
rect 6932 15706 7052 15722
rect 6920 15700 7052 15706
rect 6972 15694 7052 15700
rect 6920 15642 6972 15648
rect 6920 15564 6972 15570
rect 6920 15506 6972 15512
rect 6828 15360 6880 15366
rect 6828 15302 6880 15308
rect 6644 12164 6696 12170
rect 6644 12106 6696 12112
rect 6460 12096 6512 12102
rect 6460 12038 6512 12044
rect 5538 11384 5594 11393
rect 5448 11348 5500 11354
rect 5538 11319 5594 11328
rect 5448 11290 5500 11296
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5736 10130 5764 10406
rect 6472 10130 6500 12038
rect 6656 11218 6684 12106
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 6552 11008 6604 11014
rect 6552 10950 6604 10956
rect 6564 10606 6592 10950
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 5724 10124 5776 10130
rect 5724 10066 5776 10072
rect 6460 10124 6512 10130
rect 6460 10066 6512 10072
rect 6368 10056 6420 10062
rect 6368 9998 6420 10004
rect 6380 9722 6408 9998
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6472 9382 6500 10066
rect 6656 10062 6684 10610
rect 6644 10056 6696 10062
rect 6644 9998 6696 10004
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5460 8634 5488 8910
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 5552 8265 5580 8434
rect 5538 8256 5594 8265
rect 5538 8191 5594 8200
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5460 6866 5488 7346
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5460 5642 5488 6802
rect 5552 6458 5580 8191
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5644 6390 5672 7278
rect 5736 7002 5764 7822
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5724 6996 5776 7002
rect 5724 6938 5776 6944
rect 5632 6384 5684 6390
rect 5632 6326 5684 6332
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5552 5778 5580 6054
rect 5736 5846 5764 6054
rect 5724 5840 5776 5846
rect 5724 5782 5776 5788
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 5448 5636 5500 5642
rect 5448 5578 5500 5584
rect 4908 5358 5396 5386
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 4421 4380 4717 4400
rect 4477 4378 4501 4380
rect 4557 4378 4581 4380
rect 4637 4378 4661 4380
rect 4499 4326 4501 4378
rect 4563 4326 4575 4378
rect 4637 4326 4639 4378
rect 4477 4324 4501 4326
rect 4557 4324 4581 4326
rect 4637 4324 4661 4326
rect 4421 4304 4717 4324
rect 4816 4146 4844 4422
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4908 4026 4936 5358
rect 5724 5228 5776 5234
rect 5724 5170 5776 5176
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 4816 3998 4936 4026
rect 5356 4004 5408 4010
rect 4421 3292 4717 3312
rect 4477 3290 4501 3292
rect 4557 3290 4581 3292
rect 4637 3290 4661 3292
rect 4499 3238 4501 3290
rect 4563 3238 4575 3290
rect 4637 3238 4639 3290
rect 4477 3236 4501 3238
rect 4557 3236 4581 3238
rect 4637 3236 4661 3238
rect 4421 3216 4717 3236
rect 4421 2204 4717 2224
rect 4477 2202 4501 2204
rect 4557 2202 4581 2204
rect 4637 2202 4661 2204
rect 4499 2150 4501 2202
rect 4563 2150 4575 2202
rect 4637 2150 4639 2202
rect 4477 2148 4501 2150
rect 4557 2148 4581 2150
rect 4637 2148 4661 2150
rect 4421 2128 4717 2148
rect 4816 1170 4844 3998
rect 5356 3946 5408 3952
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 4908 2650 4936 3878
rect 5264 3732 5316 3738
rect 5264 3674 5316 3680
rect 5276 2650 5304 3674
rect 4896 2644 4948 2650
rect 4896 2586 4948 2592
rect 5264 2644 5316 2650
rect 5264 2586 5316 2592
rect 5368 1442 5396 3946
rect 5460 3534 5488 4082
rect 5552 4078 5580 4966
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 5644 3754 5672 4762
rect 5736 4622 5764 5170
rect 5724 4616 5776 4622
rect 5724 4558 5776 4564
rect 5552 3726 5672 3754
rect 5552 3670 5580 3726
rect 5540 3664 5592 3670
rect 5540 3606 5592 3612
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5460 3194 5488 3470
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 5540 3120 5592 3126
rect 5540 3062 5592 3068
rect 4264 870 4384 898
rect 4724 1142 4844 1170
rect 5092 1414 5396 1442
rect 4264 800 4292 870
rect 4724 800 4752 1142
rect 5092 800 5120 1414
rect 5552 800 5580 3062
rect 5736 2990 5764 4558
rect 5828 4554 5856 7142
rect 6092 6112 6144 6118
rect 6092 6054 6144 6060
rect 6104 5914 6132 6054
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 6196 5794 6224 8434
rect 6276 6860 6328 6866
rect 6276 6802 6328 6808
rect 6288 6322 6316 6802
rect 6472 6474 6500 9318
rect 6550 9208 6606 9217
rect 6550 9143 6606 9152
rect 6564 9042 6592 9143
rect 6552 9036 6604 9042
rect 6552 8978 6604 8984
rect 6380 6446 6500 6474
rect 6276 6316 6328 6322
rect 6276 6258 6328 6264
rect 6276 6180 6328 6186
rect 6276 6122 6328 6128
rect 6104 5766 6224 5794
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 5816 4548 5868 4554
rect 5816 4490 5868 4496
rect 5908 4480 5960 4486
rect 5908 4422 5960 4428
rect 5920 3738 5948 4422
rect 6012 4146 6040 5102
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 5908 3732 5960 3738
rect 5908 3674 5960 3680
rect 5816 3664 5868 3670
rect 5816 3606 5868 3612
rect 5724 2984 5776 2990
rect 5724 2926 5776 2932
rect 5828 2650 5856 3606
rect 6104 3398 6132 5766
rect 6288 5710 6316 6122
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 6288 5574 6316 5646
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 6092 3392 6144 3398
rect 6092 3334 6144 3340
rect 6288 2990 6316 5510
rect 5908 2984 5960 2990
rect 5908 2926 5960 2932
rect 6276 2984 6328 2990
rect 6276 2926 6328 2932
rect 5816 2644 5868 2650
rect 5816 2586 5868 2592
rect 5920 2106 5948 2926
rect 6288 2446 6316 2926
rect 6276 2440 6328 2446
rect 6276 2382 6328 2388
rect 5908 2100 5960 2106
rect 5908 2042 5960 2048
rect 6288 2038 6316 2382
rect 6276 2032 6328 2038
rect 6276 1974 6328 1980
rect 6000 1556 6052 1562
rect 6000 1498 6052 1504
rect 6012 800 6040 1498
rect 2318 640 2374 649
rect 2318 575 2374 584
rect 2410 0 2466 800
rect 2870 0 2926 800
rect 3330 0 3386 800
rect 3790 0 3846 800
rect 4250 0 4306 800
rect 4710 0 4766 800
rect 5078 0 5134 800
rect 5538 0 5594 800
rect 5998 0 6054 800
rect 6380 241 6408 6446
rect 6460 6384 6512 6390
rect 6460 6326 6512 6332
rect 6472 5302 6500 6326
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6460 5296 6512 5302
rect 6460 5238 6512 5244
rect 6472 5030 6500 5238
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6460 4072 6512 4078
rect 6460 4014 6512 4020
rect 6472 800 6500 4014
rect 6564 2582 6592 5714
rect 6748 5522 6776 12038
rect 6840 11150 6868 15302
rect 6932 14890 6960 15506
rect 6920 14884 6972 14890
rect 6920 14826 6972 14832
rect 6932 13530 6960 14826
rect 7024 13938 7052 15694
rect 7104 14408 7156 14414
rect 7104 14350 7156 14356
rect 7116 14074 7144 14350
rect 7104 14068 7156 14074
rect 7104 14010 7156 14016
rect 7012 13932 7064 13938
rect 7012 13874 7064 13880
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 7012 13456 7064 13462
rect 7012 13398 7064 13404
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6932 11354 6960 11698
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 6932 10538 6960 10950
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 6920 9988 6972 9994
rect 6920 9930 6972 9936
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 6840 8634 6868 9318
rect 6932 8974 6960 9930
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 6932 7750 6960 8230
rect 6828 7744 6880 7750
rect 6828 7686 6880 7692
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6840 5914 6868 7686
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6656 5494 6776 5522
rect 6656 3126 6684 5494
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 6644 3120 6696 3126
rect 6644 3062 6696 3068
rect 6552 2576 6604 2582
rect 6552 2518 6604 2524
rect 6748 2446 6776 3334
rect 6828 2984 6880 2990
rect 6828 2926 6880 2932
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 6748 2106 6776 2382
rect 6840 2310 6868 2926
rect 6828 2304 6880 2310
rect 6828 2246 6880 2252
rect 6736 2100 6788 2106
rect 6736 2042 6788 2048
rect 6932 800 6960 7686
rect 7024 3210 7052 13398
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 7116 11898 7144 13330
rect 7196 13320 7248 13326
rect 7196 13262 7248 13268
rect 7208 12442 7236 13262
rect 7196 12436 7248 12442
rect 7196 12378 7248 12384
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 7104 11892 7156 11898
rect 7104 11834 7156 11840
rect 7208 11694 7236 12174
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 7104 11552 7156 11558
rect 7104 11494 7156 11500
rect 7116 6866 7144 11494
rect 7300 11200 7328 15982
rect 7380 15972 7432 15978
rect 7380 15914 7432 15920
rect 7392 15434 7420 15914
rect 7380 15428 7432 15434
rect 7380 15370 7432 15376
rect 7472 15360 7524 15366
rect 7472 15302 7524 15308
rect 7484 14890 7512 15302
rect 7472 14884 7524 14890
rect 7472 14826 7524 14832
rect 7380 14544 7432 14550
rect 7380 14486 7432 14492
rect 7392 12986 7420 14486
rect 7484 14414 7512 14826
rect 7472 14408 7524 14414
rect 7472 14350 7524 14356
rect 7484 13326 7512 14350
rect 7472 13320 7524 13326
rect 7472 13262 7524 13268
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 7484 11370 7512 12786
rect 7576 11558 7604 16730
rect 7668 14618 7696 20402
rect 10048 20392 10100 20398
rect 10048 20334 10100 20340
rect 7886 20156 8182 20176
rect 7942 20154 7966 20156
rect 8022 20154 8046 20156
rect 8102 20154 8126 20156
rect 7964 20102 7966 20154
rect 8028 20102 8040 20154
rect 8102 20102 8104 20154
rect 7942 20100 7966 20102
rect 8022 20100 8046 20102
rect 8102 20100 8126 20102
rect 7886 20080 8182 20100
rect 8392 19848 8444 19854
rect 8392 19790 8444 19796
rect 8404 19310 8432 19790
rect 9496 19508 9548 19514
rect 9496 19450 9548 19456
rect 8116 19304 8168 19310
rect 8392 19304 8444 19310
rect 8168 19252 8248 19258
rect 8116 19246 8248 19252
rect 8392 19246 8444 19252
rect 8128 19230 8248 19246
rect 7886 19068 8182 19088
rect 7942 19066 7966 19068
rect 8022 19066 8046 19068
rect 8102 19066 8126 19068
rect 7964 19014 7966 19066
rect 8028 19014 8040 19066
rect 8102 19014 8104 19066
rect 7942 19012 7966 19014
rect 8022 19012 8046 19014
rect 8102 19012 8126 19014
rect 7886 18992 8182 19012
rect 8220 18902 8248 19230
rect 8404 18970 8432 19246
rect 9508 19174 9536 19450
rect 9496 19168 9548 19174
rect 9496 19110 9548 19116
rect 9508 18970 9536 19110
rect 8392 18964 8444 18970
rect 8392 18906 8444 18912
rect 9496 18964 9548 18970
rect 9496 18906 9548 18912
rect 8208 18896 8260 18902
rect 8208 18838 8260 18844
rect 8404 18290 8432 18906
rect 8944 18828 8996 18834
rect 8944 18770 8996 18776
rect 8392 18284 8444 18290
rect 8392 18226 8444 18232
rect 8208 18080 8260 18086
rect 8208 18022 8260 18028
rect 8484 18080 8536 18086
rect 8484 18022 8536 18028
rect 8576 18080 8628 18086
rect 8576 18022 8628 18028
rect 7886 17980 8182 18000
rect 7942 17978 7966 17980
rect 8022 17978 8046 17980
rect 8102 17978 8126 17980
rect 7964 17926 7966 17978
rect 8028 17926 8040 17978
rect 8102 17926 8104 17978
rect 7942 17924 7966 17926
rect 8022 17924 8046 17926
rect 8102 17924 8126 17926
rect 7886 17904 8182 17924
rect 8220 17814 8248 18022
rect 8208 17808 8260 17814
rect 8208 17750 8260 17756
rect 8300 17740 8352 17746
rect 8300 17682 8352 17688
rect 8208 17060 8260 17066
rect 8208 17002 8260 17008
rect 7886 16892 8182 16912
rect 7942 16890 7966 16892
rect 8022 16890 8046 16892
rect 8102 16890 8126 16892
rect 7964 16838 7966 16890
rect 8028 16838 8040 16890
rect 8102 16838 8104 16890
rect 7942 16836 7966 16838
rect 8022 16836 8046 16838
rect 8102 16836 8126 16838
rect 7886 16816 8182 16836
rect 8220 16794 8248 17002
rect 8208 16788 8260 16794
rect 8208 16730 8260 16736
rect 7886 15804 8182 15824
rect 7942 15802 7966 15804
rect 8022 15802 8046 15804
rect 8102 15802 8126 15804
rect 7964 15750 7966 15802
rect 8028 15750 8040 15802
rect 8102 15750 8104 15802
rect 7942 15748 7966 15750
rect 8022 15748 8046 15750
rect 8102 15748 8126 15750
rect 7886 15728 8182 15748
rect 7886 14716 8182 14736
rect 7942 14714 7966 14716
rect 8022 14714 8046 14716
rect 8102 14714 8126 14716
rect 7964 14662 7966 14714
rect 8028 14662 8040 14714
rect 8102 14662 8104 14714
rect 7942 14660 7966 14662
rect 8022 14660 8046 14662
rect 8102 14660 8126 14662
rect 7886 14640 8182 14660
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 7668 13734 7696 14554
rect 8312 14074 8340 17682
rect 8496 17338 8524 18022
rect 8588 17882 8616 18022
rect 8576 17876 8628 17882
rect 8576 17818 8628 17824
rect 8760 17740 8812 17746
rect 8760 17682 8812 17688
rect 8484 17332 8536 17338
rect 8484 17274 8536 17280
rect 8392 17196 8444 17202
rect 8392 17138 8444 17144
rect 8404 16250 8432 17138
rect 8772 16998 8800 17682
rect 8956 17678 8984 18770
rect 9588 18148 9640 18154
rect 9588 18090 9640 18096
rect 9220 18080 9272 18086
rect 9220 18022 9272 18028
rect 9232 17814 9260 18022
rect 9600 17864 9628 18090
rect 9600 17836 9904 17864
rect 9220 17808 9272 17814
rect 9220 17750 9272 17756
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 9772 17740 9824 17746
rect 9772 17682 9824 17688
rect 8944 17672 8996 17678
rect 8944 17614 8996 17620
rect 8956 17202 8984 17614
rect 9496 17604 9548 17610
rect 9496 17546 9548 17552
rect 9508 17338 9536 17546
rect 9496 17332 9548 17338
rect 9496 17274 9548 17280
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 8760 16992 8812 16998
rect 8760 16934 8812 16940
rect 9312 16992 9364 16998
rect 9312 16934 9364 16940
rect 9036 16516 9088 16522
rect 9036 16458 9088 16464
rect 8392 16244 8444 16250
rect 8392 16186 8444 16192
rect 8404 16114 8432 16186
rect 8392 16108 8444 16114
rect 8392 16050 8444 16056
rect 8484 16040 8536 16046
rect 8484 15982 8536 15988
rect 8496 15706 8524 15982
rect 8852 15972 8904 15978
rect 8852 15914 8904 15920
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 8496 15026 8524 15642
rect 8864 15162 8892 15914
rect 8852 15156 8904 15162
rect 8852 15098 8904 15104
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 8864 13938 8892 15098
rect 8208 13932 8260 13938
rect 8208 13874 8260 13880
rect 8852 13932 8904 13938
rect 8852 13874 8904 13880
rect 7656 13728 7708 13734
rect 7656 13670 7708 13676
rect 7668 13190 7696 13670
rect 7886 13628 8182 13648
rect 7942 13626 7966 13628
rect 8022 13626 8046 13628
rect 8102 13626 8126 13628
rect 7964 13574 7966 13626
rect 8028 13574 8040 13626
rect 8102 13574 8104 13626
rect 7942 13572 7966 13574
rect 8022 13572 8046 13574
rect 8102 13572 8126 13574
rect 7886 13552 8182 13572
rect 8220 13512 8248 13874
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 8128 13484 8248 13512
rect 7656 13184 7708 13190
rect 7656 13126 7708 13132
rect 8128 12850 8156 13484
rect 8312 13394 8340 13806
rect 8668 13728 8720 13734
rect 8668 13670 8720 13676
rect 8208 13388 8260 13394
rect 8208 13330 8260 13336
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 8128 12714 8156 12786
rect 7656 12708 7708 12714
rect 7656 12650 7708 12656
rect 8116 12708 8168 12714
rect 8116 12650 8168 12656
rect 7668 12322 7696 12650
rect 7886 12540 8182 12560
rect 7942 12538 7966 12540
rect 8022 12538 8046 12540
rect 8102 12538 8126 12540
rect 7964 12486 7966 12538
rect 8028 12486 8040 12538
rect 8102 12486 8104 12538
rect 7942 12484 7966 12486
rect 8022 12484 8046 12486
rect 8102 12484 8126 12486
rect 7886 12464 8182 12484
rect 7668 12294 7788 12322
rect 7760 12238 7788 12294
rect 7748 12232 7800 12238
rect 7748 12174 7800 12180
rect 7760 11762 7788 12174
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7886 11452 8182 11472
rect 7942 11450 7966 11452
rect 8022 11450 8046 11452
rect 8102 11450 8126 11452
rect 7964 11398 7966 11450
rect 8028 11398 8040 11450
rect 8102 11398 8104 11450
rect 7942 11396 7966 11398
rect 8022 11396 8046 11398
rect 8102 11396 8126 11398
rect 7886 11376 8182 11396
rect 7484 11342 7696 11370
rect 7300 11172 7604 11200
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 7300 10606 7328 11018
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 7300 9994 7328 10542
rect 7288 9988 7340 9994
rect 7288 9930 7340 9936
rect 7300 9586 7328 9930
rect 7288 9580 7340 9586
rect 7288 9522 7340 9528
rect 7196 9172 7248 9178
rect 7300 9160 7328 9522
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 7392 9178 7420 9318
rect 7248 9132 7328 9160
rect 7380 9172 7432 9178
rect 7196 9114 7248 9120
rect 7380 9114 7432 9120
rect 7472 9104 7524 9110
rect 7472 9046 7524 9052
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 7300 8634 7328 8978
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 7392 8378 7420 8910
rect 7484 8498 7512 9046
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7392 8350 7512 8378
rect 7104 6860 7156 6866
rect 7104 6802 7156 6808
rect 7116 6118 7144 6802
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 7208 4826 7236 6190
rect 7392 5710 7420 6258
rect 7484 5817 7512 8350
rect 7470 5808 7526 5817
rect 7470 5743 7526 5752
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 7484 4758 7512 5743
rect 7472 4752 7524 4758
rect 7472 4694 7524 4700
rect 7484 4282 7512 4694
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7288 3936 7340 3942
rect 7340 3896 7420 3924
rect 7288 3878 7340 3884
rect 7392 3466 7420 3896
rect 7380 3460 7432 3466
rect 7380 3402 7432 3408
rect 7024 3182 7420 3210
rect 7392 800 7420 3182
rect 7576 2122 7604 11172
rect 7668 4146 7696 11342
rect 7748 11212 7800 11218
rect 7748 11154 7800 11160
rect 7760 10266 7788 11154
rect 8024 11144 8076 11150
rect 8024 11086 8076 11092
rect 8036 10742 8064 11086
rect 8220 11082 8248 13330
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 8312 11694 8340 13126
rect 8680 12986 8708 13670
rect 8760 13388 8812 13394
rect 8760 13330 8812 13336
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8576 12776 8628 12782
rect 8576 12718 8628 12724
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 8496 11898 8524 12582
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 8300 11688 8352 11694
rect 8300 11630 8352 11636
rect 8208 11076 8260 11082
rect 8208 11018 8260 11024
rect 8024 10736 8076 10742
rect 8024 10678 8076 10684
rect 7886 10364 8182 10384
rect 7942 10362 7966 10364
rect 8022 10362 8046 10364
rect 8102 10362 8126 10364
rect 7964 10310 7966 10362
rect 8028 10310 8040 10362
rect 8102 10310 8104 10362
rect 7942 10308 7966 10310
rect 8022 10308 8046 10310
rect 8102 10308 8126 10310
rect 7886 10288 8182 10308
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 8220 9518 8248 11018
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8312 10130 8340 10406
rect 8300 10124 8352 10130
rect 8300 10066 8352 10072
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 7886 9276 8182 9296
rect 7942 9274 7966 9276
rect 8022 9274 8046 9276
rect 8102 9274 8126 9276
rect 7964 9222 7966 9274
rect 8028 9222 8040 9274
rect 8102 9222 8104 9274
rect 7942 9220 7966 9222
rect 8022 9220 8046 9222
rect 8102 9220 8126 9222
rect 7886 9200 8182 9220
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7760 7818 7788 9114
rect 8220 8430 8248 9318
rect 8312 8498 8340 10066
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8404 8974 8432 9318
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 7886 8188 8182 8208
rect 7942 8186 7966 8188
rect 8022 8186 8046 8188
rect 8102 8186 8126 8188
rect 7964 8134 7966 8186
rect 8028 8134 8040 8186
rect 8102 8134 8104 8186
rect 7942 8132 7966 8134
rect 8022 8132 8046 8134
rect 8102 8132 8126 8134
rect 7886 8112 8182 8132
rect 8220 7954 8248 8366
rect 8312 8090 8340 8434
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 7748 7812 7800 7818
rect 7748 7754 7800 7760
rect 8312 7698 8340 8026
rect 8220 7670 8340 7698
rect 8220 7546 8248 7670
rect 8588 7562 8616 12718
rect 8668 8968 8720 8974
rect 8668 8910 8720 8916
rect 8680 8566 8708 8910
rect 8772 8906 8800 13330
rect 8852 11552 8904 11558
rect 8852 11494 8904 11500
rect 8864 11354 8892 11494
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8852 9172 8904 9178
rect 8852 9114 8904 9120
rect 8760 8900 8812 8906
rect 8760 8842 8812 8848
rect 8668 8560 8720 8566
rect 8668 8502 8720 8508
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8312 7534 8616 7562
rect 7748 7268 7800 7274
rect 7748 7210 7800 7216
rect 7760 7002 7788 7210
rect 7886 7100 8182 7120
rect 7942 7098 7966 7100
rect 8022 7098 8046 7100
rect 8102 7098 8126 7100
rect 7964 7046 7966 7098
rect 8028 7046 8040 7098
rect 8102 7046 8104 7098
rect 7942 7044 7966 7046
rect 8022 7044 8046 7046
rect 8102 7044 8126 7046
rect 7886 7024 8182 7044
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7760 5710 7788 6938
rect 8114 6760 8170 6769
rect 8220 6730 8248 7482
rect 8114 6695 8170 6704
rect 8208 6724 8260 6730
rect 8128 6390 8156 6695
rect 8208 6666 8260 6672
rect 8116 6384 8168 6390
rect 8116 6326 8168 6332
rect 8220 6322 8248 6666
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 7886 6012 8182 6032
rect 7942 6010 7966 6012
rect 8022 6010 8046 6012
rect 8102 6010 8126 6012
rect 7964 5958 7966 6010
rect 8028 5958 8040 6010
rect 8102 5958 8104 6010
rect 7942 5956 7966 5958
rect 8022 5956 8046 5958
rect 8102 5956 8126 5958
rect 7886 5936 8182 5956
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 8208 5092 8260 5098
rect 8208 5034 8260 5040
rect 7886 4924 8182 4944
rect 7942 4922 7966 4924
rect 8022 4922 8046 4924
rect 8102 4922 8126 4924
rect 7964 4870 7966 4922
rect 8028 4870 8040 4922
rect 8102 4870 8104 4922
rect 7942 4868 7966 4870
rect 8022 4868 8046 4870
rect 8102 4868 8126 4870
rect 7886 4848 8182 4868
rect 8220 4826 8248 5034
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 7840 4480 7892 4486
rect 7840 4422 7892 4428
rect 7748 4208 7800 4214
rect 7748 4150 7800 4156
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 7668 2650 7696 3878
rect 7760 3534 7788 4150
rect 7852 4146 7880 4422
rect 7840 4140 7892 4146
rect 7840 4082 7892 4088
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 7886 3836 8182 3856
rect 7942 3834 7966 3836
rect 8022 3834 8046 3836
rect 8102 3834 8126 3836
rect 7964 3782 7966 3834
rect 8028 3782 8040 3834
rect 8102 3782 8104 3834
rect 7942 3780 7966 3782
rect 8022 3780 8046 3782
rect 8102 3780 8126 3782
rect 7886 3760 8182 3780
rect 8220 3738 8248 3878
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 7748 3528 7800 3534
rect 7748 3470 7800 3476
rect 7760 3126 7788 3470
rect 8116 3460 8168 3466
rect 8116 3402 8168 3408
rect 7748 3120 7800 3126
rect 7748 3062 7800 3068
rect 8128 3058 8156 3402
rect 8116 3052 8168 3058
rect 8116 2994 8168 3000
rect 7886 2748 8182 2768
rect 7942 2746 7966 2748
rect 8022 2746 8046 2748
rect 8102 2746 8126 2748
rect 7964 2694 7966 2746
rect 8028 2694 8040 2746
rect 8102 2694 8104 2746
rect 7942 2692 7966 2694
rect 8022 2692 8046 2694
rect 8102 2692 8126 2694
rect 7886 2672 8182 2692
rect 7656 2644 7708 2650
rect 7656 2586 7708 2592
rect 7576 2094 7880 2122
rect 7852 800 7880 2094
rect 8312 800 8340 7534
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 8588 5574 8616 5646
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 8588 4758 8616 5510
rect 8864 4842 8892 9114
rect 9048 7002 9076 16458
rect 9324 16164 9352 16934
rect 9496 16176 9548 16182
rect 9324 16136 9496 16164
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 9140 11082 9168 11494
rect 9128 11076 9180 11082
rect 9128 11018 9180 11024
rect 9036 6996 9088 7002
rect 9036 6938 9088 6944
rect 8680 4814 8892 4842
rect 8576 4752 8628 4758
rect 8576 4694 8628 4700
rect 8588 4282 8616 4694
rect 8576 4276 8628 4282
rect 8576 4218 8628 4224
rect 8392 4208 8444 4214
rect 8392 4150 8444 4156
rect 8404 2922 8432 4150
rect 8484 4072 8536 4078
rect 8484 4014 8536 4020
rect 8496 3466 8524 4014
rect 8484 3460 8536 3466
rect 8484 3402 8536 3408
rect 8392 2916 8444 2922
rect 8392 2858 8444 2864
rect 8680 1562 8708 4814
rect 8944 4616 8996 4622
rect 8944 4558 8996 4564
rect 8852 4548 8904 4554
rect 8852 4490 8904 4496
rect 8864 4010 8892 4490
rect 8852 4004 8904 4010
rect 8852 3946 8904 3952
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8772 3534 8800 3878
rect 8864 3534 8892 3946
rect 8956 3738 8984 4558
rect 8944 3732 8996 3738
rect 8944 3674 8996 3680
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 8852 3528 8904 3534
rect 8852 3470 8904 3476
rect 8668 1556 8720 1562
rect 8668 1498 8720 1504
rect 9140 1442 9168 11018
rect 9324 9178 9352 16136
rect 9496 16118 9548 16124
rect 9692 16046 9720 17682
rect 9784 16590 9812 17682
rect 9772 16584 9824 16590
rect 9772 16526 9824 16532
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9692 15026 9720 15982
rect 9876 15978 9904 17836
rect 9956 16992 10008 16998
rect 9956 16934 10008 16940
rect 9968 16561 9996 16934
rect 9954 16552 10010 16561
rect 9954 16487 10010 16496
rect 9968 16454 9996 16487
rect 9956 16448 10008 16454
rect 9956 16390 10008 16396
rect 9864 15972 9916 15978
rect 9864 15914 9916 15920
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 9692 14482 9720 14962
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 9876 14278 9904 14894
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9876 13938 9904 14214
rect 9864 13932 9916 13938
rect 9864 13874 9916 13880
rect 9680 13728 9732 13734
rect 9680 13670 9732 13676
rect 9772 13728 9824 13734
rect 9772 13670 9824 13676
rect 9692 13138 9720 13670
rect 9784 13530 9812 13670
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 9692 13110 9812 13138
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9692 12442 9720 12582
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9494 12200 9550 12209
rect 9494 12135 9550 12144
rect 9508 9654 9536 12135
rect 9784 11898 9812 13110
rect 9876 12850 9904 13874
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 9968 12730 9996 16390
rect 10060 13394 10088 20334
rect 14817 20156 15113 20176
rect 14873 20154 14897 20156
rect 14953 20154 14977 20156
rect 15033 20154 15057 20156
rect 14895 20102 14897 20154
rect 14959 20102 14971 20154
rect 15033 20102 15035 20154
rect 14873 20100 14897 20102
rect 14953 20100 14977 20102
rect 15033 20100 15057 20102
rect 14817 20080 15113 20100
rect 11352 19612 11648 19632
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11430 19558 11432 19610
rect 11494 19558 11506 19610
rect 11568 19558 11570 19610
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11352 19536 11648 19556
rect 10416 19304 10468 19310
rect 10416 19246 10468 19252
rect 11980 19304 12032 19310
rect 11980 19246 12032 19252
rect 10428 18902 10456 19246
rect 11796 19168 11848 19174
rect 11796 19110 11848 19116
rect 10416 18896 10468 18902
rect 10416 18838 10468 18844
rect 10428 18290 10456 18838
rect 11808 18834 11836 19110
rect 11796 18828 11848 18834
rect 11796 18770 11848 18776
rect 11992 18766 12020 19246
rect 13360 19236 13412 19242
rect 13360 19178 13412 19184
rect 11980 18760 12032 18766
rect 11980 18702 12032 18708
rect 11352 18524 11648 18544
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11430 18470 11432 18522
rect 11494 18470 11506 18522
rect 11568 18470 11570 18522
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11352 18448 11648 18468
rect 10416 18284 10468 18290
rect 10416 18226 10468 18232
rect 10428 17814 10456 18226
rect 10968 18148 11020 18154
rect 10968 18090 11020 18096
rect 10508 18080 10560 18086
rect 10508 18022 10560 18028
rect 10520 17814 10548 18022
rect 10416 17808 10468 17814
rect 10416 17750 10468 17756
rect 10508 17808 10560 17814
rect 10508 17750 10560 17756
rect 10692 17672 10744 17678
rect 10692 17614 10744 17620
rect 10140 17332 10192 17338
rect 10140 17274 10192 17280
rect 10048 13388 10100 13394
rect 10048 13330 10100 13336
rect 10152 13326 10180 17274
rect 10324 17128 10376 17134
rect 10324 17070 10376 17076
rect 10232 16992 10284 16998
rect 10232 16934 10284 16940
rect 10244 16726 10272 16934
rect 10232 16720 10284 16726
rect 10232 16662 10284 16668
rect 10336 16454 10364 17070
rect 10508 16652 10560 16658
rect 10508 16594 10560 16600
rect 10324 16448 10376 16454
rect 10324 16390 10376 16396
rect 10336 16250 10364 16390
rect 10324 16244 10376 16250
rect 10324 16186 10376 16192
rect 10232 14816 10284 14822
rect 10232 14758 10284 14764
rect 10244 14482 10272 14758
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 10244 13326 10272 14418
rect 10324 13932 10376 13938
rect 10324 13874 10376 13880
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 10232 13320 10284 13326
rect 10232 13262 10284 13268
rect 10152 12850 10180 13262
rect 10140 12844 10192 12850
rect 10140 12786 10192 12792
rect 9876 12702 9996 12730
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 9496 9648 9548 9654
rect 9496 9590 9548 9596
rect 9588 9512 9640 9518
rect 9640 9460 9720 9466
rect 9588 9454 9720 9460
rect 9600 9438 9720 9454
rect 9692 9432 9720 9438
rect 9772 9444 9824 9450
rect 9692 9404 9772 9432
rect 9772 9386 9824 9392
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 9312 8900 9364 8906
rect 9312 8842 9364 8848
rect 9324 8430 9352 8842
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 8772 1414 9168 1442
rect 8772 800 8800 1414
rect 9232 800 9260 7686
rect 9324 7546 9352 8366
rect 9312 7540 9364 7546
rect 9416 7528 9444 9318
rect 9876 9042 9904 12702
rect 9956 12640 10008 12646
rect 9956 12582 10008 12588
rect 9968 12170 9996 12582
rect 10244 12238 10272 13262
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 9956 12164 10008 12170
rect 9956 12106 10008 12112
rect 9968 11558 9996 12106
rect 10244 11762 10272 12174
rect 10232 11756 10284 11762
rect 10232 11698 10284 11704
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 10152 10112 10180 10610
rect 10232 10124 10284 10130
rect 10152 10084 10232 10112
rect 10152 9586 10180 10084
rect 10232 10066 10284 10072
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 9968 9466 9996 9522
rect 9968 9438 10088 9466
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 9968 9178 9996 9318
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 10060 9042 10088 9438
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9864 9036 9916 9042
rect 9864 8978 9916 8984
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 9508 7750 9536 8978
rect 10060 8945 10088 8978
rect 10046 8936 10102 8945
rect 9968 8894 10046 8922
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9784 7546 9812 8570
rect 9864 8016 9916 8022
rect 9864 7958 9916 7964
rect 9496 7540 9548 7546
rect 9416 7500 9496 7528
rect 9312 7482 9364 7488
rect 9496 7482 9548 7488
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9508 6866 9536 7482
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 9324 6186 9352 6734
rect 9312 6180 9364 6186
rect 9312 6122 9364 6128
rect 9324 5710 9352 6122
rect 9312 5704 9364 5710
rect 9310 5672 9312 5681
rect 9364 5672 9366 5681
rect 9310 5607 9366 5616
rect 9404 5296 9456 5302
rect 9404 5238 9456 5244
rect 9416 2292 9444 5238
rect 9508 3738 9536 6802
rect 9588 6656 9640 6662
rect 9588 6598 9640 6604
rect 9600 6322 9628 6598
rect 9876 6458 9904 7958
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 9588 5840 9640 5846
rect 9588 5782 9640 5788
rect 9600 5574 9628 5782
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 9600 5302 9628 5510
rect 9968 5370 9996 8894
rect 10046 8871 10102 8880
rect 10152 8634 10180 9522
rect 10336 9450 10364 13874
rect 10416 13864 10468 13870
rect 10416 13806 10468 13812
rect 10428 12918 10456 13806
rect 10416 12912 10468 12918
rect 10416 12854 10468 12860
rect 10324 9444 10376 9450
rect 10324 9386 10376 9392
rect 10324 9172 10376 9178
rect 10324 9114 10376 9120
rect 10336 9042 10364 9114
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 9588 5296 9640 5302
rect 9588 5238 9640 5244
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9496 3732 9548 3738
rect 9496 3674 9548 3680
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 9508 3194 9536 3538
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 9508 3074 9536 3130
rect 9508 3046 9628 3074
rect 9692 3058 9720 3334
rect 9600 2446 9628 3046
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9680 2916 9732 2922
rect 9680 2858 9732 2864
rect 9588 2440 9640 2446
rect 9588 2382 9640 2388
rect 9692 2378 9720 2858
rect 9784 2854 9812 3878
rect 9968 3602 9996 5306
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 9772 2848 9824 2854
rect 9772 2790 9824 2796
rect 9784 2446 9812 2790
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 9680 2372 9732 2378
rect 9680 2314 9732 2320
rect 9416 2264 9628 2292
rect 9600 800 9628 2264
rect 10060 800 10088 7686
rect 10322 6896 10378 6905
rect 10322 6831 10324 6840
rect 10376 6831 10378 6840
rect 10324 6802 10376 6808
rect 10140 6724 10192 6730
rect 10140 6666 10192 6672
rect 10152 5234 10180 6666
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10244 5914 10272 6054
rect 10232 5908 10284 5914
rect 10232 5850 10284 5856
rect 10324 5636 10376 5642
rect 10324 5578 10376 5584
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 10152 4282 10180 5170
rect 10140 4276 10192 4282
rect 10140 4218 10192 4224
rect 10336 3466 10364 5578
rect 10324 3460 10376 3466
rect 10324 3402 10376 3408
rect 10140 3392 10192 3398
rect 10140 3334 10192 3340
rect 10152 2514 10180 3334
rect 10232 2848 10284 2854
rect 10232 2790 10284 2796
rect 10244 2650 10272 2790
rect 10232 2644 10284 2650
rect 10232 2586 10284 2592
rect 10140 2508 10192 2514
rect 10140 2450 10192 2456
rect 10428 898 10456 12854
rect 10520 7342 10548 16594
rect 10600 12708 10652 12714
rect 10600 12650 10652 12656
rect 10612 8634 10640 12650
rect 10704 12442 10732 17614
rect 10980 17542 11008 18090
rect 11888 17808 11940 17814
rect 11888 17750 11940 17756
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 10968 17536 11020 17542
rect 10968 17478 11020 17484
rect 11152 17536 11204 17542
rect 11152 17478 11204 17484
rect 10784 17264 10836 17270
rect 10836 17224 10916 17252
rect 10784 17206 10836 17212
rect 10888 16590 10916 17224
rect 10980 17202 11008 17478
rect 10968 17196 11020 17202
rect 10968 17138 11020 17144
rect 11164 17134 11192 17478
rect 11352 17436 11648 17456
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11430 17382 11432 17434
rect 11494 17382 11506 17434
rect 11568 17382 11570 17434
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11352 17360 11648 17380
rect 11152 17128 11204 17134
rect 11152 17070 11204 17076
rect 10968 16992 11020 16998
rect 10968 16934 11020 16940
rect 11244 16992 11296 16998
rect 11244 16934 11296 16940
rect 10980 16794 11008 16934
rect 11256 16794 11284 16934
rect 10968 16788 11020 16794
rect 10968 16730 11020 16736
rect 11244 16788 11296 16794
rect 11244 16730 11296 16736
rect 11716 16590 11744 17682
rect 10876 16584 10928 16590
rect 10876 16526 10928 16532
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 10888 15910 10916 16526
rect 11352 16348 11648 16368
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11430 16294 11432 16346
rect 11494 16294 11506 16346
rect 11568 16294 11570 16346
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11352 16272 11648 16292
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 10876 15904 10928 15910
rect 10876 15846 10928 15852
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10784 10736 10836 10742
rect 10784 10678 10836 10684
rect 10690 9616 10746 9625
rect 10690 9551 10746 9560
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10612 8430 10640 8570
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10598 7984 10654 7993
rect 10598 7919 10654 7928
rect 10508 7336 10560 7342
rect 10508 7278 10560 7284
rect 10612 7274 10640 7919
rect 10600 7268 10652 7274
rect 10600 7210 10652 7216
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10520 6322 10548 6938
rect 10600 6384 10652 6390
rect 10600 6326 10652 6332
rect 10508 6316 10560 6322
rect 10508 6258 10560 6264
rect 10612 5710 10640 6326
rect 10704 6118 10732 9551
rect 10796 9382 10824 10678
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10782 7440 10838 7449
rect 10782 7375 10838 7384
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 10692 5772 10744 5778
rect 10692 5714 10744 5720
rect 10600 5704 10652 5710
rect 10600 5646 10652 5652
rect 10508 3664 10560 3670
rect 10508 3606 10560 3612
rect 10520 2854 10548 3606
rect 10704 3058 10732 5714
rect 10796 4826 10824 7375
rect 10888 4842 10916 15846
rect 11352 15260 11648 15280
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11430 15206 11432 15258
rect 11494 15206 11506 15258
rect 11568 15206 11570 15258
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11352 15184 11648 15204
rect 11352 14172 11648 14192
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11430 14118 11432 14170
rect 11494 14118 11506 14170
rect 11568 14118 11570 14170
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11352 14096 11648 14116
rect 11716 13870 11744 16050
rect 11900 14362 11928 17750
rect 11992 15570 12020 18702
rect 13372 18698 13400 19178
rect 14740 19168 14792 19174
rect 14740 19110 14792 19116
rect 15568 19168 15620 19174
rect 15568 19110 15620 19116
rect 14648 18828 14700 18834
rect 14648 18770 14700 18776
rect 13360 18692 13412 18698
rect 13360 18634 13412 18640
rect 12164 18080 12216 18086
rect 12164 18022 12216 18028
rect 12072 17128 12124 17134
rect 12072 17070 12124 17076
rect 12084 16658 12112 17070
rect 12072 16652 12124 16658
rect 12072 16594 12124 16600
rect 12176 16590 12204 18022
rect 13372 17898 13400 18634
rect 14188 18624 14240 18630
rect 14188 18566 14240 18572
rect 14200 18222 14228 18566
rect 14188 18216 14240 18222
rect 14188 18158 14240 18164
rect 13544 18080 13596 18086
rect 13544 18022 13596 18028
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 12440 17876 12492 17882
rect 13372 17870 13492 17898
rect 12440 17818 12492 17824
rect 12256 17672 12308 17678
rect 12254 17640 12256 17649
rect 12308 17640 12310 17649
rect 12254 17575 12310 17584
rect 12452 17202 12480 17818
rect 13464 17814 13492 17870
rect 13452 17808 13504 17814
rect 13266 17776 13322 17785
rect 13452 17750 13504 17756
rect 13266 17711 13268 17720
rect 13320 17711 13322 17720
rect 13268 17682 13320 17688
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 12992 16992 13044 16998
rect 12992 16934 13044 16940
rect 12164 16584 12216 16590
rect 13004 16561 13032 16934
rect 12164 16526 12216 16532
rect 12990 16552 13046 16561
rect 12176 15638 12204 16526
rect 12990 16487 12992 16496
rect 13044 16487 13046 16496
rect 12992 16458 13044 16464
rect 12164 15632 12216 15638
rect 12164 15574 12216 15580
rect 11980 15564 12032 15570
rect 11980 15506 12032 15512
rect 11992 15162 12020 15506
rect 12348 15428 12400 15434
rect 12348 15370 12400 15376
rect 11980 15156 12032 15162
rect 11980 15098 12032 15104
rect 11992 14482 12020 15098
rect 12360 14550 12388 15370
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12348 14544 12400 14550
rect 12348 14486 12400 14492
rect 11980 14476 12032 14482
rect 11980 14418 12032 14424
rect 11900 14334 12112 14362
rect 11796 13932 11848 13938
rect 11796 13874 11848 13880
rect 11704 13864 11756 13870
rect 11704 13806 11756 13812
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 11164 13326 11192 13670
rect 11244 13388 11296 13394
rect 11244 13330 11296 13336
rect 11152 13320 11204 13326
rect 11152 13262 11204 13268
rect 11164 12918 11192 13262
rect 11256 12918 11284 13330
rect 11808 13326 11836 13874
rect 11888 13796 11940 13802
rect 11888 13738 11940 13744
rect 11796 13320 11848 13326
rect 11796 13262 11848 13268
rect 11900 13258 11928 13738
rect 11888 13252 11940 13258
rect 11888 13194 11940 13200
rect 11352 13084 11648 13104
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11430 13030 11432 13082
rect 11494 13030 11506 13082
rect 11568 13030 11570 13082
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11352 13008 11648 13028
rect 11152 12912 11204 12918
rect 11152 12854 11204 12860
rect 11244 12912 11296 12918
rect 11244 12854 11296 12860
rect 11888 12708 11940 12714
rect 11888 12650 11940 12656
rect 11072 12396 11652 12424
rect 10968 12368 11020 12374
rect 11072 12356 11100 12396
rect 11020 12328 11100 12356
rect 10968 12310 11020 12316
rect 11624 12306 11652 12396
rect 11152 12300 11204 12306
rect 11152 12242 11204 12248
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 11164 11762 11192 12242
rect 11352 11996 11648 12016
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11430 11942 11432 11994
rect 11494 11942 11506 11994
rect 11568 11942 11570 11994
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11352 11920 11648 11940
rect 11900 11898 11928 12650
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 11980 11688 12032 11694
rect 11980 11630 12032 11636
rect 11796 11620 11848 11626
rect 11796 11562 11848 11568
rect 11352 10908 11648 10928
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11430 10854 11432 10906
rect 11494 10854 11506 10906
rect 11568 10854 11570 10906
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11352 10832 11648 10852
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 10980 8974 11008 9862
rect 11256 9586 11284 10066
rect 11352 9820 11648 9840
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11430 9766 11432 9818
rect 11494 9766 11506 9818
rect 11568 9766 11570 9818
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11352 9744 11648 9764
rect 11808 9602 11836 11562
rect 11992 11558 12020 11630
rect 11888 11552 11940 11558
rect 11888 11494 11940 11500
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 11900 11393 11928 11494
rect 11886 11384 11942 11393
rect 11886 11319 11942 11328
rect 11244 9580 11296 9586
rect 11808 9574 11928 9602
rect 11244 9522 11296 9528
rect 11796 9444 11848 9450
rect 11796 9386 11848 9392
rect 11808 9042 11836 9386
rect 11152 9036 11204 9042
rect 11428 9036 11480 9042
rect 11204 8996 11428 9024
rect 11152 8978 11204 8984
rect 11428 8978 11480 8984
rect 11796 9036 11848 9042
rect 11796 8978 11848 8984
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 10980 7750 11008 8910
rect 11164 7886 11192 8978
rect 11702 8936 11758 8945
rect 11702 8871 11758 8880
rect 11352 8732 11648 8752
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11430 8678 11432 8730
rect 11494 8678 11506 8730
rect 11568 8678 11570 8730
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11352 8656 11648 8676
rect 11716 8634 11744 8871
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11428 8560 11480 8566
rect 11428 8502 11480 8508
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 11256 7886 11284 8434
rect 11440 8294 11468 8502
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11428 8288 11480 8294
rect 11428 8230 11480 8236
rect 11348 8090 11376 8230
rect 11900 8106 11928 9574
rect 12084 8537 12112 14334
rect 12360 13938 12388 14486
rect 12348 13932 12400 13938
rect 12348 13874 12400 13880
rect 12624 13456 12676 13462
rect 12624 13398 12676 13404
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12164 12164 12216 12170
rect 12164 12106 12216 12112
rect 12176 11914 12204 12106
rect 12256 12096 12308 12102
rect 12452 12084 12480 12582
rect 12308 12056 12480 12084
rect 12256 12038 12308 12044
rect 12176 11886 12296 11914
rect 12164 11620 12216 11626
rect 12164 11562 12216 11568
rect 12070 8528 12126 8537
rect 11336 8084 11388 8090
rect 11336 8026 11388 8032
rect 11808 8078 11928 8106
rect 11992 8486 12070 8514
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 11244 7880 11296 7886
rect 11244 7822 11296 7828
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 11256 7342 11284 7822
rect 11704 7744 11756 7750
rect 11704 7686 11756 7692
rect 11352 7644 11648 7664
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11430 7590 11432 7642
rect 11494 7590 11506 7642
rect 11568 7590 11570 7642
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11352 7568 11648 7588
rect 11244 7336 11296 7342
rect 11244 7278 11296 7284
rect 11716 7002 11744 7686
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11808 6769 11836 8078
rect 11794 6760 11850 6769
rect 11794 6695 11850 6704
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 10980 5642 11008 6598
rect 11352 6556 11648 6576
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11430 6502 11432 6554
rect 11494 6502 11506 6554
rect 11568 6502 11570 6554
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11352 6480 11648 6500
rect 11428 6112 11480 6118
rect 11428 6054 11480 6060
rect 11440 5710 11468 6054
rect 11796 5908 11848 5914
rect 11796 5850 11848 5856
rect 11428 5704 11480 5710
rect 11428 5646 11480 5652
rect 10968 5636 11020 5642
rect 10968 5578 11020 5584
rect 10980 5166 11008 5578
rect 11808 5574 11836 5850
rect 11244 5568 11296 5574
rect 11244 5510 11296 5516
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 10968 5160 11020 5166
rect 10968 5102 11020 5108
rect 10784 4820 10836 4826
rect 10888 4814 11008 4842
rect 10784 4762 10836 4768
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 10796 3058 10824 3470
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 10784 3052 10836 3058
rect 10784 2994 10836 3000
rect 10508 2848 10560 2854
rect 10508 2790 10560 2796
rect 10428 870 10548 898
rect 10520 800 10548 870
rect 10980 800 11008 4814
rect 11164 1306 11192 5306
rect 11256 4758 11284 5510
rect 11352 5468 11648 5488
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11430 5414 11432 5466
rect 11494 5414 11506 5466
rect 11568 5414 11570 5466
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11352 5392 11648 5412
rect 11612 5024 11664 5030
rect 11612 4966 11664 4972
rect 11244 4752 11296 4758
rect 11244 4694 11296 4700
rect 11624 4622 11652 4966
rect 11716 4826 11744 5510
rect 11704 4820 11756 4826
rect 11704 4762 11756 4768
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11704 4480 11756 4486
rect 11704 4422 11756 4428
rect 11352 4380 11648 4400
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11430 4326 11432 4378
rect 11494 4326 11506 4378
rect 11568 4326 11570 4378
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11352 4304 11648 4324
rect 11244 4276 11296 4282
rect 11244 4218 11296 4224
rect 11256 3738 11284 4218
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 11716 3602 11744 4422
rect 11704 3596 11756 3602
rect 11704 3538 11756 3544
rect 11352 3292 11648 3312
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11430 3238 11432 3290
rect 11494 3238 11506 3290
rect 11568 3238 11570 3290
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11352 3216 11648 3236
rect 11900 2990 11928 6598
rect 11992 6458 12020 8486
rect 12070 8463 12126 8472
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 12084 6866 12112 7142
rect 12072 6860 12124 6866
rect 12072 6802 12124 6808
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 11992 5914 12020 6394
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 11992 4826 12020 5714
rect 11980 4820 12032 4826
rect 11980 4762 12032 4768
rect 11888 2984 11940 2990
rect 11888 2926 11940 2932
rect 11796 2916 11848 2922
rect 11796 2858 11848 2864
rect 11808 2514 11836 2858
rect 11796 2508 11848 2514
rect 11796 2450 11848 2456
rect 11352 2204 11648 2224
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11430 2150 11432 2202
rect 11494 2150 11506 2202
rect 11568 2150 11570 2202
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11352 2128 11648 2148
rect 12176 1986 12204 11562
rect 12268 11506 12296 11886
rect 12452 11642 12480 12056
rect 12636 11898 12664 13398
rect 12728 12374 12756 14962
rect 13280 13462 13308 17682
rect 13464 17202 13492 17750
rect 13556 17660 13584 18022
rect 13726 17776 13782 17785
rect 13726 17711 13728 17720
rect 13780 17711 13782 17720
rect 13728 17682 13780 17688
rect 13636 17672 13688 17678
rect 13556 17632 13636 17660
rect 13452 17196 13504 17202
rect 13452 17138 13504 17144
rect 13452 16992 13504 16998
rect 13452 16934 13504 16940
rect 13464 16794 13492 16934
rect 13452 16788 13504 16794
rect 13452 16730 13504 16736
rect 13556 16250 13584 17632
rect 13636 17614 13688 17620
rect 13832 17338 13860 18022
rect 14660 17882 14688 18770
rect 14752 18766 14780 19110
rect 14817 19068 15113 19088
rect 14873 19066 14897 19068
rect 14953 19066 14977 19068
rect 15033 19066 15057 19068
rect 14895 19014 14897 19066
rect 14959 19014 14971 19066
rect 15033 19014 15035 19066
rect 14873 19012 14897 19014
rect 14953 19012 14977 19014
rect 15033 19012 15057 19014
rect 14817 18992 15113 19012
rect 15292 18896 15344 18902
rect 15292 18838 15344 18844
rect 14740 18760 14792 18766
rect 14740 18702 14792 18708
rect 14752 18290 14780 18702
rect 15200 18692 15252 18698
rect 15200 18634 15252 18640
rect 14740 18284 14792 18290
rect 14740 18226 14792 18232
rect 14740 18148 14792 18154
rect 14740 18090 14792 18096
rect 14648 17876 14700 17882
rect 14648 17818 14700 17824
rect 14004 17808 14056 17814
rect 14004 17750 14056 17756
rect 13820 17332 13872 17338
rect 13820 17274 13872 17280
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 13544 16244 13596 16250
rect 13544 16186 13596 16192
rect 13452 14884 13504 14890
rect 13452 14826 13504 14832
rect 13464 14346 13492 14826
rect 13452 14340 13504 14346
rect 13452 14282 13504 14288
rect 13268 13456 13320 13462
rect 13268 13398 13320 13404
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12716 12368 12768 12374
rect 12716 12310 12768 12316
rect 12728 12170 12756 12310
rect 12716 12164 12768 12170
rect 12716 12106 12768 12112
rect 12624 11892 12676 11898
rect 12624 11834 12676 11840
rect 12532 11824 12584 11830
rect 12532 11766 12584 11772
rect 12360 11626 12480 11642
rect 12348 11620 12480 11626
rect 12400 11614 12480 11620
rect 12348 11562 12400 11568
rect 12268 11478 12388 11506
rect 12256 8288 12308 8294
rect 12256 8230 12308 8236
rect 12268 6934 12296 8230
rect 12256 6928 12308 6934
rect 12256 6870 12308 6876
rect 12360 5370 12388 11478
rect 12544 11218 12572 11766
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 12452 10606 12480 11154
rect 12820 11014 12848 13330
rect 12900 13320 12952 13326
rect 12900 13262 12952 13268
rect 12912 12918 12940 13262
rect 12900 12912 12952 12918
rect 12900 12854 12952 12860
rect 12912 12442 12940 12854
rect 13084 12844 13136 12850
rect 13084 12786 13136 12792
rect 12900 12436 12952 12442
rect 12900 12378 12952 12384
rect 12912 12306 12940 12378
rect 13096 12322 13124 12786
rect 12900 12300 12952 12306
rect 13096 12294 13216 12322
rect 12900 12242 12952 12248
rect 13082 11384 13138 11393
rect 13082 11319 13138 11328
rect 13096 11286 13124 11319
rect 13084 11280 13136 11286
rect 13084 11222 13136 11228
rect 12808 11008 12860 11014
rect 12808 10950 12860 10956
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12544 9722 12572 10746
rect 13084 10124 13136 10130
rect 13084 10066 13136 10072
rect 12992 10056 13044 10062
rect 12992 9998 13044 10004
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12532 9716 12584 9722
rect 12532 9658 12584 9664
rect 12624 9376 12676 9382
rect 12624 9318 12676 9324
rect 12532 8356 12584 8362
rect 12532 8298 12584 8304
rect 12544 6934 12572 8298
rect 12532 6928 12584 6934
rect 12532 6870 12584 6876
rect 12532 5840 12584 5846
rect 12530 5808 12532 5817
rect 12584 5808 12586 5817
rect 12440 5772 12492 5778
rect 12530 5743 12586 5752
rect 12440 5714 12492 5720
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12452 5166 12480 5714
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 11900 1958 12204 1986
rect 11164 1278 11468 1306
rect 11440 800 11468 1278
rect 11900 800 11928 1958
rect 12360 800 12388 4762
rect 12452 4146 12480 5102
rect 12440 4140 12492 4146
rect 12440 4082 12492 4088
rect 12636 2514 12664 9318
rect 12728 8498 12756 9862
rect 13004 9518 13032 9998
rect 12992 9512 13044 9518
rect 12992 9454 13044 9460
rect 13096 8974 13124 10066
rect 13084 8968 13136 8974
rect 13084 8910 13136 8916
rect 13084 8832 13136 8838
rect 13084 8774 13136 8780
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 12716 8288 12768 8294
rect 12716 8230 12768 8236
rect 12728 8090 12756 8230
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 13004 8022 13032 8434
rect 13096 8362 13124 8774
rect 13188 8430 13216 12294
rect 13176 8424 13228 8430
rect 13176 8366 13228 8372
rect 13084 8356 13136 8362
rect 13084 8298 13136 8304
rect 12992 8016 13044 8022
rect 12992 7958 13044 7964
rect 12808 7948 12860 7954
rect 12860 7908 12940 7936
rect 12808 7890 12860 7896
rect 12912 7342 12940 7908
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 12716 7268 12768 7274
rect 12716 7210 12768 7216
rect 12728 6254 12756 7210
rect 12808 6996 12860 7002
rect 12808 6938 12860 6944
rect 12716 6248 12768 6254
rect 12716 6190 12768 6196
rect 12820 5710 12848 6938
rect 12912 5778 12940 7278
rect 13096 7274 13124 8298
rect 13188 8090 13216 8366
rect 13176 8084 13228 8090
rect 13176 8026 13228 8032
rect 13084 7268 13136 7274
rect 13084 7210 13136 7216
rect 12900 5772 12952 5778
rect 12900 5714 12952 5720
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 13280 4214 13308 13398
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 13372 12442 13400 12718
rect 13360 12436 13412 12442
rect 13360 12378 13412 12384
rect 13360 11144 13412 11150
rect 13360 11086 13412 11092
rect 13372 10810 13400 11086
rect 13360 10804 13412 10810
rect 13360 10746 13412 10752
rect 13556 4826 13584 16186
rect 13832 16182 13860 16594
rect 14016 16454 14044 17750
rect 14280 17672 14332 17678
rect 14280 17614 14332 17620
rect 14292 17542 14320 17614
rect 14280 17536 14332 17542
rect 14280 17478 14332 17484
rect 14004 16448 14056 16454
rect 14004 16390 14056 16396
rect 13820 16176 13872 16182
rect 13820 16118 13872 16124
rect 13820 16040 13872 16046
rect 13820 15982 13872 15988
rect 13832 15706 13860 15982
rect 13820 15700 13872 15706
rect 13820 15642 13872 15648
rect 14188 15564 14240 15570
rect 14188 15506 14240 15512
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 13832 14006 13860 15438
rect 13912 14816 13964 14822
rect 13912 14758 13964 14764
rect 13924 14006 13952 14758
rect 14200 14618 14228 15506
rect 14188 14612 14240 14618
rect 14188 14554 14240 14560
rect 14096 14408 14148 14414
rect 14096 14350 14148 14356
rect 14108 14074 14136 14350
rect 14096 14068 14148 14074
rect 14096 14010 14148 14016
rect 13820 14000 13872 14006
rect 13820 13942 13872 13948
rect 13912 14000 13964 14006
rect 13912 13942 13964 13948
rect 13924 13258 13952 13942
rect 14188 13728 14240 13734
rect 14188 13670 14240 13676
rect 14200 13530 14228 13670
rect 14188 13524 14240 13530
rect 14188 13466 14240 13472
rect 14096 13388 14148 13394
rect 14096 13330 14148 13336
rect 13912 13252 13964 13258
rect 13912 13194 13964 13200
rect 13636 13184 13688 13190
rect 13636 13126 13688 13132
rect 13648 12730 13676 13126
rect 13820 12776 13872 12782
rect 13648 12702 13768 12730
rect 13820 12718 13872 12724
rect 13740 11694 13768 12702
rect 13832 12374 13860 12718
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 13820 12368 13872 12374
rect 13820 12310 13872 12316
rect 13924 11762 13952 12582
rect 13912 11756 13964 11762
rect 13912 11698 13964 11704
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13636 11620 13688 11626
rect 13636 11562 13688 11568
rect 13648 11150 13676 11562
rect 13636 11144 13688 11150
rect 13636 11086 13688 11092
rect 14108 10742 14136 13330
rect 14188 12708 14240 12714
rect 14188 12650 14240 12656
rect 14200 12442 14228 12650
rect 14188 12436 14240 12442
rect 14188 12378 14240 12384
rect 14200 11762 14228 12378
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 14096 10736 14148 10742
rect 14096 10678 14148 10684
rect 13820 10532 13872 10538
rect 13820 10474 13872 10480
rect 13728 9444 13780 9450
rect 13728 9386 13780 9392
rect 13740 8838 13768 9386
rect 13832 8906 13860 10474
rect 14004 10464 14056 10470
rect 14004 10406 14056 10412
rect 13820 8900 13872 8906
rect 13820 8842 13872 8848
rect 13728 8832 13780 8838
rect 13728 8774 13780 8780
rect 13740 8362 13768 8774
rect 14016 8430 14044 10406
rect 14108 9586 14136 10678
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14004 8424 14056 8430
rect 14004 8366 14056 8372
rect 14186 8392 14242 8401
rect 13728 8356 13780 8362
rect 14186 8327 14242 8336
rect 13728 8298 13780 8304
rect 13740 7342 13768 8298
rect 14200 8294 14228 8327
rect 14188 8288 14240 8294
rect 14188 8230 14240 8236
rect 13728 7336 13780 7342
rect 13728 7278 13780 7284
rect 14292 6934 14320 17478
rect 14752 17338 14780 18090
rect 14817 17980 15113 18000
rect 14873 17978 14897 17980
rect 14953 17978 14977 17980
rect 15033 17978 15057 17980
rect 14895 17926 14897 17978
rect 14959 17926 14971 17978
rect 15033 17926 15035 17978
rect 14873 17924 14897 17926
rect 14953 17924 14977 17926
rect 15033 17924 15057 17926
rect 14817 17904 15113 17924
rect 14740 17332 14792 17338
rect 14740 17274 14792 17280
rect 14817 16892 15113 16912
rect 14873 16890 14897 16892
rect 14953 16890 14977 16892
rect 15033 16890 15057 16892
rect 14895 16838 14897 16890
rect 14959 16838 14971 16890
rect 15033 16838 15035 16890
rect 14873 16836 14897 16838
rect 14953 16836 14977 16838
rect 15033 16836 15057 16838
rect 14817 16816 15113 16836
rect 15212 16590 15240 18634
rect 15304 17882 15332 18838
rect 15580 18834 15608 19110
rect 17236 18970 17264 22200
rect 18282 20700 18578 20720
rect 18338 20698 18362 20700
rect 18418 20698 18442 20700
rect 18498 20698 18522 20700
rect 18360 20646 18362 20698
rect 18424 20646 18436 20698
rect 18498 20646 18500 20698
rect 18338 20644 18362 20646
rect 18418 20644 18442 20646
rect 18498 20644 18522 20646
rect 18282 20624 18578 20644
rect 18282 19612 18578 19632
rect 18338 19610 18362 19612
rect 18418 19610 18442 19612
rect 18498 19610 18522 19612
rect 18360 19558 18362 19610
rect 18424 19558 18436 19610
rect 18498 19558 18500 19610
rect 18338 19556 18362 19558
rect 18418 19556 18442 19558
rect 18498 19556 18522 19558
rect 18282 19536 18578 19556
rect 17224 18964 17276 18970
rect 17224 18906 17276 18912
rect 17408 18896 17460 18902
rect 17408 18838 17460 18844
rect 15568 18828 15620 18834
rect 15568 18770 15620 18776
rect 16028 18624 16080 18630
rect 16028 18566 16080 18572
rect 16040 18290 16068 18566
rect 16028 18284 16080 18290
rect 16028 18226 16080 18232
rect 15292 17876 15344 17882
rect 15292 17818 15344 17824
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15856 17202 15884 17614
rect 15844 17196 15896 17202
rect 15844 17138 15896 17144
rect 15568 16992 15620 16998
rect 15568 16934 15620 16940
rect 15580 16794 15608 16934
rect 15568 16788 15620 16794
rect 15568 16730 15620 16736
rect 15200 16584 15252 16590
rect 15200 16526 15252 16532
rect 14817 15804 15113 15824
rect 14873 15802 14897 15804
rect 14953 15802 14977 15804
rect 15033 15802 15057 15804
rect 14895 15750 14897 15802
rect 14959 15750 14971 15802
rect 15033 15750 15035 15802
rect 14873 15748 14897 15750
rect 14953 15748 14977 15750
rect 15033 15748 15057 15750
rect 14817 15728 15113 15748
rect 15384 15700 15436 15706
rect 15384 15642 15436 15648
rect 14556 15496 14608 15502
rect 14556 15438 14608 15444
rect 14568 14822 14596 15438
rect 15200 15428 15252 15434
rect 15200 15370 15252 15376
rect 15212 15026 15240 15370
rect 15200 15020 15252 15026
rect 15200 14962 15252 14968
rect 15396 14958 15424 15642
rect 16040 15638 16068 18226
rect 17040 18148 17092 18154
rect 17040 18090 17092 18096
rect 17052 17882 17080 18090
rect 17132 18080 17184 18086
rect 17132 18022 17184 18028
rect 17040 17876 17092 17882
rect 17040 17818 17092 17824
rect 16856 17672 16908 17678
rect 16856 17614 16908 17620
rect 16396 17536 16448 17542
rect 16396 17478 16448 17484
rect 16408 17134 16436 17478
rect 16488 17196 16540 17202
rect 16488 17138 16540 17144
rect 16396 17128 16448 17134
rect 16396 17070 16448 17076
rect 16500 16522 16528 17138
rect 16868 16794 16896 17614
rect 16856 16788 16908 16794
rect 16856 16730 16908 16736
rect 16856 16652 16908 16658
rect 16856 16594 16908 16600
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 16488 16516 16540 16522
rect 16488 16458 16540 16464
rect 16684 16250 16712 16526
rect 16672 16244 16724 16250
rect 16672 16186 16724 16192
rect 16396 15972 16448 15978
rect 16396 15914 16448 15920
rect 16028 15632 16080 15638
rect 16028 15574 16080 15580
rect 15660 15564 15712 15570
rect 15712 15524 15792 15552
rect 15660 15506 15712 15512
rect 15384 14952 15436 14958
rect 15384 14894 15436 14900
rect 14556 14816 14608 14822
rect 14556 14758 14608 14764
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 15200 14816 15252 14822
rect 15200 14758 15252 14764
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 14384 13938 14412 14350
rect 14372 13932 14424 13938
rect 14372 13874 14424 13880
rect 14568 11286 14596 14758
rect 14752 14550 14780 14758
rect 14817 14716 15113 14736
rect 14873 14714 14897 14716
rect 14953 14714 14977 14716
rect 15033 14714 15057 14716
rect 14895 14662 14897 14714
rect 14959 14662 14971 14714
rect 15033 14662 15035 14714
rect 14873 14660 14897 14662
rect 14953 14660 14977 14662
rect 15033 14660 15057 14662
rect 14817 14640 15113 14660
rect 15212 14618 15240 14758
rect 15200 14612 15252 14618
rect 15200 14554 15252 14560
rect 14740 14544 14792 14550
rect 14740 14486 14792 14492
rect 15396 14482 15424 14894
rect 15200 14476 15252 14482
rect 15200 14418 15252 14424
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 14817 13628 15113 13648
rect 14873 13626 14897 13628
rect 14953 13626 14977 13628
rect 15033 13626 15057 13628
rect 14895 13574 14897 13626
rect 14959 13574 14971 13626
rect 15033 13574 15035 13626
rect 14873 13572 14897 13574
rect 14953 13572 14977 13574
rect 15033 13572 15057 13574
rect 14817 13552 15113 13572
rect 14817 12540 15113 12560
rect 14873 12538 14897 12540
rect 14953 12538 14977 12540
rect 15033 12538 15057 12540
rect 14895 12486 14897 12538
rect 14959 12486 14971 12538
rect 15033 12486 15035 12538
rect 14873 12484 14897 12486
rect 14953 12484 14977 12486
rect 15033 12484 15057 12486
rect 14817 12464 15113 12484
rect 14648 12096 14700 12102
rect 14648 12038 14700 12044
rect 14660 11898 14688 12038
rect 14648 11892 14700 11898
rect 14648 11834 14700 11840
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14752 11354 14780 11834
rect 14817 11452 15113 11472
rect 14873 11450 14897 11452
rect 14953 11450 14977 11452
rect 15033 11450 15057 11452
rect 14895 11398 14897 11450
rect 14959 11398 14971 11450
rect 15033 11398 15035 11450
rect 14873 11396 14897 11398
rect 14953 11396 14977 11398
rect 15033 11396 15057 11398
rect 14817 11376 15113 11396
rect 15212 11354 15240 14418
rect 15292 13864 15344 13870
rect 15292 13806 15344 13812
rect 15304 13530 15332 13806
rect 15476 13796 15528 13802
rect 15476 13738 15528 13744
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 14740 11348 14792 11354
rect 14740 11290 14792 11296
rect 15200 11348 15252 11354
rect 15200 11290 15252 11296
rect 14556 11280 14608 11286
rect 14556 11222 14608 11228
rect 15212 11218 15240 11290
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 14648 11076 14700 11082
rect 14648 11018 14700 11024
rect 14556 10600 14608 10606
rect 14556 10542 14608 10548
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 14384 10266 14412 10406
rect 14372 10260 14424 10266
rect 14372 10202 14424 10208
rect 14568 10198 14596 10542
rect 14660 10198 14688 11018
rect 15488 11014 15516 13738
rect 15672 13274 15700 14418
rect 15764 14414 15792 15524
rect 15936 15020 15988 15026
rect 15936 14962 15988 14968
rect 15844 14816 15896 14822
rect 15844 14758 15896 14764
rect 15752 14408 15804 14414
rect 15752 14350 15804 14356
rect 15764 14278 15792 14350
rect 15752 14272 15804 14278
rect 15752 14214 15804 14220
rect 15764 13716 15792 14214
rect 15856 14074 15884 14758
rect 15844 14068 15896 14074
rect 15844 14010 15896 14016
rect 15844 13728 15896 13734
rect 15764 13688 15844 13716
rect 15844 13670 15896 13676
rect 15580 13258 15700 13274
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 15568 13252 15700 13258
rect 15620 13246 15700 13252
rect 15568 13194 15620 13200
rect 15672 12986 15700 13246
rect 15660 12980 15712 12986
rect 15660 12922 15712 12928
rect 15672 12170 15700 12922
rect 15764 12918 15792 13262
rect 15752 12912 15804 12918
rect 15752 12854 15804 12860
rect 15856 12288 15884 13670
rect 15948 13326 15976 14962
rect 16212 13728 16264 13734
rect 16212 13670 16264 13676
rect 16304 13728 16356 13734
rect 16304 13670 16356 13676
rect 15936 13320 15988 13326
rect 15936 13262 15988 13268
rect 16224 12442 16252 13670
rect 16316 13530 16344 13670
rect 16304 13524 16356 13530
rect 16304 13466 16356 13472
rect 16212 12436 16264 12442
rect 16212 12378 16264 12384
rect 15936 12300 15988 12306
rect 15856 12260 15936 12288
rect 15936 12242 15988 12248
rect 15660 12164 15712 12170
rect 15660 12106 15712 12112
rect 15948 11218 15976 12242
rect 16408 11393 16436 15914
rect 16868 15910 16896 16594
rect 17052 16454 17080 17818
rect 17144 17202 17172 18022
rect 17420 17746 17448 18838
rect 18282 18524 18578 18544
rect 18338 18522 18362 18524
rect 18418 18522 18442 18524
rect 18498 18522 18522 18524
rect 18360 18470 18362 18522
rect 18424 18470 18436 18522
rect 18498 18470 18500 18522
rect 18338 18468 18362 18470
rect 18418 18468 18442 18470
rect 18498 18468 18522 18470
rect 18282 18448 18578 18468
rect 17500 17876 17552 17882
rect 17500 17818 17552 17824
rect 17512 17746 17540 17818
rect 17408 17740 17460 17746
rect 17408 17682 17460 17688
rect 17500 17740 17552 17746
rect 17500 17682 17552 17688
rect 17684 17740 17736 17746
rect 17684 17682 17736 17688
rect 17960 17740 18012 17746
rect 17960 17682 18012 17688
rect 17132 17196 17184 17202
rect 17132 17138 17184 17144
rect 17420 17134 17448 17682
rect 17498 17640 17554 17649
rect 17498 17575 17554 17584
rect 17512 17270 17540 17575
rect 17500 17264 17552 17270
rect 17500 17206 17552 17212
rect 17408 17128 17460 17134
rect 17408 17070 17460 17076
rect 17224 16992 17276 16998
rect 17224 16934 17276 16940
rect 17236 16658 17264 16934
rect 17224 16652 17276 16658
rect 17224 16594 17276 16600
rect 17040 16448 17092 16454
rect 17040 16390 17092 16396
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16764 14340 16816 14346
rect 16764 14282 16816 14288
rect 16776 13938 16804 14282
rect 16764 13932 16816 13938
rect 16764 13874 16816 13880
rect 16672 13388 16724 13394
rect 16672 13330 16724 13336
rect 16488 13252 16540 13258
rect 16488 13194 16540 13200
rect 16500 12850 16528 13194
rect 16488 12844 16540 12850
rect 16488 12786 16540 12792
rect 16684 12782 16712 13330
rect 16672 12776 16724 12782
rect 16672 12718 16724 12724
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 16776 11626 16804 12378
rect 16764 11620 16816 11626
rect 16764 11562 16816 11568
rect 16394 11384 16450 11393
rect 16394 11319 16450 11328
rect 15936 11212 15988 11218
rect 15936 11154 15988 11160
rect 15476 11008 15528 11014
rect 15476 10950 15528 10956
rect 16408 10962 16436 11319
rect 16868 11082 16896 15846
rect 16948 15360 17000 15366
rect 16948 15302 17000 15308
rect 16960 12374 16988 15302
rect 17052 13716 17080 16390
rect 17224 13728 17276 13734
rect 17052 13688 17224 13716
rect 17224 13670 17276 13676
rect 17236 13530 17264 13670
rect 17224 13524 17276 13530
rect 17224 13466 17276 13472
rect 17132 12844 17184 12850
rect 17132 12786 17184 12792
rect 17144 12442 17172 12786
rect 17132 12436 17184 12442
rect 17132 12378 17184 12384
rect 16948 12368 17000 12374
rect 16948 12310 17000 12316
rect 17236 11642 17264 13466
rect 17408 13456 17460 13462
rect 17408 13398 17460 13404
rect 17420 11762 17448 13398
rect 17408 11756 17460 11762
rect 17408 11698 17460 11704
rect 17236 11614 17448 11642
rect 16672 11076 16724 11082
rect 16672 11018 16724 11024
rect 16856 11076 16908 11082
rect 16856 11018 16908 11024
rect 16408 10934 16528 10962
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 14740 10668 14792 10674
rect 14740 10610 14792 10616
rect 14556 10192 14608 10198
rect 14556 10134 14608 10140
rect 14648 10192 14700 10198
rect 14648 10134 14700 10140
rect 14752 9926 14780 10610
rect 14817 10364 15113 10384
rect 14873 10362 14897 10364
rect 14953 10362 14977 10364
rect 15033 10362 15057 10364
rect 14895 10310 14897 10362
rect 14959 10310 14971 10362
rect 15033 10310 15035 10362
rect 14873 10308 14897 10310
rect 14953 10308 14977 10310
rect 15033 10308 15057 10310
rect 14817 10288 15113 10308
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 14752 9518 14780 9862
rect 15672 9586 15700 10066
rect 15660 9580 15712 9586
rect 15660 9522 15712 9528
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 14556 9376 14608 9382
rect 14556 9318 14608 9324
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14476 8498 14504 8774
rect 14464 8492 14516 8498
rect 14464 8434 14516 8440
rect 14568 8378 14596 9318
rect 14752 8974 14780 9454
rect 15200 9376 15252 9382
rect 15200 9318 15252 9324
rect 15660 9376 15712 9382
rect 15660 9318 15712 9324
rect 14817 9276 15113 9296
rect 14873 9274 14897 9276
rect 14953 9274 14977 9276
rect 15033 9274 15057 9276
rect 14895 9222 14897 9274
rect 14959 9222 14971 9274
rect 15033 9222 15035 9274
rect 14873 9220 14897 9222
rect 14953 9220 14977 9222
rect 15033 9220 15057 9222
rect 14817 9200 15113 9220
rect 15212 9042 15240 9318
rect 15672 9178 15700 9318
rect 15660 9172 15712 9178
rect 15660 9114 15712 9120
rect 15200 9036 15252 9042
rect 15200 8978 15252 8984
rect 14740 8968 14792 8974
rect 14740 8910 14792 8916
rect 14832 8492 14884 8498
rect 14832 8434 14884 8440
rect 14844 8378 14872 8434
rect 14568 8350 14872 8378
rect 14568 7342 14596 8350
rect 14648 8288 14700 8294
rect 14648 8230 14700 8236
rect 14660 8090 14688 8230
rect 14817 8188 15113 8208
rect 14873 8186 14897 8188
rect 14953 8186 14977 8188
rect 15033 8186 15057 8188
rect 14895 8134 14897 8186
rect 14959 8134 14971 8186
rect 15033 8134 15035 8186
rect 14873 8132 14897 8134
rect 14953 8132 14977 8134
rect 15033 8132 15057 8134
rect 14817 8112 15113 8132
rect 14648 8084 14700 8090
rect 14648 8026 14700 8032
rect 14832 7744 14884 7750
rect 14832 7686 14884 7692
rect 15568 7744 15620 7750
rect 15568 7686 15620 7692
rect 14844 7449 14872 7686
rect 14830 7440 14886 7449
rect 15580 7410 15608 7686
rect 14830 7375 14886 7384
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 14556 7336 14608 7342
rect 14556 7278 14608 7284
rect 15384 7200 15436 7206
rect 15384 7142 15436 7148
rect 14817 7100 15113 7120
rect 14873 7098 14897 7100
rect 14953 7098 14977 7100
rect 15033 7098 15057 7100
rect 14895 7046 14897 7098
rect 14959 7046 14971 7098
rect 15033 7046 15035 7098
rect 14873 7044 14897 7046
rect 14953 7044 14977 7046
rect 15033 7044 15057 7046
rect 14817 7024 15113 7044
rect 14280 6928 14332 6934
rect 14280 6870 14332 6876
rect 14648 6928 14700 6934
rect 14648 6870 14700 6876
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 13648 6322 13676 6734
rect 14372 6384 14424 6390
rect 14372 6326 14424 6332
rect 13636 6316 13688 6322
rect 13636 6258 13688 6264
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 13832 5794 13860 6258
rect 14188 6112 14240 6118
rect 14188 6054 14240 6060
rect 13740 5778 13860 5794
rect 13728 5772 13860 5778
rect 13780 5766 13860 5772
rect 13728 5714 13780 5720
rect 13832 5370 13860 5766
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 14200 5166 14228 6054
rect 14280 5568 14332 5574
rect 14280 5510 14332 5516
rect 14292 5234 14320 5510
rect 14280 5228 14332 5234
rect 14280 5170 14332 5176
rect 14188 5160 14240 5166
rect 14188 5102 14240 5108
rect 13912 5024 13964 5030
rect 13912 4966 13964 4972
rect 13544 4820 13596 4826
rect 13544 4762 13596 4768
rect 13268 4208 13320 4214
rect 13268 4150 13320 4156
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 13452 3596 13504 3602
rect 13452 3538 13504 3544
rect 12820 2582 12848 3538
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13268 3392 13320 3398
rect 13268 3334 13320 3340
rect 13280 3058 13308 3334
rect 13268 3052 13320 3058
rect 13268 2994 13320 3000
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 12808 2576 12860 2582
rect 12808 2518 12860 2524
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 12808 2304 12860 2310
rect 12808 2246 12860 2252
rect 12820 800 12848 2246
rect 13280 800 13308 2790
rect 13372 2514 13400 3470
rect 13464 2582 13492 3538
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13452 2576 13504 2582
rect 13452 2518 13504 2524
rect 13360 2508 13412 2514
rect 13360 2450 13412 2456
rect 13740 800 13768 3334
rect 13924 2990 13952 4966
rect 14292 4078 14320 5170
rect 14384 5098 14412 6326
rect 14660 6118 14688 6870
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 14556 6112 14608 6118
rect 14556 6054 14608 6060
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14568 5914 14596 6054
rect 14817 6012 15113 6032
rect 14873 6010 14897 6012
rect 14953 6010 14977 6012
rect 15033 6010 15057 6012
rect 14895 5958 14897 6010
rect 14959 5958 14971 6010
rect 15033 5958 15035 6010
rect 14873 5956 14897 5958
rect 14953 5956 14977 5958
rect 15033 5956 15057 5958
rect 14817 5936 15113 5956
rect 14556 5908 14608 5914
rect 14556 5850 14608 5856
rect 15304 5302 15332 6734
rect 15396 5710 15424 7142
rect 15752 6112 15804 6118
rect 15752 6054 15804 6060
rect 15764 5778 15792 6054
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 15292 5296 15344 5302
rect 15292 5238 15344 5244
rect 14372 5092 14424 5098
rect 14372 5034 14424 5040
rect 14817 4924 15113 4944
rect 14873 4922 14897 4924
rect 14953 4922 14977 4924
rect 15033 4922 15057 4924
rect 14895 4870 14897 4922
rect 14959 4870 14971 4922
rect 15033 4870 15035 4922
rect 14873 4868 14897 4870
rect 14953 4868 14977 4870
rect 15033 4868 15057 4870
rect 14817 4848 15113 4868
rect 15304 4622 15332 5238
rect 15396 5234 15424 5646
rect 15476 5636 15528 5642
rect 15476 5578 15528 5584
rect 15384 5228 15436 5234
rect 15384 5170 15436 5176
rect 15488 5166 15516 5578
rect 16040 5370 16068 10746
rect 16212 9988 16264 9994
rect 16212 9930 16264 9936
rect 16224 9586 16252 9930
rect 16212 9580 16264 9586
rect 16212 9522 16264 9528
rect 16396 8900 16448 8906
rect 16396 8842 16448 8848
rect 16212 8356 16264 8362
rect 16212 8298 16264 8304
rect 16224 7886 16252 8298
rect 16212 7880 16264 7886
rect 16212 7822 16264 7828
rect 16408 7546 16436 8842
rect 16500 8566 16528 10934
rect 16580 10124 16632 10130
rect 16580 10066 16632 10072
rect 16592 8838 16620 10066
rect 16684 9926 16712 11018
rect 16764 10124 16816 10130
rect 16764 10066 16816 10072
rect 16672 9920 16724 9926
rect 16672 9862 16724 9868
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16672 8832 16724 8838
rect 16672 8774 16724 8780
rect 16488 8560 16540 8566
rect 16488 8502 16540 8508
rect 16500 8090 16528 8502
rect 16592 8090 16620 8774
rect 16684 8634 16712 8774
rect 16776 8634 16804 10066
rect 16868 9654 16896 11018
rect 17132 10464 17184 10470
rect 17132 10406 17184 10412
rect 16856 9648 16908 9654
rect 16908 9608 16988 9636
rect 16856 9590 16908 9596
rect 16868 9382 16896 9590
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16672 8628 16724 8634
rect 16672 8570 16724 8576
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 16670 8392 16726 8401
rect 16670 8327 16672 8336
rect 16724 8327 16726 8336
rect 16672 8298 16724 8304
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16580 8084 16632 8090
rect 16580 8026 16632 8032
rect 16592 7886 16620 8026
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16212 6860 16264 6866
rect 16212 6802 16264 6808
rect 16224 6746 16252 6802
rect 16224 6718 16344 6746
rect 16316 6322 16344 6718
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 16408 5370 16436 7482
rect 16592 7290 16620 7822
rect 16776 7478 16804 8570
rect 16856 7948 16908 7954
rect 16856 7890 16908 7896
rect 16764 7472 16816 7478
rect 16764 7414 16816 7420
rect 16500 7262 16620 7290
rect 16500 6662 16528 7262
rect 16580 7200 16632 7206
rect 16580 7142 16632 7148
rect 16488 6656 16540 6662
rect 16488 6598 16540 6604
rect 16488 6112 16540 6118
rect 16488 6054 16540 6060
rect 16500 5914 16528 6054
rect 16488 5908 16540 5914
rect 16488 5850 16540 5856
rect 16028 5364 16080 5370
rect 16028 5306 16080 5312
rect 16396 5364 16448 5370
rect 16396 5306 16448 5312
rect 15476 5160 15528 5166
rect 15476 5102 15528 5108
rect 15568 5024 15620 5030
rect 15568 4966 15620 4972
rect 15580 4690 15608 4966
rect 15568 4684 15620 4690
rect 15568 4626 15620 4632
rect 15292 4616 15344 4622
rect 15292 4558 15344 4564
rect 14280 4072 14332 4078
rect 14280 4014 14332 4020
rect 15200 3936 15252 3942
rect 15200 3878 15252 3884
rect 14817 3836 15113 3856
rect 14873 3834 14897 3836
rect 14953 3834 14977 3836
rect 15033 3834 15057 3836
rect 14895 3782 14897 3834
rect 14959 3782 14971 3834
rect 15033 3782 15035 3834
rect 14873 3780 14897 3782
rect 14953 3780 14977 3782
rect 15033 3780 15057 3782
rect 14817 3760 15113 3780
rect 14556 3392 14608 3398
rect 14556 3334 14608 3340
rect 13912 2984 13964 2990
rect 13912 2926 13964 2932
rect 13820 2916 13872 2922
rect 13820 2858 13872 2864
rect 13832 2514 13860 2858
rect 13820 2508 13872 2514
rect 13820 2450 13872 2456
rect 14004 2304 14056 2310
rect 14004 2246 14056 2252
rect 14016 1170 14044 2246
rect 14016 1142 14136 1170
rect 14108 800 14136 1142
rect 14568 800 14596 3334
rect 15212 3058 15240 3878
rect 15304 3602 15332 4558
rect 15476 4480 15528 4486
rect 15476 4422 15528 4428
rect 15488 3942 15516 4422
rect 15568 4140 15620 4146
rect 15568 4082 15620 4088
rect 15476 3936 15528 3942
rect 15476 3878 15528 3884
rect 15292 3596 15344 3602
rect 15292 3538 15344 3544
rect 15488 3126 15516 3878
rect 15580 3670 15608 4082
rect 16040 4010 16068 5306
rect 16408 4078 16436 5306
rect 16488 4684 16540 4690
rect 16488 4626 16540 4632
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16028 4004 16080 4010
rect 16028 3946 16080 3952
rect 15844 3936 15896 3942
rect 15844 3878 15896 3884
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 15568 3664 15620 3670
rect 15568 3606 15620 3612
rect 15476 3120 15528 3126
rect 15476 3062 15528 3068
rect 15200 3052 15252 3058
rect 15200 2994 15252 3000
rect 15856 2922 15884 3878
rect 16316 3738 16344 3878
rect 16500 3738 16528 4626
rect 16304 3732 16356 3738
rect 16304 3674 16356 3680
rect 16488 3732 16540 3738
rect 16488 3674 16540 3680
rect 16500 3126 16528 3674
rect 16592 3602 16620 7142
rect 16868 7002 16896 7890
rect 16856 6996 16908 7002
rect 16856 6938 16908 6944
rect 16868 5710 16896 6938
rect 16856 5704 16908 5710
rect 16856 5646 16908 5652
rect 16580 3596 16632 3602
rect 16580 3538 16632 3544
rect 16488 3120 16540 3126
rect 16488 3062 16540 3068
rect 14740 2916 14792 2922
rect 14740 2858 14792 2864
rect 15844 2916 15896 2922
rect 15844 2858 15896 2864
rect 16580 2916 16632 2922
rect 16580 2858 16632 2864
rect 16856 2916 16908 2922
rect 16856 2858 16908 2864
rect 14752 2514 14780 2858
rect 15384 2848 15436 2854
rect 15384 2790 15436 2796
rect 14817 2748 15113 2768
rect 14873 2746 14897 2748
rect 14953 2746 14977 2748
rect 15033 2746 15057 2748
rect 14895 2694 14897 2746
rect 14959 2694 14971 2746
rect 15033 2694 15035 2746
rect 14873 2692 14897 2694
rect 14953 2692 14977 2694
rect 15033 2692 15057 2694
rect 14817 2672 15113 2692
rect 14740 2508 14792 2514
rect 14740 2450 14792 2456
rect 15016 2372 15068 2378
rect 15016 2314 15068 2320
rect 15028 800 15056 2314
rect 15396 898 15424 2790
rect 16592 2514 16620 2858
rect 16868 2514 16896 2858
rect 16580 2508 16632 2514
rect 16580 2450 16632 2456
rect 16856 2508 16908 2514
rect 16856 2450 16908 2456
rect 15936 2304 15988 2310
rect 15936 2246 15988 2252
rect 16396 2304 16448 2310
rect 16396 2246 16448 2252
rect 16856 2304 16908 2310
rect 16856 2246 16908 2252
rect 15396 870 15516 898
rect 15488 800 15516 870
rect 15948 800 15976 2246
rect 16408 800 16436 2246
rect 16868 800 16896 2246
rect 6366 232 6422 241
rect 6366 167 6422 176
rect 6458 0 6514 800
rect 6918 0 6974 800
rect 7378 0 7434 800
rect 7838 0 7894 800
rect 8298 0 8354 800
rect 8758 0 8814 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 10046 0 10102 800
rect 10506 0 10562 800
rect 10966 0 11022 800
rect 11426 0 11482 800
rect 11886 0 11942 800
rect 12346 0 12402 800
rect 12806 0 12862 800
rect 13266 0 13322 800
rect 13726 0 13782 800
rect 14094 0 14150 800
rect 14554 0 14610 800
rect 15014 0 15070 800
rect 15474 0 15530 800
rect 15934 0 15990 800
rect 16394 0 16450 800
rect 16854 0 16910 800
rect 16960 649 16988 9608
rect 17144 7993 17172 10406
rect 17130 7984 17186 7993
rect 17130 7919 17186 7928
rect 17132 6792 17184 6798
rect 17132 6734 17184 6740
rect 17144 6254 17172 6734
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 17224 6248 17276 6254
rect 17224 6190 17276 6196
rect 17236 5914 17264 6190
rect 17224 5908 17276 5914
rect 17224 5850 17276 5856
rect 17040 5568 17092 5574
rect 17040 5510 17092 5516
rect 17052 2990 17080 5510
rect 17328 4826 17356 6258
rect 17316 4820 17368 4826
rect 17316 4762 17368 4768
rect 17224 3528 17276 3534
rect 17420 3505 17448 11614
rect 17512 8634 17540 17206
rect 17696 16998 17724 17682
rect 17972 17270 18000 17682
rect 18282 17436 18578 17456
rect 18338 17434 18362 17436
rect 18418 17434 18442 17436
rect 18498 17434 18522 17436
rect 18360 17382 18362 17434
rect 18424 17382 18436 17434
rect 18498 17382 18500 17434
rect 18338 17380 18362 17382
rect 18418 17380 18442 17382
rect 18498 17380 18522 17382
rect 18282 17360 18578 17380
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 17776 17128 17828 17134
rect 17776 17070 17828 17076
rect 17684 16992 17736 16998
rect 17684 16934 17736 16940
rect 17696 16522 17724 16934
rect 17684 16516 17736 16522
rect 17684 16458 17736 16464
rect 17788 15570 17816 17070
rect 18052 17060 18104 17066
rect 18052 17002 18104 17008
rect 17868 16584 17920 16590
rect 17920 16532 18000 16538
rect 17868 16526 18000 16532
rect 17880 16510 18000 16526
rect 17972 16250 18000 16510
rect 17960 16244 18012 16250
rect 17960 16186 18012 16192
rect 17776 15564 17828 15570
rect 17776 15506 17828 15512
rect 17960 15564 18012 15570
rect 17960 15506 18012 15512
rect 17972 15026 18000 15506
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 17960 14544 18012 14550
rect 17960 14486 18012 14492
rect 17972 12866 18000 14486
rect 18064 14074 18092 17002
rect 18282 16348 18578 16368
rect 18338 16346 18362 16348
rect 18418 16346 18442 16348
rect 18498 16346 18522 16348
rect 18360 16294 18362 16346
rect 18424 16294 18436 16346
rect 18498 16294 18500 16346
rect 18338 16292 18362 16294
rect 18418 16292 18442 16294
rect 18498 16292 18522 16294
rect 18282 16272 18578 16292
rect 18708 16250 18736 22607
rect 20626 22264 20682 22273
rect 20626 22199 20682 22208
rect 19154 21720 19210 21729
rect 19154 21655 19210 21664
rect 18880 19304 18932 19310
rect 18880 19246 18932 19252
rect 18144 16244 18196 16250
rect 18144 16186 18196 16192
rect 18696 16244 18748 16250
rect 18696 16186 18748 16192
rect 18052 14068 18104 14074
rect 18052 14010 18104 14016
rect 17880 12838 18000 12866
rect 18064 12850 18092 14010
rect 18156 14006 18184 16186
rect 18892 15706 18920 19246
rect 19168 19174 19196 21655
rect 19246 21312 19302 21321
rect 19246 21247 19302 21256
rect 19260 19242 19288 21247
rect 20442 20768 20498 20777
rect 20442 20703 20498 20712
rect 19984 20392 20036 20398
rect 19984 20334 20036 20340
rect 19892 19712 19944 19718
rect 19892 19654 19944 19660
rect 19904 19378 19932 19654
rect 19892 19372 19944 19378
rect 19892 19314 19944 19320
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 19248 19236 19300 19242
rect 19248 19178 19300 19184
rect 19156 19168 19208 19174
rect 19156 19110 19208 19116
rect 19352 18630 19380 19246
rect 19340 18624 19392 18630
rect 19340 18566 19392 18572
rect 19352 17746 19380 18566
rect 19800 18080 19852 18086
rect 19800 18022 19852 18028
rect 19340 17740 19392 17746
rect 19340 17682 19392 17688
rect 19616 17740 19668 17746
rect 19616 17682 19668 17688
rect 19246 17504 19302 17513
rect 19246 17439 19302 17448
rect 19064 17060 19116 17066
rect 19064 17002 19116 17008
rect 18972 16652 19024 16658
rect 18972 16594 19024 16600
rect 18984 16454 19012 16594
rect 18972 16448 19024 16454
rect 18972 16390 19024 16396
rect 18984 16114 19012 16390
rect 18972 16108 19024 16114
rect 18972 16050 19024 16056
rect 19076 15706 19104 17002
rect 19260 16794 19288 17439
rect 19248 16788 19300 16794
rect 19248 16730 19300 16736
rect 19524 16652 19576 16658
rect 19524 16594 19576 16600
rect 18880 15700 18932 15706
rect 18880 15642 18932 15648
rect 19064 15700 19116 15706
rect 19064 15642 19116 15648
rect 18282 15260 18578 15280
rect 18338 15258 18362 15260
rect 18418 15258 18442 15260
rect 18498 15258 18522 15260
rect 18360 15206 18362 15258
rect 18424 15206 18436 15258
rect 18498 15206 18500 15258
rect 18338 15204 18362 15206
rect 18418 15204 18442 15206
rect 18498 15204 18522 15206
rect 18282 15184 18578 15204
rect 19076 15094 19104 15642
rect 19340 15496 19392 15502
rect 19340 15438 19392 15444
rect 19064 15088 19116 15094
rect 19064 15030 19116 15036
rect 18788 15020 18840 15026
rect 18788 14962 18840 14968
rect 19248 15020 19300 15026
rect 19248 14962 19300 14968
rect 18800 14278 18828 14962
rect 19260 14482 19288 14962
rect 19352 14890 19380 15438
rect 19340 14884 19392 14890
rect 19340 14826 19392 14832
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 19444 14618 19472 14758
rect 19432 14612 19484 14618
rect 19432 14554 19484 14560
rect 19248 14476 19300 14482
rect 19248 14418 19300 14424
rect 18788 14272 18840 14278
rect 18788 14214 18840 14220
rect 18282 14172 18578 14192
rect 18338 14170 18362 14172
rect 18418 14170 18442 14172
rect 18498 14170 18522 14172
rect 18360 14118 18362 14170
rect 18424 14118 18436 14170
rect 18498 14118 18500 14170
rect 18338 14116 18362 14118
rect 18418 14116 18442 14118
rect 18498 14116 18522 14118
rect 18282 14096 18578 14116
rect 18144 14000 18196 14006
rect 18144 13942 18196 13948
rect 18800 13870 18828 14214
rect 19260 13938 19288 14418
rect 18972 13932 19024 13938
rect 19248 13932 19300 13938
rect 18972 13874 19024 13880
rect 19168 13892 19248 13920
rect 18788 13864 18840 13870
rect 18788 13806 18840 13812
rect 18788 13388 18840 13394
rect 18788 13330 18840 13336
rect 18604 13320 18656 13326
rect 18604 13262 18656 13268
rect 18144 13184 18196 13190
rect 18144 13126 18196 13132
rect 18052 12844 18104 12850
rect 17684 12708 17736 12714
rect 17684 12650 17736 12656
rect 17696 11558 17724 12650
rect 17776 11688 17828 11694
rect 17774 11656 17776 11665
rect 17828 11656 17830 11665
rect 17774 11591 17830 11600
rect 17684 11552 17736 11558
rect 17684 11494 17736 11500
rect 17592 11348 17644 11354
rect 17592 11290 17644 11296
rect 17604 9518 17632 11290
rect 17880 10826 17908 12838
rect 18052 12786 18104 12792
rect 18156 12646 18184 13126
rect 18282 13084 18578 13104
rect 18338 13082 18362 13084
rect 18418 13082 18442 13084
rect 18498 13082 18522 13084
rect 18360 13030 18362 13082
rect 18424 13030 18436 13082
rect 18498 13030 18500 13082
rect 18338 13028 18362 13030
rect 18418 13028 18442 13030
rect 18498 13028 18522 13030
rect 18282 13008 18578 13028
rect 18616 12918 18644 13262
rect 18696 13252 18748 13258
rect 18696 13194 18748 13200
rect 18604 12912 18656 12918
rect 18604 12854 18656 12860
rect 18052 12640 18104 12646
rect 18052 12582 18104 12588
rect 18144 12640 18196 12646
rect 18144 12582 18196 12588
rect 18064 12442 18092 12582
rect 18616 12442 18644 12854
rect 18708 12782 18736 13194
rect 18800 12986 18828 13330
rect 18880 13320 18932 13326
rect 18880 13262 18932 13268
rect 18892 12986 18920 13262
rect 18984 13258 19012 13874
rect 19168 13326 19196 13892
rect 19248 13874 19300 13880
rect 19432 13796 19484 13802
rect 19432 13738 19484 13744
rect 19340 13728 19392 13734
rect 19340 13670 19392 13676
rect 19352 13530 19380 13670
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 19156 13320 19208 13326
rect 19156 13262 19208 13268
rect 18972 13252 19024 13258
rect 18972 13194 19024 13200
rect 18788 12980 18840 12986
rect 18788 12922 18840 12928
rect 18880 12980 18932 12986
rect 18880 12922 18932 12928
rect 19156 12912 19208 12918
rect 19156 12854 19208 12860
rect 18696 12776 18748 12782
rect 18696 12718 18748 12724
rect 18052 12436 18104 12442
rect 18052 12378 18104 12384
rect 18604 12436 18656 12442
rect 18604 12378 18656 12384
rect 18144 12300 18196 12306
rect 18144 12242 18196 12248
rect 18156 11880 18184 12242
rect 18604 12232 18656 12238
rect 18604 12174 18656 12180
rect 18282 11996 18578 12016
rect 18338 11994 18362 11996
rect 18418 11994 18442 11996
rect 18498 11994 18522 11996
rect 18360 11942 18362 11994
rect 18424 11942 18436 11994
rect 18498 11942 18500 11994
rect 18338 11940 18362 11942
rect 18418 11940 18442 11942
rect 18498 11940 18522 11942
rect 18282 11920 18578 11940
rect 18156 11852 18552 11880
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 18236 11756 18288 11762
rect 18236 11698 18288 11704
rect 17972 11540 18000 11698
rect 18248 11626 18276 11698
rect 18524 11694 18552 11852
rect 18616 11762 18644 12174
rect 18604 11756 18656 11762
rect 18604 11698 18656 11704
rect 18420 11688 18472 11694
rect 18418 11656 18420 11665
rect 18512 11688 18564 11694
rect 18472 11656 18474 11665
rect 18236 11620 18288 11626
rect 18512 11630 18564 11636
rect 18418 11591 18474 11600
rect 18236 11562 18288 11568
rect 18144 11552 18196 11558
rect 17972 11512 18144 11540
rect 18144 11494 18196 11500
rect 18432 11506 18460 11591
rect 18708 11506 18736 12718
rect 18972 12436 19024 12442
rect 18972 12378 19024 12384
rect 18984 11558 19012 12378
rect 19062 11928 19118 11937
rect 19062 11863 19118 11872
rect 19076 11830 19104 11863
rect 19064 11824 19116 11830
rect 19064 11766 19116 11772
rect 18432 11478 18736 11506
rect 18972 11552 19024 11558
rect 18972 11494 19024 11500
rect 18052 11212 18104 11218
rect 18052 11154 18104 11160
rect 17960 11144 18012 11150
rect 17960 11086 18012 11092
rect 17696 10798 17908 10826
rect 17696 10606 17724 10798
rect 17684 10600 17736 10606
rect 17684 10542 17736 10548
rect 17868 10600 17920 10606
rect 17868 10542 17920 10548
rect 17592 9512 17644 9518
rect 17592 9454 17644 9460
rect 17500 8628 17552 8634
rect 17500 8570 17552 8576
rect 17696 6254 17724 10542
rect 17880 10198 17908 10542
rect 17868 10192 17920 10198
rect 17868 10134 17920 10140
rect 17880 9722 17908 10134
rect 17868 9716 17920 9722
rect 17868 9658 17920 9664
rect 17776 8288 17828 8294
rect 17776 8230 17828 8236
rect 17788 8129 17816 8230
rect 17774 8120 17830 8129
rect 17774 8055 17830 8064
rect 17868 8084 17920 8090
rect 17868 8026 17920 8032
rect 17880 7954 17908 8026
rect 17868 7948 17920 7954
rect 17868 7890 17920 7896
rect 17972 7018 18000 11086
rect 18064 9654 18092 11154
rect 18144 11144 18196 11150
rect 18144 11086 18196 11092
rect 18156 10674 18184 11086
rect 18282 10908 18578 10928
rect 18338 10906 18362 10908
rect 18418 10906 18442 10908
rect 18498 10906 18522 10908
rect 18360 10854 18362 10906
rect 18424 10854 18436 10906
rect 18498 10854 18500 10906
rect 18338 10852 18362 10854
rect 18418 10852 18442 10854
rect 18498 10852 18522 10854
rect 18282 10832 18578 10852
rect 18144 10668 18196 10674
rect 18144 10610 18196 10616
rect 18604 10668 18656 10674
rect 18604 10610 18656 10616
rect 18144 10464 18196 10470
rect 18144 10406 18196 10412
rect 18052 9648 18104 9654
rect 18052 9590 18104 9596
rect 18156 9518 18184 10406
rect 18616 10198 18644 10610
rect 18604 10192 18656 10198
rect 18604 10134 18656 10140
rect 18282 9820 18578 9840
rect 18338 9818 18362 9820
rect 18418 9818 18442 9820
rect 18498 9818 18522 9820
rect 18360 9766 18362 9818
rect 18424 9766 18436 9818
rect 18498 9766 18500 9818
rect 18338 9764 18362 9766
rect 18418 9764 18442 9766
rect 18498 9764 18522 9766
rect 18282 9744 18578 9764
rect 18326 9616 18382 9625
rect 18616 9586 18644 10134
rect 18326 9551 18328 9560
rect 18380 9551 18382 9560
rect 18604 9580 18656 9586
rect 18328 9522 18380 9528
rect 18604 9522 18656 9528
rect 18144 9512 18196 9518
rect 18144 9454 18196 9460
rect 18602 9480 18658 9489
rect 18602 9415 18658 9424
rect 18282 8732 18578 8752
rect 18338 8730 18362 8732
rect 18418 8730 18442 8732
rect 18498 8730 18522 8732
rect 18360 8678 18362 8730
rect 18424 8678 18436 8730
rect 18498 8678 18500 8730
rect 18338 8676 18362 8678
rect 18418 8676 18442 8678
rect 18498 8676 18522 8678
rect 18282 8656 18578 8676
rect 18144 8492 18196 8498
rect 18144 8434 18196 8440
rect 18052 8288 18104 8294
rect 18052 8230 18104 8236
rect 18064 7342 18092 8230
rect 18156 8090 18184 8434
rect 18420 8288 18472 8294
rect 18420 8230 18472 8236
rect 18432 8090 18460 8230
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 18420 8084 18472 8090
rect 18420 8026 18472 8032
rect 18282 7644 18578 7664
rect 18338 7642 18362 7644
rect 18418 7642 18442 7644
rect 18498 7642 18522 7644
rect 18360 7590 18362 7642
rect 18424 7590 18436 7642
rect 18498 7590 18500 7642
rect 18338 7588 18362 7590
rect 18418 7588 18442 7590
rect 18498 7588 18522 7590
rect 18282 7568 18578 7588
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 17972 6990 18092 7018
rect 17684 6248 17736 6254
rect 17684 6190 17736 6196
rect 17960 5840 18012 5846
rect 17958 5808 17960 5817
rect 18012 5808 18014 5817
rect 17958 5743 18014 5752
rect 17868 5296 17920 5302
rect 17868 5238 17920 5244
rect 17880 4690 17908 5238
rect 17958 4856 18014 4865
rect 17958 4791 18014 4800
rect 17868 4684 17920 4690
rect 17868 4626 17920 4632
rect 17972 4282 18000 4791
rect 17960 4276 18012 4282
rect 17960 4218 18012 4224
rect 17224 3470 17276 3476
rect 17406 3496 17462 3505
rect 17040 2984 17092 2990
rect 17040 2926 17092 2932
rect 17236 2514 17264 3470
rect 17406 3431 17462 3440
rect 17776 3392 17828 3398
rect 17776 3334 17828 3340
rect 17224 2508 17276 2514
rect 17224 2450 17276 2456
rect 17316 2304 17368 2310
rect 17316 2246 17368 2252
rect 17328 800 17356 2246
rect 17788 800 17816 3334
rect 18064 2990 18092 6990
rect 18616 6866 18644 9415
rect 18604 6860 18656 6866
rect 18604 6802 18656 6808
rect 18144 6792 18196 6798
rect 18144 6734 18196 6740
rect 18156 6458 18184 6734
rect 18282 6556 18578 6576
rect 18338 6554 18362 6556
rect 18418 6554 18442 6556
rect 18498 6554 18522 6556
rect 18360 6502 18362 6554
rect 18424 6502 18436 6554
rect 18498 6502 18500 6554
rect 18338 6500 18362 6502
rect 18418 6500 18442 6502
rect 18498 6500 18522 6502
rect 18282 6480 18578 6500
rect 18144 6452 18196 6458
rect 18144 6394 18196 6400
rect 18708 6118 18736 11478
rect 18788 11280 18840 11286
rect 18788 11222 18840 11228
rect 18800 9382 18828 11222
rect 18880 11008 18932 11014
rect 18880 10950 18932 10956
rect 18892 10441 18920 10950
rect 18878 10432 18934 10441
rect 18878 10367 18934 10376
rect 18788 9376 18840 9382
rect 18788 9318 18840 9324
rect 18696 6112 18748 6118
rect 18696 6054 18748 6060
rect 18708 5914 18736 6054
rect 18696 5908 18748 5914
rect 18696 5850 18748 5856
rect 18604 5704 18656 5710
rect 18604 5646 18656 5652
rect 18282 5468 18578 5488
rect 18338 5466 18362 5468
rect 18418 5466 18442 5468
rect 18498 5466 18522 5468
rect 18360 5414 18362 5466
rect 18424 5414 18436 5466
rect 18498 5414 18500 5466
rect 18338 5412 18362 5414
rect 18418 5412 18442 5414
rect 18498 5412 18522 5414
rect 18282 5392 18578 5412
rect 18616 5098 18644 5646
rect 18604 5092 18656 5098
rect 18604 5034 18656 5040
rect 18282 4380 18578 4400
rect 18338 4378 18362 4380
rect 18418 4378 18442 4380
rect 18498 4378 18522 4380
rect 18360 4326 18362 4378
rect 18424 4326 18436 4378
rect 18498 4326 18500 4378
rect 18338 4324 18362 4326
rect 18418 4324 18442 4326
rect 18498 4324 18522 4326
rect 18282 4304 18578 4324
rect 18144 3596 18196 3602
rect 18144 3538 18196 3544
rect 18156 3058 18184 3538
rect 18282 3292 18578 3312
rect 18338 3290 18362 3292
rect 18418 3290 18442 3292
rect 18498 3290 18522 3292
rect 18360 3238 18362 3290
rect 18424 3238 18436 3290
rect 18498 3238 18500 3290
rect 18338 3236 18362 3238
rect 18418 3236 18442 3238
rect 18498 3236 18522 3238
rect 18282 3216 18578 3236
rect 18144 3052 18196 3058
rect 18144 2994 18196 3000
rect 18052 2984 18104 2990
rect 18708 2961 18736 5850
rect 18052 2926 18104 2932
rect 18694 2952 18750 2961
rect 18512 2916 18564 2922
rect 18694 2887 18750 2896
rect 18512 2858 18564 2864
rect 18524 2514 18552 2858
rect 18604 2848 18656 2854
rect 18604 2790 18656 2796
rect 18512 2508 18564 2514
rect 18512 2450 18564 2456
rect 18144 2304 18196 2310
rect 18144 2246 18196 2252
rect 18156 1170 18184 2246
rect 18282 2204 18578 2224
rect 18338 2202 18362 2204
rect 18418 2202 18442 2204
rect 18498 2202 18522 2204
rect 18360 2150 18362 2202
rect 18424 2150 18436 2202
rect 18498 2150 18500 2202
rect 18338 2148 18362 2150
rect 18418 2148 18442 2150
rect 18498 2148 18522 2150
rect 18282 2128 18578 2148
rect 18156 1142 18276 1170
rect 18248 800 18276 1142
rect 18616 800 18644 2790
rect 18800 2553 18828 9318
rect 18892 6798 18920 10367
rect 18880 6792 18932 6798
rect 18880 6734 18932 6740
rect 18880 6656 18932 6662
rect 18880 6598 18932 6604
rect 18892 3602 18920 6598
rect 18880 3596 18932 3602
rect 18880 3538 18932 3544
rect 18786 2544 18842 2553
rect 18786 2479 18842 2488
rect 16946 640 17002 649
rect 16946 575 17002 584
rect 17314 0 17370 800
rect 17774 0 17830 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 18984 241 19012 11494
rect 19076 11354 19104 11766
rect 19064 11348 19116 11354
rect 19064 11290 19116 11296
rect 19076 10606 19104 11290
rect 19168 11286 19196 12854
rect 19248 12640 19300 12646
rect 19248 12582 19300 12588
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 19260 12374 19288 12582
rect 19248 12368 19300 12374
rect 19248 12310 19300 12316
rect 19248 12164 19300 12170
rect 19248 12106 19300 12112
rect 19260 11558 19288 12106
rect 19352 11762 19380 12582
rect 19444 12442 19472 13738
rect 19536 12714 19564 16594
rect 19524 12708 19576 12714
rect 19524 12650 19576 12656
rect 19432 12436 19484 12442
rect 19432 12378 19484 12384
rect 19340 11756 19392 11762
rect 19340 11698 19392 11704
rect 19248 11552 19300 11558
rect 19248 11494 19300 11500
rect 19156 11280 19208 11286
rect 19156 11222 19208 11228
rect 19156 11144 19208 11150
rect 19156 11086 19208 11092
rect 19064 10600 19116 10606
rect 19064 10542 19116 10548
rect 19168 10538 19196 11086
rect 19260 11082 19288 11494
rect 19536 11082 19564 12650
rect 19248 11076 19300 11082
rect 19248 11018 19300 11024
rect 19524 11076 19576 11082
rect 19524 11018 19576 11024
rect 19156 10532 19208 10538
rect 19156 10474 19208 10480
rect 19168 10266 19196 10474
rect 19156 10260 19208 10266
rect 19156 10202 19208 10208
rect 19062 10024 19118 10033
rect 19062 9959 19118 9968
rect 19076 8906 19104 9959
rect 19156 9104 19208 9110
rect 19156 9046 19208 9052
rect 19064 8900 19116 8906
rect 19064 8842 19116 8848
rect 19168 7721 19196 9046
rect 19154 7712 19210 7721
rect 19154 7647 19210 7656
rect 19260 7290 19288 11018
rect 19524 8560 19576 8566
rect 19524 8502 19576 8508
rect 19432 7948 19484 7954
rect 19432 7890 19484 7896
rect 19444 7410 19472 7890
rect 19432 7404 19484 7410
rect 19432 7346 19484 7352
rect 19076 7262 19288 7290
rect 19076 5778 19104 7262
rect 19156 7200 19208 7206
rect 19156 7142 19208 7148
rect 19246 7168 19302 7177
rect 19168 7002 19196 7142
rect 19246 7103 19302 7112
rect 19156 6996 19208 7002
rect 19156 6938 19208 6944
rect 19064 5772 19116 5778
rect 19064 5714 19116 5720
rect 19076 5574 19104 5714
rect 19156 5636 19208 5642
rect 19156 5578 19208 5584
rect 19064 5568 19116 5574
rect 19064 5510 19116 5516
rect 19076 3482 19104 5510
rect 19168 5234 19196 5578
rect 19156 5228 19208 5234
rect 19156 5170 19208 5176
rect 19260 4146 19288 7103
rect 19444 6254 19472 7346
rect 19340 6248 19392 6254
rect 19338 6216 19340 6225
rect 19432 6248 19484 6254
rect 19392 6216 19394 6225
rect 19432 6190 19484 6196
rect 19338 6151 19394 6160
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 19432 6112 19484 6118
rect 19432 6054 19484 6060
rect 19352 5914 19380 6054
rect 19340 5908 19392 5914
rect 19340 5850 19392 5856
rect 19444 5370 19472 6054
rect 19432 5364 19484 5370
rect 19432 5306 19484 5312
rect 19432 5024 19484 5030
rect 19432 4966 19484 4972
rect 19444 4758 19472 4966
rect 19432 4752 19484 4758
rect 19432 4694 19484 4700
rect 19340 4684 19392 4690
rect 19340 4626 19392 4632
rect 19352 4146 19380 4626
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 19340 4140 19392 4146
rect 19340 4082 19392 4088
rect 19260 3602 19288 4082
rect 19536 3618 19564 8502
rect 19628 8362 19656 17682
rect 19708 17332 19760 17338
rect 19708 17274 19760 17280
rect 19720 16658 19748 17274
rect 19708 16652 19760 16658
rect 19708 16594 19760 16600
rect 19708 15904 19760 15910
rect 19708 15846 19760 15852
rect 19720 15570 19748 15846
rect 19708 15564 19760 15570
rect 19708 15506 19760 15512
rect 19708 14476 19760 14482
rect 19708 14418 19760 14424
rect 19720 12850 19748 14418
rect 19708 12844 19760 12850
rect 19708 12786 19760 12792
rect 19708 12164 19760 12170
rect 19708 12106 19760 12112
rect 19720 11218 19748 12106
rect 19708 11212 19760 11218
rect 19708 11154 19760 11160
rect 19708 9920 19760 9926
rect 19708 9862 19760 9868
rect 19720 8430 19748 9862
rect 19812 9625 19840 18022
rect 19904 17882 19932 19314
rect 19892 17876 19944 17882
rect 19892 17818 19944 17824
rect 19892 17536 19944 17542
rect 19892 17478 19944 17484
rect 19904 17134 19932 17478
rect 19892 17128 19944 17134
rect 19892 17070 19944 17076
rect 19892 15360 19944 15366
rect 19892 15302 19944 15308
rect 19904 12102 19932 15302
rect 19996 13802 20024 20334
rect 20260 20256 20312 20262
rect 20260 20198 20312 20204
rect 20168 19916 20220 19922
rect 20168 19858 20220 19864
rect 20180 18902 20208 19858
rect 20272 19310 20300 20198
rect 20456 20058 20484 20703
rect 20640 20602 20668 22199
rect 20628 20596 20680 20602
rect 20628 20538 20680 20544
rect 21086 20360 21142 20369
rect 21086 20295 21142 20304
rect 20812 20256 20864 20262
rect 20812 20198 20864 20204
rect 20444 20052 20496 20058
rect 20444 19994 20496 20000
rect 20824 19922 20852 20198
rect 21100 20058 21128 20295
rect 21088 20052 21140 20058
rect 21088 19994 21140 20000
rect 20812 19916 20864 19922
rect 20812 19858 20864 19864
rect 20442 19816 20498 19825
rect 20442 19751 20498 19760
rect 20456 19514 20484 19751
rect 20444 19508 20496 19514
rect 20444 19450 20496 19456
rect 20260 19304 20312 19310
rect 20260 19246 20312 19252
rect 20168 18896 20220 18902
rect 20168 18838 20220 18844
rect 20076 18828 20128 18834
rect 20076 18770 20128 18776
rect 20088 17814 20116 18770
rect 20272 17898 20300 19246
rect 20352 18760 20404 18766
rect 20352 18702 20404 18708
rect 20180 17870 20300 17898
rect 20076 17808 20128 17814
rect 20076 17750 20128 17756
rect 20076 14816 20128 14822
rect 20076 14758 20128 14764
rect 20088 14482 20116 14758
rect 20076 14476 20128 14482
rect 20076 14418 20128 14424
rect 20180 14362 20208 17870
rect 20260 17740 20312 17746
rect 20260 17682 20312 17688
rect 20272 16114 20300 17682
rect 20260 16108 20312 16114
rect 20260 16050 20312 16056
rect 20260 14816 20312 14822
rect 20260 14758 20312 14764
rect 20088 14334 20208 14362
rect 19984 13796 20036 13802
rect 19984 13738 20036 13744
rect 19984 13320 20036 13326
rect 19984 13262 20036 13268
rect 19996 12850 20024 13262
rect 19984 12844 20036 12850
rect 19984 12786 20036 12792
rect 19996 12238 20024 12786
rect 19984 12232 20036 12238
rect 19984 12174 20036 12180
rect 19892 12096 19944 12102
rect 19892 12038 19944 12044
rect 19892 11756 19944 11762
rect 19892 11698 19944 11704
rect 19904 11150 19932 11698
rect 20088 11234 20116 14334
rect 20168 14272 20220 14278
rect 20168 14214 20220 14220
rect 19996 11206 20116 11234
rect 19892 11144 19944 11150
rect 19892 11086 19944 11092
rect 19798 9616 19854 9625
rect 19798 9551 19854 9560
rect 19800 8832 19852 8838
rect 19800 8774 19852 8780
rect 19812 8498 19840 8774
rect 19800 8492 19852 8498
rect 19800 8434 19852 8440
rect 19708 8424 19760 8430
rect 19708 8366 19760 8372
rect 19616 8356 19668 8362
rect 19616 8298 19668 8304
rect 19708 6860 19760 6866
rect 19708 6802 19760 6808
rect 19720 5846 19748 6802
rect 19904 6474 19932 11086
rect 19996 10810 20024 11206
rect 20076 11076 20128 11082
rect 20076 11018 20128 11024
rect 19984 10804 20036 10810
rect 19984 10746 20036 10752
rect 19984 9376 20036 9382
rect 19984 9318 20036 9324
rect 19996 8498 20024 9318
rect 20088 9110 20116 11018
rect 20076 9104 20128 9110
rect 20076 9046 20128 9052
rect 19984 8492 20036 8498
rect 19984 8434 20036 8440
rect 19996 8022 20024 8434
rect 19984 8016 20036 8022
rect 20180 7993 20208 14214
rect 20272 14074 20300 14758
rect 20260 14068 20312 14074
rect 20260 14010 20312 14016
rect 20260 13728 20312 13734
rect 20260 13670 20312 13676
rect 20272 13190 20300 13670
rect 20260 13184 20312 13190
rect 20260 13126 20312 13132
rect 20260 12844 20312 12850
rect 20260 12786 20312 12792
rect 20272 11626 20300 12786
rect 20260 11620 20312 11626
rect 20260 11562 20312 11568
rect 20260 11144 20312 11150
rect 20260 11086 20312 11092
rect 20272 10198 20300 11086
rect 20260 10192 20312 10198
rect 20260 10134 20312 10140
rect 19984 7958 20036 7964
rect 20166 7984 20222 7993
rect 20166 7919 20222 7928
rect 20168 7744 20220 7750
rect 20168 7686 20220 7692
rect 20180 7342 20208 7686
rect 20168 7336 20220 7342
rect 20168 7278 20220 7284
rect 20180 6798 20208 7278
rect 20260 7200 20312 7206
rect 20260 7142 20312 7148
rect 20168 6792 20220 6798
rect 20168 6734 20220 6740
rect 20272 6730 20300 7142
rect 20260 6724 20312 6730
rect 20260 6666 20312 6672
rect 19904 6446 20116 6474
rect 19892 6316 19944 6322
rect 19892 6258 19944 6264
rect 19798 6216 19854 6225
rect 19798 6151 19800 6160
rect 19852 6151 19854 6160
rect 19800 6122 19852 6128
rect 19708 5840 19760 5846
rect 19708 5782 19760 5788
rect 19904 4554 19932 6258
rect 19984 5772 20036 5778
rect 19984 5714 20036 5720
rect 19996 4826 20024 5714
rect 19984 4820 20036 4826
rect 19984 4762 20036 4768
rect 19892 4548 19944 4554
rect 19892 4490 19944 4496
rect 19904 4078 19932 4490
rect 19984 4480 20036 4486
rect 19984 4422 20036 4428
rect 19892 4072 19944 4078
rect 19892 4014 19944 4020
rect 19800 3732 19852 3738
rect 19800 3674 19852 3680
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 19444 3590 19564 3618
rect 19076 3454 19288 3482
rect 19064 3188 19116 3194
rect 19064 3130 19116 3136
rect 19076 2650 19104 3130
rect 19064 2644 19116 2650
rect 19064 2586 19116 2592
rect 19156 2304 19208 2310
rect 19156 2246 19208 2252
rect 19168 1170 19196 2246
rect 19076 1142 19196 1170
rect 19076 800 19104 1142
rect 19260 1057 19288 3454
rect 19444 3058 19472 3590
rect 19524 3528 19576 3534
rect 19524 3470 19576 3476
rect 19432 3052 19484 3058
rect 19432 2994 19484 3000
rect 19536 2990 19564 3470
rect 19616 3392 19668 3398
rect 19616 3334 19668 3340
rect 19524 2984 19576 2990
rect 19524 2926 19576 2932
rect 19246 1048 19302 1057
rect 19246 983 19302 992
rect 19628 898 19656 3334
rect 19812 2514 19840 3674
rect 19800 2508 19852 2514
rect 19800 2450 19852 2456
rect 19536 870 19656 898
rect 19536 800 19564 870
rect 19996 800 20024 4422
rect 20088 2009 20116 6446
rect 20272 6254 20300 6666
rect 20364 6458 20392 18702
rect 20442 18456 20498 18465
rect 20442 18391 20444 18400
rect 20496 18391 20498 18400
rect 20444 18362 20496 18368
rect 20536 18216 20588 18222
rect 20536 18158 20588 18164
rect 20442 16144 20498 16153
rect 20442 16079 20498 16088
rect 20456 15706 20484 16079
rect 20444 15700 20496 15706
rect 20444 15642 20496 15648
rect 20444 15564 20496 15570
rect 20444 15506 20496 15512
rect 20456 14278 20484 15506
rect 20548 15042 20576 18158
rect 20628 16992 20680 16998
rect 20628 16934 20680 16940
rect 20640 16561 20668 16934
rect 20720 16652 20772 16658
rect 20720 16594 20772 16600
rect 20626 16552 20682 16561
rect 20626 16487 20682 16496
rect 20732 16046 20760 16594
rect 20720 16040 20772 16046
rect 20720 15982 20772 15988
rect 20628 15904 20680 15910
rect 20824 15858 20852 19858
rect 20994 19408 21050 19417
rect 20994 19343 21050 19352
rect 21008 19174 21036 19343
rect 20996 19168 21048 19174
rect 20996 19110 21048 19116
rect 21088 18964 21140 18970
rect 21088 18906 21140 18912
rect 21100 18873 21128 18906
rect 21086 18864 21142 18873
rect 21086 18799 21142 18808
rect 20996 18080 21048 18086
rect 20994 18048 20996 18057
rect 21048 18048 21050 18057
rect 20994 17983 21050 17992
rect 21088 17536 21140 17542
rect 21088 17478 21140 17484
rect 21100 17105 21128 17478
rect 21086 17096 21142 17105
rect 20904 17060 20956 17066
rect 21086 17031 21142 17040
rect 20904 17002 20956 17008
rect 20916 16658 20944 17002
rect 21272 16788 21324 16794
rect 21272 16730 21324 16736
rect 20904 16652 20956 16658
rect 20904 16594 20956 16600
rect 20628 15846 20680 15852
rect 20640 15201 20668 15846
rect 20732 15830 20852 15858
rect 20626 15192 20682 15201
rect 20626 15127 20682 15136
rect 20548 15014 20668 15042
rect 20444 14272 20496 14278
rect 20444 14214 20496 14220
rect 20444 13796 20496 13802
rect 20444 13738 20496 13744
rect 20456 11150 20484 13738
rect 20536 12640 20588 12646
rect 20536 12582 20588 12588
rect 20444 11144 20496 11150
rect 20444 11086 20496 11092
rect 20442 10976 20498 10985
rect 20442 10911 20498 10920
rect 20456 7546 20484 10911
rect 20548 9178 20576 12582
rect 20640 11778 20668 15014
rect 20732 14550 20760 15830
rect 21088 15700 21140 15706
rect 21088 15642 21140 15648
rect 21100 15609 21128 15642
rect 21086 15600 21142 15609
rect 21086 15535 21142 15544
rect 20812 14952 20864 14958
rect 20812 14894 20864 14900
rect 20824 14550 20852 14894
rect 20996 14816 21048 14822
rect 20996 14758 21048 14764
rect 20720 14544 20772 14550
rect 20720 14486 20772 14492
rect 20812 14544 20864 14550
rect 20812 14486 20864 14492
rect 21008 14249 21036 14758
rect 21086 14648 21142 14657
rect 21086 14583 21142 14592
rect 20994 14240 21050 14249
rect 20994 14175 21050 14184
rect 21100 14074 21128 14583
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 20812 13864 20864 13870
rect 20812 13806 20864 13812
rect 21178 13832 21234 13841
rect 20824 13462 20852 13806
rect 21178 13767 21234 13776
rect 20812 13456 20864 13462
rect 20812 13398 20864 13404
rect 20720 13388 20772 13394
rect 20720 13330 20772 13336
rect 20732 12102 20760 13330
rect 21088 13320 21140 13326
rect 21088 13262 21140 13268
rect 20902 12880 20958 12889
rect 20902 12815 20958 12824
rect 20916 12646 20944 12815
rect 20996 12776 21048 12782
rect 20996 12718 21048 12724
rect 20904 12640 20956 12646
rect 20904 12582 20956 12588
rect 20720 12096 20772 12102
rect 20720 12038 20772 12044
rect 20732 11898 20852 11914
rect 20720 11892 20852 11898
rect 20772 11886 20852 11892
rect 20720 11834 20772 11840
rect 20640 11750 20760 11778
rect 20628 11620 20680 11626
rect 20628 11562 20680 11568
rect 20640 10810 20668 11562
rect 20628 10804 20680 10810
rect 20628 10746 20680 10752
rect 20732 10690 20760 11750
rect 20640 10662 20760 10690
rect 20536 9172 20588 9178
rect 20536 9114 20588 9120
rect 20534 9072 20590 9081
rect 20534 9007 20590 9016
rect 20444 7540 20496 7546
rect 20444 7482 20496 7488
rect 20456 6866 20484 7482
rect 20444 6860 20496 6866
rect 20444 6802 20496 6808
rect 20352 6452 20404 6458
rect 20352 6394 20404 6400
rect 20260 6248 20312 6254
rect 20260 6190 20312 6196
rect 20260 5704 20312 5710
rect 20260 5646 20312 5652
rect 20272 5234 20300 5646
rect 20260 5228 20312 5234
rect 20260 5170 20312 5176
rect 20444 5024 20496 5030
rect 20444 4966 20496 4972
rect 20074 2000 20130 2009
rect 20074 1935 20130 1944
rect 20456 800 20484 4966
rect 20548 3738 20576 9007
rect 20640 5914 20668 10662
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 20732 9518 20760 9998
rect 20720 9512 20772 9518
rect 20720 9454 20772 9460
rect 20732 8974 20760 9454
rect 20720 8968 20772 8974
rect 20720 8910 20772 8916
rect 20628 5908 20680 5914
rect 20628 5850 20680 5856
rect 20626 5264 20682 5273
rect 20626 5199 20682 5208
rect 20640 4690 20668 5199
rect 20628 4684 20680 4690
rect 20628 4626 20680 4632
rect 20640 4282 20668 4626
rect 20628 4276 20680 4282
rect 20628 4218 20680 4224
rect 20720 4004 20772 4010
rect 20720 3946 20772 3952
rect 20626 3904 20682 3913
rect 20626 3839 20682 3848
rect 20536 3732 20588 3738
rect 20536 3674 20588 3680
rect 20640 2514 20668 3839
rect 20732 2990 20760 3946
rect 20824 3058 20852 11886
rect 20916 11354 20944 12582
rect 21008 12345 21036 12718
rect 20994 12336 21050 12345
rect 21100 12306 21128 13262
rect 21192 12442 21220 13767
rect 21284 13297 21312 16730
rect 21270 13288 21326 13297
rect 21270 13223 21326 13232
rect 21180 12436 21232 12442
rect 21180 12378 21232 12384
rect 20994 12271 21050 12280
rect 21088 12300 21140 12306
rect 21088 12242 21140 12248
rect 20996 12096 21048 12102
rect 20996 12038 21048 12044
rect 21008 11694 21036 12038
rect 20996 11688 21048 11694
rect 20996 11630 21048 11636
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 20904 11348 20956 11354
rect 20904 11290 20956 11296
rect 20904 10124 20956 10130
rect 20904 10066 20956 10072
rect 20916 9178 20944 10066
rect 21376 10062 21404 11494
rect 21364 10056 21416 10062
rect 21364 9998 21416 10004
rect 20904 9172 20956 9178
rect 20904 9114 20956 9120
rect 21180 9104 21232 9110
rect 21180 9046 21232 9052
rect 20812 3052 20864 3058
rect 20812 2994 20864 3000
rect 20720 2984 20772 2990
rect 20720 2926 20772 2932
rect 20628 2508 20680 2514
rect 20628 2450 20680 2456
rect 20904 2304 20956 2310
rect 20904 2246 20956 2252
rect 20916 800 20944 2246
rect 21192 1601 21220 9046
rect 21364 6112 21416 6118
rect 21364 6054 21416 6060
rect 21376 5681 21404 6054
rect 21362 5672 21418 5681
rect 21362 5607 21418 5616
rect 21272 5568 21324 5574
rect 21272 5510 21324 5516
rect 21284 5166 21312 5510
rect 21272 5160 21324 5166
rect 21272 5102 21324 5108
rect 21284 4457 21312 5102
rect 21270 4448 21326 4457
rect 21270 4383 21326 4392
rect 21824 3936 21876 3942
rect 21824 3878 21876 3884
rect 21836 3602 21864 3878
rect 21824 3596 21876 3602
rect 21824 3538 21876 3544
rect 21364 2372 21416 2378
rect 21364 2314 21416 2320
rect 21178 1592 21234 1601
rect 21178 1527 21234 1536
rect 21376 800 21404 2314
rect 21836 800 21864 3538
rect 22284 3392 22336 3398
rect 22284 3334 22336 3340
rect 22296 800 22324 3334
rect 22744 2984 22796 2990
rect 22744 2926 22796 2932
rect 22756 800 22784 2926
rect 18970 232 19026 241
rect 18970 167 19026 176
rect 19062 0 19118 800
rect 19522 0 19578 800
rect 19982 0 20038 800
rect 20442 0 20498 800
rect 20902 0 20958 800
rect 21362 0 21418 800
rect 21822 0 21878 800
rect 22282 0 22338 800
rect 22742 0 22798 800
<< via2 >>
rect 3330 22616 3386 22672
rect 2870 22208 2926 22264
rect 2778 21664 2834 21720
rect 1950 21256 2006 21312
rect 3054 20712 3110 20768
rect 2962 20304 3018 20360
rect 1950 19760 2006 19816
rect 2778 19352 2834 19408
rect 1950 18808 2006 18864
rect 1950 18420 2006 18456
rect 1950 18400 1952 18420
rect 1952 18400 2004 18420
rect 2004 18400 2006 18420
rect 1674 17992 1730 18048
rect 1950 17040 2006 17096
rect 1674 16124 1676 16144
rect 1676 16124 1728 16144
rect 1728 16124 1730 16144
rect 1674 16088 1730 16124
rect 1950 15544 2006 15600
rect 1858 15136 1914 15192
rect 1858 14592 1914 14648
rect 1950 14184 2006 14240
rect 2778 17448 2834 17504
rect 18694 22616 18750 22672
rect 4421 20698 4477 20700
rect 4501 20698 4557 20700
rect 4581 20698 4637 20700
rect 4661 20698 4717 20700
rect 4421 20646 4447 20698
rect 4447 20646 4477 20698
rect 4501 20646 4511 20698
rect 4511 20646 4557 20698
rect 4581 20646 4627 20698
rect 4627 20646 4637 20698
rect 4661 20646 4691 20698
rect 4691 20646 4717 20698
rect 4421 20644 4477 20646
rect 4501 20644 4557 20646
rect 4581 20644 4637 20646
rect 4661 20644 4717 20646
rect 2502 16516 2558 16552
rect 2502 16496 2504 16516
rect 2504 16496 2556 16516
rect 2556 16496 2558 16516
rect 2134 12144 2190 12200
rect 2870 13776 2926 13832
rect 2778 13232 2834 13288
rect 4421 19610 4477 19612
rect 4501 19610 4557 19612
rect 4581 19610 4637 19612
rect 4661 19610 4717 19612
rect 4421 19558 4447 19610
rect 4447 19558 4477 19610
rect 4501 19558 4511 19610
rect 4511 19558 4557 19610
rect 4581 19558 4627 19610
rect 4627 19558 4637 19610
rect 4661 19558 4691 19610
rect 4691 19558 4717 19610
rect 4421 19556 4477 19558
rect 4501 19556 4557 19558
rect 4581 19556 4637 19558
rect 4661 19556 4717 19558
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11378 20698
rect 11378 20646 11408 20698
rect 11432 20646 11442 20698
rect 11442 20646 11488 20698
rect 11512 20646 11558 20698
rect 11558 20646 11568 20698
rect 11592 20646 11622 20698
rect 11622 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 4421 18522 4477 18524
rect 4501 18522 4557 18524
rect 4581 18522 4637 18524
rect 4661 18522 4717 18524
rect 4421 18470 4447 18522
rect 4447 18470 4477 18522
rect 4501 18470 4511 18522
rect 4511 18470 4557 18522
rect 4581 18470 4627 18522
rect 4627 18470 4637 18522
rect 4661 18470 4691 18522
rect 4691 18470 4717 18522
rect 4421 18468 4477 18470
rect 4501 18468 4557 18470
rect 4581 18468 4637 18470
rect 4661 18468 4717 18470
rect 4421 17434 4477 17436
rect 4501 17434 4557 17436
rect 4581 17434 4637 17436
rect 4661 17434 4717 17436
rect 4421 17382 4447 17434
rect 4447 17382 4477 17434
rect 4501 17382 4511 17434
rect 4511 17382 4557 17434
rect 4581 17382 4627 17434
rect 4627 17382 4637 17434
rect 4661 17382 4691 17434
rect 4691 17382 4717 17434
rect 4421 17380 4477 17382
rect 4501 17380 4557 17382
rect 4581 17380 4637 17382
rect 4661 17380 4717 17382
rect 2042 9152 2098 9208
rect 1398 7148 1400 7168
rect 1400 7148 1452 7168
rect 1452 7148 1454 7168
rect 1398 7112 1454 7148
rect 1950 3596 2006 3632
rect 1950 3576 1952 3596
rect 1952 3576 2004 3596
rect 2004 3576 2006 3596
rect 2042 3440 2098 3496
rect 1674 2488 1730 2544
rect 1306 1536 1362 1592
rect 3054 8200 3110 8256
rect 4421 16346 4477 16348
rect 4501 16346 4557 16348
rect 4581 16346 4637 16348
rect 4661 16346 4717 16348
rect 4421 16294 4447 16346
rect 4447 16294 4477 16346
rect 4501 16294 4511 16346
rect 4511 16294 4557 16346
rect 4581 16294 4627 16346
rect 4627 16294 4637 16346
rect 4661 16294 4691 16346
rect 4691 16294 4717 16346
rect 4421 16292 4477 16294
rect 4501 16292 4557 16294
rect 4581 16292 4637 16294
rect 4661 16292 4717 16294
rect 3146 6296 3202 6352
rect 4421 15258 4477 15260
rect 4501 15258 4557 15260
rect 4581 15258 4637 15260
rect 4661 15258 4717 15260
rect 4421 15206 4447 15258
rect 4447 15206 4477 15258
rect 4501 15206 4511 15258
rect 4511 15206 4557 15258
rect 4581 15206 4627 15258
rect 4627 15206 4637 15258
rect 4661 15206 4691 15258
rect 4691 15206 4717 15258
rect 4421 15204 4477 15206
rect 4501 15204 4557 15206
rect 4581 15204 4637 15206
rect 4661 15204 4717 15206
rect 4421 14170 4477 14172
rect 4501 14170 4557 14172
rect 4581 14170 4637 14172
rect 4661 14170 4717 14172
rect 4421 14118 4447 14170
rect 4447 14118 4477 14170
rect 4501 14118 4511 14170
rect 4511 14118 4557 14170
rect 4581 14118 4627 14170
rect 4627 14118 4637 14170
rect 4661 14118 4691 14170
rect 4691 14118 4717 14170
rect 4421 14116 4477 14118
rect 4501 14116 4557 14118
rect 4581 14116 4637 14118
rect 4661 14116 4717 14118
rect 4421 13082 4477 13084
rect 4501 13082 4557 13084
rect 4581 13082 4637 13084
rect 4661 13082 4717 13084
rect 4421 13030 4447 13082
rect 4447 13030 4477 13082
rect 4501 13030 4511 13082
rect 4511 13030 4557 13082
rect 4581 13030 4627 13082
rect 4627 13030 4637 13082
rect 4661 13030 4691 13082
rect 4691 13030 4717 13082
rect 4421 13028 4477 13030
rect 4501 13028 4557 13030
rect 4581 13028 4637 13030
rect 4661 13028 4717 13030
rect 4066 12824 4122 12880
rect 3882 12280 3938 12336
rect 4066 11872 4122 11928
rect 4421 11994 4477 11996
rect 4501 11994 4557 11996
rect 4581 11994 4637 11996
rect 4661 11994 4717 11996
rect 4421 11942 4447 11994
rect 4447 11942 4477 11994
rect 4501 11942 4511 11994
rect 4511 11942 4557 11994
rect 4581 11942 4627 11994
rect 4627 11942 4637 11994
rect 4661 11942 4691 11994
rect 4691 11942 4717 11994
rect 4421 11940 4477 11942
rect 4501 11940 4557 11942
rect 4581 11940 4637 11942
rect 4661 11940 4717 11942
rect 4066 10920 4122 10976
rect 4421 10906 4477 10908
rect 4501 10906 4557 10908
rect 4581 10906 4637 10908
rect 4661 10906 4717 10908
rect 4421 10854 4447 10906
rect 4447 10854 4477 10906
rect 4501 10854 4511 10906
rect 4511 10854 4557 10906
rect 4581 10854 4627 10906
rect 4627 10854 4637 10906
rect 4661 10854 4691 10906
rect 4691 10854 4717 10906
rect 4421 10852 4477 10854
rect 4501 10852 4557 10854
rect 4581 10852 4637 10854
rect 4661 10852 4717 10854
rect 4066 10376 4122 10432
rect 4066 9968 4122 10024
rect 4066 9016 4122 9072
rect 4421 9818 4477 9820
rect 4501 9818 4557 9820
rect 4581 9818 4637 9820
rect 4661 9818 4717 9820
rect 4421 9766 4447 9818
rect 4447 9766 4477 9818
rect 4501 9766 4511 9818
rect 4511 9766 4557 9818
rect 4581 9766 4627 9818
rect 4627 9766 4637 9818
rect 4661 9766 4691 9818
rect 4691 9766 4717 9818
rect 4421 9764 4477 9766
rect 4501 9764 4557 9766
rect 4581 9764 4637 9766
rect 4661 9764 4717 9766
rect 4250 9560 4306 9616
rect 4421 8730 4477 8732
rect 4501 8730 4557 8732
rect 4581 8730 4637 8732
rect 4661 8730 4717 8732
rect 4421 8678 4447 8730
rect 4447 8678 4477 8730
rect 4501 8678 4511 8730
rect 4511 8678 4557 8730
rect 4581 8678 4627 8730
rect 4627 8678 4637 8730
rect 4661 8678 4691 8730
rect 4691 8678 4717 8730
rect 4421 8676 4477 8678
rect 4501 8676 4557 8678
rect 4581 8676 4637 8678
rect 4661 8676 4717 8678
rect 4250 8608 4306 8664
rect 4066 8064 4122 8120
rect 3974 7656 4030 7712
rect 4421 7642 4477 7644
rect 4501 7642 4557 7644
rect 4581 7642 4637 7644
rect 4661 7642 4717 7644
rect 4421 7590 4447 7642
rect 4447 7590 4477 7642
rect 4501 7590 4511 7642
rect 4511 7590 4557 7642
rect 4581 7590 4627 7642
rect 4627 7590 4637 7642
rect 4661 7590 4691 7642
rect 4691 7590 4717 7642
rect 4421 7588 4477 7590
rect 4501 7588 4557 7590
rect 4581 7588 4637 7590
rect 4661 7588 4717 7590
rect 5078 9424 5134 9480
rect 3974 6704 4030 6760
rect 4158 6160 4214 6216
rect 3882 5752 3938 5808
rect 3974 5208 4030 5264
rect 3882 4800 3938 4856
rect 4066 4392 4122 4448
rect 3882 3848 3938 3904
rect 3698 2896 3754 2952
rect 3606 1944 3662 2000
rect 4158 3576 4214 3632
rect 3974 992 4030 1048
rect 4421 6554 4477 6556
rect 4501 6554 4557 6556
rect 4581 6554 4637 6556
rect 4661 6554 4717 6556
rect 4421 6502 4447 6554
rect 4447 6502 4477 6554
rect 4501 6502 4511 6554
rect 4511 6502 4557 6554
rect 4581 6502 4627 6554
rect 4627 6502 4637 6554
rect 4661 6502 4691 6554
rect 4691 6502 4717 6554
rect 4421 6500 4477 6502
rect 4501 6500 4557 6502
rect 4581 6500 4637 6502
rect 4661 6500 4717 6502
rect 5170 6024 5226 6080
rect 4421 5466 4477 5468
rect 4501 5466 4557 5468
rect 4581 5466 4637 5468
rect 4661 5466 4717 5468
rect 4421 5414 4447 5466
rect 4447 5414 4477 5466
rect 4501 5414 4511 5466
rect 4511 5414 4557 5466
rect 4581 5414 4627 5466
rect 4627 5414 4637 5466
rect 4661 5414 4691 5466
rect 4691 5414 4717 5466
rect 4421 5412 4477 5414
rect 4501 5412 4557 5414
rect 4581 5412 4637 5414
rect 4661 5412 4717 5414
rect 5538 11328 5594 11384
rect 5538 8200 5594 8256
rect 4421 4378 4477 4380
rect 4501 4378 4557 4380
rect 4581 4378 4637 4380
rect 4661 4378 4717 4380
rect 4421 4326 4447 4378
rect 4447 4326 4477 4378
rect 4501 4326 4511 4378
rect 4511 4326 4557 4378
rect 4581 4326 4627 4378
rect 4627 4326 4637 4378
rect 4661 4326 4691 4378
rect 4691 4326 4717 4378
rect 4421 4324 4477 4326
rect 4501 4324 4557 4326
rect 4581 4324 4637 4326
rect 4661 4324 4717 4326
rect 4421 3290 4477 3292
rect 4501 3290 4557 3292
rect 4581 3290 4637 3292
rect 4661 3290 4717 3292
rect 4421 3238 4447 3290
rect 4447 3238 4477 3290
rect 4501 3238 4511 3290
rect 4511 3238 4557 3290
rect 4581 3238 4627 3290
rect 4627 3238 4637 3290
rect 4661 3238 4691 3290
rect 4691 3238 4717 3290
rect 4421 3236 4477 3238
rect 4501 3236 4557 3238
rect 4581 3236 4637 3238
rect 4661 3236 4717 3238
rect 4421 2202 4477 2204
rect 4501 2202 4557 2204
rect 4581 2202 4637 2204
rect 4661 2202 4717 2204
rect 4421 2150 4447 2202
rect 4447 2150 4477 2202
rect 4501 2150 4511 2202
rect 4511 2150 4557 2202
rect 4581 2150 4627 2202
rect 4627 2150 4637 2202
rect 4661 2150 4691 2202
rect 4691 2150 4717 2202
rect 4421 2148 4477 2150
rect 4501 2148 4557 2150
rect 4581 2148 4637 2150
rect 4661 2148 4717 2150
rect 6550 9152 6606 9208
rect 2318 584 2374 640
rect 7886 20154 7942 20156
rect 7966 20154 8022 20156
rect 8046 20154 8102 20156
rect 8126 20154 8182 20156
rect 7886 20102 7912 20154
rect 7912 20102 7942 20154
rect 7966 20102 7976 20154
rect 7976 20102 8022 20154
rect 8046 20102 8092 20154
rect 8092 20102 8102 20154
rect 8126 20102 8156 20154
rect 8156 20102 8182 20154
rect 7886 20100 7942 20102
rect 7966 20100 8022 20102
rect 8046 20100 8102 20102
rect 8126 20100 8182 20102
rect 7886 19066 7942 19068
rect 7966 19066 8022 19068
rect 8046 19066 8102 19068
rect 8126 19066 8182 19068
rect 7886 19014 7912 19066
rect 7912 19014 7942 19066
rect 7966 19014 7976 19066
rect 7976 19014 8022 19066
rect 8046 19014 8092 19066
rect 8092 19014 8102 19066
rect 8126 19014 8156 19066
rect 8156 19014 8182 19066
rect 7886 19012 7942 19014
rect 7966 19012 8022 19014
rect 8046 19012 8102 19014
rect 8126 19012 8182 19014
rect 7886 17978 7942 17980
rect 7966 17978 8022 17980
rect 8046 17978 8102 17980
rect 8126 17978 8182 17980
rect 7886 17926 7912 17978
rect 7912 17926 7942 17978
rect 7966 17926 7976 17978
rect 7976 17926 8022 17978
rect 8046 17926 8092 17978
rect 8092 17926 8102 17978
rect 8126 17926 8156 17978
rect 8156 17926 8182 17978
rect 7886 17924 7942 17926
rect 7966 17924 8022 17926
rect 8046 17924 8102 17926
rect 8126 17924 8182 17926
rect 7886 16890 7942 16892
rect 7966 16890 8022 16892
rect 8046 16890 8102 16892
rect 8126 16890 8182 16892
rect 7886 16838 7912 16890
rect 7912 16838 7942 16890
rect 7966 16838 7976 16890
rect 7976 16838 8022 16890
rect 8046 16838 8092 16890
rect 8092 16838 8102 16890
rect 8126 16838 8156 16890
rect 8156 16838 8182 16890
rect 7886 16836 7942 16838
rect 7966 16836 8022 16838
rect 8046 16836 8102 16838
rect 8126 16836 8182 16838
rect 7886 15802 7942 15804
rect 7966 15802 8022 15804
rect 8046 15802 8102 15804
rect 8126 15802 8182 15804
rect 7886 15750 7912 15802
rect 7912 15750 7942 15802
rect 7966 15750 7976 15802
rect 7976 15750 8022 15802
rect 8046 15750 8092 15802
rect 8092 15750 8102 15802
rect 8126 15750 8156 15802
rect 8156 15750 8182 15802
rect 7886 15748 7942 15750
rect 7966 15748 8022 15750
rect 8046 15748 8102 15750
rect 8126 15748 8182 15750
rect 7886 14714 7942 14716
rect 7966 14714 8022 14716
rect 8046 14714 8102 14716
rect 8126 14714 8182 14716
rect 7886 14662 7912 14714
rect 7912 14662 7942 14714
rect 7966 14662 7976 14714
rect 7976 14662 8022 14714
rect 8046 14662 8092 14714
rect 8092 14662 8102 14714
rect 8126 14662 8156 14714
rect 8156 14662 8182 14714
rect 7886 14660 7942 14662
rect 7966 14660 8022 14662
rect 8046 14660 8102 14662
rect 8126 14660 8182 14662
rect 7886 13626 7942 13628
rect 7966 13626 8022 13628
rect 8046 13626 8102 13628
rect 8126 13626 8182 13628
rect 7886 13574 7912 13626
rect 7912 13574 7942 13626
rect 7966 13574 7976 13626
rect 7976 13574 8022 13626
rect 8046 13574 8092 13626
rect 8092 13574 8102 13626
rect 8126 13574 8156 13626
rect 8156 13574 8182 13626
rect 7886 13572 7942 13574
rect 7966 13572 8022 13574
rect 8046 13572 8102 13574
rect 8126 13572 8182 13574
rect 7886 12538 7942 12540
rect 7966 12538 8022 12540
rect 8046 12538 8102 12540
rect 8126 12538 8182 12540
rect 7886 12486 7912 12538
rect 7912 12486 7942 12538
rect 7966 12486 7976 12538
rect 7976 12486 8022 12538
rect 8046 12486 8092 12538
rect 8092 12486 8102 12538
rect 8126 12486 8156 12538
rect 8156 12486 8182 12538
rect 7886 12484 7942 12486
rect 7966 12484 8022 12486
rect 8046 12484 8102 12486
rect 8126 12484 8182 12486
rect 7886 11450 7942 11452
rect 7966 11450 8022 11452
rect 8046 11450 8102 11452
rect 8126 11450 8182 11452
rect 7886 11398 7912 11450
rect 7912 11398 7942 11450
rect 7966 11398 7976 11450
rect 7976 11398 8022 11450
rect 8046 11398 8092 11450
rect 8092 11398 8102 11450
rect 8126 11398 8156 11450
rect 8156 11398 8182 11450
rect 7886 11396 7942 11398
rect 7966 11396 8022 11398
rect 8046 11396 8102 11398
rect 8126 11396 8182 11398
rect 7470 5752 7526 5808
rect 7886 10362 7942 10364
rect 7966 10362 8022 10364
rect 8046 10362 8102 10364
rect 8126 10362 8182 10364
rect 7886 10310 7912 10362
rect 7912 10310 7942 10362
rect 7966 10310 7976 10362
rect 7976 10310 8022 10362
rect 8046 10310 8092 10362
rect 8092 10310 8102 10362
rect 8126 10310 8156 10362
rect 8156 10310 8182 10362
rect 7886 10308 7942 10310
rect 7966 10308 8022 10310
rect 8046 10308 8102 10310
rect 8126 10308 8182 10310
rect 7886 9274 7942 9276
rect 7966 9274 8022 9276
rect 8046 9274 8102 9276
rect 8126 9274 8182 9276
rect 7886 9222 7912 9274
rect 7912 9222 7942 9274
rect 7966 9222 7976 9274
rect 7976 9222 8022 9274
rect 8046 9222 8092 9274
rect 8092 9222 8102 9274
rect 8126 9222 8156 9274
rect 8156 9222 8182 9274
rect 7886 9220 7942 9222
rect 7966 9220 8022 9222
rect 8046 9220 8102 9222
rect 8126 9220 8182 9222
rect 7886 8186 7942 8188
rect 7966 8186 8022 8188
rect 8046 8186 8102 8188
rect 8126 8186 8182 8188
rect 7886 8134 7912 8186
rect 7912 8134 7942 8186
rect 7966 8134 7976 8186
rect 7976 8134 8022 8186
rect 8046 8134 8092 8186
rect 8092 8134 8102 8186
rect 8126 8134 8156 8186
rect 8156 8134 8182 8186
rect 7886 8132 7942 8134
rect 7966 8132 8022 8134
rect 8046 8132 8102 8134
rect 8126 8132 8182 8134
rect 7886 7098 7942 7100
rect 7966 7098 8022 7100
rect 8046 7098 8102 7100
rect 8126 7098 8182 7100
rect 7886 7046 7912 7098
rect 7912 7046 7942 7098
rect 7966 7046 7976 7098
rect 7976 7046 8022 7098
rect 8046 7046 8092 7098
rect 8092 7046 8102 7098
rect 8126 7046 8156 7098
rect 8156 7046 8182 7098
rect 7886 7044 7942 7046
rect 7966 7044 8022 7046
rect 8046 7044 8102 7046
rect 8126 7044 8182 7046
rect 8114 6704 8170 6760
rect 7886 6010 7942 6012
rect 7966 6010 8022 6012
rect 8046 6010 8102 6012
rect 8126 6010 8182 6012
rect 7886 5958 7912 6010
rect 7912 5958 7942 6010
rect 7966 5958 7976 6010
rect 7976 5958 8022 6010
rect 8046 5958 8092 6010
rect 8092 5958 8102 6010
rect 8126 5958 8156 6010
rect 8156 5958 8182 6010
rect 7886 5956 7942 5958
rect 7966 5956 8022 5958
rect 8046 5956 8102 5958
rect 8126 5956 8182 5958
rect 7886 4922 7942 4924
rect 7966 4922 8022 4924
rect 8046 4922 8102 4924
rect 8126 4922 8182 4924
rect 7886 4870 7912 4922
rect 7912 4870 7942 4922
rect 7966 4870 7976 4922
rect 7976 4870 8022 4922
rect 8046 4870 8092 4922
rect 8092 4870 8102 4922
rect 8126 4870 8156 4922
rect 8156 4870 8182 4922
rect 7886 4868 7942 4870
rect 7966 4868 8022 4870
rect 8046 4868 8102 4870
rect 8126 4868 8182 4870
rect 7886 3834 7942 3836
rect 7966 3834 8022 3836
rect 8046 3834 8102 3836
rect 8126 3834 8182 3836
rect 7886 3782 7912 3834
rect 7912 3782 7942 3834
rect 7966 3782 7976 3834
rect 7976 3782 8022 3834
rect 8046 3782 8092 3834
rect 8092 3782 8102 3834
rect 8126 3782 8156 3834
rect 8156 3782 8182 3834
rect 7886 3780 7942 3782
rect 7966 3780 8022 3782
rect 8046 3780 8102 3782
rect 8126 3780 8182 3782
rect 7886 2746 7942 2748
rect 7966 2746 8022 2748
rect 8046 2746 8102 2748
rect 8126 2746 8182 2748
rect 7886 2694 7912 2746
rect 7912 2694 7942 2746
rect 7966 2694 7976 2746
rect 7976 2694 8022 2746
rect 8046 2694 8092 2746
rect 8092 2694 8102 2746
rect 8126 2694 8156 2746
rect 8156 2694 8182 2746
rect 7886 2692 7942 2694
rect 7966 2692 8022 2694
rect 8046 2692 8102 2694
rect 8126 2692 8182 2694
rect 9954 16496 10010 16552
rect 9494 12144 9550 12200
rect 14817 20154 14873 20156
rect 14897 20154 14953 20156
rect 14977 20154 15033 20156
rect 15057 20154 15113 20156
rect 14817 20102 14843 20154
rect 14843 20102 14873 20154
rect 14897 20102 14907 20154
rect 14907 20102 14953 20154
rect 14977 20102 15023 20154
rect 15023 20102 15033 20154
rect 15057 20102 15087 20154
rect 15087 20102 15113 20154
rect 14817 20100 14873 20102
rect 14897 20100 14953 20102
rect 14977 20100 15033 20102
rect 15057 20100 15113 20102
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11378 19610
rect 11378 19558 11408 19610
rect 11432 19558 11442 19610
rect 11442 19558 11488 19610
rect 11512 19558 11558 19610
rect 11558 19558 11568 19610
rect 11592 19558 11622 19610
rect 11622 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11378 18522
rect 11378 18470 11408 18522
rect 11432 18470 11442 18522
rect 11442 18470 11488 18522
rect 11512 18470 11558 18522
rect 11558 18470 11568 18522
rect 11592 18470 11622 18522
rect 11622 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 9310 5652 9312 5672
rect 9312 5652 9364 5672
rect 9364 5652 9366 5672
rect 9310 5616 9366 5652
rect 10046 8880 10102 8936
rect 10322 6860 10378 6896
rect 10322 6840 10324 6860
rect 10324 6840 10376 6860
rect 10376 6840 10378 6860
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11378 17434
rect 11378 17382 11408 17434
rect 11432 17382 11442 17434
rect 11442 17382 11488 17434
rect 11512 17382 11558 17434
rect 11558 17382 11568 17434
rect 11592 17382 11622 17434
rect 11622 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11378 16346
rect 11378 16294 11408 16346
rect 11432 16294 11442 16346
rect 11442 16294 11488 16346
rect 11512 16294 11558 16346
rect 11558 16294 11568 16346
rect 11592 16294 11622 16346
rect 11622 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 10690 9560 10746 9616
rect 10598 7928 10654 7984
rect 10782 7384 10838 7440
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11378 15258
rect 11378 15206 11408 15258
rect 11432 15206 11442 15258
rect 11442 15206 11488 15258
rect 11512 15206 11558 15258
rect 11558 15206 11568 15258
rect 11592 15206 11622 15258
rect 11622 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11378 14170
rect 11378 14118 11408 14170
rect 11432 14118 11442 14170
rect 11442 14118 11488 14170
rect 11512 14118 11558 14170
rect 11558 14118 11568 14170
rect 11592 14118 11622 14170
rect 11622 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 12254 17620 12256 17640
rect 12256 17620 12308 17640
rect 12308 17620 12310 17640
rect 12254 17584 12310 17620
rect 13266 17740 13322 17776
rect 13266 17720 13268 17740
rect 13268 17720 13320 17740
rect 13320 17720 13322 17740
rect 12990 16516 13046 16552
rect 12990 16496 12992 16516
rect 12992 16496 13044 16516
rect 13044 16496 13046 16516
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11378 13082
rect 11378 13030 11408 13082
rect 11432 13030 11442 13082
rect 11442 13030 11488 13082
rect 11512 13030 11558 13082
rect 11558 13030 11568 13082
rect 11592 13030 11622 13082
rect 11622 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11378 11994
rect 11378 11942 11408 11994
rect 11432 11942 11442 11994
rect 11442 11942 11488 11994
rect 11512 11942 11558 11994
rect 11558 11942 11568 11994
rect 11592 11942 11622 11994
rect 11622 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11378 10906
rect 11378 10854 11408 10906
rect 11432 10854 11442 10906
rect 11442 10854 11488 10906
rect 11512 10854 11558 10906
rect 11558 10854 11568 10906
rect 11592 10854 11622 10906
rect 11622 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11378 9818
rect 11378 9766 11408 9818
rect 11432 9766 11442 9818
rect 11442 9766 11488 9818
rect 11512 9766 11558 9818
rect 11558 9766 11568 9818
rect 11592 9766 11622 9818
rect 11622 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11886 11328 11942 11384
rect 11702 8880 11758 8936
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11378 8730
rect 11378 8678 11408 8730
rect 11432 8678 11442 8730
rect 11442 8678 11488 8730
rect 11512 8678 11558 8730
rect 11558 8678 11568 8730
rect 11592 8678 11622 8730
rect 11622 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11378 7642
rect 11378 7590 11408 7642
rect 11432 7590 11442 7642
rect 11442 7590 11488 7642
rect 11512 7590 11558 7642
rect 11558 7590 11568 7642
rect 11592 7590 11622 7642
rect 11622 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11794 6704 11850 6760
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11378 6554
rect 11378 6502 11408 6554
rect 11432 6502 11442 6554
rect 11442 6502 11488 6554
rect 11512 6502 11558 6554
rect 11558 6502 11568 6554
rect 11592 6502 11622 6554
rect 11622 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11378 5466
rect 11378 5414 11408 5466
rect 11432 5414 11442 5466
rect 11442 5414 11488 5466
rect 11512 5414 11558 5466
rect 11558 5414 11568 5466
rect 11592 5414 11622 5466
rect 11622 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11378 4378
rect 11378 4326 11408 4378
rect 11432 4326 11442 4378
rect 11442 4326 11488 4378
rect 11512 4326 11558 4378
rect 11558 4326 11568 4378
rect 11592 4326 11622 4378
rect 11622 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11378 3290
rect 11378 3238 11408 3290
rect 11432 3238 11442 3290
rect 11442 3238 11488 3290
rect 11512 3238 11558 3290
rect 11558 3238 11568 3290
rect 11592 3238 11622 3290
rect 11622 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 12070 8472 12126 8528
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11378 2202
rect 11378 2150 11408 2202
rect 11432 2150 11442 2202
rect 11442 2150 11488 2202
rect 11512 2150 11558 2202
rect 11558 2150 11568 2202
rect 11592 2150 11622 2202
rect 11622 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 13726 17740 13782 17776
rect 13726 17720 13728 17740
rect 13728 17720 13780 17740
rect 13780 17720 13782 17740
rect 14817 19066 14873 19068
rect 14897 19066 14953 19068
rect 14977 19066 15033 19068
rect 15057 19066 15113 19068
rect 14817 19014 14843 19066
rect 14843 19014 14873 19066
rect 14897 19014 14907 19066
rect 14907 19014 14953 19066
rect 14977 19014 15023 19066
rect 15023 19014 15033 19066
rect 15057 19014 15087 19066
rect 15087 19014 15113 19066
rect 14817 19012 14873 19014
rect 14897 19012 14953 19014
rect 14977 19012 15033 19014
rect 15057 19012 15113 19014
rect 13082 11328 13138 11384
rect 12530 5788 12532 5808
rect 12532 5788 12584 5808
rect 12584 5788 12586 5808
rect 12530 5752 12586 5788
rect 14186 8336 14242 8392
rect 14817 17978 14873 17980
rect 14897 17978 14953 17980
rect 14977 17978 15033 17980
rect 15057 17978 15113 17980
rect 14817 17926 14843 17978
rect 14843 17926 14873 17978
rect 14897 17926 14907 17978
rect 14907 17926 14953 17978
rect 14977 17926 15023 17978
rect 15023 17926 15033 17978
rect 15057 17926 15087 17978
rect 15087 17926 15113 17978
rect 14817 17924 14873 17926
rect 14897 17924 14953 17926
rect 14977 17924 15033 17926
rect 15057 17924 15113 17926
rect 14817 16890 14873 16892
rect 14897 16890 14953 16892
rect 14977 16890 15033 16892
rect 15057 16890 15113 16892
rect 14817 16838 14843 16890
rect 14843 16838 14873 16890
rect 14897 16838 14907 16890
rect 14907 16838 14953 16890
rect 14977 16838 15023 16890
rect 15023 16838 15033 16890
rect 15057 16838 15087 16890
rect 15087 16838 15113 16890
rect 14817 16836 14873 16838
rect 14897 16836 14953 16838
rect 14977 16836 15033 16838
rect 15057 16836 15113 16838
rect 18282 20698 18338 20700
rect 18362 20698 18418 20700
rect 18442 20698 18498 20700
rect 18522 20698 18578 20700
rect 18282 20646 18308 20698
rect 18308 20646 18338 20698
rect 18362 20646 18372 20698
rect 18372 20646 18418 20698
rect 18442 20646 18488 20698
rect 18488 20646 18498 20698
rect 18522 20646 18552 20698
rect 18552 20646 18578 20698
rect 18282 20644 18338 20646
rect 18362 20644 18418 20646
rect 18442 20644 18498 20646
rect 18522 20644 18578 20646
rect 18282 19610 18338 19612
rect 18362 19610 18418 19612
rect 18442 19610 18498 19612
rect 18522 19610 18578 19612
rect 18282 19558 18308 19610
rect 18308 19558 18338 19610
rect 18362 19558 18372 19610
rect 18372 19558 18418 19610
rect 18442 19558 18488 19610
rect 18488 19558 18498 19610
rect 18522 19558 18552 19610
rect 18552 19558 18578 19610
rect 18282 19556 18338 19558
rect 18362 19556 18418 19558
rect 18442 19556 18498 19558
rect 18522 19556 18578 19558
rect 14817 15802 14873 15804
rect 14897 15802 14953 15804
rect 14977 15802 15033 15804
rect 15057 15802 15113 15804
rect 14817 15750 14843 15802
rect 14843 15750 14873 15802
rect 14897 15750 14907 15802
rect 14907 15750 14953 15802
rect 14977 15750 15023 15802
rect 15023 15750 15033 15802
rect 15057 15750 15087 15802
rect 15087 15750 15113 15802
rect 14817 15748 14873 15750
rect 14897 15748 14953 15750
rect 14977 15748 15033 15750
rect 15057 15748 15113 15750
rect 14817 14714 14873 14716
rect 14897 14714 14953 14716
rect 14977 14714 15033 14716
rect 15057 14714 15113 14716
rect 14817 14662 14843 14714
rect 14843 14662 14873 14714
rect 14897 14662 14907 14714
rect 14907 14662 14953 14714
rect 14977 14662 15023 14714
rect 15023 14662 15033 14714
rect 15057 14662 15087 14714
rect 15087 14662 15113 14714
rect 14817 14660 14873 14662
rect 14897 14660 14953 14662
rect 14977 14660 15033 14662
rect 15057 14660 15113 14662
rect 14817 13626 14873 13628
rect 14897 13626 14953 13628
rect 14977 13626 15033 13628
rect 15057 13626 15113 13628
rect 14817 13574 14843 13626
rect 14843 13574 14873 13626
rect 14897 13574 14907 13626
rect 14907 13574 14953 13626
rect 14977 13574 15023 13626
rect 15023 13574 15033 13626
rect 15057 13574 15087 13626
rect 15087 13574 15113 13626
rect 14817 13572 14873 13574
rect 14897 13572 14953 13574
rect 14977 13572 15033 13574
rect 15057 13572 15113 13574
rect 14817 12538 14873 12540
rect 14897 12538 14953 12540
rect 14977 12538 15033 12540
rect 15057 12538 15113 12540
rect 14817 12486 14843 12538
rect 14843 12486 14873 12538
rect 14897 12486 14907 12538
rect 14907 12486 14953 12538
rect 14977 12486 15023 12538
rect 15023 12486 15033 12538
rect 15057 12486 15087 12538
rect 15087 12486 15113 12538
rect 14817 12484 14873 12486
rect 14897 12484 14953 12486
rect 14977 12484 15033 12486
rect 15057 12484 15113 12486
rect 14817 11450 14873 11452
rect 14897 11450 14953 11452
rect 14977 11450 15033 11452
rect 15057 11450 15113 11452
rect 14817 11398 14843 11450
rect 14843 11398 14873 11450
rect 14897 11398 14907 11450
rect 14907 11398 14953 11450
rect 14977 11398 15023 11450
rect 15023 11398 15033 11450
rect 15057 11398 15087 11450
rect 15087 11398 15113 11450
rect 14817 11396 14873 11398
rect 14897 11396 14953 11398
rect 14977 11396 15033 11398
rect 15057 11396 15113 11398
rect 18282 18522 18338 18524
rect 18362 18522 18418 18524
rect 18442 18522 18498 18524
rect 18522 18522 18578 18524
rect 18282 18470 18308 18522
rect 18308 18470 18338 18522
rect 18362 18470 18372 18522
rect 18372 18470 18418 18522
rect 18442 18470 18488 18522
rect 18488 18470 18498 18522
rect 18522 18470 18552 18522
rect 18552 18470 18578 18522
rect 18282 18468 18338 18470
rect 18362 18468 18418 18470
rect 18442 18468 18498 18470
rect 18522 18468 18578 18470
rect 17498 17584 17554 17640
rect 16394 11328 16450 11384
rect 14817 10362 14873 10364
rect 14897 10362 14953 10364
rect 14977 10362 15033 10364
rect 15057 10362 15113 10364
rect 14817 10310 14843 10362
rect 14843 10310 14873 10362
rect 14897 10310 14907 10362
rect 14907 10310 14953 10362
rect 14977 10310 15023 10362
rect 15023 10310 15033 10362
rect 15057 10310 15087 10362
rect 15087 10310 15113 10362
rect 14817 10308 14873 10310
rect 14897 10308 14953 10310
rect 14977 10308 15033 10310
rect 15057 10308 15113 10310
rect 14817 9274 14873 9276
rect 14897 9274 14953 9276
rect 14977 9274 15033 9276
rect 15057 9274 15113 9276
rect 14817 9222 14843 9274
rect 14843 9222 14873 9274
rect 14897 9222 14907 9274
rect 14907 9222 14953 9274
rect 14977 9222 15023 9274
rect 15023 9222 15033 9274
rect 15057 9222 15087 9274
rect 15087 9222 15113 9274
rect 14817 9220 14873 9222
rect 14897 9220 14953 9222
rect 14977 9220 15033 9222
rect 15057 9220 15113 9222
rect 14817 8186 14873 8188
rect 14897 8186 14953 8188
rect 14977 8186 15033 8188
rect 15057 8186 15113 8188
rect 14817 8134 14843 8186
rect 14843 8134 14873 8186
rect 14897 8134 14907 8186
rect 14907 8134 14953 8186
rect 14977 8134 15023 8186
rect 15023 8134 15033 8186
rect 15057 8134 15087 8186
rect 15087 8134 15113 8186
rect 14817 8132 14873 8134
rect 14897 8132 14953 8134
rect 14977 8132 15033 8134
rect 15057 8132 15113 8134
rect 14830 7384 14886 7440
rect 14817 7098 14873 7100
rect 14897 7098 14953 7100
rect 14977 7098 15033 7100
rect 15057 7098 15113 7100
rect 14817 7046 14843 7098
rect 14843 7046 14873 7098
rect 14897 7046 14907 7098
rect 14907 7046 14953 7098
rect 14977 7046 15023 7098
rect 15023 7046 15033 7098
rect 15057 7046 15087 7098
rect 15087 7046 15113 7098
rect 14817 7044 14873 7046
rect 14897 7044 14953 7046
rect 14977 7044 15033 7046
rect 15057 7044 15113 7046
rect 14817 6010 14873 6012
rect 14897 6010 14953 6012
rect 14977 6010 15033 6012
rect 15057 6010 15113 6012
rect 14817 5958 14843 6010
rect 14843 5958 14873 6010
rect 14897 5958 14907 6010
rect 14907 5958 14953 6010
rect 14977 5958 15023 6010
rect 15023 5958 15033 6010
rect 15057 5958 15087 6010
rect 15087 5958 15113 6010
rect 14817 5956 14873 5958
rect 14897 5956 14953 5958
rect 14977 5956 15033 5958
rect 15057 5956 15113 5958
rect 14817 4922 14873 4924
rect 14897 4922 14953 4924
rect 14977 4922 15033 4924
rect 15057 4922 15113 4924
rect 14817 4870 14843 4922
rect 14843 4870 14873 4922
rect 14897 4870 14907 4922
rect 14907 4870 14953 4922
rect 14977 4870 15023 4922
rect 15023 4870 15033 4922
rect 15057 4870 15087 4922
rect 15087 4870 15113 4922
rect 14817 4868 14873 4870
rect 14897 4868 14953 4870
rect 14977 4868 15033 4870
rect 15057 4868 15113 4870
rect 16670 8356 16726 8392
rect 16670 8336 16672 8356
rect 16672 8336 16724 8356
rect 16724 8336 16726 8356
rect 14817 3834 14873 3836
rect 14897 3834 14953 3836
rect 14977 3834 15033 3836
rect 15057 3834 15113 3836
rect 14817 3782 14843 3834
rect 14843 3782 14873 3834
rect 14897 3782 14907 3834
rect 14907 3782 14953 3834
rect 14977 3782 15023 3834
rect 15023 3782 15033 3834
rect 15057 3782 15087 3834
rect 15087 3782 15113 3834
rect 14817 3780 14873 3782
rect 14897 3780 14953 3782
rect 14977 3780 15033 3782
rect 15057 3780 15113 3782
rect 14817 2746 14873 2748
rect 14897 2746 14953 2748
rect 14977 2746 15033 2748
rect 15057 2746 15113 2748
rect 14817 2694 14843 2746
rect 14843 2694 14873 2746
rect 14897 2694 14907 2746
rect 14907 2694 14953 2746
rect 14977 2694 15023 2746
rect 15023 2694 15033 2746
rect 15057 2694 15087 2746
rect 15087 2694 15113 2746
rect 14817 2692 14873 2694
rect 14897 2692 14953 2694
rect 14977 2692 15033 2694
rect 15057 2692 15113 2694
rect 6366 176 6422 232
rect 17130 7928 17186 7984
rect 18282 17434 18338 17436
rect 18362 17434 18418 17436
rect 18442 17434 18498 17436
rect 18522 17434 18578 17436
rect 18282 17382 18308 17434
rect 18308 17382 18338 17434
rect 18362 17382 18372 17434
rect 18372 17382 18418 17434
rect 18442 17382 18488 17434
rect 18488 17382 18498 17434
rect 18522 17382 18552 17434
rect 18552 17382 18578 17434
rect 18282 17380 18338 17382
rect 18362 17380 18418 17382
rect 18442 17380 18498 17382
rect 18522 17380 18578 17382
rect 18282 16346 18338 16348
rect 18362 16346 18418 16348
rect 18442 16346 18498 16348
rect 18522 16346 18578 16348
rect 18282 16294 18308 16346
rect 18308 16294 18338 16346
rect 18362 16294 18372 16346
rect 18372 16294 18418 16346
rect 18442 16294 18488 16346
rect 18488 16294 18498 16346
rect 18522 16294 18552 16346
rect 18552 16294 18578 16346
rect 18282 16292 18338 16294
rect 18362 16292 18418 16294
rect 18442 16292 18498 16294
rect 18522 16292 18578 16294
rect 20626 22208 20682 22264
rect 19154 21664 19210 21720
rect 19246 21256 19302 21312
rect 20442 20712 20498 20768
rect 19246 17448 19302 17504
rect 18282 15258 18338 15260
rect 18362 15258 18418 15260
rect 18442 15258 18498 15260
rect 18522 15258 18578 15260
rect 18282 15206 18308 15258
rect 18308 15206 18338 15258
rect 18362 15206 18372 15258
rect 18372 15206 18418 15258
rect 18442 15206 18488 15258
rect 18488 15206 18498 15258
rect 18522 15206 18552 15258
rect 18552 15206 18578 15258
rect 18282 15204 18338 15206
rect 18362 15204 18418 15206
rect 18442 15204 18498 15206
rect 18522 15204 18578 15206
rect 18282 14170 18338 14172
rect 18362 14170 18418 14172
rect 18442 14170 18498 14172
rect 18522 14170 18578 14172
rect 18282 14118 18308 14170
rect 18308 14118 18338 14170
rect 18362 14118 18372 14170
rect 18372 14118 18418 14170
rect 18442 14118 18488 14170
rect 18488 14118 18498 14170
rect 18522 14118 18552 14170
rect 18552 14118 18578 14170
rect 18282 14116 18338 14118
rect 18362 14116 18418 14118
rect 18442 14116 18498 14118
rect 18522 14116 18578 14118
rect 17774 11636 17776 11656
rect 17776 11636 17828 11656
rect 17828 11636 17830 11656
rect 17774 11600 17830 11636
rect 18282 13082 18338 13084
rect 18362 13082 18418 13084
rect 18442 13082 18498 13084
rect 18522 13082 18578 13084
rect 18282 13030 18308 13082
rect 18308 13030 18338 13082
rect 18362 13030 18372 13082
rect 18372 13030 18418 13082
rect 18442 13030 18488 13082
rect 18488 13030 18498 13082
rect 18522 13030 18552 13082
rect 18552 13030 18578 13082
rect 18282 13028 18338 13030
rect 18362 13028 18418 13030
rect 18442 13028 18498 13030
rect 18522 13028 18578 13030
rect 18282 11994 18338 11996
rect 18362 11994 18418 11996
rect 18442 11994 18498 11996
rect 18522 11994 18578 11996
rect 18282 11942 18308 11994
rect 18308 11942 18338 11994
rect 18362 11942 18372 11994
rect 18372 11942 18418 11994
rect 18442 11942 18488 11994
rect 18488 11942 18498 11994
rect 18522 11942 18552 11994
rect 18552 11942 18578 11994
rect 18282 11940 18338 11942
rect 18362 11940 18418 11942
rect 18442 11940 18498 11942
rect 18522 11940 18578 11942
rect 18418 11636 18420 11656
rect 18420 11636 18472 11656
rect 18472 11636 18474 11656
rect 18418 11600 18474 11636
rect 19062 11872 19118 11928
rect 17774 8064 17830 8120
rect 18282 10906 18338 10908
rect 18362 10906 18418 10908
rect 18442 10906 18498 10908
rect 18522 10906 18578 10908
rect 18282 10854 18308 10906
rect 18308 10854 18338 10906
rect 18362 10854 18372 10906
rect 18372 10854 18418 10906
rect 18442 10854 18488 10906
rect 18488 10854 18498 10906
rect 18522 10854 18552 10906
rect 18552 10854 18578 10906
rect 18282 10852 18338 10854
rect 18362 10852 18418 10854
rect 18442 10852 18498 10854
rect 18522 10852 18578 10854
rect 18282 9818 18338 9820
rect 18362 9818 18418 9820
rect 18442 9818 18498 9820
rect 18522 9818 18578 9820
rect 18282 9766 18308 9818
rect 18308 9766 18338 9818
rect 18362 9766 18372 9818
rect 18372 9766 18418 9818
rect 18442 9766 18488 9818
rect 18488 9766 18498 9818
rect 18522 9766 18552 9818
rect 18552 9766 18578 9818
rect 18282 9764 18338 9766
rect 18362 9764 18418 9766
rect 18442 9764 18498 9766
rect 18522 9764 18578 9766
rect 18326 9580 18382 9616
rect 18326 9560 18328 9580
rect 18328 9560 18380 9580
rect 18380 9560 18382 9580
rect 18602 9424 18658 9480
rect 18282 8730 18338 8732
rect 18362 8730 18418 8732
rect 18442 8730 18498 8732
rect 18522 8730 18578 8732
rect 18282 8678 18308 8730
rect 18308 8678 18338 8730
rect 18362 8678 18372 8730
rect 18372 8678 18418 8730
rect 18442 8678 18488 8730
rect 18488 8678 18498 8730
rect 18522 8678 18552 8730
rect 18552 8678 18578 8730
rect 18282 8676 18338 8678
rect 18362 8676 18418 8678
rect 18442 8676 18498 8678
rect 18522 8676 18578 8678
rect 18282 7642 18338 7644
rect 18362 7642 18418 7644
rect 18442 7642 18498 7644
rect 18522 7642 18578 7644
rect 18282 7590 18308 7642
rect 18308 7590 18338 7642
rect 18362 7590 18372 7642
rect 18372 7590 18418 7642
rect 18442 7590 18488 7642
rect 18488 7590 18498 7642
rect 18522 7590 18552 7642
rect 18552 7590 18578 7642
rect 18282 7588 18338 7590
rect 18362 7588 18418 7590
rect 18442 7588 18498 7590
rect 18522 7588 18578 7590
rect 17958 5788 17960 5808
rect 17960 5788 18012 5808
rect 18012 5788 18014 5808
rect 17958 5752 18014 5788
rect 17958 4800 18014 4856
rect 17406 3440 17462 3496
rect 18282 6554 18338 6556
rect 18362 6554 18418 6556
rect 18442 6554 18498 6556
rect 18522 6554 18578 6556
rect 18282 6502 18308 6554
rect 18308 6502 18338 6554
rect 18362 6502 18372 6554
rect 18372 6502 18418 6554
rect 18442 6502 18488 6554
rect 18488 6502 18498 6554
rect 18522 6502 18552 6554
rect 18552 6502 18578 6554
rect 18282 6500 18338 6502
rect 18362 6500 18418 6502
rect 18442 6500 18498 6502
rect 18522 6500 18578 6502
rect 18878 10376 18934 10432
rect 18282 5466 18338 5468
rect 18362 5466 18418 5468
rect 18442 5466 18498 5468
rect 18522 5466 18578 5468
rect 18282 5414 18308 5466
rect 18308 5414 18338 5466
rect 18362 5414 18372 5466
rect 18372 5414 18418 5466
rect 18442 5414 18488 5466
rect 18488 5414 18498 5466
rect 18522 5414 18552 5466
rect 18552 5414 18578 5466
rect 18282 5412 18338 5414
rect 18362 5412 18418 5414
rect 18442 5412 18498 5414
rect 18522 5412 18578 5414
rect 18282 4378 18338 4380
rect 18362 4378 18418 4380
rect 18442 4378 18498 4380
rect 18522 4378 18578 4380
rect 18282 4326 18308 4378
rect 18308 4326 18338 4378
rect 18362 4326 18372 4378
rect 18372 4326 18418 4378
rect 18442 4326 18488 4378
rect 18488 4326 18498 4378
rect 18522 4326 18552 4378
rect 18552 4326 18578 4378
rect 18282 4324 18338 4326
rect 18362 4324 18418 4326
rect 18442 4324 18498 4326
rect 18522 4324 18578 4326
rect 18282 3290 18338 3292
rect 18362 3290 18418 3292
rect 18442 3290 18498 3292
rect 18522 3290 18578 3292
rect 18282 3238 18308 3290
rect 18308 3238 18338 3290
rect 18362 3238 18372 3290
rect 18372 3238 18418 3290
rect 18442 3238 18488 3290
rect 18488 3238 18498 3290
rect 18522 3238 18552 3290
rect 18552 3238 18578 3290
rect 18282 3236 18338 3238
rect 18362 3236 18418 3238
rect 18442 3236 18498 3238
rect 18522 3236 18578 3238
rect 18694 2896 18750 2952
rect 18282 2202 18338 2204
rect 18362 2202 18418 2204
rect 18442 2202 18498 2204
rect 18522 2202 18578 2204
rect 18282 2150 18308 2202
rect 18308 2150 18338 2202
rect 18362 2150 18372 2202
rect 18372 2150 18418 2202
rect 18442 2150 18488 2202
rect 18488 2150 18498 2202
rect 18522 2150 18552 2202
rect 18552 2150 18578 2202
rect 18282 2148 18338 2150
rect 18362 2148 18418 2150
rect 18442 2148 18498 2150
rect 18522 2148 18578 2150
rect 18786 2488 18842 2544
rect 16946 584 17002 640
rect 19062 9968 19118 10024
rect 19154 7656 19210 7712
rect 19246 7112 19302 7168
rect 19338 6196 19340 6216
rect 19340 6196 19392 6216
rect 19392 6196 19394 6216
rect 19338 6160 19394 6196
rect 21086 20304 21142 20360
rect 20442 19760 20498 19816
rect 19798 9560 19854 9616
rect 20166 7928 20222 7984
rect 19798 6180 19854 6216
rect 19798 6160 19800 6180
rect 19800 6160 19852 6180
rect 19852 6160 19854 6180
rect 19246 992 19302 1048
rect 20442 18420 20498 18456
rect 20442 18400 20444 18420
rect 20444 18400 20496 18420
rect 20496 18400 20498 18420
rect 20442 16088 20498 16144
rect 20626 16496 20682 16552
rect 20994 19352 21050 19408
rect 21086 18808 21142 18864
rect 20994 18028 20996 18048
rect 20996 18028 21048 18048
rect 21048 18028 21050 18048
rect 20994 17992 21050 18028
rect 21086 17040 21142 17096
rect 20626 15136 20682 15192
rect 20442 10920 20498 10976
rect 21086 15544 21142 15600
rect 21086 14592 21142 14648
rect 20994 14184 21050 14240
rect 21178 13776 21234 13832
rect 20902 12824 20958 12880
rect 20534 9016 20590 9072
rect 20074 1944 20130 2000
rect 20626 5208 20682 5264
rect 20626 3848 20682 3904
rect 20994 12280 21050 12336
rect 21270 13232 21326 13288
rect 21362 5616 21418 5672
rect 21270 4392 21326 4448
rect 21178 1536 21234 1592
rect 18970 176 19026 232
<< metal3 >>
rect 0 22674 800 22704
rect 3325 22674 3391 22677
rect 0 22672 3391 22674
rect 0 22616 3330 22672
rect 3386 22616 3391 22672
rect 0 22614 3391 22616
rect 0 22584 800 22614
rect 3325 22611 3391 22614
rect 18689 22674 18755 22677
rect 22200 22674 23000 22704
rect 18689 22672 23000 22674
rect 18689 22616 18694 22672
rect 18750 22616 23000 22672
rect 18689 22614 23000 22616
rect 18689 22611 18755 22614
rect 22200 22584 23000 22614
rect 0 22266 800 22296
rect 2865 22266 2931 22269
rect 0 22264 2931 22266
rect 0 22208 2870 22264
rect 2926 22208 2931 22264
rect 0 22206 2931 22208
rect 0 22176 800 22206
rect 2865 22203 2931 22206
rect 20621 22266 20687 22269
rect 22200 22266 23000 22296
rect 20621 22264 23000 22266
rect 20621 22208 20626 22264
rect 20682 22208 23000 22264
rect 20621 22206 23000 22208
rect 20621 22203 20687 22206
rect 22200 22176 23000 22206
rect 0 21722 800 21752
rect 2773 21722 2839 21725
rect 0 21720 2839 21722
rect 0 21664 2778 21720
rect 2834 21664 2839 21720
rect 0 21662 2839 21664
rect 0 21632 800 21662
rect 2773 21659 2839 21662
rect 19149 21722 19215 21725
rect 22200 21722 23000 21752
rect 19149 21720 23000 21722
rect 19149 21664 19154 21720
rect 19210 21664 23000 21720
rect 19149 21662 23000 21664
rect 19149 21659 19215 21662
rect 22200 21632 23000 21662
rect 0 21314 800 21344
rect 1945 21314 2011 21317
rect 0 21312 2011 21314
rect 0 21256 1950 21312
rect 2006 21256 2011 21312
rect 0 21254 2011 21256
rect 0 21224 800 21254
rect 1945 21251 2011 21254
rect 19241 21314 19307 21317
rect 22200 21314 23000 21344
rect 19241 21312 23000 21314
rect 19241 21256 19246 21312
rect 19302 21256 23000 21312
rect 19241 21254 23000 21256
rect 19241 21251 19307 21254
rect 22200 21224 23000 21254
rect 0 20770 800 20800
rect 3049 20770 3115 20773
rect 0 20768 3115 20770
rect 0 20712 3054 20768
rect 3110 20712 3115 20768
rect 0 20710 3115 20712
rect 0 20680 800 20710
rect 3049 20707 3115 20710
rect 20437 20770 20503 20773
rect 22200 20770 23000 20800
rect 20437 20768 23000 20770
rect 20437 20712 20442 20768
rect 20498 20712 23000 20768
rect 20437 20710 23000 20712
rect 20437 20707 20503 20710
rect 4409 20704 4729 20705
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 20639 4729 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 18270 20704 18590 20705
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 22200 20680 23000 20710
rect 18270 20639 18590 20640
rect 0 20362 800 20392
rect 2957 20362 3023 20365
rect 0 20360 3023 20362
rect 0 20304 2962 20360
rect 3018 20304 3023 20360
rect 0 20302 3023 20304
rect 0 20272 800 20302
rect 2957 20299 3023 20302
rect 21081 20362 21147 20365
rect 22200 20362 23000 20392
rect 21081 20360 23000 20362
rect 21081 20304 21086 20360
rect 21142 20304 23000 20360
rect 21081 20302 23000 20304
rect 21081 20299 21147 20302
rect 22200 20272 23000 20302
rect 7874 20160 8194 20161
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8194 20160
rect 7874 20095 8194 20096
rect 14805 20160 15125 20161
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 20095 15125 20096
rect 0 19818 800 19848
rect 1945 19818 2011 19821
rect 0 19816 2011 19818
rect 0 19760 1950 19816
rect 2006 19760 2011 19816
rect 0 19758 2011 19760
rect 0 19728 800 19758
rect 1945 19755 2011 19758
rect 20437 19818 20503 19821
rect 22200 19818 23000 19848
rect 20437 19816 23000 19818
rect 20437 19760 20442 19816
rect 20498 19760 23000 19816
rect 20437 19758 23000 19760
rect 20437 19755 20503 19758
rect 22200 19728 23000 19758
rect 4409 19616 4729 19617
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 19551 4729 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 18270 19616 18590 19617
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 19551 18590 19552
rect 0 19410 800 19440
rect 2773 19410 2839 19413
rect 0 19408 2839 19410
rect 0 19352 2778 19408
rect 2834 19352 2839 19408
rect 0 19350 2839 19352
rect 0 19320 800 19350
rect 2773 19347 2839 19350
rect 20989 19410 21055 19413
rect 22200 19410 23000 19440
rect 20989 19408 23000 19410
rect 20989 19352 20994 19408
rect 21050 19352 23000 19408
rect 20989 19350 23000 19352
rect 20989 19347 21055 19350
rect 22200 19320 23000 19350
rect 7874 19072 8194 19073
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8194 19072
rect 7874 19007 8194 19008
rect 14805 19072 15125 19073
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 19007 15125 19008
rect 0 18866 800 18896
rect 1945 18866 2011 18869
rect 0 18864 2011 18866
rect 0 18808 1950 18864
rect 2006 18808 2011 18864
rect 0 18806 2011 18808
rect 0 18776 800 18806
rect 1945 18803 2011 18806
rect 21081 18866 21147 18869
rect 22200 18866 23000 18896
rect 21081 18864 23000 18866
rect 21081 18808 21086 18864
rect 21142 18808 23000 18864
rect 21081 18806 23000 18808
rect 21081 18803 21147 18806
rect 22200 18776 23000 18806
rect 4409 18528 4729 18529
rect 0 18458 800 18488
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 18463 4729 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 18270 18528 18590 18529
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 18270 18463 18590 18464
rect 1945 18458 2011 18461
rect 0 18456 2011 18458
rect 0 18400 1950 18456
rect 2006 18400 2011 18456
rect 0 18398 2011 18400
rect 0 18368 800 18398
rect 1945 18395 2011 18398
rect 20437 18458 20503 18461
rect 22200 18458 23000 18488
rect 20437 18456 23000 18458
rect 20437 18400 20442 18456
rect 20498 18400 23000 18456
rect 20437 18398 23000 18400
rect 20437 18395 20503 18398
rect 22200 18368 23000 18398
rect 0 18050 800 18080
rect 1669 18050 1735 18053
rect 0 18048 1735 18050
rect 0 17992 1674 18048
rect 1730 17992 1735 18048
rect 0 17990 1735 17992
rect 0 17960 800 17990
rect 1669 17987 1735 17990
rect 20989 18050 21055 18053
rect 22200 18050 23000 18080
rect 20989 18048 23000 18050
rect 20989 17992 20994 18048
rect 21050 17992 23000 18048
rect 20989 17990 23000 17992
rect 20989 17987 21055 17990
rect 7874 17984 8194 17985
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8194 17984
rect 7874 17919 8194 17920
rect 14805 17984 15125 17985
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 22200 17960 23000 17990
rect 14805 17919 15125 17920
rect 13261 17778 13327 17781
rect 13721 17778 13787 17781
rect 13261 17776 13787 17778
rect 13261 17720 13266 17776
rect 13322 17720 13726 17776
rect 13782 17720 13787 17776
rect 13261 17718 13787 17720
rect 13261 17715 13327 17718
rect 13721 17715 13787 17718
rect 12249 17642 12315 17645
rect 17493 17642 17559 17645
rect 12249 17640 17559 17642
rect 12249 17584 12254 17640
rect 12310 17584 17498 17640
rect 17554 17584 17559 17640
rect 12249 17582 17559 17584
rect 12249 17579 12315 17582
rect 17493 17579 17559 17582
rect 0 17506 800 17536
rect 2773 17506 2839 17509
rect 0 17504 2839 17506
rect 0 17448 2778 17504
rect 2834 17448 2839 17504
rect 0 17446 2839 17448
rect 0 17416 800 17446
rect 2773 17443 2839 17446
rect 19241 17506 19307 17509
rect 22200 17506 23000 17536
rect 19241 17504 23000 17506
rect 19241 17448 19246 17504
rect 19302 17448 23000 17504
rect 19241 17446 23000 17448
rect 19241 17443 19307 17446
rect 4409 17440 4729 17441
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 17375 4729 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 18270 17440 18590 17441
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 22200 17416 23000 17446
rect 18270 17375 18590 17376
rect 0 17098 800 17128
rect 1945 17098 2011 17101
rect 0 17096 2011 17098
rect 0 17040 1950 17096
rect 2006 17040 2011 17096
rect 0 17038 2011 17040
rect 0 17008 800 17038
rect 1945 17035 2011 17038
rect 21081 17098 21147 17101
rect 22200 17098 23000 17128
rect 21081 17096 23000 17098
rect 21081 17040 21086 17096
rect 21142 17040 23000 17096
rect 21081 17038 23000 17040
rect 21081 17035 21147 17038
rect 22200 17008 23000 17038
rect 7874 16896 8194 16897
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8194 16896
rect 7874 16831 8194 16832
rect 14805 16896 15125 16897
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 16831 15125 16832
rect 0 16554 800 16584
rect 2497 16554 2563 16557
rect 0 16552 2563 16554
rect 0 16496 2502 16552
rect 2558 16496 2563 16552
rect 0 16494 2563 16496
rect 0 16464 800 16494
rect 2497 16491 2563 16494
rect 9949 16554 10015 16557
rect 12985 16554 13051 16557
rect 9949 16552 13051 16554
rect 9949 16496 9954 16552
rect 10010 16496 12990 16552
rect 13046 16496 13051 16552
rect 9949 16494 13051 16496
rect 9949 16491 10015 16494
rect 12985 16491 13051 16494
rect 20621 16554 20687 16557
rect 22200 16554 23000 16584
rect 20621 16552 23000 16554
rect 20621 16496 20626 16552
rect 20682 16496 23000 16552
rect 20621 16494 23000 16496
rect 20621 16491 20687 16494
rect 22200 16464 23000 16494
rect 4409 16352 4729 16353
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 16287 4729 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 18270 16352 18590 16353
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 16287 18590 16288
rect 0 16146 800 16176
rect 1669 16146 1735 16149
rect 0 16144 1735 16146
rect 0 16088 1674 16144
rect 1730 16088 1735 16144
rect 0 16086 1735 16088
rect 0 16056 800 16086
rect 1669 16083 1735 16086
rect 20437 16146 20503 16149
rect 22200 16146 23000 16176
rect 20437 16144 23000 16146
rect 20437 16088 20442 16144
rect 20498 16088 23000 16144
rect 20437 16086 23000 16088
rect 20437 16083 20503 16086
rect 22200 16056 23000 16086
rect 7874 15808 8194 15809
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8194 15808
rect 7874 15743 8194 15744
rect 14805 15808 15125 15809
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 15743 15125 15744
rect 0 15602 800 15632
rect 1945 15602 2011 15605
rect 0 15600 2011 15602
rect 0 15544 1950 15600
rect 2006 15544 2011 15600
rect 0 15542 2011 15544
rect 0 15512 800 15542
rect 1945 15539 2011 15542
rect 21081 15602 21147 15605
rect 22200 15602 23000 15632
rect 21081 15600 23000 15602
rect 21081 15544 21086 15600
rect 21142 15544 23000 15600
rect 21081 15542 23000 15544
rect 21081 15539 21147 15542
rect 22200 15512 23000 15542
rect 4409 15264 4729 15265
rect 0 15194 800 15224
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 15199 4729 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 18270 15264 18590 15265
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 18270 15199 18590 15200
rect 1853 15194 1919 15197
rect 0 15192 1919 15194
rect 0 15136 1858 15192
rect 1914 15136 1919 15192
rect 0 15134 1919 15136
rect 0 15104 800 15134
rect 1853 15131 1919 15134
rect 20621 15194 20687 15197
rect 22200 15194 23000 15224
rect 20621 15192 23000 15194
rect 20621 15136 20626 15192
rect 20682 15136 23000 15192
rect 20621 15134 23000 15136
rect 20621 15131 20687 15134
rect 22200 15104 23000 15134
rect 7874 14720 8194 14721
rect 0 14650 800 14680
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8194 14720
rect 7874 14655 8194 14656
rect 14805 14720 15125 14721
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 14655 15125 14656
rect 1853 14650 1919 14653
rect 0 14648 1919 14650
rect 0 14592 1858 14648
rect 1914 14592 1919 14648
rect 0 14590 1919 14592
rect 0 14560 800 14590
rect 1853 14587 1919 14590
rect 21081 14650 21147 14653
rect 22200 14650 23000 14680
rect 21081 14648 23000 14650
rect 21081 14592 21086 14648
rect 21142 14592 23000 14648
rect 21081 14590 23000 14592
rect 21081 14587 21147 14590
rect 22200 14560 23000 14590
rect 0 14242 800 14272
rect 1945 14242 2011 14245
rect 0 14240 2011 14242
rect 0 14184 1950 14240
rect 2006 14184 2011 14240
rect 0 14182 2011 14184
rect 0 14152 800 14182
rect 1945 14179 2011 14182
rect 20989 14242 21055 14245
rect 22200 14242 23000 14272
rect 20989 14240 23000 14242
rect 20989 14184 20994 14240
rect 21050 14184 23000 14240
rect 20989 14182 23000 14184
rect 20989 14179 21055 14182
rect 4409 14176 4729 14177
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 14111 4729 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 18270 14176 18590 14177
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 22200 14152 23000 14182
rect 18270 14111 18590 14112
rect 0 13834 800 13864
rect 2865 13834 2931 13837
rect 0 13832 2931 13834
rect 0 13776 2870 13832
rect 2926 13776 2931 13832
rect 0 13774 2931 13776
rect 0 13744 800 13774
rect 2865 13771 2931 13774
rect 21173 13834 21239 13837
rect 22200 13834 23000 13864
rect 21173 13832 23000 13834
rect 21173 13776 21178 13832
rect 21234 13776 23000 13832
rect 21173 13774 23000 13776
rect 21173 13771 21239 13774
rect 22200 13744 23000 13774
rect 7874 13632 8194 13633
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8194 13632
rect 7874 13567 8194 13568
rect 14805 13632 15125 13633
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 13567 15125 13568
rect 0 13290 800 13320
rect 2773 13290 2839 13293
rect 0 13288 2839 13290
rect 0 13232 2778 13288
rect 2834 13232 2839 13288
rect 0 13230 2839 13232
rect 0 13200 800 13230
rect 2773 13227 2839 13230
rect 21265 13290 21331 13293
rect 22200 13290 23000 13320
rect 21265 13288 23000 13290
rect 21265 13232 21270 13288
rect 21326 13232 23000 13288
rect 21265 13230 23000 13232
rect 21265 13227 21331 13230
rect 22200 13200 23000 13230
rect 4409 13088 4729 13089
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 13023 4729 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 18270 13088 18590 13089
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 13023 18590 13024
rect 0 12882 800 12912
rect 4061 12882 4127 12885
rect 0 12880 4127 12882
rect 0 12824 4066 12880
rect 4122 12824 4127 12880
rect 0 12822 4127 12824
rect 0 12792 800 12822
rect 4061 12819 4127 12822
rect 20897 12882 20963 12885
rect 22200 12882 23000 12912
rect 20897 12880 23000 12882
rect 20897 12824 20902 12880
rect 20958 12824 23000 12880
rect 20897 12822 23000 12824
rect 20897 12819 20963 12822
rect 22200 12792 23000 12822
rect 7874 12544 8194 12545
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8194 12544
rect 7874 12479 8194 12480
rect 14805 12544 15125 12545
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 12479 15125 12480
rect 0 12338 800 12368
rect 3877 12338 3943 12341
rect 0 12336 3943 12338
rect 0 12280 3882 12336
rect 3938 12280 3943 12336
rect 0 12278 3943 12280
rect 0 12248 800 12278
rect 3877 12275 3943 12278
rect 20989 12338 21055 12341
rect 22200 12338 23000 12368
rect 20989 12336 23000 12338
rect 20989 12280 20994 12336
rect 21050 12280 23000 12336
rect 20989 12278 23000 12280
rect 20989 12275 21055 12278
rect 22200 12248 23000 12278
rect 2129 12202 2195 12205
rect 9489 12202 9555 12205
rect 2129 12200 9555 12202
rect 2129 12144 2134 12200
rect 2190 12144 9494 12200
rect 9550 12144 9555 12200
rect 2129 12142 9555 12144
rect 2129 12139 2195 12142
rect 9489 12139 9555 12142
rect 4409 12000 4729 12001
rect 0 11930 800 11960
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 11935 4729 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 18270 12000 18590 12001
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 18270 11935 18590 11936
rect 4061 11930 4127 11933
rect 0 11928 4127 11930
rect 0 11872 4066 11928
rect 4122 11872 4127 11928
rect 0 11870 4127 11872
rect 0 11840 800 11870
rect 4061 11867 4127 11870
rect 19057 11930 19123 11933
rect 22200 11930 23000 11960
rect 19057 11928 23000 11930
rect 19057 11872 19062 11928
rect 19118 11872 23000 11928
rect 19057 11870 23000 11872
rect 19057 11867 19123 11870
rect 22200 11840 23000 11870
rect 17769 11658 17835 11661
rect 18413 11658 18479 11661
rect 17769 11656 18479 11658
rect 17769 11600 17774 11656
rect 17830 11600 18418 11656
rect 18474 11600 18479 11656
rect 17769 11598 18479 11600
rect 17769 11595 17835 11598
rect 18413 11595 18479 11598
rect 7874 11456 8194 11457
rect 0 11386 800 11416
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8194 11456
rect 7874 11391 8194 11392
rect 14805 11456 15125 11457
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 11391 15125 11392
rect 5533 11386 5599 11389
rect 0 11384 5599 11386
rect 0 11328 5538 11384
rect 5594 11328 5599 11384
rect 0 11326 5599 11328
rect 0 11296 800 11326
rect 5533 11323 5599 11326
rect 11881 11386 11947 11389
rect 13077 11386 13143 11389
rect 11881 11384 13143 11386
rect 11881 11328 11886 11384
rect 11942 11328 13082 11384
rect 13138 11328 13143 11384
rect 11881 11326 13143 11328
rect 11881 11323 11947 11326
rect 13077 11323 13143 11326
rect 16389 11386 16455 11389
rect 22200 11386 23000 11416
rect 16389 11384 23000 11386
rect 16389 11328 16394 11384
rect 16450 11328 23000 11384
rect 16389 11326 23000 11328
rect 16389 11323 16455 11326
rect 22200 11296 23000 11326
rect 0 10978 800 11008
rect 4061 10978 4127 10981
rect 0 10976 4127 10978
rect 0 10920 4066 10976
rect 4122 10920 4127 10976
rect 0 10918 4127 10920
rect 0 10888 800 10918
rect 4061 10915 4127 10918
rect 20437 10978 20503 10981
rect 22200 10978 23000 11008
rect 20437 10976 23000 10978
rect 20437 10920 20442 10976
rect 20498 10920 23000 10976
rect 20437 10918 23000 10920
rect 20437 10915 20503 10918
rect 4409 10912 4729 10913
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 10847 4729 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 18270 10912 18590 10913
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 22200 10888 23000 10918
rect 18270 10847 18590 10848
rect 0 10434 800 10464
rect 4061 10434 4127 10437
rect 0 10432 4127 10434
rect 0 10376 4066 10432
rect 4122 10376 4127 10432
rect 0 10374 4127 10376
rect 0 10344 800 10374
rect 4061 10371 4127 10374
rect 18873 10434 18939 10437
rect 22200 10434 23000 10464
rect 18873 10432 23000 10434
rect 18873 10376 18878 10432
rect 18934 10376 23000 10432
rect 18873 10374 23000 10376
rect 18873 10371 18939 10374
rect 7874 10368 8194 10369
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8194 10368
rect 7874 10303 8194 10304
rect 14805 10368 15125 10369
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 22200 10344 23000 10374
rect 14805 10303 15125 10304
rect 0 10026 800 10056
rect 4061 10026 4127 10029
rect 0 10024 4127 10026
rect 0 9968 4066 10024
rect 4122 9968 4127 10024
rect 0 9966 4127 9968
rect 0 9936 800 9966
rect 4061 9963 4127 9966
rect 19057 10026 19123 10029
rect 22200 10026 23000 10056
rect 19057 10024 23000 10026
rect 19057 9968 19062 10024
rect 19118 9968 23000 10024
rect 19057 9966 23000 9968
rect 19057 9963 19123 9966
rect 22200 9936 23000 9966
rect 4409 9824 4729 9825
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 9759 4729 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 18270 9824 18590 9825
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 9759 18590 9760
rect 4245 9618 4311 9621
rect 10685 9618 10751 9621
rect 4245 9616 10751 9618
rect 4245 9560 4250 9616
rect 4306 9560 10690 9616
rect 10746 9560 10751 9616
rect 4245 9558 10751 9560
rect 4245 9555 4311 9558
rect 10685 9555 10751 9558
rect 18321 9618 18387 9621
rect 19793 9618 19859 9621
rect 18321 9616 19859 9618
rect 18321 9560 18326 9616
rect 18382 9560 19798 9616
rect 19854 9560 19859 9616
rect 18321 9558 19859 9560
rect 18321 9555 18387 9558
rect 19793 9555 19859 9558
rect 0 9482 800 9512
rect 5073 9482 5139 9485
rect 0 9480 5139 9482
rect 0 9424 5078 9480
rect 5134 9424 5139 9480
rect 0 9422 5139 9424
rect 0 9392 800 9422
rect 5073 9419 5139 9422
rect 18597 9482 18663 9485
rect 22200 9482 23000 9512
rect 18597 9480 23000 9482
rect 18597 9424 18602 9480
rect 18658 9424 23000 9480
rect 18597 9422 23000 9424
rect 18597 9419 18663 9422
rect 22200 9392 23000 9422
rect 7874 9280 8194 9281
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8194 9280
rect 7874 9215 8194 9216
rect 14805 9280 15125 9281
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 9215 15125 9216
rect 2037 9210 2103 9213
rect 6545 9210 6611 9213
rect 2037 9208 6611 9210
rect 2037 9152 2042 9208
rect 2098 9152 6550 9208
rect 6606 9152 6611 9208
rect 2037 9150 6611 9152
rect 2037 9147 2103 9150
rect 6545 9147 6611 9150
rect 0 9074 800 9104
rect 4061 9074 4127 9077
rect 0 9072 4127 9074
rect 0 9016 4066 9072
rect 4122 9016 4127 9072
rect 0 9014 4127 9016
rect 0 8984 800 9014
rect 4061 9011 4127 9014
rect 20529 9074 20595 9077
rect 22200 9074 23000 9104
rect 20529 9072 23000 9074
rect 20529 9016 20534 9072
rect 20590 9016 23000 9072
rect 20529 9014 23000 9016
rect 20529 9011 20595 9014
rect 22200 8984 23000 9014
rect 10041 8938 10107 8941
rect 11697 8938 11763 8941
rect 10041 8936 11763 8938
rect 10041 8880 10046 8936
rect 10102 8880 11702 8936
rect 11758 8880 11763 8936
rect 10041 8878 11763 8880
rect 10041 8875 10107 8878
rect 11697 8875 11763 8878
rect 17902 8876 17908 8940
rect 17972 8938 17978 8940
rect 17972 8878 18890 8938
rect 17972 8876 17978 8878
rect 18830 8802 18890 8878
rect 18830 8742 22202 8802
rect 4409 8736 4729 8737
rect 0 8666 800 8696
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 8671 4729 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 18270 8736 18590 8737
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 8671 18590 8672
rect 22142 8696 22202 8742
rect 4245 8666 4311 8669
rect 0 8664 4311 8666
rect 0 8608 4250 8664
rect 4306 8608 4311 8664
rect 0 8606 4311 8608
rect 22142 8606 23000 8696
rect 0 8576 800 8606
rect 4245 8603 4311 8606
rect 22200 8576 23000 8606
rect 12065 8530 12131 8533
rect 17902 8530 17908 8532
rect 12065 8528 17908 8530
rect 12065 8472 12070 8528
rect 12126 8472 17908 8528
rect 12065 8470 17908 8472
rect 12065 8467 12131 8470
rect 17902 8468 17908 8470
rect 17972 8468 17978 8532
rect 14181 8394 14247 8397
rect 16665 8394 16731 8397
rect 14181 8392 16731 8394
rect 14181 8336 14186 8392
rect 14242 8336 16670 8392
rect 16726 8336 16731 8392
rect 14181 8334 16731 8336
rect 14181 8331 14247 8334
rect 16665 8331 16731 8334
rect 3049 8258 3115 8261
rect 5533 8258 5599 8261
rect 3049 8256 5599 8258
rect 3049 8200 3054 8256
rect 3110 8200 5538 8256
rect 5594 8200 5599 8256
rect 3049 8198 5599 8200
rect 3049 8195 3115 8198
rect 5533 8195 5599 8198
rect 7874 8192 8194 8193
rect 0 8122 800 8152
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8194 8192
rect 7874 8127 8194 8128
rect 14805 8192 15125 8193
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 8127 15125 8128
rect 4061 8122 4127 8125
rect 0 8120 4127 8122
rect 0 8064 4066 8120
rect 4122 8064 4127 8120
rect 0 8062 4127 8064
rect 0 8032 800 8062
rect 4061 8059 4127 8062
rect 17769 8122 17835 8125
rect 22200 8122 23000 8152
rect 17769 8120 23000 8122
rect 17769 8064 17774 8120
rect 17830 8064 23000 8120
rect 17769 8062 23000 8064
rect 17769 8059 17835 8062
rect 22200 8032 23000 8062
rect 10593 7986 10659 7989
rect 17125 7986 17191 7989
rect 10593 7984 17191 7986
rect 10593 7928 10598 7984
rect 10654 7928 17130 7984
rect 17186 7928 17191 7984
rect 10593 7926 17191 7928
rect 10593 7923 10659 7926
rect 17125 7923 17191 7926
rect 19374 7924 19380 7988
rect 19444 7986 19450 7988
rect 20161 7986 20227 7989
rect 19444 7984 20227 7986
rect 19444 7928 20166 7984
rect 20222 7928 20227 7984
rect 19444 7926 20227 7928
rect 19444 7924 19450 7926
rect 20161 7923 20227 7926
rect 0 7714 800 7744
rect 3969 7714 4035 7717
rect 0 7712 4035 7714
rect 0 7656 3974 7712
rect 4030 7656 4035 7712
rect 0 7654 4035 7656
rect 0 7624 800 7654
rect 3969 7651 4035 7654
rect 19149 7714 19215 7717
rect 22200 7714 23000 7744
rect 19149 7712 23000 7714
rect 19149 7656 19154 7712
rect 19210 7656 23000 7712
rect 19149 7654 23000 7656
rect 19149 7651 19215 7654
rect 4409 7648 4729 7649
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 7583 4729 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 18270 7648 18590 7649
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 22200 7624 23000 7654
rect 18270 7583 18590 7584
rect 10777 7442 10843 7445
rect 14825 7442 14891 7445
rect 10777 7440 14891 7442
rect 10777 7384 10782 7440
rect 10838 7384 14830 7440
rect 14886 7384 14891 7440
rect 10777 7382 14891 7384
rect 10777 7379 10843 7382
rect 14825 7379 14891 7382
rect 0 7170 800 7200
rect 1393 7170 1459 7173
rect 0 7168 1459 7170
rect 0 7112 1398 7168
rect 1454 7112 1459 7168
rect 0 7110 1459 7112
rect 0 7080 800 7110
rect 1393 7107 1459 7110
rect 19241 7170 19307 7173
rect 22200 7170 23000 7200
rect 19241 7168 23000 7170
rect 19241 7112 19246 7168
rect 19302 7112 23000 7168
rect 19241 7110 23000 7112
rect 19241 7107 19307 7110
rect 7874 7104 8194 7105
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8194 7104
rect 7874 7039 8194 7040
rect 14805 7104 15125 7105
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 22200 7080 23000 7110
rect 14805 7039 15125 7040
rect 10317 6898 10383 6901
rect 10317 6896 12082 6898
rect 10317 6840 10322 6896
rect 10378 6840 12082 6896
rect 10317 6838 12082 6840
rect 10317 6835 10383 6838
rect 0 6762 800 6792
rect 3969 6762 4035 6765
rect 0 6760 4035 6762
rect 0 6704 3974 6760
rect 4030 6704 4035 6760
rect 0 6702 4035 6704
rect 0 6672 800 6702
rect 3969 6699 4035 6702
rect 8109 6762 8175 6765
rect 11789 6762 11855 6765
rect 8109 6760 11855 6762
rect 8109 6704 8114 6760
rect 8170 6704 11794 6760
rect 11850 6704 11855 6760
rect 8109 6702 11855 6704
rect 12022 6762 12082 6838
rect 22200 6762 23000 6792
rect 12022 6702 23000 6762
rect 8109 6699 8175 6702
rect 11789 6699 11855 6702
rect 22200 6672 23000 6702
rect 4409 6560 4729 6561
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 6495 4729 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 18270 6560 18590 6561
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 18270 6495 18590 6496
rect 3141 6354 3207 6357
rect 19374 6354 19380 6356
rect 3006 6352 19380 6354
rect 3006 6296 3146 6352
rect 3202 6296 19380 6352
rect 3006 6294 19380 6296
rect 0 6218 800 6248
rect 3006 6218 3066 6294
rect 3141 6291 3207 6294
rect 19374 6292 19380 6294
rect 19444 6292 19450 6356
rect 0 6158 3066 6218
rect 4153 6218 4219 6221
rect 19333 6218 19399 6221
rect 4153 6216 8402 6218
rect 4153 6160 4158 6216
rect 4214 6160 8402 6216
rect 4153 6158 8402 6160
rect 0 6128 800 6158
rect 4153 6155 4219 6158
rect 5214 6085 5274 6158
rect 5165 6080 5274 6085
rect 5165 6024 5170 6080
rect 5226 6024 5274 6080
rect 5165 6022 5274 6024
rect 8342 6082 8402 6158
rect 14414 6216 19399 6218
rect 14414 6160 19338 6216
rect 19394 6160 19399 6216
rect 14414 6158 19399 6160
rect 14414 6082 14474 6158
rect 19333 6155 19399 6158
rect 19793 6218 19859 6221
rect 22200 6218 23000 6248
rect 19793 6216 23000 6218
rect 19793 6160 19798 6216
rect 19854 6160 23000 6216
rect 19793 6158 23000 6160
rect 19793 6155 19859 6158
rect 22200 6128 23000 6158
rect 8342 6022 14474 6082
rect 5165 6019 5231 6022
rect 7874 6016 8194 6017
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8194 6016
rect 7874 5951 8194 5952
rect 14805 6016 15125 6017
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 5951 15125 5952
rect 0 5810 800 5840
rect 3877 5810 3943 5813
rect 0 5808 3943 5810
rect 0 5752 3882 5808
rect 3938 5752 3943 5808
rect 0 5750 3943 5752
rect 0 5720 800 5750
rect 3877 5747 3943 5750
rect 7465 5810 7531 5813
rect 12525 5810 12591 5813
rect 7465 5808 12591 5810
rect 7465 5752 7470 5808
rect 7526 5752 12530 5808
rect 12586 5752 12591 5808
rect 7465 5750 12591 5752
rect 7465 5747 7531 5750
rect 12525 5747 12591 5750
rect 17953 5810 18019 5813
rect 22200 5810 23000 5840
rect 17953 5808 23000 5810
rect 17953 5752 17958 5808
rect 18014 5752 23000 5808
rect 17953 5750 23000 5752
rect 17953 5747 18019 5750
rect 22200 5720 23000 5750
rect 9305 5674 9371 5677
rect 21357 5674 21423 5677
rect 9305 5672 21423 5674
rect 9305 5616 9310 5672
rect 9366 5616 21362 5672
rect 21418 5616 21423 5672
rect 9305 5614 21423 5616
rect 9305 5611 9371 5614
rect 21357 5611 21423 5614
rect 4409 5472 4729 5473
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 5407 4729 5408
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 18270 5472 18590 5473
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 5407 18590 5408
rect 0 5266 800 5296
rect 3969 5266 4035 5269
rect 0 5264 4035 5266
rect 0 5208 3974 5264
rect 4030 5208 4035 5264
rect 0 5206 4035 5208
rect 0 5176 800 5206
rect 3969 5203 4035 5206
rect 20621 5266 20687 5269
rect 22200 5266 23000 5296
rect 20621 5264 23000 5266
rect 20621 5208 20626 5264
rect 20682 5208 23000 5264
rect 20621 5206 23000 5208
rect 20621 5203 20687 5206
rect 22200 5176 23000 5206
rect 7874 4928 8194 4929
rect 0 4858 800 4888
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8194 4928
rect 7874 4863 8194 4864
rect 14805 4928 15125 4929
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 4863 15125 4864
rect 3877 4858 3943 4861
rect 0 4856 3943 4858
rect 0 4800 3882 4856
rect 3938 4800 3943 4856
rect 0 4798 3943 4800
rect 0 4768 800 4798
rect 3877 4795 3943 4798
rect 17953 4858 18019 4861
rect 22200 4858 23000 4888
rect 17953 4856 23000 4858
rect 17953 4800 17958 4856
rect 18014 4800 23000 4856
rect 17953 4798 23000 4800
rect 17953 4795 18019 4798
rect 22200 4768 23000 4798
rect 0 4450 800 4480
rect 4061 4450 4127 4453
rect 0 4448 4127 4450
rect 0 4392 4066 4448
rect 4122 4392 4127 4448
rect 0 4390 4127 4392
rect 0 4360 800 4390
rect 4061 4387 4127 4390
rect 21265 4450 21331 4453
rect 22200 4450 23000 4480
rect 21265 4448 23000 4450
rect 21265 4392 21270 4448
rect 21326 4392 23000 4448
rect 21265 4390 23000 4392
rect 21265 4387 21331 4390
rect 4409 4384 4729 4385
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 4319 4729 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 18270 4384 18590 4385
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 22200 4360 23000 4390
rect 18270 4319 18590 4320
rect 0 3906 800 3936
rect 3877 3906 3943 3909
rect 0 3904 3943 3906
rect 0 3848 3882 3904
rect 3938 3848 3943 3904
rect 0 3846 3943 3848
rect 0 3816 800 3846
rect 3877 3843 3943 3846
rect 20621 3906 20687 3909
rect 22200 3906 23000 3936
rect 20621 3904 23000 3906
rect 20621 3848 20626 3904
rect 20682 3848 23000 3904
rect 20621 3846 23000 3848
rect 20621 3843 20687 3846
rect 7874 3840 8194 3841
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8194 3840
rect 7874 3775 8194 3776
rect 14805 3840 15125 3841
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 22200 3816 23000 3846
rect 14805 3775 15125 3776
rect 1945 3634 2011 3637
rect 4153 3634 4219 3637
rect 1945 3632 4219 3634
rect 1945 3576 1950 3632
rect 2006 3576 4158 3632
rect 4214 3576 4219 3632
rect 1945 3574 4219 3576
rect 1945 3571 2011 3574
rect 4153 3571 4219 3574
rect 0 3498 800 3528
rect 2037 3498 2103 3501
rect 0 3496 2103 3498
rect 0 3440 2042 3496
rect 2098 3440 2103 3496
rect 0 3438 2103 3440
rect 0 3408 800 3438
rect 2037 3435 2103 3438
rect 17401 3498 17467 3501
rect 22200 3498 23000 3528
rect 17401 3496 23000 3498
rect 17401 3440 17406 3496
rect 17462 3440 23000 3496
rect 17401 3438 23000 3440
rect 17401 3435 17467 3438
rect 22200 3408 23000 3438
rect 4409 3296 4729 3297
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 3231 4729 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 18270 3296 18590 3297
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 18270 3231 18590 3232
rect 0 2954 800 2984
rect 3693 2954 3759 2957
rect 0 2952 3759 2954
rect 0 2896 3698 2952
rect 3754 2896 3759 2952
rect 0 2894 3759 2896
rect 0 2864 800 2894
rect 3693 2891 3759 2894
rect 18689 2954 18755 2957
rect 22200 2954 23000 2984
rect 18689 2952 23000 2954
rect 18689 2896 18694 2952
rect 18750 2896 23000 2952
rect 18689 2894 23000 2896
rect 18689 2891 18755 2894
rect 22200 2864 23000 2894
rect 7874 2752 8194 2753
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8194 2752
rect 7874 2687 8194 2688
rect 14805 2752 15125 2753
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2687 15125 2688
rect 0 2546 800 2576
rect 1669 2546 1735 2549
rect 0 2544 1735 2546
rect 0 2488 1674 2544
rect 1730 2488 1735 2544
rect 0 2486 1735 2488
rect 0 2456 800 2486
rect 1669 2483 1735 2486
rect 18781 2546 18847 2549
rect 22200 2546 23000 2576
rect 18781 2544 23000 2546
rect 18781 2488 18786 2544
rect 18842 2488 23000 2544
rect 18781 2486 23000 2488
rect 18781 2483 18847 2486
rect 22200 2456 23000 2486
rect 4409 2208 4729 2209
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2143 4729 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 18270 2208 18590 2209
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2143 18590 2144
rect 0 2002 800 2032
rect 3601 2002 3667 2005
rect 0 2000 3667 2002
rect 0 1944 3606 2000
rect 3662 1944 3667 2000
rect 0 1942 3667 1944
rect 0 1912 800 1942
rect 3601 1939 3667 1942
rect 20069 2002 20135 2005
rect 22200 2002 23000 2032
rect 20069 2000 23000 2002
rect 20069 1944 20074 2000
rect 20130 1944 23000 2000
rect 20069 1942 23000 1944
rect 20069 1939 20135 1942
rect 22200 1912 23000 1942
rect 0 1594 800 1624
rect 1301 1594 1367 1597
rect 0 1592 1367 1594
rect 0 1536 1306 1592
rect 1362 1536 1367 1592
rect 0 1534 1367 1536
rect 0 1504 800 1534
rect 1301 1531 1367 1534
rect 21173 1594 21239 1597
rect 22200 1594 23000 1624
rect 21173 1592 23000 1594
rect 21173 1536 21178 1592
rect 21234 1536 23000 1592
rect 21173 1534 23000 1536
rect 21173 1531 21239 1534
rect 22200 1504 23000 1534
rect 0 1050 800 1080
rect 3969 1050 4035 1053
rect 0 1048 4035 1050
rect 0 992 3974 1048
rect 4030 992 4035 1048
rect 0 990 4035 992
rect 0 960 800 990
rect 3969 987 4035 990
rect 19241 1050 19307 1053
rect 22200 1050 23000 1080
rect 19241 1048 23000 1050
rect 19241 992 19246 1048
rect 19302 992 23000 1048
rect 19241 990 23000 992
rect 19241 987 19307 990
rect 22200 960 23000 990
rect 0 642 800 672
rect 2313 642 2379 645
rect 0 640 2379 642
rect 0 584 2318 640
rect 2374 584 2379 640
rect 0 582 2379 584
rect 0 552 800 582
rect 2313 579 2379 582
rect 16941 642 17007 645
rect 22200 642 23000 672
rect 16941 640 23000 642
rect 16941 584 16946 640
rect 17002 584 23000 640
rect 16941 582 23000 584
rect 16941 579 17007 582
rect 22200 552 23000 582
rect 0 234 800 264
rect 6361 234 6427 237
rect 0 232 6427 234
rect 0 176 6366 232
rect 6422 176 6427 232
rect 0 174 6427 176
rect 0 144 800 174
rect 6361 171 6427 174
rect 18965 234 19031 237
rect 22200 234 23000 264
rect 18965 232 23000 234
rect 18965 176 18970 232
rect 19026 176 23000 232
rect 18965 174 23000 176
rect 18965 171 19031 174
rect 22200 144 23000 174
<< via3 >>
rect 4417 20700 4481 20704
rect 4417 20644 4421 20700
rect 4421 20644 4477 20700
rect 4477 20644 4481 20700
rect 4417 20640 4481 20644
rect 4497 20700 4561 20704
rect 4497 20644 4501 20700
rect 4501 20644 4557 20700
rect 4557 20644 4561 20700
rect 4497 20640 4561 20644
rect 4577 20700 4641 20704
rect 4577 20644 4581 20700
rect 4581 20644 4637 20700
rect 4637 20644 4641 20700
rect 4577 20640 4641 20644
rect 4657 20700 4721 20704
rect 4657 20644 4661 20700
rect 4661 20644 4717 20700
rect 4717 20644 4721 20700
rect 4657 20640 4721 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 18278 20700 18342 20704
rect 18278 20644 18282 20700
rect 18282 20644 18338 20700
rect 18338 20644 18342 20700
rect 18278 20640 18342 20644
rect 18358 20700 18422 20704
rect 18358 20644 18362 20700
rect 18362 20644 18418 20700
rect 18418 20644 18422 20700
rect 18358 20640 18422 20644
rect 18438 20700 18502 20704
rect 18438 20644 18442 20700
rect 18442 20644 18498 20700
rect 18498 20644 18502 20700
rect 18438 20640 18502 20644
rect 18518 20700 18582 20704
rect 18518 20644 18522 20700
rect 18522 20644 18578 20700
rect 18578 20644 18582 20700
rect 18518 20640 18582 20644
rect 7882 20156 7946 20160
rect 7882 20100 7886 20156
rect 7886 20100 7942 20156
rect 7942 20100 7946 20156
rect 7882 20096 7946 20100
rect 7962 20156 8026 20160
rect 7962 20100 7966 20156
rect 7966 20100 8022 20156
rect 8022 20100 8026 20156
rect 7962 20096 8026 20100
rect 8042 20156 8106 20160
rect 8042 20100 8046 20156
rect 8046 20100 8102 20156
rect 8102 20100 8106 20156
rect 8042 20096 8106 20100
rect 8122 20156 8186 20160
rect 8122 20100 8126 20156
rect 8126 20100 8182 20156
rect 8182 20100 8186 20156
rect 8122 20096 8186 20100
rect 14813 20156 14877 20160
rect 14813 20100 14817 20156
rect 14817 20100 14873 20156
rect 14873 20100 14877 20156
rect 14813 20096 14877 20100
rect 14893 20156 14957 20160
rect 14893 20100 14897 20156
rect 14897 20100 14953 20156
rect 14953 20100 14957 20156
rect 14893 20096 14957 20100
rect 14973 20156 15037 20160
rect 14973 20100 14977 20156
rect 14977 20100 15033 20156
rect 15033 20100 15037 20156
rect 14973 20096 15037 20100
rect 15053 20156 15117 20160
rect 15053 20100 15057 20156
rect 15057 20100 15113 20156
rect 15113 20100 15117 20156
rect 15053 20096 15117 20100
rect 4417 19612 4481 19616
rect 4417 19556 4421 19612
rect 4421 19556 4477 19612
rect 4477 19556 4481 19612
rect 4417 19552 4481 19556
rect 4497 19612 4561 19616
rect 4497 19556 4501 19612
rect 4501 19556 4557 19612
rect 4557 19556 4561 19612
rect 4497 19552 4561 19556
rect 4577 19612 4641 19616
rect 4577 19556 4581 19612
rect 4581 19556 4637 19612
rect 4637 19556 4641 19612
rect 4577 19552 4641 19556
rect 4657 19612 4721 19616
rect 4657 19556 4661 19612
rect 4661 19556 4717 19612
rect 4717 19556 4721 19612
rect 4657 19552 4721 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 18278 19612 18342 19616
rect 18278 19556 18282 19612
rect 18282 19556 18338 19612
rect 18338 19556 18342 19612
rect 18278 19552 18342 19556
rect 18358 19612 18422 19616
rect 18358 19556 18362 19612
rect 18362 19556 18418 19612
rect 18418 19556 18422 19612
rect 18358 19552 18422 19556
rect 18438 19612 18502 19616
rect 18438 19556 18442 19612
rect 18442 19556 18498 19612
rect 18498 19556 18502 19612
rect 18438 19552 18502 19556
rect 18518 19612 18582 19616
rect 18518 19556 18522 19612
rect 18522 19556 18578 19612
rect 18578 19556 18582 19612
rect 18518 19552 18582 19556
rect 7882 19068 7946 19072
rect 7882 19012 7886 19068
rect 7886 19012 7942 19068
rect 7942 19012 7946 19068
rect 7882 19008 7946 19012
rect 7962 19068 8026 19072
rect 7962 19012 7966 19068
rect 7966 19012 8022 19068
rect 8022 19012 8026 19068
rect 7962 19008 8026 19012
rect 8042 19068 8106 19072
rect 8042 19012 8046 19068
rect 8046 19012 8102 19068
rect 8102 19012 8106 19068
rect 8042 19008 8106 19012
rect 8122 19068 8186 19072
rect 8122 19012 8126 19068
rect 8126 19012 8182 19068
rect 8182 19012 8186 19068
rect 8122 19008 8186 19012
rect 14813 19068 14877 19072
rect 14813 19012 14817 19068
rect 14817 19012 14873 19068
rect 14873 19012 14877 19068
rect 14813 19008 14877 19012
rect 14893 19068 14957 19072
rect 14893 19012 14897 19068
rect 14897 19012 14953 19068
rect 14953 19012 14957 19068
rect 14893 19008 14957 19012
rect 14973 19068 15037 19072
rect 14973 19012 14977 19068
rect 14977 19012 15033 19068
rect 15033 19012 15037 19068
rect 14973 19008 15037 19012
rect 15053 19068 15117 19072
rect 15053 19012 15057 19068
rect 15057 19012 15113 19068
rect 15113 19012 15117 19068
rect 15053 19008 15117 19012
rect 4417 18524 4481 18528
rect 4417 18468 4421 18524
rect 4421 18468 4477 18524
rect 4477 18468 4481 18524
rect 4417 18464 4481 18468
rect 4497 18524 4561 18528
rect 4497 18468 4501 18524
rect 4501 18468 4557 18524
rect 4557 18468 4561 18524
rect 4497 18464 4561 18468
rect 4577 18524 4641 18528
rect 4577 18468 4581 18524
rect 4581 18468 4637 18524
rect 4637 18468 4641 18524
rect 4577 18464 4641 18468
rect 4657 18524 4721 18528
rect 4657 18468 4661 18524
rect 4661 18468 4717 18524
rect 4717 18468 4721 18524
rect 4657 18464 4721 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 18278 18524 18342 18528
rect 18278 18468 18282 18524
rect 18282 18468 18338 18524
rect 18338 18468 18342 18524
rect 18278 18464 18342 18468
rect 18358 18524 18422 18528
rect 18358 18468 18362 18524
rect 18362 18468 18418 18524
rect 18418 18468 18422 18524
rect 18358 18464 18422 18468
rect 18438 18524 18502 18528
rect 18438 18468 18442 18524
rect 18442 18468 18498 18524
rect 18498 18468 18502 18524
rect 18438 18464 18502 18468
rect 18518 18524 18582 18528
rect 18518 18468 18522 18524
rect 18522 18468 18578 18524
rect 18578 18468 18582 18524
rect 18518 18464 18582 18468
rect 7882 17980 7946 17984
rect 7882 17924 7886 17980
rect 7886 17924 7942 17980
rect 7942 17924 7946 17980
rect 7882 17920 7946 17924
rect 7962 17980 8026 17984
rect 7962 17924 7966 17980
rect 7966 17924 8022 17980
rect 8022 17924 8026 17980
rect 7962 17920 8026 17924
rect 8042 17980 8106 17984
rect 8042 17924 8046 17980
rect 8046 17924 8102 17980
rect 8102 17924 8106 17980
rect 8042 17920 8106 17924
rect 8122 17980 8186 17984
rect 8122 17924 8126 17980
rect 8126 17924 8182 17980
rect 8182 17924 8186 17980
rect 8122 17920 8186 17924
rect 14813 17980 14877 17984
rect 14813 17924 14817 17980
rect 14817 17924 14873 17980
rect 14873 17924 14877 17980
rect 14813 17920 14877 17924
rect 14893 17980 14957 17984
rect 14893 17924 14897 17980
rect 14897 17924 14953 17980
rect 14953 17924 14957 17980
rect 14893 17920 14957 17924
rect 14973 17980 15037 17984
rect 14973 17924 14977 17980
rect 14977 17924 15033 17980
rect 15033 17924 15037 17980
rect 14973 17920 15037 17924
rect 15053 17980 15117 17984
rect 15053 17924 15057 17980
rect 15057 17924 15113 17980
rect 15113 17924 15117 17980
rect 15053 17920 15117 17924
rect 4417 17436 4481 17440
rect 4417 17380 4421 17436
rect 4421 17380 4477 17436
rect 4477 17380 4481 17436
rect 4417 17376 4481 17380
rect 4497 17436 4561 17440
rect 4497 17380 4501 17436
rect 4501 17380 4557 17436
rect 4557 17380 4561 17436
rect 4497 17376 4561 17380
rect 4577 17436 4641 17440
rect 4577 17380 4581 17436
rect 4581 17380 4637 17436
rect 4637 17380 4641 17436
rect 4577 17376 4641 17380
rect 4657 17436 4721 17440
rect 4657 17380 4661 17436
rect 4661 17380 4717 17436
rect 4717 17380 4721 17436
rect 4657 17376 4721 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 18278 17436 18342 17440
rect 18278 17380 18282 17436
rect 18282 17380 18338 17436
rect 18338 17380 18342 17436
rect 18278 17376 18342 17380
rect 18358 17436 18422 17440
rect 18358 17380 18362 17436
rect 18362 17380 18418 17436
rect 18418 17380 18422 17436
rect 18358 17376 18422 17380
rect 18438 17436 18502 17440
rect 18438 17380 18442 17436
rect 18442 17380 18498 17436
rect 18498 17380 18502 17436
rect 18438 17376 18502 17380
rect 18518 17436 18582 17440
rect 18518 17380 18522 17436
rect 18522 17380 18578 17436
rect 18578 17380 18582 17436
rect 18518 17376 18582 17380
rect 7882 16892 7946 16896
rect 7882 16836 7886 16892
rect 7886 16836 7942 16892
rect 7942 16836 7946 16892
rect 7882 16832 7946 16836
rect 7962 16892 8026 16896
rect 7962 16836 7966 16892
rect 7966 16836 8022 16892
rect 8022 16836 8026 16892
rect 7962 16832 8026 16836
rect 8042 16892 8106 16896
rect 8042 16836 8046 16892
rect 8046 16836 8102 16892
rect 8102 16836 8106 16892
rect 8042 16832 8106 16836
rect 8122 16892 8186 16896
rect 8122 16836 8126 16892
rect 8126 16836 8182 16892
rect 8182 16836 8186 16892
rect 8122 16832 8186 16836
rect 14813 16892 14877 16896
rect 14813 16836 14817 16892
rect 14817 16836 14873 16892
rect 14873 16836 14877 16892
rect 14813 16832 14877 16836
rect 14893 16892 14957 16896
rect 14893 16836 14897 16892
rect 14897 16836 14953 16892
rect 14953 16836 14957 16892
rect 14893 16832 14957 16836
rect 14973 16892 15037 16896
rect 14973 16836 14977 16892
rect 14977 16836 15033 16892
rect 15033 16836 15037 16892
rect 14973 16832 15037 16836
rect 15053 16892 15117 16896
rect 15053 16836 15057 16892
rect 15057 16836 15113 16892
rect 15113 16836 15117 16892
rect 15053 16832 15117 16836
rect 4417 16348 4481 16352
rect 4417 16292 4421 16348
rect 4421 16292 4477 16348
rect 4477 16292 4481 16348
rect 4417 16288 4481 16292
rect 4497 16348 4561 16352
rect 4497 16292 4501 16348
rect 4501 16292 4557 16348
rect 4557 16292 4561 16348
rect 4497 16288 4561 16292
rect 4577 16348 4641 16352
rect 4577 16292 4581 16348
rect 4581 16292 4637 16348
rect 4637 16292 4641 16348
rect 4577 16288 4641 16292
rect 4657 16348 4721 16352
rect 4657 16292 4661 16348
rect 4661 16292 4717 16348
rect 4717 16292 4721 16348
rect 4657 16288 4721 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 18278 16348 18342 16352
rect 18278 16292 18282 16348
rect 18282 16292 18338 16348
rect 18338 16292 18342 16348
rect 18278 16288 18342 16292
rect 18358 16348 18422 16352
rect 18358 16292 18362 16348
rect 18362 16292 18418 16348
rect 18418 16292 18422 16348
rect 18358 16288 18422 16292
rect 18438 16348 18502 16352
rect 18438 16292 18442 16348
rect 18442 16292 18498 16348
rect 18498 16292 18502 16348
rect 18438 16288 18502 16292
rect 18518 16348 18582 16352
rect 18518 16292 18522 16348
rect 18522 16292 18578 16348
rect 18578 16292 18582 16348
rect 18518 16288 18582 16292
rect 7882 15804 7946 15808
rect 7882 15748 7886 15804
rect 7886 15748 7942 15804
rect 7942 15748 7946 15804
rect 7882 15744 7946 15748
rect 7962 15804 8026 15808
rect 7962 15748 7966 15804
rect 7966 15748 8022 15804
rect 8022 15748 8026 15804
rect 7962 15744 8026 15748
rect 8042 15804 8106 15808
rect 8042 15748 8046 15804
rect 8046 15748 8102 15804
rect 8102 15748 8106 15804
rect 8042 15744 8106 15748
rect 8122 15804 8186 15808
rect 8122 15748 8126 15804
rect 8126 15748 8182 15804
rect 8182 15748 8186 15804
rect 8122 15744 8186 15748
rect 14813 15804 14877 15808
rect 14813 15748 14817 15804
rect 14817 15748 14873 15804
rect 14873 15748 14877 15804
rect 14813 15744 14877 15748
rect 14893 15804 14957 15808
rect 14893 15748 14897 15804
rect 14897 15748 14953 15804
rect 14953 15748 14957 15804
rect 14893 15744 14957 15748
rect 14973 15804 15037 15808
rect 14973 15748 14977 15804
rect 14977 15748 15033 15804
rect 15033 15748 15037 15804
rect 14973 15744 15037 15748
rect 15053 15804 15117 15808
rect 15053 15748 15057 15804
rect 15057 15748 15113 15804
rect 15113 15748 15117 15804
rect 15053 15744 15117 15748
rect 4417 15260 4481 15264
rect 4417 15204 4421 15260
rect 4421 15204 4477 15260
rect 4477 15204 4481 15260
rect 4417 15200 4481 15204
rect 4497 15260 4561 15264
rect 4497 15204 4501 15260
rect 4501 15204 4557 15260
rect 4557 15204 4561 15260
rect 4497 15200 4561 15204
rect 4577 15260 4641 15264
rect 4577 15204 4581 15260
rect 4581 15204 4637 15260
rect 4637 15204 4641 15260
rect 4577 15200 4641 15204
rect 4657 15260 4721 15264
rect 4657 15204 4661 15260
rect 4661 15204 4717 15260
rect 4717 15204 4721 15260
rect 4657 15200 4721 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 18278 15260 18342 15264
rect 18278 15204 18282 15260
rect 18282 15204 18338 15260
rect 18338 15204 18342 15260
rect 18278 15200 18342 15204
rect 18358 15260 18422 15264
rect 18358 15204 18362 15260
rect 18362 15204 18418 15260
rect 18418 15204 18422 15260
rect 18358 15200 18422 15204
rect 18438 15260 18502 15264
rect 18438 15204 18442 15260
rect 18442 15204 18498 15260
rect 18498 15204 18502 15260
rect 18438 15200 18502 15204
rect 18518 15260 18582 15264
rect 18518 15204 18522 15260
rect 18522 15204 18578 15260
rect 18578 15204 18582 15260
rect 18518 15200 18582 15204
rect 7882 14716 7946 14720
rect 7882 14660 7886 14716
rect 7886 14660 7942 14716
rect 7942 14660 7946 14716
rect 7882 14656 7946 14660
rect 7962 14716 8026 14720
rect 7962 14660 7966 14716
rect 7966 14660 8022 14716
rect 8022 14660 8026 14716
rect 7962 14656 8026 14660
rect 8042 14716 8106 14720
rect 8042 14660 8046 14716
rect 8046 14660 8102 14716
rect 8102 14660 8106 14716
rect 8042 14656 8106 14660
rect 8122 14716 8186 14720
rect 8122 14660 8126 14716
rect 8126 14660 8182 14716
rect 8182 14660 8186 14716
rect 8122 14656 8186 14660
rect 14813 14716 14877 14720
rect 14813 14660 14817 14716
rect 14817 14660 14873 14716
rect 14873 14660 14877 14716
rect 14813 14656 14877 14660
rect 14893 14716 14957 14720
rect 14893 14660 14897 14716
rect 14897 14660 14953 14716
rect 14953 14660 14957 14716
rect 14893 14656 14957 14660
rect 14973 14716 15037 14720
rect 14973 14660 14977 14716
rect 14977 14660 15033 14716
rect 15033 14660 15037 14716
rect 14973 14656 15037 14660
rect 15053 14716 15117 14720
rect 15053 14660 15057 14716
rect 15057 14660 15113 14716
rect 15113 14660 15117 14716
rect 15053 14656 15117 14660
rect 4417 14172 4481 14176
rect 4417 14116 4421 14172
rect 4421 14116 4477 14172
rect 4477 14116 4481 14172
rect 4417 14112 4481 14116
rect 4497 14172 4561 14176
rect 4497 14116 4501 14172
rect 4501 14116 4557 14172
rect 4557 14116 4561 14172
rect 4497 14112 4561 14116
rect 4577 14172 4641 14176
rect 4577 14116 4581 14172
rect 4581 14116 4637 14172
rect 4637 14116 4641 14172
rect 4577 14112 4641 14116
rect 4657 14172 4721 14176
rect 4657 14116 4661 14172
rect 4661 14116 4717 14172
rect 4717 14116 4721 14172
rect 4657 14112 4721 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 18278 14172 18342 14176
rect 18278 14116 18282 14172
rect 18282 14116 18338 14172
rect 18338 14116 18342 14172
rect 18278 14112 18342 14116
rect 18358 14172 18422 14176
rect 18358 14116 18362 14172
rect 18362 14116 18418 14172
rect 18418 14116 18422 14172
rect 18358 14112 18422 14116
rect 18438 14172 18502 14176
rect 18438 14116 18442 14172
rect 18442 14116 18498 14172
rect 18498 14116 18502 14172
rect 18438 14112 18502 14116
rect 18518 14172 18582 14176
rect 18518 14116 18522 14172
rect 18522 14116 18578 14172
rect 18578 14116 18582 14172
rect 18518 14112 18582 14116
rect 7882 13628 7946 13632
rect 7882 13572 7886 13628
rect 7886 13572 7942 13628
rect 7942 13572 7946 13628
rect 7882 13568 7946 13572
rect 7962 13628 8026 13632
rect 7962 13572 7966 13628
rect 7966 13572 8022 13628
rect 8022 13572 8026 13628
rect 7962 13568 8026 13572
rect 8042 13628 8106 13632
rect 8042 13572 8046 13628
rect 8046 13572 8102 13628
rect 8102 13572 8106 13628
rect 8042 13568 8106 13572
rect 8122 13628 8186 13632
rect 8122 13572 8126 13628
rect 8126 13572 8182 13628
rect 8182 13572 8186 13628
rect 8122 13568 8186 13572
rect 14813 13628 14877 13632
rect 14813 13572 14817 13628
rect 14817 13572 14873 13628
rect 14873 13572 14877 13628
rect 14813 13568 14877 13572
rect 14893 13628 14957 13632
rect 14893 13572 14897 13628
rect 14897 13572 14953 13628
rect 14953 13572 14957 13628
rect 14893 13568 14957 13572
rect 14973 13628 15037 13632
rect 14973 13572 14977 13628
rect 14977 13572 15033 13628
rect 15033 13572 15037 13628
rect 14973 13568 15037 13572
rect 15053 13628 15117 13632
rect 15053 13572 15057 13628
rect 15057 13572 15113 13628
rect 15113 13572 15117 13628
rect 15053 13568 15117 13572
rect 4417 13084 4481 13088
rect 4417 13028 4421 13084
rect 4421 13028 4477 13084
rect 4477 13028 4481 13084
rect 4417 13024 4481 13028
rect 4497 13084 4561 13088
rect 4497 13028 4501 13084
rect 4501 13028 4557 13084
rect 4557 13028 4561 13084
rect 4497 13024 4561 13028
rect 4577 13084 4641 13088
rect 4577 13028 4581 13084
rect 4581 13028 4637 13084
rect 4637 13028 4641 13084
rect 4577 13024 4641 13028
rect 4657 13084 4721 13088
rect 4657 13028 4661 13084
rect 4661 13028 4717 13084
rect 4717 13028 4721 13084
rect 4657 13024 4721 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 18278 13084 18342 13088
rect 18278 13028 18282 13084
rect 18282 13028 18338 13084
rect 18338 13028 18342 13084
rect 18278 13024 18342 13028
rect 18358 13084 18422 13088
rect 18358 13028 18362 13084
rect 18362 13028 18418 13084
rect 18418 13028 18422 13084
rect 18358 13024 18422 13028
rect 18438 13084 18502 13088
rect 18438 13028 18442 13084
rect 18442 13028 18498 13084
rect 18498 13028 18502 13084
rect 18438 13024 18502 13028
rect 18518 13084 18582 13088
rect 18518 13028 18522 13084
rect 18522 13028 18578 13084
rect 18578 13028 18582 13084
rect 18518 13024 18582 13028
rect 7882 12540 7946 12544
rect 7882 12484 7886 12540
rect 7886 12484 7942 12540
rect 7942 12484 7946 12540
rect 7882 12480 7946 12484
rect 7962 12540 8026 12544
rect 7962 12484 7966 12540
rect 7966 12484 8022 12540
rect 8022 12484 8026 12540
rect 7962 12480 8026 12484
rect 8042 12540 8106 12544
rect 8042 12484 8046 12540
rect 8046 12484 8102 12540
rect 8102 12484 8106 12540
rect 8042 12480 8106 12484
rect 8122 12540 8186 12544
rect 8122 12484 8126 12540
rect 8126 12484 8182 12540
rect 8182 12484 8186 12540
rect 8122 12480 8186 12484
rect 14813 12540 14877 12544
rect 14813 12484 14817 12540
rect 14817 12484 14873 12540
rect 14873 12484 14877 12540
rect 14813 12480 14877 12484
rect 14893 12540 14957 12544
rect 14893 12484 14897 12540
rect 14897 12484 14953 12540
rect 14953 12484 14957 12540
rect 14893 12480 14957 12484
rect 14973 12540 15037 12544
rect 14973 12484 14977 12540
rect 14977 12484 15033 12540
rect 15033 12484 15037 12540
rect 14973 12480 15037 12484
rect 15053 12540 15117 12544
rect 15053 12484 15057 12540
rect 15057 12484 15113 12540
rect 15113 12484 15117 12540
rect 15053 12480 15117 12484
rect 4417 11996 4481 12000
rect 4417 11940 4421 11996
rect 4421 11940 4477 11996
rect 4477 11940 4481 11996
rect 4417 11936 4481 11940
rect 4497 11996 4561 12000
rect 4497 11940 4501 11996
rect 4501 11940 4557 11996
rect 4557 11940 4561 11996
rect 4497 11936 4561 11940
rect 4577 11996 4641 12000
rect 4577 11940 4581 11996
rect 4581 11940 4637 11996
rect 4637 11940 4641 11996
rect 4577 11936 4641 11940
rect 4657 11996 4721 12000
rect 4657 11940 4661 11996
rect 4661 11940 4717 11996
rect 4717 11940 4721 11996
rect 4657 11936 4721 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 18278 11996 18342 12000
rect 18278 11940 18282 11996
rect 18282 11940 18338 11996
rect 18338 11940 18342 11996
rect 18278 11936 18342 11940
rect 18358 11996 18422 12000
rect 18358 11940 18362 11996
rect 18362 11940 18418 11996
rect 18418 11940 18422 11996
rect 18358 11936 18422 11940
rect 18438 11996 18502 12000
rect 18438 11940 18442 11996
rect 18442 11940 18498 11996
rect 18498 11940 18502 11996
rect 18438 11936 18502 11940
rect 18518 11996 18582 12000
rect 18518 11940 18522 11996
rect 18522 11940 18578 11996
rect 18578 11940 18582 11996
rect 18518 11936 18582 11940
rect 7882 11452 7946 11456
rect 7882 11396 7886 11452
rect 7886 11396 7942 11452
rect 7942 11396 7946 11452
rect 7882 11392 7946 11396
rect 7962 11452 8026 11456
rect 7962 11396 7966 11452
rect 7966 11396 8022 11452
rect 8022 11396 8026 11452
rect 7962 11392 8026 11396
rect 8042 11452 8106 11456
rect 8042 11396 8046 11452
rect 8046 11396 8102 11452
rect 8102 11396 8106 11452
rect 8042 11392 8106 11396
rect 8122 11452 8186 11456
rect 8122 11396 8126 11452
rect 8126 11396 8182 11452
rect 8182 11396 8186 11452
rect 8122 11392 8186 11396
rect 14813 11452 14877 11456
rect 14813 11396 14817 11452
rect 14817 11396 14873 11452
rect 14873 11396 14877 11452
rect 14813 11392 14877 11396
rect 14893 11452 14957 11456
rect 14893 11396 14897 11452
rect 14897 11396 14953 11452
rect 14953 11396 14957 11452
rect 14893 11392 14957 11396
rect 14973 11452 15037 11456
rect 14973 11396 14977 11452
rect 14977 11396 15033 11452
rect 15033 11396 15037 11452
rect 14973 11392 15037 11396
rect 15053 11452 15117 11456
rect 15053 11396 15057 11452
rect 15057 11396 15113 11452
rect 15113 11396 15117 11452
rect 15053 11392 15117 11396
rect 4417 10908 4481 10912
rect 4417 10852 4421 10908
rect 4421 10852 4477 10908
rect 4477 10852 4481 10908
rect 4417 10848 4481 10852
rect 4497 10908 4561 10912
rect 4497 10852 4501 10908
rect 4501 10852 4557 10908
rect 4557 10852 4561 10908
rect 4497 10848 4561 10852
rect 4577 10908 4641 10912
rect 4577 10852 4581 10908
rect 4581 10852 4637 10908
rect 4637 10852 4641 10908
rect 4577 10848 4641 10852
rect 4657 10908 4721 10912
rect 4657 10852 4661 10908
rect 4661 10852 4717 10908
rect 4717 10852 4721 10908
rect 4657 10848 4721 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 18278 10908 18342 10912
rect 18278 10852 18282 10908
rect 18282 10852 18338 10908
rect 18338 10852 18342 10908
rect 18278 10848 18342 10852
rect 18358 10908 18422 10912
rect 18358 10852 18362 10908
rect 18362 10852 18418 10908
rect 18418 10852 18422 10908
rect 18358 10848 18422 10852
rect 18438 10908 18502 10912
rect 18438 10852 18442 10908
rect 18442 10852 18498 10908
rect 18498 10852 18502 10908
rect 18438 10848 18502 10852
rect 18518 10908 18582 10912
rect 18518 10852 18522 10908
rect 18522 10852 18578 10908
rect 18578 10852 18582 10908
rect 18518 10848 18582 10852
rect 7882 10364 7946 10368
rect 7882 10308 7886 10364
rect 7886 10308 7942 10364
rect 7942 10308 7946 10364
rect 7882 10304 7946 10308
rect 7962 10364 8026 10368
rect 7962 10308 7966 10364
rect 7966 10308 8022 10364
rect 8022 10308 8026 10364
rect 7962 10304 8026 10308
rect 8042 10364 8106 10368
rect 8042 10308 8046 10364
rect 8046 10308 8102 10364
rect 8102 10308 8106 10364
rect 8042 10304 8106 10308
rect 8122 10364 8186 10368
rect 8122 10308 8126 10364
rect 8126 10308 8182 10364
rect 8182 10308 8186 10364
rect 8122 10304 8186 10308
rect 14813 10364 14877 10368
rect 14813 10308 14817 10364
rect 14817 10308 14873 10364
rect 14873 10308 14877 10364
rect 14813 10304 14877 10308
rect 14893 10364 14957 10368
rect 14893 10308 14897 10364
rect 14897 10308 14953 10364
rect 14953 10308 14957 10364
rect 14893 10304 14957 10308
rect 14973 10364 15037 10368
rect 14973 10308 14977 10364
rect 14977 10308 15033 10364
rect 15033 10308 15037 10364
rect 14973 10304 15037 10308
rect 15053 10364 15117 10368
rect 15053 10308 15057 10364
rect 15057 10308 15113 10364
rect 15113 10308 15117 10364
rect 15053 10304 15117 10308
rect 4417 9820 4481 9824
rect 4417 9764 4421 9820
rect 4421 9764 4477 9820
rect 4477 9764 4481 9820
rect 4417 9760 4481 9764
rect 4497 9820 4561 9824
rect 4497 9764 4501 9820
rect 4501 9764 4557 9820
rect 4557 9764 4561 9820
rect 4497 9760 4561 9764
rect 4577 9820 4641 9824
rect 4577 9764 4581 9820
rect 4581 9764 4637 9820
rect 4637 9764 4641 9820
rect 4577 9760 4641 9764
rect 4657 9820 4721 9824
rect 4657 9764 4661 9820
rect 4661 9764 4717 9820
rect 4717 9764 4721 9820
rect 4657 9760 4721 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 18278 9820 18342 9824
rect 18278 9764 18282 9820
rect 18282 9764 18338 9820
rect 18338 9764 18342 9820
rect 18278 9760 18342 9764
rect 18358 9820 18422 9824
rect 18358 9764 18362 9820
rect 18362 9764 18418 9820
rect 18418 9764 18422 9820
rect 18358 9760 18422 9764
rect 18438 9820 18502 9824
rect 18438 9764 18442 9820
rect 18442 9764 18498 9820
rect 18498 9764 18502 9820
rect 18438 9760 18502 9764
rect 18518 9820 18582 9824
rect 18518 9764 18522 9820
rect 18522 9764 18578 9820
rect 18578 9764 18582 9820
rect 18518 9760 18582 9764
rect 7882 9276 7946 9280
rect 7882 9220 7886 9276
rect 7886 9220 7942 9276
rect 7942 9220 7946 9276
rect 7882 9216 7946 9220
rect 7962 9276 8026 9280
rect 7962 9220 7966 9276
rect 7966 9220 8022 9276
rect 8022 9220 8026 9276
rect 7962 9216 8026 9220
rect 8042 9276 8106 9280
rect 8042 9220 8046 9276
rect 8046 9220 8102 9276
rect 8102 9220 8106 9276
rect 8042 9216 8106 9220
rect 8122 9276 8186 9280
rect 8122 9220 8126 9276
rect 8126 9220 8182 9276
rect 8182 9220 8186 9276
rect 8122 9216 8186 9220
rect 14813 9276 14877 9280
rect 14813 9220 14817 9276
rect 14817 9220 14873 9276
rect 14873 9220 14877 9276
rect 14813 9216 14877 9220
rect 14893 9276 14957 9280
rect 14893 9220 14897 9276
rect 14897 9220 14953 9276
rect 14953 9220 14957 9276
rect 14893 9216 14957 9220
rect 14973 9276 15037 9280
rect 14973 9220 14977 9276
rect 14977 9220 15033 9276
rect 15033 9220 15037 9276
rect 14973 9216 15037 9220
rect 15053 9276 15117 9280
rect 15053 9220 15057 9276
rect 15057 9220 15113 9276
rect 15113 9220 15117 9276
rect 15053 9216 15117 9220
rect 17908 8876 17972 8940
rect 4417 8732 4481 8736
rect 4417 8676 4421 8732
rect 4421 8676 4477 8732
rect 4477 8676 4481 8732
rect 4417 8672 4481 8676
rect 4497 8732 4561 8736
rect 4497 8676 4501 8732
rect 4501 8676 4557 8732
rect 4557 8676 4561 8732
rect 4497 8672 4561 8676
rect 4577 8732 4641 8736
rect 4577 8676 4581 8732
rect 4581 8676 4637 8732
rect 4637 8676 4641 8732
rect 4577 8672 4641 8676
rect 4657 8732 4721 8736
rect 4657 8676 4661 8732
rect 4661 8676 4717 8732
rect 4717 8676 4721 8732
rect 4657 8672 4721 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 18278 8732 18342 8736
rect 18278 8676 18282 8732
rect 18282 8676 18338 8732
rect 18338 8676 18342 8732
rect 18278 8672 18342 8676
rect 18358 8732 18422 8736
rect 18358 8676 18362 8732
rect 18362 8676 18418 8732
rect 18418 8676 18422 8732
rect 18358 8672 18422 8676
rect 18438 8732 18502 8736
rect 18438 8676 18442 8732
rect 18442 8676 18498 8732
rect 18498 8676 18502 8732
rect 18438 8672 18502 8676
rect 18518 8732 18582 8736
rect 18518 8676 18522 8732
rect 18522 8676 18578 8732
rect 18578 8676 18582 8732
rect 18518 8672 18582 8676
rect 17908 8468 17972 8532
rect 7882 8188 7946 8192
rect 7882 8132 7886 8188
rect 7886 8132 7942 8188
rect 7942 8132 7946 8188
rect 7882 8128 7946 8132
rect 7962 8188 8026 8192
rect 7962 8132 7966 8188
rect 7966 8132 8022 8188
rect 8022 8132 8026 8188
rect 7962 8128 8026 8132
rect 8042 8188 8106 8192
rect 8042 8132 8046 8188
rect 8046 8132 8102 8188
rect 8102 8132 8106 8188
rect 8042 8128 8106 8132
rect 8122 8188 8186 8192
rect 8122 8132 8126 8188
rect 8126 8132 8182 8188
rect 8182 8132 8186 8188
rect 8122 8128 8186 8132
rect 14813 8188 14877 8192
rect 14813 8132 14817 8188
rect 14817 8132 14873 8188
rect 14873 8132 14877 8188
rect 14813 8128 14877 8132
rect 14893 8188 14957 8192
rect 14893 8132 14897 8188
rect 14897 8132 14953 8188
rect 14953 8132 14957 8188
rect 14893 8128 14957 8132
rect 14973 8188 15037 8192
rect 14973 8132 14977 8188
rect 14977 8132 15033 8188
rect 15033 8132 15037 8188
rect 14973 8128 15037 8132
rect 15053 8188 15117 8192
rect 15053 8132 15057 8188
rect 15057 8132 15113 8188
rect 15113 8132 15117 8188
rect 15053 8128 15117 8132
rect 19380 7924 19444 7988
rect 4417 7644 4481 7648
rect 4417 7588 4421 7644
rect 4421 7588 4477 7644
rect 4477 7588 4481 7644
rect 4417 7584 4481 7588
rect 4497 7644 4561 7648
rect 4497 7588 4501 7644
rect 4501 7588 4557 7644
rect 4557 7588 4561 7644
rect 4497 7584 4561 7588
rect 4577 7644 4641 7648
rect 4577 7588 4581 7644
rect 4581 7588 4637 7644
rect 4637 7588 4641 7644
rect 4577 7584 4641 7588
rect 4657 7644 4721 7648
rect 4657 7588 4661 7644
rect 4661 7588 4717 7644
rect 4717 7588 4721 7644
rect 4657 7584 4721 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 18278 7644 18342 7648
rect 18278 7588 18282 7644
rect 18282 7588 18338 7644
rect 18338 7588 18342 7644
rect 18278 7584 18342 7588
rect 18358 7644 18422 7648
rect 18358 7588 18362 7644
rect 18362 7588 18418 7644
rect 18418 7588 18422 7644
rect 18358 7584 18422 7588
rect 18438 7644 18502 7648
rect 18438 7588 18442 7644
rect 18442 7588 18498 7644
rect 18498 7588 18502 7644
rect 18438 7584 18502 7588
rect 18518 7644 18582 7648
rect 18518 7588 18522 7644
rect 18522 7588 18578 7644
rect 18578 7588 18582 7644
rect 18518 7584 18582 7588
rect 7882 7100 7946 7104
rect 7882 7044 7886 7100
rect 7886 7044 7942 7100
rect 7942 7044 7946 7100
rect 7882 7040 7946 7044
rect 7962 7100 8026 7104
rect 7962 7044 7966 7100
rect 7966 7044 8022 7100
rect 8022 7044 8026 7100
rect 7962 7040 8026 7044
rect 8042 7100 8106 7104
rect 8042 7044 8046 7100
rect 8046 7044 8102 7100
rect 8102 7044 8106 7100
rect 8042 7040 8106 7044
rect 8122 7100 8186 7104
rect 8122 7044 8126 7100
rect 8126 7044 8182 7100
rect 8182 7044 8186 7100
rect 8122 7040 8186 7044
rect 14813 7100 14877 7104
rect 14813 7044 14817 7100
rect 14817 7044 14873 7100
rect 14873 7044 14877 7100
rect 14813 7040 14877 7044
rect 14893 7100 14957 7104
rect 14893 7044 14897 7100
rect 14897 7044 14953 7100
rect 14953 7044 14957 7100
rect 14893 7040 14957 7044
rect 14973 7100 15037 7104
rect 14973 7044 14977 7100
rect 14977 7044 15033 7100
rect 15033 7044 15037 7100
rect 14973 7040 15037 7044
rect 15053 7100 15117 7104
rect 15053 7044 15057 7100
rect 15057 7044 15113 7100
rect 15113 7044 15117 7100
rect 15053 7040 15117 7044
rect 4417 6556 4481 6560
rect 4417 6500 4421 6556
rect 4421 6500 4477 6556
rect 4477 6500 4481 6556
rect 4417 6496 4481 6500
rect 4497 6556 4561 6560
rect 4497 6500 4501 6556
rect 4501 6500 4557 6556
rect 4557 6500 4561 6556
rect 4497 6496 4561 6500
rect 4577 6556 4641 6560
rect 4577 6500 4581 6556
rect 4581 6500 4637 6556
rect 4637 6500 4641 6556
rect 4577 6496 4641 6500
rect 4657 6556 4721 6560
rect 4657 6500 4661 6556
rect 4661 6500 4717 6556
rect 4717 6500 4721 6556
rect 4657 6496 4721 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 18278 6556 18342 6560
rect 18278 6500 18282 6556
rect 18282 6500 18338 6556
rect 18338 6500 18342 6556
rect 18278 6496 18342 6500
rect 18358 6556 18422 6560
rect 18358 6500 18362 6556
rect 18362 6500 18418 6556
rect 18418 6500 18422 6556
rect 18358 6496 18422 6500
rect 18438 6556 18502 6560
rect 18438 6500 18442 6556
rect 18442 6500 18498 6556
rect 18498 6500 18502 6556
rect 18438 6496 18502 6500
rect 18518 6556 18582 6560
rect 18518 6500 18522 6556
rect 18522 6500 18578 6556
rect 18578 6500 18582 6556
rect 18518 6496 18582 6500
rect 19380 6292 19444 6356
rect 7882 6012 7946 6016
rect 7882 5956 7886 6012
rect 7886 5956 7942 6012
rect 7942 5956 7946 6012
rect 7882 5952 7946 5956
rect 7962 6012 8026 6016
rect 7962 5956 7966 6012
rect 7966 5956 8022 6012
rect 8022 5956 8026 6012
rect 7962 5952 8026 5956
rect 8042 6012 8106 6016
rect 8042 5956 8046 6012
rect 8046 5956 8102 6012
rect 8102 5956 8106 6012
rect 8042 5952 8106 5956
rect 8122 6012 8186 6016
rect 8122 5956 8126 6012
rect 8126 5956 8182 6012
rect 8182 5956 8186 6012
rect 8122 5952 8186 5956
rect 14813 6012 14877 6016
rect 14813 5956 14817 6012
rect 14817 5956 14873 6012
rect 14873 5956 14877 6012
rect 14813 5952 14877 5956
rect 14893 6012 14957 6016
rect 14893 5956 14897 6012
rect 14897 5956 14953 6012
rect 14953 5956 14957 6012
rect 14893 5952 14957 5956
rect 14973 6012 15037 6016
rect 14973 5956 14977 6012
rect 14977 5956 15033 6012
rect 15033 5956 15037 6012
rect 14973 5952 15037 5956
rect 15053 6012 15117 6016
rect 15053 5956 15057 6012
rect 15057 5956 15113 6012
rect 15113 5956 15117 6012
rect 15053 5952 15117 5956
rect 4417 5468 4481 5472
rect 4417 5412 4421 5468
rect 4421 5412 4477 5468
rect 4477 5412 4481 5468
rect 4417 5408 4481 5412
rect 4497 5468 4561 5472
rect 4497 5412 4501 5468
rect 4501 5412 4557 5468
rect 4557 5412 4561 5468
rect 4497 5408 4561 5412
rect 4577 5468 4641 5472
rect 4577 5412 4581 5468
rect 4581 5412 4637 5468
rect 4637 5412 4641 5468
rect 4577 5408 4641 5412
rect 4657 5468 4721 5472
rect 4657 5412 4661 5468
rect 4661 5412 4717 5468
rect 4717 5412 4721 5468
rect 4657 5408 4721 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 18278 5468 18342 5472
rect 18278 5412 18282 5468
rect 18282 5412 18338 5468
rect 18338 5412 18342 5468
rect 18278 5408 18342 5412
rect 18358 5468 18422 5472
rect 18358 5412 18362 5468
rect 18362 5412 18418 5468
rect 18418 5412 18422 5468
rect 18358 5408 18422 5412
rect 18438 5468 18502 5472
rect 18438 5412 18442 5468
rect 18442 5412 18498 5468
rect 18498 5412 18502 5468
rect 18438 5408 18502 5412
rect 18518 5468 18582 5472
rect 18518 5412 18522 5468
rect 18522 5412 18578 5468
rect 18578 5412 18582 5468
rect 18518 5408 18582 5412
rect 7882 4924 7946 4928
rect 7882 4868 7886 4924
rect 7886 4868 7942 4924
rect 7942 4868 7946 4924
rect 7882 4864 7946 4868
rect 7962 4924 8026 4928
rect 7962 4868 7966 4924
rect 7966 4868 8022 4924
rect 8022 4868 8026 4924
rect 7962 4864 8026 4868
rect 8042 4924 8106 4928
rect 8042 4868 8046 4924
rect 8046 4868 8102 4924
rect 8102 4868 8106 4924
rect 8042 4864 8106 4868
rect 8122 4924 8186 4928
rect 8122 4868 8126 4924
rect 8126 4868 8182 4924
rect 8182 4868 8186 4924
rect 8122 4864 8186 4868
rect 14813 4924 14877 4928
rect 14813 4868 14817 4924
rect 14817 4868 14873 4924
rect 14873 4868 14877 4924
rect 14813 4864 14877 4868
rect 14893 4924 14957 4928
rect 14893 4868 14897 4924
rect 14897 4868 14953 4924
rect 14953 4868 14957 4924
rect 14893 4864 14957 4868
rect 14973 4924 15037 4928
rect 14973 4868 14977 4924
rect 14977 4868 15033 4924
rect 15033 4868 15037 4924
rect 14973 4864 15037 4868
rect 15053 4924 15117 4928
rect 15053 4868 15057 4924
rect 15057 4868 15113 4924
rect 15113 4868 15117 4924
rect 15053 4864 15117 4868
rect 4417 4380 4481 4384
rect 4417 4324 4421 4380
rect 4421 4324 4477 4380
rect 4477 4324 4481 4380
rect 4417 4320 4481 4324
rect 4497 4380 4561 4384
rect 4497 4324 4501 4380
rect 4501 4324 4557 4380
rect 4557 4324 4561 4380
rect 4497 4320 4561 4324
rect 4577 4380 4641 4384
rect 4577 4324 4581 4380
rect 4581 4324 4637 4380
rect 4637 4324 4641 4380
rect 4577 4320 4641 4324
rect 4657 4380 4721 4384
rect 4657 4324 4661 4380
rect 4661 4324 4717 4380
rect 4717 4324 4721 4380
rect 4657 4320 4721 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 18278 4380 18342 4384
rect 18278 4324 18282 4380
rect 18282 4324 18338 4380
rect 18338 4324 18342 4380
rect 18278 4320 18342 4324
rect 18358 4380 18422 4384
rect 18358 4324 18362 4380
rect 18362 4324 18418 4380
rect 18418 4324 18422 4380
rect 18358 4320 18422 4324
rect 18438 4380 18502 4384
rect 18438 4324 18442 4380
rect 18442 4324 18498 4380
rect 18498 4324 18502 4380
rect 18438 4320 18502 4324
rect 18518 4380 18582 4384
rect 18518 4324 18522 4380
rect 18522 4324 18578 4380
rect 18578 4324 18582 4380
rect 18518 4320 18582 4324
rect 7882 3836 7946 3840
rect 7882 3780 7886 3836
rect 7886 3780 7942 3836
rect 7942 3780 7946 3836
rect 7882 3776 7946 3780
rect 7962 3836 8026 3840
rect 7962 3780 7966 3836
rect 7966 3780 8022 3836
rect 8022 3780 8026 3836
rect 7962 3776 8026 3780
rect 8042 3836 8106 3840
rect 8042 3780 8046 3836
rect 8046 3780 8102 3836
rect 8102 3780 8106 3836
rect 8042 3776 8106 3780
rect 8122 3836 8186 3840
rect 8122 3780 8126 3836
rect 8126 3780 8182 3836
rect 8182 3780 8186 3836
rect 8122 3776 8186 3780
rect 14813 3836 14877 3840
rect 14813 3780 14817 3836
rect 14817 3780 14873 3836
rect 14873 3780 14877 3836
rect 14813 3776 14877 3780
rect 14893 3836 14957 3840
rect 14893 3780 14897 3836
rect 14897 3780 14953 3836
rect 14953 3780 14957 3836
rect 14893 3776 14957 3780
rect 14973 3836 15037 3840
rect 14973 3780 14977 3836
rect 14977 3780 15033 3836
rect 15033 3780 15037 3836
rect 14973 3776 15037 3780
rect 15053 3836 15117 3840
rect 15053 3780 15057 3836
rect 15057 3780 15113 3836
rect 15113 3780 15117 3836
rect 15053 3776 15117 3780
rect 4417 3292 4481 3296
rect 4417 3236 4421 3292
rect 4421 3236 4477 3292
rect 4477 3236 4481 3292
rect 4417 3232 4481 3236
rect 4497 3292 4561 3296
rect 4497 3236 4501 3292
rect 4501 3236 4557 3292
rect 4557 3236 4561 3292
rect 4497 3232 4561 3236
rect 4577 3292 4641 3296
rect 4577 3236 4581 3292
rect 4581 3236 4637 3292
rect 4637 3236 4641 3292
rect 4577 3232 4641 3236
rect 4657 3292 4721 3296
rect 4657 3236 4661 3292
rect 4661 3236 4717 3292
rect 4717 3236 4721 3292
rect 4657 3232 4721 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 18278 3292 18342 3296
rect 18278 3236 18282 3292
rect 18282 3236 18338 3292
rect 18338 3236 18342 3292
rect 18278 3232 18342 3236
rect 18358 3292 18422 3296
rect 18358 3236 18362 3292
rect 18362 3236 18418 3292
rect 18418 3236 18422 3292
rect 18358 3232 18422 3236
rect 18438 3292 18502 3296
rect 18438 3236 18442 3292
rect 18442 3236 18498 3292
rect 18498 3236 18502 3292
rect 18438 3232 18502 3236
rect 18518 3292 18582 3296
rect 18518 3236 18522 3292
rect 18522 3236 18578 3292
rect 18578 3236 18582 3292
rect 18518 3232 18582 3236
rect 7882 2748 7946 2752
rect 7882 2692 7886 2748
rect 7886 2692 7942 2748
rect 7942 2692 7946 2748
rect 7882 2688 7946 2692
rect 7962 2748 8026 2752
rect 7962 2692 7966 2748
rect 7966 2692 8022 2748
rect 8022 2692 8026 2748
rect 7962 2688 8026 2692
rect 8042 2748 8106 2752
rect 8042 2692 8046 2748
rect 8046 2692 8102 2748
rect 8102 2692 8106 2748
rect 8042 2688 8106 2692
rect 8122 2748 8186 2752
rect 8122 2692 8126 2748
rect 8126 2692 8182 2748
rect 8182 2692 8186 2748
rect 8122 2688 8186 2692
rect 14813 2748 14877 2752
rect 14813 2692 14817 2748
rect 14817 2692 14873 2748
rect 14873 2692 14877 2748
rect 14813 2688 14877 2692
rect 14893 2748 14957 2752
rect 14893 2692 14897 2748
rect 14897 2692 14953 2748
rect 14953 2692 14957 2748
rect 14893 2688 14957 2692
rect 14973 2748 15037 2752
rect 14973 2692 14977 2748
rect 14977 2692 15033 2748
rect 15033 2692 15037 2748
rect 14973 2688 15037 2692
rect 15053 2748 15117 2752
rect 15053 2692 15057 2748
rect 15057 2692 15113 2748
rect 15113 2692 15117 2748
rect 15053 2688 15117 2692
rect 4417 2204 4481 2208
rect 4417 2148 4421 2204
rect 4421 2148 4477 2204
rect 4477 2148 4481 2204
rect 4417 2144 4481 2148
rect 4497 2204 4561 2208
rect 4497 2148 4501 2204
rect 4501 2148 4557 2204
rect 4557 2148 4561 2204
rect 4497 2144 4561 2148
rect 4577 2204 4641 2208
rect 4577 2148 4581 2204
rect 4581 2148 4637 2204
rect 4637 2148 4641 2204
rect 4577 2144 4641 2148
rect 4657 2204 4721 2208
rect 4657 2148 4661 2204
rect 4661 2148 4717 2204
rect 4717 2148 4721 2204
rect 4657 2144 4721 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 18278 2204 18342 2208
rect 18278 2148 18282 2204
rect 18282 2148 18338 2204
rect 18338 2148 18342 2204
rect 18278 2144 18342 2148
rect 18358 2204 18422 2208
rect 18358 2148 18362 2204
rect 18362 2148 18418 2204
rect 18418 2148 18422 2204
rect 18358 2144 18422 2148
rect 18438 2204 18502 2208
rect 18438 2148 18442 2204
rect 18442 2148 18498 2204
rect 18498 2148 18502 2204
rect 18438 2144 18502 2148
rect 18518 2204 18582 2208
rect 18518 2148 18522 2204
rect 18522 2148 18578 2204
rect 18578 2148 18582 2204
rect 18518 2144 18582 2148
<< metal4 >>
rect 4409 20704 4729 20720
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 19616 4729 20640
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 18528 4729 19552
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 17440 4729 18464
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 16352 4729 17376
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 15264 4729 16288
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 14176 4729 15200
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 13088 4729 14112
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 12000 4729 13024
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 10912 4729 11936
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 9824 4729 10848
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 8736 4729 9760
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 7648 4729 8672
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 6560 4729 7584
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 5472 4729 6496
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 4384 4729 5408
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 3296 4729 4320
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 2208 4729 3232
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2128 4729 2144
rect 7874 20160 8195 20720
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8195 20160
rect 7874 19072 8195 20096
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8195 19072
rect 7874 17984 8195 19008
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8195 17984
rect 7874 16896 8195 17920
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8195 16896
rect 7874 15808 8195 16832
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8195 15808
rect 7874 14720 8195 15744
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8195 14720
rect 7874 13632 8195 14656
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8195 13632
rect 7874 12544 8195 13568
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8195 12544
rect 7874 11456 8195 12480
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8195 11456
rect 7874 10368 8195 11392
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8195 10368
rect 7874 9280 8195 10304
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8195 9280
rect 7874 8192 8195 9216
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8195 8192
rect 7874 7104 8195 8128
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8195 7104
rect 7874 6016 8195 7040
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8195 6016
rect 7874 4928 8195 5952
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8195 4928
rect 7874 3840 8195 4864
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8195 3840
rect 7874 2752 8195 3776
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8195 2752
rect 7874 2128 8195 2688
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 14805 20160 15125 20720
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 19072 15125 20096
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 17984 15125 19008
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 16896 15125 17920
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 15808 15125 16832
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 14720 15125 15744
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 13632 15125 14656
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 12544 15125 13568
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 11456 15125 12480
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 10368 15125 11392
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 9280 15125 10304
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 8192 15125 9216
rect 18270 20704 18591 20720
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18591 20704
rect 18270 19616 18591 20640
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18591 19616
rect 18270 18528 18591 19552
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18591 18528
rect 18270 17440 18591 18464
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18591 17440
rect 18270 16352 18591 17376
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18591 16352
rect 18270 15264 18591 16288
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18591 15264
rect 18270 14176 18591 15200
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18591 14176
rect 18270 13088 18591 14112
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18591 13088
rect 18270 12000 18591 13024
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18591 12000
rect 18270 10912 18591 11936
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18591 10912
rect 18270 9824 18591 10848
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18591 9824
rect 17907 8940 17973 8941
rect 17907 8876 17908 8940
rect 17972 8876 17973 8940
rect 17907 8875 17973 8876
rect 17910 8533 17970 8875
rect 18270 8736 18591 9760
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18591 8736
rect 17907 8532 17973 8533
rect 17907 8468 17908 8532
rect 17972 8468 17973 8532
rect 17907 8467 17973 8468
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 7104 15125 8128
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 6016 15125 7040
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 4928 15125 5952
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 3840 15125 4864
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 2752 15125 3776
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2128 15125 2688
rect 18270 7648 18591 8672
rect 19379 7988 19445 7989
rect 19379 7924 19380 7988
rect 19444 7924 19445 7988
rect 19379 7923 19445 7924
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18591 7648
rect 18270 6560 18591 7584
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18591 6560
rect 18270 5472 18591 6496
rect 19382 6357 19442 7923
rect 19379 6356 19445 6357
rect 19379 6292 19380 6356
rect 19444 6292 19445 6356
rect 19379 6291 19445 6292
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18591 5472
rect 18270 4384 18591 5408
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18591 4384
rect 18270 3296 18591 4320
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18591 3296
rect 18270 2208 18591 3232
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18591 2208
rect 18270 2128 18591 2144
use sky130_fd_sc_hd__decap_3  FILLER_1_15 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 2484 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15
timestamp 1608910539
transform 1 0 2484 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1608910539
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1608910539
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608910539
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 2760 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 2760 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_1_34 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 4232 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 4600 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 4048 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30
timestamp 1608910539
transform 1 0 3864 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24
timestamp 1608910539
transform 1 0 3312 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 4692 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 4416 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48
timestamp 1608910539
transform 1 0 5520 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1608910539
transform 1 0 5796 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_60
timestamp 1608910539
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 6256 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_52
timestamp 1608910539
transform 1 0 5888 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60
timestamp 1608910539
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 6072 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608910539
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608910539
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 6808 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_74
timestamp 1608910539
transform 1 0 7912 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_68
timestamp 1608910539
transform 1 0 7360 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81
timestamp 1608910539
transform 1 0 8556 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77
timestamp 1608910539
transform 1 0 8188 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_65
timestamp 1608910539
transform 1 0 7084 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 7728 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 6900 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1608910539
transform 1 0 8648 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 8096 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_1_97
timestamp 1608910539
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_92
timestamp 1608910539
transform 1 0 9568 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_103
timestamp 1608910539
transform 1 0 10580 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1608910539
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 9844 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608910539
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1608910539
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1608910539
transform 1 0 10212 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_108
timestamp 1608910539
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 11224 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_116
timestamp 1608910539
transform 1 0 11776 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115
timestamp 1608910539
transform 1 0 11684 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _097_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 11776 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120
timestamp 1608910539
transform 1 0 12144 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608910539
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608910539
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 12420 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 12604 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_129
timestamp 1608910539
transform 1 0 12972 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_131
timestamp 1608910539
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1608910539
transform 1 0 13156 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_135
timestamp 1608910539
transform 1 0 13524 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_137
timestamp 1608910539
transform 1 0 13708 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1608910539
transform 1 0 13340 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_145
timestamp 1608910539
transform 1 0 14444 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_143
timestamp 1608910539
transform 1 0 14260 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 13892 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1608910539
transform 1 0 13892 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_155
timestamp 1608910539
transform 1 0 15364 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_151
timestamp 1608910539
transform 1 0 14996 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_152
timestamp 1608910539
transform 1 0 15088 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_147
timestamp 1608910539
transform 1 0 14628 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608910539
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1608910539
transform 1 0 14720 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1608910539
transform 1 0 14628 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_165
timestamp 1608910539
transform 1 0 16284 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_162
timestamp 1608910539
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_156
timestamp 1608910539
transform 1 0 15456 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1608910539
transform 1 0 15456 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1608910539
transform 1 0 16100 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_173
timestamp 1608910539
transform 1 0 17020 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_173
timestamp 1608910539
transform 1 0 17020 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_167
timestamp 1608910539
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 16468 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1608910539
transform 1 0 16652 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_179
timestamp 1608910539
transform 1 0 17572 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 17204 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1608910539
transform 1 0 17204 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1608910539
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_187
timestamp 1608910539
transform 1 0 18308 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_185
timestamp 1608910539
transform 1 0 18124 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608910539
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608910539
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 18032 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_190
timestamp 1608910539
transform 1 0 18584 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1608910539
transform 1 0 19228 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_193
timestamp 1608910539
transform 1 0 18860 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1608910539
transform 1 0 19044 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 18768 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1608910539
transform 1 0 18492 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_204
timestamp 1608910539
transform 1 0 19872 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_198
timestamp 1608910539
transform 1 0 19320 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_203
timestamp 1608910539
transform 1 0 19780 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1608910539
transform 1 0 19964 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1608910539
transform 1 0 19412 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1608910539
transform 1 0 19504 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 20148 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_219
timestamp 1608910539
transform 1 0 21252 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_220
timestamp 1608910539
transform 1 0 21344 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1608910539
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_209
timestamp 1608910539
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1608910539
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608910539
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608910539
transform -1 0 21896 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608910539
transform -1 0 21896 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1608910539
transform 1 0 20516 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp 1608910539
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608910539
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 1656 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1608910539
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_30
timestamp 1608910539
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_26
timestamp 1608910539
transform 1 0 3496 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_22
timestamp 1608910539
transform 1 0 3128 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 3312 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608910539
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_54
timestamp 1608910539
transform 1 0 6072 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_44
timestamp 1608910539
transform 1 0 5152 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1608910539
transform 1 0 5244 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 6348 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_73
timestamp 1608910539
transform 1 0 7820 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_3_
timestamp 1608910539
transform 1 0 8188 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_97
timestamp 1608910539
transform 1 0 10028 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_93
timestamp 1608910539
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1608910539
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_86
timestamp 1608910539
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9844 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608910539
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10212 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_121
timestamp 1608910539
transform 1 0 12236 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_112
timestamp 1608910539
transform 1 0 11408 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_108
timestamp 1608910539
transform 1 0 11040 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 11224 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 12420 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 11684 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1608910539
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_135
timestamp 1608910539
transform 1 0 13524 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_129
timestamp 1608910539
transform 1 0 12972 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1608910539
transform 1 0 13708 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1608910539
transform 1 0 13156 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608910539
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 15272 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_180
timestamp 1608910539
transform 1 0 17664 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_170
timestamp 1608910539
transform 1 0 16744 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 17112 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1608910539
transform 1 0 18032 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_208
timestamp 1608910539
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_203
timestamp 1608910539
transform 1 0 19780 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_199
timestamp 1608910539
transform 1 0 19412 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_192
timestamp 1608910539
transform 1 0 18768 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_188
timestamp 1608910539
transform 1 0 18400 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 18860 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1608910539
transform 1 0 19872 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_219
timestamp 1608910539
transform 1 0 21252 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_212
timestamp 1608910539
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1608910539
transform 1 0 20424 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608910539
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608910539
transform -1 0 21896 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _056_
timestamp 1608910539
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_20
timestamp 1608910539
transform 1 0 2944 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1608910539
transform 1 0 1380 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608910539
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 1472 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_39
timestamp 1608910539
transform 1 0 4692 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_31 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3956 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1608910539
transform 1 0 3128 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1608910539
transform 1 0 4876 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_60
timestamp 1608910539
transform 1 0 6624 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_56
timestamp 1608910539
transform 1 0 6256 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_50
timestamp 1608910539
transform 1 0 5704 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 6808 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608910539
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _054_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 5980 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_77
timestamp 1608910539
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_64
timestamp 1608910539
transform 1 0 6992 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1608910539
transform 1 0 7360 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 8372 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_3_95
timestamp 1608910539
transform 1 0 9844 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1608910539
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_119
timestamp 1608910539
transform 1 0 12052 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_107
timestamp 1608910539
transform 1 0 10948 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608910539
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 13524 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_162
timestamp 1608910539
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_151
timestamp 1608910539
transform 1 0 14996 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1608910539
transform 1 0 16192 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1608910539
transform 1 0 15180 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_184
timestamp 1608910539
transform 1 0 18032 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_182
timestamp 1608910539
transform 1 0 17848 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_178
timestamp 1608910539
transform 1 0 17480 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_173
timestamp 1608910539
transform 1 0 17020 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608910539
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1608910539
transform 1 0 17204 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_199
timestamp 1608910539
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_195
timestamp 1608910539
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_191
timestamp 1608910539
transform 1 0 18676 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_188
timestamp 1608910539
transform 1 0 18400 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1608910539
transform 1 0 18492 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1608910539
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1608910539
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 19596 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_221
timestamp 1608910539
transform 1 0 21436 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_217
timestamp 1608910539
transform 1 0 21068 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__056__A
timestamp 1608910539
transform 1 0 21252 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608910539
transform -1 0 21896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_11
timestamp 1608910539
transform 1 0 2116 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_3
timestamp 1608910539
transform 1 0 1380 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608910539
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1608910539
transform 1 0 2208 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_38
timestamp 1608910539
transform 1 0 4600 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_34
timestamp 1608910539
transform 1 0 4232 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_25
timestamp 1608910539
transform 1 0 3404 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_21
timestamp 1608910539
transform 1 0 3036 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 4416 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608910539
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1608910539
transform 1 0 4784 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_61
timestamp 1608910539
transform 1 0 6716 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_49
timestamp 1608910539
transform 1 0 5612 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1608910539
transform 1 0 5888 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_83
timestamp 1608910539
transform 1 0 8740 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_72
timestamp 1608910539
transform 1 0 7728 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_69
timestamp 1608910539
transform 1 0 7452 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_65
timestamp 1608910539
transform 1 0 7084 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 7544 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6900 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1608910539
transform 1 0 7912 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1608910539
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_88
timestamp 1608910539
transform 1 0 9200 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608910539
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1608910539
transform 1 0 8924 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1608910539
transform 1 0 12236 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_116
timestamp 1608910539
transform 1 0 11776 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_105
timestamp 1608910539
transform 1 0 10764 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l2_in_0_
timestamp 1608910539
transform 1 0 10948 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1608910539
transform 1 0 11960 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_145
timestamp 1608910539
transform 1 0 14444 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_133
timestamp 1608910539
transform 1 0 13340 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_156
timestamp 1608910539
transform 1 0 15456 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_150
timestamp 1608910539
transform 1 0 14904 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 14720 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 15272 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608910539
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15732 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_187
timestamp 1608910539
transform 1 0 18308 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_175
timestamp 1608910539
transform 1 0 17204 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_207
timestamp 1608910539
transform 1 0 20148 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 18676 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_219
timestamp 1608910539
transform 1 0 21252 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_212
timestamp 1608910539
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608910539
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608910539
transform -1 0 21896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1608910539
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1608910539
transform 1 0 20332 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_13
timestamp 1608910539
transform 1 0 2300 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3
timestamp 1608910539
transform 1 0 1380 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608910539
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1608910539
transform 1 0 1472 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1608910539
transform 1 0 2484 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_5_32
timestamp 1608910539
transform 1 0 4048 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_28
timestamp 1608910539
transform 1 0 3680 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_24
timestamp 1608910539
transform 1 0 3312 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 3864 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 3496 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_62
timestamp 1608910539
transform 1 0 6808 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1608910539
transform 1 0 6348 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_46
timestamp 1608910539
transform 1 0 5336 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 5152 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608910539
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1608910539
transform 1 0 5520 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_5_72
timestamp 1608910539
transform 1 0 7728 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 7544 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_100
timestamp 1608910539
transform 1 0 10304 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_96
timestamp 1608910539
transform 1 0 9936 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_84
timestamp 1608910539
transform 1 0 8832 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 10396 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_5_121
timestamp 1608910539
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_117
timestamp 1608910539
transform 1 0 11868 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608910539
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 12420 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_139
timestamp 1608910539
transform 1 0 13892 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l2_in_0_
timestamp 1608910539
transform 1 0 14076 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_165
timestamp 1608910539
transform 1 0 16284 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_161
timestamp 1608910539
transform 1 0 15916 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_150
timestamp 1608910539
transform 1 0 14904 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 16100 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1608910539
transform 1 0 15088 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_181
timestamp 1608910539
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1608910539
transform 1 0 16652 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 16468 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608910539
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 18032 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_200
timestamp 1608910539
transform 1 0 19504 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1608910539
transform 1 0 19688 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_222
timestamp 1608910539
transform 1 0 21528 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_218
timestamp 1608910539
transform 1 0 21160 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_211
timestamp 1608910539
transform 1 0 20516 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608910539
transform -1 0 21896 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1608910539
transform 1 0 20792 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1608910539
transform 1 0 1380 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp 1608910539
transform 1 0 1748 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1608910539
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608910539
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608910539
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1608910539
transform 1 0 1472 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1608910539
transform 1 0 1840 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_13
timestamp 1608910539
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_11
timestamp 1608910539
transform 1 0 2116 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1608910539
transform 1 0 2484 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 2300 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_7_40
timestamp 1608910539
transform 1 0 4784 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_28
timestamp 1608910539
transform 1 0 3680 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_24
timestamp 1608910539
transform 1 0 3312 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1608910539
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 4876 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 3496 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608910539
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4048 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_48
timestamp 1608910539
transform 1 0 5520 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_43
timestamp 1608910539
transform 1 0 5060 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_48
timestamp 1608910539
transform 1 0 5520 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 5336 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 5796 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_0_
timestamp 1608910539
transform 1 0 5704 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1608910539
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_53
timestamp 1608910539
transform 1 0 5980 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608910539
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_1_
timestamp 1608910539
transform 1 0 6164 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_0_
timestamp 1608910539
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_71
timestamp 1608910539
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_64
timestamp 1608910539
transform 1 0 6992 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l3_in_0_
timestamp 1608910539
transform 1 0 7176 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_75
timestamp 1608910539
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_79
timestamp 1608910539
transform 1 0 8372 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_75
timestamp 1608910539
transform 1 0 8004 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 8188 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1608910539
transform 1 0 8556 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 8188 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_93
timestamp 1608910539
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1608910539
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608910539
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_101
timestamp 1608910539
transform 1 0 10396 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_95
timestamp 1608910539
transform 1 0 9844 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 10212 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1608910539
transform 1 0 9844 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10580 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_7_104
timestamp 1608910539
transform 1 0 10672 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_123
timestamp 1608910539
transform 1 0 12420 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_118
timestamp 1608910539
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_114
timestamp 1608910539
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_123
timestamp 1608910539
transform 1 0 12420 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_112
timestamp 1608910539
transform 1 0 11408 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608910539
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_1_
timestamp 1608910539
transform 1 0 11592 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_140
timestamp 1608910539
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_129
timestamp 1608910539
transform 1 0 12972 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_144
timestamp 1608910539
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_127
timestamp 1608910539
transform 1 0 12788 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 12788 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_1_
timestamp 1608910539
transform 1 0 14168 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_0_
timestamp 1608910539
transform 1 0 13156 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 12880 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_7_151
timestamp 1608910539
transform 1 0 14996 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_149
timestamp 1608910539
transform 1 0 14812 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 15272 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608910539
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1608910539
transform 1 0 14536 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_157
timestamp 1608910539
transform 1 0 15548 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_162
timestamp 1608910539
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_156
timestamp 1608910539
transform 1 0 15456 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l2_in_0_
timestamp 1608910539
transform 1 0 16100 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_0_
timestamp 1608910539
transform 1 0 15732 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_168
timestamp 1608910539
transform 1 0 16560 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_176
timestamp 1608910539
transform 1 0 17296 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_172
timestamp 1608910539
transform 1 0 16928 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 17112 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_1_
timestamp 1608910539
transform 1 0 16744 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_7_186
timestamp 1608910539
transform 1 0 18216 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_179
timestamp 1608910539
transform 1 0 17572 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 18032 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608910539
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1608910539
transform 1 0 17848 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_192
timestamp 1608910539
transform 1 0 18768 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_195
timestamp 1608910539
transform 1 0 19044 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_191
timestamp 1608910539
transform 1 0 18676 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 18584 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 18860 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 19228 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1608910539
transform 1 0 18952 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_203
timestamp 1608910539
transform 1 0 19780 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_199
timestamp 1608910539
transform 1 0 19412 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1608910539
transform 1 0 19596 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 19964 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_221
timestamp 1608910539
transform 1 0 21436 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_220
timestamp 1608910539
transform 1 0 21344 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_215
timestamp 1608910539
transform 1 0 20884 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_210
timestamp 1608910539
transform 1 0 20424 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1608910539
transform 1 0 21160 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608910539
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608910539
transform -1 0 21896 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608910539
transform -1 0 21896 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_18
timestamp 1608910539
transform 1 0 2760 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_14
timestamp 1608910539
transform 1 0 2392 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1608910539
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 2576 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608910539
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_3_
timestamp 1608910539
transform 1 0 1564 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_34
timestamp 1608910539
transform 1 0 4232 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_30
timestamp 1608910539
transform 1 0 3864 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608910539
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 4416 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_8_56
timestamp 1608910539
transform 1 0 6256 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_52
timestamp 1608910539
transform 1 0 5888 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 6348 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_77
timestamp 1608910539
transform 1 0 8188 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_73
timestamp 1608910539
transform 1 0 7820 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8004 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8556 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_95
timestamp 1608910539
transform 1 0 9844 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1608910539
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608910539
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 10212 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_115
timestamp 1608910539
transform 1 0 11684 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l3_in_0_
timestamp 1608910539
transform 1 0 11868 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_142
timestamp 1608910539
transform 1 0 14168 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1608910539
transform 1 0 13800 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_126
timestamp 1608910539
transform 1 0 12696 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 14352 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_154
timestamp 1608910539
transform 1 0 15272 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_152
timestamp 1608910539
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_146
timestamp 1608910539
transform 1 0 14536 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608910539
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 15364 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_8_176
timestamp 1608910539
transform 1 0 17296 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_171
timestamp 1608910539
transform 1 0 16836 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1608910539
transform 1 0 17020 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_199
timestamp 1608910539
transform 1 0 19412 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_188
timestamp 1608910539
transform 1 0 18400 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l2_in_0_
timestamp 1608910539
transform 1 0 18584 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l1_in_0_
timestamp 1608910539
transform 1 0 19596 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_222
timestamp 1608910539
transform 1 0 21528 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_218
timestamp 1608910539
transform 1 0 21160 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_210
timestamp 1608910539
transform 1 0 20424 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608910539
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608910539
transform -1 0 21896 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1608910539
transform 1 0 20884 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_12
timestamp 1608910539
transform 1 0 2208 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_9
timestamp 1608910539
transform 1 0 1932 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_5
timestamp 1608910539
transform 1 0 1564 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 2024 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608910539
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1608910539
transform 1 0 2392 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_32
timestamp 1608910539
transform 1 0 4048 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_23
timestamp 1608910539
transform 1 0 3220 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_3_
timestamp 1608910539
transform 1 0 4232 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1608910539
transform 1 0 3772 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_62
timestamp 1608910539
transform 1 0 6808 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_58
timestamp 1608910539
transform 1 0 6440 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1608910539
transform 1 0 6072 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_43
timestamp 1608910539
transform 1 0 5060 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 6256 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608910539
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_2_
timestamp 1608910539
transform 1 0 5244 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_9_70
timestamp 1608910539
transform 1 0 7544 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 7820 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_102
timestamp 1608910539
transform 1 0 10488 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_94
timestamp 1608910539
transform 1 0 9752 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_89
timestamp 1608910539
transform 1 0 9292 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9568 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 10672 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1608910539
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1608910539
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608910539
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_139
timestamp 1608910539
transform 1 0 13892 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_135
timestamp 1608910539
transform 1 0 13524 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 13984 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_9_156
timestamp 1608910539
transform 1 0 15456 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_184
timestamp 1608910539
transform 1 0 18032 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_9_177
timestamp 1608910539
transform 1 0 17388 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608910539
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l2_in_0_
timestamp 1608910539
transform 1 0 16560 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_197
timestamp 1608910539
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_192
timestamp 1608910539
transform 1 0 18768 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 19412 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_219
timestamp 1608910539
transform 1 0 21252 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_215
timestamp 1608910539
transform 1 0 20884 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 21068 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608910539
transform -1 0 21896 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_12
timestamp 1608910539
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_8
timestamp 1608910539
transform 1 0 1840 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 1608910539
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 1656 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608910539
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1608910539
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_41
timestamp 1608910539
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_28
timestamp 1608910539
transform 1 0 3680 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_23
timestamp 1608910539
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608910539
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1608910539
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1608910539
transform 1 0 3404 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_52
timestamp 1608910539
transform 1 0 5888 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_1_
timestamp 1608910539
transform 1 0 5060 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_82
timestamp 1608910539
transform 1 0 8648 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_78
timestamp 1608910539
transform 1 0 8280 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_73
timestamp 1608910539
transform 1 0 7820 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_70
timestamp 1608910539
transform 1 0 7544 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_64
timestamp 1608910539
transform 1 0 6992 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 8464 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 8004 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_103
timestamp 1608910539
transform 1 0 10580 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_93
timestamp 1608910539
transform 1 0 9660 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1608910539
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 10396 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608910539
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_124
timestamp 1608910539
transform 1 0 12512 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_113
timestamp 1608910539
transform 1 0 11500 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_108
timestamp 1608910539
transform 1 0 11040 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 10856 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_0_
timestamp 1608910539
transform 1 0 11684 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1608910539
transform 1 0 11224 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_142
timestamp 1608910539
transform 1 0 14168 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 14352 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 12696 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_166
timestamp 1608910539
transform 1 0 16376 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_154
timestamp 1608910539
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1608910539
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_146
timestamp 1608910539
transform 1 0 14536 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608910539
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_0_
timestamp 1608910539
transform 1 0 15548 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_184
timestamp 1608910539
transform 1 0 18032 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 16560 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1608910539
transform 1 0 18216 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_208
timestamp 1608910539
transform 1 0 20240 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_10_189
timestamp 1608910539
transform 1 0 18492 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 18768 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_10_215
timestamp 1608910539
transform 1 0 20884 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608910539
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608910539
transform -1 0 21896 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_7
timestamp 1608910539
transform 1 0 1748 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1608910539
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608910539
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 1840 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_11_39
timestamp 1608910539
transform 1 0 4692 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_28
timestamp 1608910539
transform 1 0 3680 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_24
timestamp 1608910539
transform 1 0 3312 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 3496 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1608910539
transform 1 0 3864 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1608910539
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_53
timestamp 1608910539
transform 1 0 5980 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_47
timestamp 1608910539
transform 1 0 5428 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 5704 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608910539
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1608910539
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_79
timestamp 1608910539
transform 1 0 8372 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_75
timestamp 1608910539
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_71
timestamp 1608910539
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 8740 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_99
timestamp 1608910539
transform 1 0 10212 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_123
timestamp 1608910539
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_116
timestamp 1608910539
transform 1 0 11776 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_105
timestamp 1608910539
transform 1 0 10764 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608910539
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_1_
timestamp 1608910539
transform 1 0 10948 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_139
timestamp 1608910539
transform 1 0 13892 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_135
timestamp 1608910539
transform 1 0 13524 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1608910539
transform 1 0 13984 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l1_in_0_
timestamp 1608910539
transform 1 0 12696 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_155
timestamp 1608910539
transform 1 0 15364 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_149
timestamp 1608910539
transform 1 0 14812 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 15456 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_181
timestamp 1608910539
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_176
timestamp 1608910539
transform 1 0 17296 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_172
timestamp 1608910539
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608910539
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_1_
timestamp 1608910539
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_11_207
timestamp 1608910539
transform 1 0 20148 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_197
timestamp 1608910539
transform 1 0 19228 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_193
timestamp 1608910539
transform 1 0 18860 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1608910539
transform 1 0 19320 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_219
timestamp 1608910539
transform 1 0 21252 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608910539
transform -1 0 21896 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_11
timestamp 1608910539
transform 1 0 2116 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3
timestamp 1608910539
transform 1 0 1380 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608910539
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1608910539
transform 1 0 2208 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_12_28
timestamp 1608910539
transform 1 0 3680 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_25
timestamp 1608910539
transform 1 0 3404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_21
timestamp 1608910539
transform 1 0 3036 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 3496 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608910539
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4048 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_48
timestamp 1608910539
transform 1 0 5520 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 5704 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_77
timestamp 1608910539
transform 1 0 8188 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_66
timestamp 1608910539
transform 1 0 7176 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1608910539
transform 1 0 8372 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1608910539
transform 1 0 7360 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_12_102
timestamp 1608910539
transform 1 0 10488 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_88
timestamp 1608910539
transform 1 0 9200 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608910539
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1608910539
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_122
timestamp 1608910539
transform 1 0 12328 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_118
timestamp 1608910539
transform 1 0 11960 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_114
timestamp 1608910539
transform 1 0 11592 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 12144 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 11776 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 12512 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1608910539
transform 1 0 10764 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_140
timestamp 1608910539
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_134
timestamp 1608910539
transform 1 0 13432 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_126
timestamp 1608910539
transform 1 0 12696 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 13708 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1608910539
transform 1 0 14168 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_12_162
timestamp 1608910539
transform 1 0 16008 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_158
timestamp 1608910539
transform 1 0 15640 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_154
timestamp 1608910539
transform 1 0 15272 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1608910539
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 15732 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608910539
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_186
timestamp 1608910539
transform 1 0 18216 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_174
timestamp 1608910539
transform 1 0 17112 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_201
timestamp 1608910539
transform 1 0 19596 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_198
timestamp 1608910539
transform 1 0 19320 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 19412 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1608910539
transform 1 0 19780 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_222
timestamp 1608910539
transform 1 0 21528 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_218
timestamp 1608910539
transform 1 0 21160 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_212
timestamp 1608910539
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608910539
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608910539
transform -1 0 21896 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1608910539
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_11
timestamp 1608910539
transform 1 0 2116 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1608910539
transform 1 0 1380 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_9
timestamp 1608910539
transform 1 0 1932 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1608910539
transform 1 0 1380 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608910539
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608910539
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1608910539
transform 1 0 2300 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 2024 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_14_40
timestamp 1608910539
transform 1 0 4784 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_32
timestamp 1608910539
transform 1 0 4048 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_30
timestamp 1608910539
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_22
timestamp 1608910539
transform 1 0 3128 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_38
timestamp 1608910539
transform 1 0 4600 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_26
timestamp 1608910539
transform 1 0 3496 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608910539
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1608910539
transform 1 0 4876 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_61
timestamp 1608910539
transform 1 0 6716 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_50
timestamp 1608910539
transform 1 0 5704 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1608910539
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_56
timestamp 1608910539
transform 1 0 6256 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_50
timestamp 1608910539
transform 1 0 5704 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608910539
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1608910539
transform 1 0 5888 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1608910539
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_72
timestamp 1608910539
transform 1 0 7728 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_71
timestamp 1608910539
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1608910539
transform 1 0 6900 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_14_81
timestamp 1608910539
transform 1 0 8556 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_77
timestamp 1608910539
transform 1 0 8188 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_81
timestamp 1608910539
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_76
timestamp 1608910539
transform 1 0 8096 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 7820 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1608910539
transform 1 0 7912 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_89
timestamp 1608910539
transform 1 0 9292 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_100
timestamp 1608910539
transform 1 0 10304 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_89
timestamp 1608910539
transform 1 0 9292 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_85
timestamp 1608910539
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9108 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1608910539
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1608910539
transform 1 0 10488 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1608910539
transform 1 0 9476 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 9660 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_14_109
timestamp 1608910539
transform 1 0 11132 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_123
timestamp 1608910539
transform 1 0 12420 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_13_119
timestamp 1608910539
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_111
timestamp 1608910539
transform 1 0 11316 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608910539
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 11316 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_14_145
timestamp 1608910539
transform 1 0 14444 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_127
timestamp 1608910539
transform 1 0 12788 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_129
timestamp 1608910539
transform 1 0 12972 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 13064 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 12972 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1608910539
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_151
timestamp 1608910539
transform 1 0 14996 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_146
timestamp 1608910539
transform 1 0 14536 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 14720 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1608910539
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_3_
timestamp 1608910539
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1608910539
transform 1 0 15180 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_163
timestamp 1608910539
transform 1 0 16100 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_156
timestamp 1608910539
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1608910539
transform 1 0 15640 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_13_175
timestamp 1608910539
transform 1 0 17204 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_171
timestamp 1608910539
transform 1 0 16836 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_167
timestamp 1608910539
transform 1 0 16468 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 17020 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 16652 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_183
timestamp 1608910539
transform 1 0 17940 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1608910539
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608910539
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_1_
timestamp 1608910539
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 18124 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 16468 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_14_201
timestamp 1608910539
transform 1 0 19596 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_193
timestamp 1608910539
transform 1 0 18860 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1608910539
transform 1 0 19780 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 19596 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_14_217
timestamp 1608910539
transform 1 0 21068 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_212
timestamp 1608910539
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1608910539
transform 1 0 21068 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 20884 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1608910539
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608910539
transform -1 0 21896 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608910539
transform -1 0 21896 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_20
timestamp 1608910539
transform 1 0 2944 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_14
timestamp 1608910539
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_6
timestamp 1608910539
transform 1 0 1656 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1608910539
transform 1 0 1380 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_5__A0
timestamp 1608910539
transform 1 0 1472 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608910539
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1840 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1608910539
transform 1 0 2576 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_28
timestamp 1608910539
transform 1 0 3680 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 3864 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_62
timestamp 1608910539
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1608910539
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_46
timestamp 1608910539
transform 1 0 5336 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1608910539
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1608910539
transform 1 0 5704 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_80
timestamp 1608910539
transform 1 0 8464 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 8648 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 6992 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_100
timestamp 1608910539
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_89
timestamp 1608910539
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_84
timestamp 1608910539
transform 1 0 8832 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 9108 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1608910539
transform 1 0 9476 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1608910539
transform 1 0 10488 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_125
timestamp 1608910539
transform 1 0 12604 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1608910539
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_117
timestamp 1608910539
transform 1 0 11868 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_105
timestamp 1608910539
transform 1 0 10764 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1608910539
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_139
timestamp 1608910539
transform 1 0 13892 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_133
timestamp 1608910539
transform 1 0 13340 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_129
timestamp 1608910539
transform 1 0 12972 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 13064 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1608910539
transform 1 0 13984 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_15_161
timestamp 1608910539
transform 1 0 15916 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1608910539
transform 1 0 14812 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1608910539
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_176
timestamp 1608910539
transform 1 0 17296 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_173
timestamp 1608910539
transform 1 0 17020 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 17112 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1608910539
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_0_
timestamp 1608910539
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1608910539
transform 1 0 17480 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_193
timestamp 1608910539
transform 1 0 18860 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 19228 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_221
timestamp 1608910539
transform 1 0 21436 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_213
timestamp 1608910539
transform 1 0 20700 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608910539
transform -1 0 21896 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_12
timestamp 1608910539
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1608910539
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608910539
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_5_
timestamp 1608910539
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1656 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_16_32
timestamp 1608910539
transform 1 0 4048 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1608910539
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_23
timestamp 1608910539
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_5__A1
timestamp 1608910539
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1608910539
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4324 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_57
timestamp 1608910539
transform 1 0 6348 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_51
timestamp 1608910539
transform 1 0 5796 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 6164 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1608910539
transform 1 0 6532 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_79
timestamp 1608910539
transform 1 0 8372 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_68
timestamp 1608910539
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 8556 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1608910539
transform 1 0 7544 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_16_102
timestamp 1608910539
transform 1 0 10488 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_96
timestamp 1608910539
transform 1 0 9936 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1608910539
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_84
timestamp 1608910539
transform 1 0 8832 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 10304 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1608910539
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1608910539
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_125
timestamp 1608910539
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 10764 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_16_140
timestamp 1608910539
transform 1 0 13984 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_136
timestamp 1608910539
transform 1 0 13616 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_mem_bottom_track_1.prog_clk_A
timestamp 1608910539
transform 1 0 13800 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1608910539
transform 1 0 12788 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1608910539
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1608910539
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15272 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_178
timestamp 1608910539
transform 1 0 17480 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_170
timestamp 1608910539
transform 1 0 16744 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l2_in_0_
timestamp 1608910539
transform 1 0 17664 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_205
timestamp 1608910539
transform 1 0 19964 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_199
timestamp 1608910539
transform 1 0 19412 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_195
timestamp 1608910539
transform 1 0 19044 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_189
timestamp 1608910539
transform 1 0 18492 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 19780 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 19228 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 20148 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 18860 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_221
timestamp 1608910539
transform 1 0 21436 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_217
timestamp 1608910539
transform 1 0 21068 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_213
timestamp 1608910539
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_209
timestamp 1608910539
transform 1 0 20332 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 20884 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 21252 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1608910539
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608910539
transform -1 0 21896 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_10
timestamp 1608910539
transform 1 0 2024 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_3
timestamp 1608910539
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608910539
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 2208 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1608910539
transform 1 0 1656 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_37
timestamp 1608910539
transform 1 0 4508 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_34
timestamp 1608910539
transform 1 0 4232 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_28
timestamp 1608910539
transform 1 0 3680 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A0
timestamp 1608910539
transform 1 0 4324 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1608910539
transform 1 0 6348 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_53
timestamp 1608910539
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_49
timestamp 1608910539
transform 1 0 5612 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1608910539
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_3_
timestamp 1608910539
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_78
timestamp 1608910539
transform 1 0 8280 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_75
timestamp 1608910539
transform 1 0 8004 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_71
timestamp 1608910539
transform 1 0 7636 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 8096 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_3_
timestamp 1608910539
transform 1 0 8464 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_100
timestamp 1608910539
transform 1 0 10304 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_89
timestamp 1608910539
transform 1 0 9292 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1608910539
transform 1 0 10488 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1608910539
transform 1 0 9476 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1608910539
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_115
timestamp 1608910539
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_111
timestamp 1608910539
transform 1 0 11316 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 11500 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1608910539
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1608910539
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1608910539
transform 1 0 11868 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_143
timestamp 1608910539
transform 1 0 14260 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_132
timestamp 1608910539
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1608910539
transform 1 0 13432 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_17_155
timestamp 1608910539
transform 1 0 15364 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1608910539
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_177
timestamp 1608910539
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_167
timestamp 1608910539
transform 1 0 16468 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1608910539
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1608910539
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_203
timestamp 1608910539
transform 1 0 19780 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_197
timestamp 1608910539
transform 1 0 19228 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_193
timestamp 1608910539
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 19596 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 19964 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_221
timestamp 1608910539
transform 1 0 21436 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608910539
transform -1 0 21896 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_12
timestamp 1608910539
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_8
timestamp 1608910539
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1608910539
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_4__A0
timestamp 1608910539
transform 1 0 1656 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_4__A1
timestamp 1608910539
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608910539
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_4_
timestamp 1608910539
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_37
timestamp 1608910539
transform 1 0 4508 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_32
timestamp 1608910539
transform 1 0 4048 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_23
timestamp 1608910539
transform 1 0 3220 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 4324 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1608910539
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1608910539
transform 1 0 4692 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_59
timestamp 1608910539
transform 1 0 6532 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_56
timestamp 1608910539
transform 1 0 6256 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_48
timestamp 1608910539
transform 1 0 5520 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 6348 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1608910539
transform 1 0 6716 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_79
timestamp 1608910539
transform 1 0 8372 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_75
timestamp 1608910539
transform 1 0 8004 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_64
timestamp 1608910539
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 8188 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1608910539
transform 1 0 7176 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_102
timestamp 1608910539
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_89
timestamp 1608910539
transform 1 0 9292 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1608910539
transform 1 0 8924 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 9108 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1608910539
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1608910539
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_18_124
timestamp 1608910539
transform 1 0 12512 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_106
timestamp 1608910539
transform 1 0 10856 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 11040 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_143
timestamp 1608910539
transform 1 0 14260 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_5__A0
timestamp 1608910539
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 12788 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_18_163
timestamp 1608910539
transform 1 0 16100 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1608910539
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_147
timestamp 1608910539
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_5__A1
timestamp 1608910539
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1608910539
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_5_
timestamp 1608910539
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 16376 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_182
timestamp 1608910539
transform 1 0 17848 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1608910539
transform 1 0 18032 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_18_207
timestamp 1608910539
transform 1 0 20148 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_197
timestamp 1608910539
transform 1 0 19228 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_193
timestamp 1608910539
transform 1 0 18860 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1608910539
transform 1 0 19320 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_219
timestamp 1608910539
transform 1 0 21252 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1608910539
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 20424 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1608910539
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608910539
transform -1 0 21896 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1608910539
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_8
timestamp 1608910539
transform 1 0 1840 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3
timestamp 1608910539
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1608910539
transform 1 0 1380 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_6__A1
timestamp 1608910539
transform 1 0 1656 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608910539
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608910539
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_12
timestamp 1608910539
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_11
timestamp 1608910539
transform 1 0 2116 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__A
timestamp 1608910539
transform 1 0 2024 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1608910539
transform 1 0 2208 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_6_
timestamp 1608910539
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1608910539
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_23
timestamp 1608910539
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_21
timestamp 1608910539
transform 1 0 3036 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_6__A0
timestamp 1608910539
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1608910539
transform 1 0 3588 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_38
timestamp 1608910539
transform 1 0 4600 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_32
timestamp 1608910539
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_36
timestamp 1608910539
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 4416 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1608910539
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1608910539
transform 1 0 4600 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1608910539
transform 1 0 4784 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_49
timestamp 1608910539
transform 1 0 5612 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1608910539
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_47
timestamp 1608910539
transform 1 0 5428 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 5612 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 5796 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_57
timestamp 1608910539
transform 1 0 6348 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_53
timestamp 1608910539
transform 1 0 5980 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1608910539
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 6164 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1608910539
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1608910539
transform 1 0 6716 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_62
timestamp 1608910539
transform 1 0 6808 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_70
timestamp 1608910539
transform 1 0 7544 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_66
timestamp 1608910539
transform 1 0 7176 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 6992 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 7728 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1608910539
transform 1 0 7360 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_75
timestamp 1608910539
transform 1 0 8004 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_81
timestamp 1608910539
transform 1 0 8556 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_77
timestamp 1608910539
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8188 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_79
timestamp 1608910539
transform 1 0 8372 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1608910539
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1608910539
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1608910539
transform 1 0 9108 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1608910539
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_102
timestamp 1608910539
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_100
timestamp 1608910539
transform 1 0 10304 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_96
timestamp 1608910539
transform 1 0 9936 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 10120 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 10672 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_106
timestamp 1608910539
transform 1 0 10856 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_114
timestamp 1608910539
transform 1 0 11592 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1608910539
transform 1 0 11224 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_106
timestamp 1608910539
transform 1 0 10856 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 11040 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1608910539
transform 1 0 11132 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_118
timestamp 1608910539
transform 1 0 11960 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1608910539
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1608910539
transform 1 0 12144 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_19_125
timestamp 1608910539
transform 1 0 12604 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_142
timestamp 1608910539
transform 1 0 14168 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_137
timestamp 1608910539
transform 1 0 13708 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_129
timestamp 1608910539
transform 1 0 12972 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_140
timestamp 1608910539
transform 1 0 13984 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 13892 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1608910539
transform 1 0 13156 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 14260 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_20_163
timestamp 1608910539
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_150
timestamp 1608910539
transform 1 0 14904 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_165
timestamp 1608910539
transform 1 0 16284 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_159
timestamp 1608910539
transform 1 0 15732 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_4__A0
timestamp 1608910539
transform 1 0 16100 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1608910539
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_4_
timestamp 1608910539
transform 1 0 16284 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1608910539
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_174
timestamp 1608910539
transform 1 0 17112 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1608910539
transform 1 0 16652 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 17296 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 16468 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1608910539
transform 1 0 16836 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_186
timestamp 1608910539
transform 1 0 18216 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_182
timestamp 1608910539
transform 1 0 17848 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_178
timestamp 1608910539
transform 1 0 17480 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_184
timestamp 1608910539
transform 1 0 18032 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_180
timestamp 1608910539
transform 1 0 17664 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A0
timestamp 1608910539
transform 1 0 17664 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 18032 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1608910539
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1608910539
transform 1 0 18308 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_208
timestamp 1608910539
transform 1 0 20240 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1608910539
transform 1 0 19228 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_207
timestamp 1608910539
transform 1 0 20148 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_196
timestamp 1608910539
transform 1 0 19136 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1608910539
transform 1 0 18400 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1608910539
transform 1 0 19320 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1608910539
transform 1 0 19412 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_221
timestamp 1608910539
transform 1 0 21436 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_212
timestamp 1608910539
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_220
timestamp 1608910539
transform 1 0 21344 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1608910539
transform 1 0 20424 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1608910539
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608910539
transform -1 0 21896 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608910539
transform -1 0 21896 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 20884 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1608910539
transform 1 0 20516 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_10
timestamp 1608910539
transform 1 0 2024 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1608910539
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608910539
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1608910539
transform 1 0 2208 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1608910539
transform 1 0 1656 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_41
timestamp 1608910539
transform 1 0 4876 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_26
timestamp 1608910539
transform 1 0 3496 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_21
timestamp 1608910539
transform 1 0 3036 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1608910539
transform 1 0 4048 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1608910539
transform 1 0 3220 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_62
timestamp 1608910539
transform 1 0 6808 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_60
timestamp 1608910539
transform 1 0 6624 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_56
timestamp 1608910539
transform 1 0 6256 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_52
timestamp 1608910539
transform 1 0 5888 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 6072 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1608910539
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1608910539
transform 1 0 5060 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_74
timestamp 1608910539
transform 1 0 7912 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1608910539
transform 1 0 8280 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1608910539
transform 1 0 7084 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_102
timestamp 1608910539
transform 1 0 10488 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_98
timestamp 1608910539
transform 1 0 10120 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_87
timestamp 1608910539
transform 1 0 9108 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1608910539
transform 1 0 9292 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1608910539
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_120
timestamp 1608910539
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_109
timestamp 1608910539
transform 1 0 11132 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_105
timestamp 1608910539
transform 1 0 10764 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 10948 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1608910539
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1608910539
transform 1 0 11316 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_21_135
timestamp 1608910539
transform 1 0 13524 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1608910539
transform 1 0 13800 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_158
timestamp 1608910539
transform 1 0 15640 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_147
timestamp 1608910539
transform 1 0 14628 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 15364 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1608910539
transform 1 0 15824 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_187
timestamp 1608910539
transform 1 0 18308 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_184
timestamp 1608910539
transform 1 0 18032 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_182
timestamp 1608910539
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_176
timestamp 1608910539
transform 1 0 17296 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_173
timestamp 1608910539
transform 1 0 17020 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_169
timestamp 1608910539
transform 1 0 16652 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 18124 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_4__A1
timestamp 1608910539
transform 1 0 17112 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1608910539
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_202
timestamp 1608910539
transform 1 0 19688 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_191
timestamp 1608910539
transform 1 0 18676 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 18492 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1608910539
transform 1 0 19872 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1608910539
transform 1 0 18860 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_219
timestamp 1608910539
transform 1 0 21252 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_213
timestamp 1608910539
transform 1 0 20700 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608910539
transform -1 0 21896 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1608910539
transform 1 0 20884 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_11
timestamp 1608910539
transform 1 0 2116 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1608910539
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608910539
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1564 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1608910539
transform 1 0 2300 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_41
timestamp 1608910539
transform 1 0 4876 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_30
timestamp 1608910539
transform 1 0 3864 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_22
timestamp 1608910539
transform 1 0 3128 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1608910539
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1608910539
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_60
timestamp 1608910539
transform 1 0 6624 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_45
timestamp 1608910539
transform 1 0 5244 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 5060 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1608910539
transform 1 0 5796 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1608910539
transform 1 0 6808 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_22_76
timestamp 1608910539
transform 1 0 8096 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_71
timestamp 1608910539
transform 1 0 7636 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 7912 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_88
timestamp 1608910539
transform 1 0 9200 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1608910539
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9660 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_22_117
timestamp 1608910539
transform 1 0 11868 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_109
timestamp 1608910539
transform 1 0 11132 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 11960 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_145
timestamp 1608910539
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_134
timestamp 1608910539
transform 1 0 13432 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1608910539
transform 1 0 13616 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_22_158
timestamp 1608910539
transform 1 0 15640 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_154
timestamp 1608910539
transform 1 0 15272 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_150
timestamp 1608910539
transform 1 0 14904 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1608910539
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 15732 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1608910539
transform 1 0 14628 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_175
timestamp 1608910539
transform 1 0 17204 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 17388 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_208
timestamp 1608910539
transform 1 0 20240 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1608910539
transform 1 0 19228 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_193
timestamp 1608910539
transform 1 0 18860 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A0
timestamp 1608910539
transform 1 0 19044 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_6_
timestamp 1608910539
transform 1 0 19412 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_221
timestamp 1608910539
transform 1 0 21436 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1608910539
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A1
timestamp 1608910539
transform 1 0 20424 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1608910539
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608910539
transform -1 0 21896 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 20884 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_11
timestamp 1608910539
transform 1 0 2116 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1608910539
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1608910539
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 2484 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1608910539
transform 1 0 1748 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_31
timestamp 1608910539
transform 1 0 3956 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1608910539
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1608910539
transform 1 0 6164 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_43
timestamp 1608910539
transform 1 0 5060 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 6256 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1608910539
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 6808 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_78
timestamp 1608910539
transform 1 0 8280 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 8464 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_96
timestamp 1608910539
transform 1 0 9936 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 10120 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_23_123
timestamp 1608910539
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_114
timestamp 1608910539
transform 1 0 11592 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1608910539
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_129
timestamp 1608910539
transform 1 0 12972 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 12696 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 13156 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_23_158
timestamp 1608910539
transform 1 0 15640 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_147
timestamp 1608910539
transform 1 0 14628 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_3_
timestamp 1608910539
transform 1 0 14812 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_23_184
timestamp 1608910539
transform 1 0 18032 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_181
timestamp 1608910539
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_170
timestamp 1608910539
transform 1 0 16744 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1608910539
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1608910539
transform 1 0 16928 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_201
timestamp 1608910539
transform 1 0 19596 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1608910539
transform 1 0 19780 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1608910539
transform 1 0 18768 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_23_222
timestamp 1608910539
transform 1 0 21528 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_218
timestamp 1608910539
transform 1 0 21160 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_212
timestamp 1608910539
transform 1 0 20608 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1608910539
transform -1 0 21896 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1608910539
transform 1 0 20792 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_15
timestamp 1608910539
transform 1 0 2484 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_11
timestamp 1608910539
transform 1 0 2116 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1608910539
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__A
timestamp 1608910539
transform 1 0 2300 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1608910539
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1608910539
transform 1 0 2668 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1608910539
transform 1 0 1748 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_30
timestamp 1608910539
transform 1 0 3864 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_26
timestamp 1608910539
transform 1 0 3496 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1608910539
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 4048 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_24_48
timestamp 1608910539
transform 1 0 5520 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 5888 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_24_81
timestamp 1608910539
transform 1 0 8556 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_24_72
timestamp 1608910539
transform 1 0 7728 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_68
timestamp 1608910539
transform 1 0 7360 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 7544 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 8280 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1608910539
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_89
timestamp 1608910539
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1608910539
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_105
timestamp 1608910539
transform 1 0 10764 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 11316 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_24_135
timestamp 1608910539
transform 1 0 13524 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_127
timestamp 1608910539
transform 1 0 12788 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1608910539
transform 1 0 13800 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_24_154
timestamp 1608910539
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_151
timestamp 1608910539
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_147
timestamp 1608910539
transform 1 0 14628 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 14812 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1608910539
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15548 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_24_179
timestamp 1608910539
transform 1 0 17572 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_173
timestamp 1608910539
transform 1 0 17020 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 17664 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_206
timestamp 1608910539
transform 1 0 20056 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_201
timestamp 1608910539
transform 1 0 19596 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_196
timestamp 1608910539
transform 1 0 19136 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1608910539
transform 1 0 19872 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1608910539
transform 1 0 20240 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1608910539
transform 1 0 19320 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_219
timestamp 1608910539
transform 1 0 21252 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_212
timestamp 1608910539
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1608910539
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1608910539
transform -1 0 21896 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1608910539
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_20
timestamp 1608910539
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_16
timestamp 1608910539
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_8
timestamp 1608910539
transform 1 0 1840 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1608910539
transform 1 0 1380 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A
timestamp 1608910539
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1608910539
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2024 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1608910539
transform 1 0 1472 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_24
timestamp 1608910539
transform 1 0 3312 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 3128 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4416 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_25_62
timestamp 1608910539
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1608910539
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_56
timestamp 1608910539
transform 1 0 6256 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1608910539
transform 1 0 5888 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1608910539
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_78
timestamp 1608910539
transform 1 0 8280 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_74
timestamp 1608910539
transform 1 0 7912 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 8096 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1608910539
transform 1 0 7084 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 8464 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_25_96
timestamp 1608910539
transform 1 0 9936 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_123
timestamp 1608910539
transform 1 0 12420 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_118
timestamp 1608910539
transform 1 0 11960 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_108
timestamp 1608910539
transform 1 0 11040 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1608910539
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_134
timestamp 1608910539
transform 1 0 13432 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_131
timestamp 1608910539
transform 1 0 13156 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_158
timestamp 1608910539
transform 1 0 15640 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_146
timestamp 1608910539
transform 1 0 14536 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_184
timestamp 1608910539
transform 1 0 18032 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_179
timestamp 1608910539
transform 1 0 17572 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_175
timestamp 1608910539
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_170
timestamp 1608910539
transform 1 0 16744 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 17020 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1608910539
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_203
timestamp 1608910539
transform 1 0 19780 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_198
timestamp 1608910539
transform 1 0 19320 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_190
timestamp 1608910539
transform 1 0 18584 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 18400 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1608910539
transform 1 0 19596 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 19964 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_222
timestamp 1608910539
transform 1 0 21528 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_218
timestamp 1608910539
transform 1 0 21160 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_211
timestamp 1608910539
transform 1 0 20516 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1608910539
transform -1 0 21896 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1608910539
transform 1 0 20792 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1608910539
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1608910539
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1608910539
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1608910539
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_5
timestamp 1608910539
transform 1 0 1564 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1608910539
transform 1 0 1748 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1608910539
transform 1 0 1748 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_11
timestamp 1608910539
transform 1 0 2116 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_11
timestamp 1608910539
transform 1 0 2116 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1608910539
transform 1 0 2300 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1608910539
transform 1 0 2300 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_17
timestamp 1608910539
transform 1 0 2668 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_17
timestamp 1608910539
transform 1 0 2668 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A
timestamp 1608910539
transform 1 0 2852 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_31
timestamp 1608910539
transform 1 0 3956 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_21
timestamp 1608910539
transform 1 0 3036 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1608910539
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_25
timestamp 1608910539
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_21
timestamp 1608910539
transform 1 0 3036 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1608910539
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1608910539
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1608910539
transform 1 0 3128 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_41
timestamp 1608910539
transform 1 0 4876 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_36
timestamp 1608910539
transform 1 0 4416 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 4692 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1608910539
transform 1 0 4140 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1608910539
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_44
timestamp 1608910539
transform 1 0 5152 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1608910539
transform 1 0 5060 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1608910539
transform 1 0 5520 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_27_60
timestamp 1608910539
transform 1 0 6624 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_52
timestamp 1608910539
transform 1 0 5888 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_61
timestamp 1608910539
transform 1 0 6716 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_57
timestamp 1608910539
transform 1 0 6348 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6532 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1608910539
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_62
timestamp 1608910539
transform 1 0 6808 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_69
timestamp 1608910539
transform 1 0 7452 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_65
timestamp 1608910539
transform 1 0 7084 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 7268 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 7636 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 6900 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1608910539
transform 1 0 6992 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_81
timestamp 1608910539
transform 1 0 8556 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_77
timestamp 1608910539
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_73
timestamp 1608910539
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_73
timestamp 1608910539
transform 1 0 7820 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1608910539
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_27_85
timestamp 1608910539
transform 1 0 8924 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_93
timestamp 1608910539
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_84
timestamp 1608910539
transform 1 0 8832 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1608910539
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1608910539
transform 1 0 9016 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_95
timestamp 1608910539
transform 1 0 9844 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_101
timestamp 1608910539
transform 1 0 10396 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_97
timestamp 1608910539
transform 1 0 10028 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 10212 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 9844 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 10580 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1608910539
transform 1 0 10212 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_27_119
timestamp 1608910539
transform 1 0 12052 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_108
timestamp 1608910539
transform 1 0 11040 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_116
timestamp 1608910539
transform 1 0 11776 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_105
timestamp 1608910539
transform 1 0 10764 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1608910539
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1608910539
transform 1 0 11960 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1608910539
transform 1 0 11224 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1608910539
transform 1 0 10948 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1608910539
transform 1 0 12420 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_130
timestamp 1608910539
transform 1 0 13064 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_126
timestamp 1608910539
transform 1 0 12696 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_131
timestamp 1608910539
transform 1 0 13156 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_127
timestamp 1608910539
transform 1 0 12788 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 12972 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1608910539
transform 1 0 13156 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1608910539
transform 1 0 13432 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_143
timestamp 1608910539
transform 1 0 14260 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 14444 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_140
timestamp 1608910539
transform 1 0 13984 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_161
timestamp 1608910539
transform 1 0 15916 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_162
timestamp 1608910539
transform 1 0 16008 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_154
timestamp 1608910539
transform 1 0 15272 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_147
timestamp 1608910539
transform 1 0 14628 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1608910539
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 15088 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1608910539
transform 1 0 16100 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 16192 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_176
timestamp 1608910539
transform 1 0 17296 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_172
timestamp 1608910539
transform 1 0 16928 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_173
timestamp 1608910539
transform 1 0 17020 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 17112 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1608910539
transform 1 0 17388 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_27_184
timestamp 1608910539
transform 1 0 18032 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_180
timestamp 1608910539
transform 1 0 17664 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_186
timestamp 1608910539
transform 1 0 18216 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 17480 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1608910539
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 18124 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_27_201
timestamp 1608910539
transform 1 0 19596 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_202
timestamp 1608910539
transform 1 0 19688 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_196
timestamp 1608910539
transform 1 0 19136 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_190
timestamp 1608910539
transform 1 0 18584 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 18400 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1608910539
transform 1 0 18952 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 19872 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 19780 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1608910539
transform 1 0 19320 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_213
timestamp 1608910539
transform 1 0 20700 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_209
timestamp 1608910539
transform 1 0 20332 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_210
timestamp 1608910539
transform 1 0 20424 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_218
timestamp 1608910539
transform 1 0 21160 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1608910539
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1608910539
transform 1 0 20792 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1608910539
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_222
timestamp 1608910539
transform 1 0 21528 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_219
timestamp 1608910539
transform 1 0 21252 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1608910539
transform -1 0 21896 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1608910539
transform -1 0 21896 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_16
timestamp 1608910539
transform 1 0 2576 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_8
timestamp 1608910539
transform 1 0 1840 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_3
timestamp 1608910539
transform 1 0 1380 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1608910539
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2024 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1608910539
transform 1 0 2944 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1608910539
transform 1 0 1472 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_34
timestamp 1608910539
transform 1 0 4232 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1608910539
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1608910539
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1608910539
transform 1 0 4508 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_46
timestamp 1608910539
transform 1 0 5336 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 5704 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_77
timestamp 1608910539
transform 1 0 8188 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_70
timestamp 1608910539
transform 1 0 7544 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_66
timestamp 1608910539
transform 1 0 7176 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8372 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 7636 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_88
timestamp 1608910539
transform 1 0 9200 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1608910539
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 9660 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_28_125
timestamp 1608910539
transform 1 0 12604 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_114
timestamp 1608910539
transform 1 0 11592 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_109
timestamp 1608910539
transform 1 0 11132 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 11408 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1608910539
transform 1 0 11776 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_142
timestamp 1608910539
transform 1 0 14168 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_131
timestamp 1608910539
transform 1 0 13156 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 12972 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 14352 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1608910539
transform 1 0 13340 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_28_163
timestamp 1608910539
transform 1 0 16100 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1608910539
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_146
timestamp 1608910539
transform 1 0 14536 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1608910539
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1608910539
transform 1 0 16376 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1608910539
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1608910539
transform 1 0 14720 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_175
timestamp 1608910539
transform 1 0 17204 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 17388 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_201
timestamp 1608910539
transform 1 0 19596 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_193
timestamp 1608910539
transform 1 0 18860 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1608910539
transform 1 0 19412 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 19780 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_219
timestamp 1608910539
transform 1 0 21252 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_213
timestamp 1608910539
transform 1 0 20700 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_209
timestamp 1608910539
transform 1 0 20332 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1608910539
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1608910539
transform -1 0 21896 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1608910539
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_15
timestamp 1608910539
transform 1 0 2484 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_11
timestamp 1608910539
transform 1 0 2116 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_5
timestamp 1608910539
transform 1 0 1564 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1608910539
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1608910539
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1608910539
transform 1 0 2576 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1608910539
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_25
timestamp 1608910539
transform 1 0 3404 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 3588 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1608910539
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_55
timestamp 1608910539
transform 1 0 6164 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_43
timestamp 1608910539
transform 1 0 5060 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1608910539
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_74
timestamp 1608910539
transform 1 0 7912 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8096 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_29_98
timestamp 1608910539
transform 1 0 10120 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_90
timestamp 1608910539
transform 1 0 9384 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_85
timestamp 1608910539
transform 1 0 8924 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9200 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 10396 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_29_123
timestamp 1608910539
transform 1 0 12420 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_121
timestamp 1608910539
transform 1 0 12236 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_117
timestamp 1608910539
transform 1 0 11868 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1608910539
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_143
timestamp 1608910539
transform 1 0 14260 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_131
timestamp 1608910539
transform 1 0 13156 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 12972 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1608910539
transform 1 0 14444 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_29_165
timestamp 1608910539
transform 1 0 16284 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_154
timestamp 1608910539
transform 1 0 15272 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1608910539
transform 1 0 15456 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1608910539
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_177
timestamp 1608910539
transform 1 0 17388 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_173
timestamp 1608910539
transform 1 0 17020 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 17204 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1608910539
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_206
timestamp 1608910539
transform 1 0 20056 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_202
timestamp 1608910539
transform 1 0 19688 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_196
timestamp 1608910539
transform 1 0 19136 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1608910539
transform 1 0 19504 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1608910539
transform 1 0 19872 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1608910539
transform 1 0 20240 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_222
timestamp 1608910539
transform 1 0 21528 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_218
timestamp 1608910539
transform 1 0 21160 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_212
timestamp 1608910539
transform 1 0 20608 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1608910539
transform -1 0 21896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1608910539
transform 1 0 20792 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_17
timestamp 1608910539
transform 1 0 2668 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_11
timestamp 1608910539
transform 1 0 2116 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1608910539
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1608910539
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1608910539
transform 1 0 2852 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1608910539
transform 1 0 2300 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1608910539
transform 1 0 1748 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_41
timestamp 1608910539
transform 1 0 4876 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1608910539
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_23
timestamp 1608910539
transform 1 0 3220 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1608910539
transform 1 0 3404 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1608910539
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1608910539
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_30_60
timestamp 1608910539
transform 1 0 6624 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 5152 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_30_82
timestamp 1608910539
transform 1 0 8648 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 7176 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1608910539
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1608910539
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1608910539
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_117
timestamp 1608910539
transform 1 0 11868 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1608910539
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 11960 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_30_134
timestamp 1608910539
transform 1 0 13432 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1608910539
transform 1 0 14168 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_151
timestamp 1608910539
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1608910539
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 15272 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_30_182
timestamp 1608910539
transform 1 0 17848 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_170
timestamp 1608910539
transform 1 0 16744 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_202
timestamp 1608910539
transform 1 0 19688 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_194
timestamp 1608910539
transform 1 0 18952 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1608910539
transform 1 0 19504 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 19872 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_219
timestamp 1608910539
transform 1 0 21252 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_210
timestamp 1608910539
transform 1 0 20424 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1608910539
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1608910539
transform -1 0 21896 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1608910539
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_17
timestamp 1608910539
transform 1 0 2668 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_11
timestamp 1608910539
transform 1 0 2116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1608910539
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1608910539
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1608910539
transform 1 0 2300 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1608910539
transform 1 0 1748 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_38
timestamp 1608910539
transform 1 0 4600 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_21
timestamp 1608910539
transform 1 0 3036 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 3128 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_31_62
timestamp 1608910539
transform 1 0 6808 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_58
timestamp 1608910539
transform 1 0 6440 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_50
timestamp 1608910539
transform 1 0 5704 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1608910539
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_74
timestamp 1608910539
transform 1 0 7912 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1608910539
transform 1 0 7084 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 8096 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_99
timestamp 1608910539
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_96
timestamp 1608910539
transform 1 0 9936 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_92
timestamp 1608910539
transform 1 0 9568 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608910539
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 10396 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_31_123
timestamp 1608910539
transform 1 0 12420 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_121
timestamp 1608910539
transform 1 0 12236 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_117
timestamp 1608910539
transform 1 0 11868 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1608910539
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_131
timestamp 1608910539
transform 1 0 13156 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 13248 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_31_160
timestamp 1608910539
transform 1 0 15824 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_148
timestamp 1608910539
transform 1 0 14720 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_184
timestamp 1608910539
transform 1 0 18032 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_180
timestamp 1608910539
transform 1 0 17664 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_172
timestamp 1608910539
transform 1 0 16928 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1608910539
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_206
timestamp 1608910539
transform 1 0 20056 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_200
timestamp 1608910539
transform 1 0 19504 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_194
timestamp 1608910539
transform 1 0 18952 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1608910539
transform 1 0 18768 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1608910539
transform 1 0 19136 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1608910539
transform 1 0 19688 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1608910539
transform 1 0 20240 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_222
timestamp 1608910539
transform 1 0 21528 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_218
timestamp 1608910539
transform 1 0 21160 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_212
timestamp 1608910539
transform 1 0 20608 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1608910539
transform -1 0 21896 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1608910539
transform 1 0 20792 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_15
timestamp 1608910539
transform 1 0 2484 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_11
timestamp 1608910539
transform 1 0 2116 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_5
timestamp 1608910539
transform 1 0 1564 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1608910539
transform 1 0 1380 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1608910539
transform 1 0 2300 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1608910539
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2760 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1608910539
transform 1 0 1748 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1608910539
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_28
timestamp 1608910539
transform 1 0 3680 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_24
timestamp 1608910539
transform 1 0 3312 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1608910539
transform 1 0 3496 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1608910539
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1608910539
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1608910539
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_79
timestamp 1608910539
transform 1 0 8372 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_68
timestamp 1608910539
transform 1 0 7360 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1608910539
transform 1 0 7544 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1608910539
transform 1 0 8556 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1608910539
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_84
timestamp 1608910539
transform 1 0 8832 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1608910539
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_117
timestamp 1608910539
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1608910539
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1608910539
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_129
timestamp 1608910539
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_166
timestamp 1608910539
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_154
timestamp 1608910539
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1608910539
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_178
timestamp 1608910539
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_206
timestamp 1608910539
transform 1 0 20056 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_202
timestamp 1608910539
transform 1 0 19688 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_190
timestamp 1608910539
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1608910539
transform 1 0 19872 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1608910539
transform 1 0 20240 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_219
timestamp 1608910539
transform 1 0 21252 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_212
timestamp 1608910539
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1608910539
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1608910539
transform -1 0 21896 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1608910539
transform 1 0 20884 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_17
timestamp 1608910539
transform 1 0 2668 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_11
timestamp 1608910539
transform 1 0 2116 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1608910539
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1608910539
transform 1 0 2852 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1608910539
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1608910539
transform 1 0 2300 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1608910539
transform 1 0 1748 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_32
timestamp 1608910539
transform 1 0 4048 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_25
timestamp 1608910539
transform 1 0 3404 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_21
timestamp 1608910539
transform 1 0 3036 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1608910539
transform 1 0 3220 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1608910539
transform 1 0 3956 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_56
timestamp 1608910539
transform 1 0 6256 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_44
timestamp 1608910539
transform 1 0 5152 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1608910539
transform 1 0 6808 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_75
timestamp 1608910539
transform 1 0 8004 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_63
timestamp 1608910539
transform 1 0 6900 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_94
timestamp 1608910539
transform 1 0 9752 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_87
timestamp 1608910539
transform 1 0 9108 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1608910539
transform 1 0 9660 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_125
timestamp 1608910539
transform 1 0 12604 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_118
timestamp 1608910539
transform 1 0 11960 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_106
timestamp 1608910539
transform 1 0 10856 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1608910539
transform 1 0 12512 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_137
timestamp 1608910539
transform 1 0 13708 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_156
timestamp 1608910539
transform 1 0 15456 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_149
timestamp 1608910539
transform 1 0 14812 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1608910539
transform 1 0 15364 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_187
timestamp 1608910539
transform 1 0 18308 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_180
timestamp 1608910539
transform 1 0 17664 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_168
timestamp 1608910539
transform 1 0 16560 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1608910539
transform 1 0 18216 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_208
timestamp 1608910539
transform 1 0 20240 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_204
timestamp 1608910539
transform 1 0 19872 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_199
timestamp 1608910539
transform 1 0 19412 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1608910539
transform 1 0 19688 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1608910539
transform 1 0 20056 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_220
timestamp 1608910539
transform 1 0 21344 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_215
timestamp 1608910539
transform 1 0 20884 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1608910539
transform 1 0 21160 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1608910539
transform 1 0 21068 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1608910539
transform -1 0 21896 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1608910539
transform 1 0 20516 0 1 20128
box -38 -48 406 592
<< labels >>
rlabel metal2 s 21822 0 21878 800 6 SC_IN_BOT
port 0 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 SC_OUT_BOT
port 1 nsew signal tristate
rlabel metal2 s 202 0 258 800 6 bottom_left_grid_pin_42_
port 2 nsew signal input
rlabel metal2 s 570 0 626 800 6 bottom_left_grid_pin_43_
port 3 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 bottom_left_grid_pin_44_
port 4 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 bottom_left_grid_pin_45_
port 5 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 bottom_left_grid_pin_46_
port 6 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 bottom_left_grid_pin_47_
port 7 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 bottom_left_grid_pin_48_
port 8 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 bottom_left_grid_pin_49_
port 9 nsew signal input
rlabel metal2 s 5722 22200 5778 23000 6 ccff_head
port 10 nsew signal input
rlabel metal2 s 17222 22200 17278 23000 6 ccff_tail
port 11 nsew signal tristate
rlabel metal3 s 0 3816 800 3936 6 chanx_left_in[0]
port 12 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 chanx_left_in[10]
port 13 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 chanx_left_in[11]
port 14 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 chanx_left_in[12]
port 15 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 chanx_left_in[13]
port 16 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 chanx_left_in[14]
port 17 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 chanx_left_in[15]
port 18 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[16]
port 19 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 chanx_left_in[17]
port 20 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[18]
port 21 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 chanx_left_in[19]
port 22 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 chanx_left_in[1]
port 23 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 chanx_left_in[2]
port 24 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 chanx_left_in[3]
port 25 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 chanx_left_in[4]
port 26 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 chanx_left_in[5]
port 27 nsew signal input
rlabel metal3 s 0 6672 800 6792 6 chanx_left_in[6]
port 28 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 chanx_left_in[7]
port 29 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 chanx_left_in[8]
port 30 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 chanx_left_in[9]
port 31 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 chanx_left_out[0]
port 32 nsew signal tristate
rlabel metal3 s 0 17960 800 18080 6 chanx_left_out[10]
port 33 nsew signal tristate
rlabel metal3 s 0 18368 800 18488 6 chanx_left_out[11]
port 34 nsew signal tristate
rlabel metal3 s 0 18776 800 18896 6 chanx_left_out[12]
port 35 nsew signal tristate
rlabel metal3 s 0 19320 800 19440 6 chanx_left_out[13]
port 36 nsew signal tristate
rlabel metal3 s 0 19728 800 19848 6 chanx_left_out[14]
port 37 nsew signal tristate
rlabel metal3 s 0 20272 800 20392 6 chanx_left_out[15]
port 38 nsew signal tristate
rlabel metal3 s 0 20680 800 20800 6 chanx_left_out[16]
port 39 nsew signal tristate
rlabel metal3 s 0 21224 800 21344 6 chanx_left_out[17]
port 40 nsew signal tristate
rlabel metal3 s 0 21632 800 21752 6 chanx_left_out[18]
port 41 nsew signal tristate
rlabel metal3 s 0 22176 800 22296 6 chanx_left_out[19]
port 42 nsew signal tristate
rlabel metal3 s 0 13744 800 13864 6 chanx_left_out[1]
port 43 nsew signal tristate
rlabel metal3 s 0 14152 800 14272 6 chanx_left_out[2]
port 44 nsew signal tristate
rlabel metal3 s 0 14560 800 14680 6 chanx_left_out[3]
port 45 nsew signal tristate
rlabel metal3 s 0 15104 800 15224 6 chanx_left_out[4]
port 46 nsew signal tristate
rlabel metal3 s 0 15512 800 15632 6 chanx_left_out[5]
port 47 nsew signal tristate
rlabel metal3 s 0 16056 800 16176 6 chanx_left_out[6]
port 48 nsew signal tristate
rlabel metal3 s 0 16464 800 16584 6 chanx_left_out[7]
port 49 nsew signal tristate
rlabel metal3 s 0 17008 800 17128 6 chanx_left_out[8]
port 50 nsew signal tristate
rlabel metal3 s 0 17416 800 17536 6 chanx_left_out[9]
port 51 nsew signal tristate
rlabel metal3 s 22200 3816 23000 3936 6 chanx_right_in[0]
port 52 nsew signal input
rlabel metal3 s 22200 8576 23000 8696 6 chanx_right_in[10]
port 53 nsew signal input
rlabel metal3 s 22200 8984 23000 9104 6 chanx_right_in[11]
port 54 nsew signal input
rlabel metal3 s 22200 9392 23000 9512 6 chanx_right_in[12]
port 55 nsew signal input
rlabel metal3 s 22200 9936 23000 10056 6 chanx_right_in[13]
port 56 nsew signal input
rlabel metal3 s 22200 10344 23000 10464 6 chanx_right_in[14]
port 57 nsew signal input
rlabel metal3 s 22200 10888 23000 11008 6 chanx_right_in[15]
port 58 nsew signal input
rlabel metal3 s 22200 11296 23000 11416 6 chanx_right_in[16]
port 59 nsew signal input
rlabel metal3 s 22200 11840 23000 11960 6 chanx_right_in[17]
port 60 nsew signal input
rlabel metal3 s 22200 12248 23000 12368 6 chanx_right_in[18]
port 61 nsew signal input
rlabel metal3 s 22200 12792 23000 12912 6 chanx_right_in[19]
port 62 nsew signal input
rlabel metal3 s 22200 4360 23000 4480 6 chanx_right_in[1]
port 63 nsew signal input
rlabel metal3 s 22200 4768 23000 4888 6 chanx_right_in[2]
port 64 nsew signal input
rlabel metal3 s 22200 5176 23000 5296 6 chanx_right_in[3]
port 65 nsew signal input
rlabel metal3 s 22200 5720 23000 5840 6 chanx_right_in[4]
port 66 nsew signal input
rlabel metal3 s 22200 6128 23000 6248 6 chanx_right_in[5]
port 67 nsew signal input
rlabel metal3 s 22200 6672 23000 6792 6 chanx_right_in[6]
port 68 nsew signal input
rlabel metal3 s 22200 7080 23000 7200 6 chanx_right_in[7]
port 69 nsew signal input
rlabel metal3 s 22200 7624 23000 7744 6 chanx_right_in[8]
port 70 nsew signal input
rlabel metal3 s 22200 8032 23000 8152 6 chanx_right_in[9]
port 71 nsew signal input
rlabel metal3 s 22200 13200 23000 13320 6 chanx_right_out[0]
port 72 nsew signal tristate
rlabel metal3 s 22200 17960 23000 18080 6 chanx_right_out[10]
port 73 nsew signal tristate
rlabel metal3 s 22200 18368 23000 18488 6 chanx_right_out[11]
port 74 nsew signal tristate
rlabel metal3 s 22200 18776 23000 18896 6 chanx_right_out[12]
port 75 nsew signal tristate
rlabel metal3 s 22200 19320 23000 19440 6 chanx_right_out[13]
port 76 nsew signal tristate
rlabel metal3 s 22200 19728 23000 19848 6 chanx_right_out[14]
port 77 nsew signal tristate
rlabel metal3 s 22200 20272 23000 20392 6 chanx_right_out[15]
port 78 nsew signal tristate
rlabel metal3 s 22200 20680 23000 20800 6 chanx_right_out[16]
port 79 nsew signal tristate
rlabel metal3 s 22200 21224 23000 21344 6 chanx_right_out[17]
port 80 nsew signal tristate
rlabel metal3 s 22200 21632 23000 21752 6 chanx_right_out[18]
port 81 nsew signal tristate
rlabel metal3 s 22200 22176 23000 22296 6 chanx_right_out[19]
port 82 nsew signal tristate
rlabel metal3 s 22200 13744 23000 13864 6 chanx_right_out[1]
port 83 nsew signal tristate
rlabel metal3 s 22200 14152 23000 14272 6 chanx_right_out[2]
port 84 nsew signal tristate
rlabel metal3 s 22200 14560 23000 14680 6 chanx_right_out[3]
port 85 nsew signal tristate
rlabel metal3 s 22200 15104 23000 15224 6 chanx_right_out[4]
port 86 nsew signal tristate
rlabel metal3 s 22200 15512 23000 15632 6 chanx_right_out[5]
port 87 nsew signal tristate
rlabel metal3 s 22200 16056 23000 16176 6 chanx_right_out[6]
port 88 nsew signal tristate
rlabel metal3 s 22200 16464 23000 16584 6 chanx_right_out[7]
port 89 nsew signal tristate
rlabel metal3 s 22200 17008 23000 17128 6 chanx_right_out[8]
port 90 nsew signal tristate
rlabel metal3 s 22200 17416 23000 17536 6 chanx_right_out[9]
port 91 nsew signal tristate
rlabel metal2 s 3790 0 3846 800 6 chany_bottom_in[0]
port 92 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 chany_bottom_in[10]
port 93 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 chany_bottom_in[11]
port 94 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 chany_bottom_in[12]
port 95 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 chany_bottom_in[13]
port 96 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 chany_bottom_in[14]
port 97 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 chany_bottom_in[15]
port 98 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 chany_bottom_in[16]
port 99 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 chany_bottom_in[17]
port 100 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 chany_bottom_in[18]
port 101 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 chany_bottom_in[19]
port 102 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 chany_bottom_in[1]
port 103 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 chany_bottom_in[2]
port 104 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 chany_bottom_in[3]
port 105 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 chany_bottom_in[4]
port 106 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 chany_bottom_in[5]
port 107 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 chany_bottom_in[6]
port 108 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 chany_bottom_in[7]
port 109 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 chany_bottom_in[8]
port 110 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 chany_bottom_in[9]
port 111 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 chany_bottom_out[0]
port 112 nsew signal tristate
rlabel metal2 s 17314 0 17370 800 6 chany_bottom_out[10]
port 113 nsew signal tristate
rlabel metal2 s 17774 0 17830 800 6 chany_bottom_out[11]
port 114 nsew signal tristate
rlabel metal2 s 18234 0 18290 800 6 chany_bottom_out[12]
port 115 nsew signal tristate
rlabel metal2 s 18602 0 18658 800 6 chany_bottom_out[13]
port 116 nsew signal tristate
rlabel metal2 s 19062 0 19118 800 6 chany_bottom_out[14]
port 117 nsew signal tristate
rlabel metal2 s 19522 0 19578 800 6 chany_bottom_out[15]
port 118 nsew signal tristate
rlabel metal2 s 19982 0 20038 800 6 chany_bottom_out[16]
port 119 nsew signal tristate
rlabel metal2 s 20442 0 20498 800 6 chany_bottom_out[17]
port 120 nsew signal tristate
rlabel metal2 s 20902 0 20958 800 6 chany_bottom_out[18]
port 121 nsew signal tristate
rlabel metal2 s 21362 0 21418 800 6 chany_bottom_out[19]
port 122 nsew signal tristate
rlabel metal2 s 13266 0 13322 800 6 chany_bottom_out[1]
port 123 nsew signal tristate
rlabel metal2 s 13726 0 13782 800 6 chany_bottom_out[2]
port 124 nsew signal tristate
rlabel metal2 s 14094 0 14150 800 6 chany_bottom_out[3]
port 125 nsew signal tristate
rlabel metal2 s 14554 0 14610 800 6 chany_bottom_out[4]
port 126 nsew signal tristate
rlabel metal2 s 15014 0 15070 800 6 chany_bottom_out[5]
port 127 nsew signal tristate
rlabel metal2 s 15474 0 15530 800 6 chany_bottom_out[6]
port 128 nsew signal tristate
rlabel metal2 s 15934 0 15990 800 6 chany_bottom_out[7]
port 129 nsew signal tristate
rlabel metal2 s 16394 0 16450 800 6 chany_bottom_out[8]
port 130 nsew signal tristate
rlabel metal2 s 16854 0 16910 800 6 chany_bottom_out[9]
port 131 nsew signal tristate
rlabel metal3 s 0 144 800 264 6 left_bottom_grid_pin_34_
port 132 nsew signal input
rlabel metal3 s 0 552 800 672 6 left_bottom_grid_pin_35_
port 133 nsew signal input
rlabel metal3 s 0 960 800 1080 6 left_bottom_grid_pin_36_
port 134 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 left_bottom_grid_pin_37_
port 135 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 left_bottom_grid_pin_38_
port 136 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 left_bottom_grid_pin_39_
port 137 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 left_bottom_grid_pin_40_
port 138 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 left_bottom_grid_pin_41_
port 139 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 left_top_grid_pin_1_
port 140 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 prog_clk_0_S_in
port 141 nsew signal input
rlabel metal3 s 22200 144 23000 264 6 right_bottom_grid_pin_34_
port 142 nsew signal input
rlabel metal3 s 22200 552 23000 672 6 right_bottom_grid_pin_35_
port 143 nsew signal input
rlabel metal3 s 22200 960 23000 1080 6 right_bottom_grid_pin_36_
port 144 nsew signal input
rlabel metal3 s 22200 1504 23000 1624 6 right_bottom_grid_pin_37_
port 145 nsew signal input
rlabel metal3 s 22200 1912 23000 2032 6 right_bottom_grid_pin_38_
port 146 nsew signal input
rlabel metal3 s 22200 2456 23000 2576 6 right_bottom_grid_pin_39_
port 147 nsew signal input
rlabel metal3 s 22200 2864 23000 2984 6 right_bottom_grid_pin_40_
port 148 nsew signal input
rlabel metal3 s 22200 3408 23000 3528 6 right_bottom_grid_pin_41_
port 149 nsew signal input
rlabel metal3 s 22200 22584 23000 22704 6 right_top_grid_pin_1_
port 150 nsew signal input
rlabel metal4 s 18271 2128 18591 20720 6 VPWR
port 151 nsew power bidirectional
rlabel metal4 s 11340 2128 11660 20720 6 VPWR
port 152 nsew power bidirectional
rlabel metal4 s 4409 2128 4729 20720 6 VPWR
port 153 nsew power bidirectional
rlabel metal4 s 14805 2128 15125 20720 6 VGND
port 154 nsew ground bidirectional
rlabel metal4 s 7875 2128 8195 20720 6 VGND
port 155 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
