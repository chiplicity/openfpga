magic
tech sky130A
magscale 1 2
timestamp 1609019112
<< locali >>
rect 2973 19159 3007 19261
rect 9045 13855 9079 14025
rect 8309 12699 8343 12937
rect 4905 12087 4939 12257
rect 4445 6103 4479 6273
rect 3893 5559 3927 5797
rect 7515 5729 7607 5763
rect 7573 5627 7607 5729
rect 7849 5015 7883 5321
rect 15485 5083 15519 5185
rect 16497 5015 16531 5321
rect 22017 4199 22051 4981
rect 9505 3587 9539 3689
rect 9505 3553 9597 3587
rect 2145 2839 2179 2941
rect 8125 2839 8159 2941
<< viali >>
rect 1961 20553 1995 20587
rect 2513 20553 2547 20587
rect 1777 20349 1811 20383
rect 2329 20349 2363 20383
rect 2605 20009 2639 20043
rect 3157 20009 3191 20043
rect 1869 19873 1903 19907
rect 2421 19873 2455 19907
rect 2973 19873 3007 19907
rect 2053 19737 2087 19771
rect 1961 19397 1995 19431
rect 2513 19329 2547 19363
rect 3249 19329 3283 19363
rect 1777 19261 1811 19295
rect 2329 19261 2363 19295
rect 2973 19261 3007 19295
rect 3065 19261 3099 19295
rect 2973 19125 3007 19159
rect 1961 18921 1995 18955
rect 10793 18921 10827 18955
rect 2605 18853 2639 18887
rect 3341 18853 3375 18887
rect 1777 18785 1811 18819
rect 2339 18785 2373 18819
rect 3065 18785 3099 18819
rect 10609 18785 10643 18819
rect 2789 18241 2823 18275
rect 11069 18241 11103 18275
rect 1777 18173 1811 18207
rect 2605 18173 2639 18207
rect 10885 18173 10919 18207
rect 1961 18037 1995 18071
rect 1869 17833 1903 17867
rect 8033 17833 8067 17867
rect 9689 17833 9723 17867
rect 11437 17833 11471 17867
rect 2513 17765 2547 17799
rect 3249 17765 3283 17799
rect 5356 17765 5390 17799
rect 1685 17697 1719 17731
rect 2226 17697 2260 17731
rect 2973 17697 3007 17731
rect 8401 17697 8435 17731
rect 10057 17697 10091 17731
rect 10701 17697 10735 17731
rect 11805 17697 11839 17731
rect 5089 17629 5123 17663
rect 8493 17629 8527 17663
rect 8677 17629 8711 17663
rect 10149 17629 10183 17663
rect 10333 17629 10367 17663
rect 11897 17629 11931 17663
rect 12081 17629 12115 17663
rect 6469 17493 6503 17527
rect 1961 17289 1995 17323
rect 6837 17289 6871 17323
rect 2605 17153 2639 17187
rect 3341 17153 3375 17187
rect 7389 17153 7423 17187
rect 8217 17153 8251 17187
rect 12449 17153 12483 17187
rect 1777 17085 1811 17119
rect 2421 17085 2455 17119
rect 3157 17085 3191 17119
rect 4169 17085 4203 17119
rect 8677 17085 8711 17119
rect 10333 17085 10367 17119
rect 4436 17017 4470 17051
rect 5825 17017 5859 17051
rect 7205 17017 7239 17051
rect 8944 17017 8978 17051
rect 10578 17017 10612 17051
rect 5549 16949 5583 16983
rect 6285 16949 6319 16983
rect 7297 16949 7331 16983
rect 7849 16949 7883 16983
rect 10057 16949 10091 16983
rect 11713 16949 11747 16983
rect 2973 16745 3007 16779
rect 5457 16745 5491 16779
rect 9321 16745 9355 16779
rect 9689 16745 9723 16779
rect 12081 16745 12115 16779
rect 13737 16745 13771 16779
rect 2329 16677 2363 16711
rect 3341 16677 3375 16711
rect 6184 16677 6218 16711
rect 10057 16677 10091 16711
rect 10946 16677 10980 16711
rect 12602 16677 12636 16711
rect 2053 16609 2087 16643
rect 4344 16609 4378 16643
rect 7573 16609 7607 16643
rect 7941 16609 7975 16643
rect 8208 16609 8242 16643
rect 12357 16609 12391 16643
rect 3433 16541 3467 16575
rect 3617 16541 3651 16575
rect 4077 16541 4111 16575
rect 5917 16541 5951 16575
rect 10149 16541 10183 16575
rect 10241 16541 10275 16575
rect 10701 16541 10735 16575
rect 7297 16405 7331 16439
rect 1961 16201 1995 16235
rect 2513 16201 2547 16235
rect 4353 16201 4387 16235
rect 5733 16201 5767 16235
rect 10149 16201 10183 16235
rect 11345 16201 11379 16235
rect 4629 16065 4663 16099
rect 6285 16065 6319 16099
rect 7757 16065 7791 16099
rect 8769 16065 8803 16099
rect 11989 16065 12023 16099
rect 1777 15997 1811 16031
rect 2329 15997 2363 16031
rect 2973 15997 3007 16031
rect 11069 15997 11103 16031
rect 11713 15997 11747 16031
rect 3240 15929 3274 15963
rect 6193 15929 6227 15963
rect 9036 15929 9070 15963
rect 10609 15929 10643 15963
rect 5089 15861 5123 15895
rect 6101 15861 6135 15895
rect 6837 15861 6871 15895
rect 7205 15861 7239 15895
rect 7573 15861 7607 15895
rect 7665 15861 7699 15895
rect 8217 15861 8251 15895
rect 11805 15861 11839 15895
rect 12449 15861 12483 15895
rect 1685 15657 1719 15691
rect 4077 15657 4111 15691
rect 8493 15657 8527 15691
rect 10057 15657 10091 15691
rect 2329 15589 2363 15623
rect 5641 15589 5675 15623
rect 5733 15589 5767 15623
rect 6828 15589 6862 15623
rect 8861 15589 8895 15623
rect 1501 15521 1535 15555
rect 2053 15521 2087 15555
rect 4445 15521 4479 15555
rect 4537 15521 4571 15555
rect 4629 15453 4663 15487
rect 5825 15453 5859 15487
rect 6561 15453 6595 15487
rect 8953 15453 8987 15487
rect 9045 15453 9079 15487
rect 9781 15385 9815 15419
rect 3709 15317 3743 15351
rect 5273 15317 5307 15351
rect 7941 15317 7975 15351
rect 1869 15113 1903 15147
rect 2973 15113 3007 15147
rect 6285 15113 6319 15147
rect 8309 15113 8343 15147
rect 9045 15113 9079 15147
rect 4629 15045 4663 15079
rect 6837 15045 6871 15079
rect 2421 14977 2455 15011
rect 3617 14977 3651 15011
rect 7297 14977 7331 15011
rect 7481 14977 7515 15011
rect 9597 14977 9631 15011
rect 1685 14909 1719 14943
rect 2247 14909 2281 14943
rect 3433 14909 3467 14943
rect 4905 14909 4939 14943
rect 3341 14841 3375 14875
rect 3985 14841 4019 14875
rect 5172 14841 5206 14875
rect 7205 14841 7239 14875
rect 7849 14841 7883 14875
rect 9413 14841 9447 14875
rect 10057 14841 10091 14875
rect 9505 14773 9539 14807
rect 3249 14569 3283 14603
rect 5825 14569 5859 14603
rect 11437 14569 11471 14603
rect 7196 14501 7230 14535
rect 1777 14433 1811 14467
rect 2339 14433 2373 14467
rect 3065 14433 3099 14467
rect 4712 14433 4746 14467
rect 6929 14433 6963 14467
rect 10057 14433 10091 14467
rect 10324 14433 10358 14467
rect 2513 14365 2547 14399
rect 4445 14365 4479 14399
rect 1961 14229 1995 14263
rect 8309 14229 8343 14263
rect 11713 14229 11747 14263
rect 3249 14025 3283 14059
rect 5365 14025 5399 14059
rect 5641 14025 5675 14059
rect 9045 14025 9079 14059
rect 10977 14025 11011 14059
rect 11253 14025 11287 14059
rect 7757 13957 7791 13991
rect 1869 13889 1903 13923
rect 6193 13889 6227 13923
rect 8309 13889 8343 13923
rect 9229 13889 9263 13923
rect 9597 13889 9631 13923
rect 11805 13889 11839 13923
rect 1593 13821 1627 13855
rect 2339 13821 2373 13855
rect 3065 13821 3099 13855
rect 3985 13821 4019 13855
rect 7389 13821 7423 13855
rect 8125 13821 8159 13855
rect 8953 13821 8987 13855
rect 9045 13821 9079 13855
rect 11621 13821 11655 13855
rect 2605 13753 2639 13787
rect 4252 13753 4286 13787
rect 6101 13753 6135 13787
rect 8217 13753 8251 13787
rect 9864 13753 9898 13787
rect 6009 13685 6043 13719
rect 8769 13685 8803 13719
rect 11713 13685 11747 13719
rect 3525 13481 3559 13515
rect 4537 13481 4571 13515
rect 11345 13481 11379 13515
rect 2145 13413 2179 13447
rect 2881 13413 2915 13447
rect 7288 13413 7322 13447
rect 1869 13345 1903 13379
rect 2605 13345 2639 13379
rect 3341 13345 3375 13379
rect 4261 13345 4295 13379
rect 5457 13345 5491 13379
rect 7021 13345 7055 13379
rect 9965 13345 9999 13379
rect 10232 13345 10266 13379
rect 5549 13277 5583 13311
rect 5641 13277 5675 13311
rect 8677 13277 8711 13311
rect 9137 13277 9171 13311
rect 5089 13209 5123 13243
rect 6101 13141 6135 13175
rect 8401 13141 8435 13175
rect 11713 13141 11747 13175
rect 2237 12937 2271 12971
rect 5549 12937 5583 12971
rect 7021 12937 7055 12971
rect 7481 12937 7515 12971
rect 8309 12937 8343 12971
rect 8493 12937 8527 12971
rect 10609 12937 10643 12971
rect 2881 12801 2915 12835
rect 3433 12801 3467 12835
rect 8125 12801 8159 12835
rect 3249 12733 3283 12767
rect 4169 12733 4203 12767
rect 6009 12733 6043 12767
rect 7205 12733 7239 12767
rect 9045 12801 9079 12835
rect 10241 12801 10275 12835
rect 11161 12801 11195 12835
rect 8953 12733 8987 12767
rect 9965 12733 9999 12767
rect 10057 12733 10091 12767
rect 11621 12733 11655 12767
rect 4436 12665 4470 12699
rect 7849 12665 7883 12699
rect 8309 12665 8343 12699
rect 8861 12665 8895 12699
rect 11069 12665 11103 12699
rect 2605 12597 2639 12631
rect 2697 12597 2731 12631
rect 5825 12597 5859 12631
rect 6469 12597 6503 12631
rect 7941 12597 7975 12631
rect 9597 12597 9631 12631
rect 10977 12597 11011 12631
rect 1593 12393 1627 12427
rect 4077 12393 4111 12427
rect 8861 12393 8895 12427
rect 11253 12393 11287 12427
rect 20269 12393 20303 12427
rect 4537 12325 4571 12359
rect 7104 12325 7138 12359
rect 1409 12257 1443 12291
rect 1961 12257 1995 12291
rect 2228 12257 2262 12291
rect 4445 12257 4479 12291
rect 4905 12257 4939 12291
rect 5089 12257 5123 12291
rect 5356 12257 5390 12291
rect 9873 12257 9907 12291
rect 10140 12257 10174 12291
rect 19717 12257 19751 12291
rect 4721 12189 4755 12223
rect 6837 12189 6871 12223
rect 3341 12053 3375 12087
rect 4905 12053 4939 12087
rect 6469 12053 6503 12087
rect 8217 12053 8251 12087
rect 9229 12053 9263 12087
rect 19901 12053 19935 12087
rect 2053 11849 2087 11883
rect 7021 11849 7055 11883
rect 10977 11849 11011 11883
rect 9597 11781 9631 11815
rect 9965 11781 9999 11815
rect 2697 11713 2731 11747
rect 4721 11713 4755 11747
rect 7665 11713 7699 11747
rect 8217 11713 8251 11747
rect 10517 11713 10551 11747
rect 11437 11713 11471 11747
rect 11529 11713 11563 11747
rect 3065 11645 3099 11679
rect 3332 11645 3366 11679
rect 8473 11645 8507 11679
rect 10425 11645 10459 11679
rect 19257 11645 19291 11679
rect 19809 11645 19843 11679
rect 1777 11577 1811 11611
rect 11345 11577 11379 11611
rect 12449 11577 12483 11611
rect 2421 11509 2455 11543
rect 2513 11509 2547 11543
rect 4445 11509 4479 11543
rect 7389 11509 7423 11543
rect 7481 11509 7515 11543
rect 10333 11509 10367 11543
rect 19441 11509 19475 11543
rect 2329 11305 2363 11339
rect 2789 11305 2823 11339
rect 3157 11305 3191 11339
rect 6009 11305 6043 11339
rect 8769 11305 8803 11339
rect 11069 11305 11103 11339
rect 2053 11237 2087 11271
rect 6653 11237 6687 11271
rect 9934 11237 9968 11271
rect 4896 11169 4930 11203
rect 6377 11169 6411 11203
rect 7380 11169 7414 11203
rect 9689 11169 9723 11203
rect 11529 11169 11563 11203
rect 18797 11169 18831 11203
rect 19349 11169 19383 11203
rect 3249 11101 3283 11135
rect 3341 11101 3375 11135
rect 4629 11101 4663 11135
rect 7113 11101 7147 11135
rect 4077 11033 4111 11067
rect 8493 11033 8527 11067
rect 9321 11033 9355 11067
rect 11345 11033 11379 11067
rect 18981 11033 19015 11067
rect 3065 10761 3099 10795
rect 5457 10761 5491 10795
rect 5733 10761 5767 10795
rect 7389 10761 7423 10795
rect 8401 10761 8435 10795
rect 9965 10761 9999 10795
rect 12909 10761 12943 10795
rect 11621 10693 11655 10727
rect 18521 10693 18555 10727
rect 6285 10625 6319 10659
rect 7849 10625 7883 10659
rect 8033 10625 8067 10659
rect 9505 10625 9539 10659
rect 1685 10557 1719 10591
rect 4077 10557 4111 10591
rect 4344 10557 4378 10591
rect 7021 10557 7055 10591
rect 7757 10557 7791 10591
rect 8585 10557 8619 10591
rect 13093 10557 13127 10591
rect 18337 10557 18371 10591
rect 18889 10557 18923 10591
rect 1952 10489 1986 10523
rect 10333 10489 10367 10523
rect 3801 10421 3835 10455
rect 6101 10421 6135 10455
rect 6193 10421 6227 10455
rect 8953 10421 8987 10455
rect 9321 10421 9355 10455
rect 9413 10421 9447 10455
rect 12541 10421 12575 10455
rect 4169 10217 4203 10251
rect 4629 10217 4663 10251
rect 7389 10217 7423 10251
rect 7849 10217 7883 10251
rect 9689 10217 9723 10251
rect 10701 10217 10735 10251
rect 2053 10149 2087 10183
rect 2789 10149 2823 10183
rect 6101 10149 6135 10183
rect 6653 10149 6687 10183
rect 8769 10149 8803 10183
rect 2697 10081 2731 10115
rect 3341 10081 3375 10115
rect 4997 10081 5031 10115
rect 5089 10081 5123 10115
rect 6009 10081 6043 10115
rect 7021 10081 7055 10115
rect 7757 10081 7791 10115
rect 8861 10081 8895 10115
rect 10057 10081 10091 10115
rect 10885 10081 10919 10115
rect 11428 10081 11462 10115
rect 2881 10013 2915 10047
rect 5181 10013 5215 10047
rect 6193 10013 6227 10047
rect 8033 10013 8067 10047
rect 9045 10013 9079 10047
rect 10149 10013 10183 10047
rect 10333 10013 10367 10047
rect 11161 10013 11195 10047
rect 5641 9945 5675 9979
rect 2329 9877 2363 9911
rect 8401 9877 8435 9911
rect 12541 9877 12575 9911
rect 2973 9605 3007 9639
rect 3249 9605 3283 9639
rect 4537 9605 4571 9639
rect 15209 9605 15243 9639
rect 3801 9537 3835 9571
rect 5181 9537 5215 9571
rect 11437 9537 11471 9571
rect 11621 9537 11655 9571
rect 13001 9537 13035 9571
rect 13829 9537 13863 9571
rect 1593 9469 1627 9503
rect 1860 9469 1894 9503
rect 3617 9469 3651 9503
rect 6837 9469 6871 9503
rect 9321 9469 9355 9503
rect 11345 9469 11379 9503
rect 4997 9401 5031 9435
rect 7104 9401 7138 9435
rect 8953 9401 8987 9435
rect 9588 9401 9622 9435
rect 12909 9401 12943 9435
rect 14096 9401 14130 9435
rect 3709 9333 3743 9367
rect 4905 9333 4939 9367
rect 5549 9333 5583 9367
rect 5917 9333 5951 9367
rect 8217 9333 8251 9367
rect 8493 9333 8527 9367
rect 10701 9333 10735 9367
rect 10977 9333 11011 9367
rect 12449 9333 12483 9367
rect 12817 9333 12851 9367
rect 2421 9129 2455 9163
rect 4537 9129 4571 9163
rect 7757 9129 7791 9163
rect 8125 9129 8159 9163
rect 8769 9129 8803 9163
rect 9689 9129 9723 9163
rect 11161 9129 11195 9163
rect 8217 9061 8251 9095
rect 11980 9061 12014 9095
rect 2789 8993 2823 9027
rect 4905 8993 4939 9027
rect 5816 8993 5850 9027
rect 7389 8993 7423 9027
rect 10057 8993 10091 9027
rect 14473 8993 14507 9027
rect 2881 8925 2915 8959
rect 3065 8925 3099 8959
rect 4997 8925 5031 8959
rect 5181 8925 5215 8959
rect 5549 8925 5583 8959
rect 8401 8925 8435 8959
rect 10149 8925 10183 8959
rect 10333 8925 10367 8959
rect 11713 8925 11747 8959
rect 14565 8925 14599 8959
rect 14657 8925 14691 8959
rect 4169 8857 4203 8891
rect 6929 8789 6963 8823
rect 7205 8789 7239 8823
rect 9229 8789 9263 8823
rect 10793 8789 10827 8823
rect 13093 8789 13127 8823
rect 14105 8789 14139 8823
rect 3341 8585 3375 8619
rect 5641 8585 5675 8619
rect 8401 8585 8435 8619
rect 11621 8585 11655 8619
rect 14841 8585 14875 8619
rect 4261 8449 4295 8483
rect 5917 8449 5951 8483
rect 7021 8449 7055 8483
rect 9505 8449 9539 8483
rect 12449 8449 12483 8483
rect 15117 8449 15151 8483
rect 1961 8381 1995 8415
rect 4528 8381 4562 8415
rect 7288 8381 7322 8415
rect 10609 8381 10643 8415
rect 11805 8381 11839 8415
rect 13461 8381 13495 8415
rect 16865 8381 16899 8415
rect 2228 8313 2262 8347
rect 13728 8313 13762 8347
rect 17141 8313 17175 8347
rect 1593 8245 1627 8279
rect 1961 8041 1995 8075
rect 2973 8041 3007 8075
rect 4445 8041 4479 8075
rect 4905 8041 4939 8075
rect 5457 8041 5491 8075
rect 7389 8041 7423 8075
rect 8953 8041 8987 8075
rect 13553 8041 13587 8075
rect 13829 8041 13863 8075
rect 5825 7973 5859 8007
rect 14197 7973 14231 8007
rect 14841 7973 14875 8007
rect 2329 7905 2363 7939
rect 3341 7905 3375 7939
rect 3433 7905 3467 7939
rect 4813 7905 4847 7939
rect 7757 7905 7791 7939
rect 8861 7905 8895 7939
rect 10517 7905 10551 7939
rect 10784 7905 10818 7939
rect 12429 7905 12463 7939
rect 15301 7905 15335 7939
rect 16589 7905 16623 7939
rect 1685 7837 1719 7871
rect 2421 7837 2455 7871
rect 2513 7837 2547 7871
rect 3617 7837 3651 7871
rect 5089 7837 5123 7871
rect 5917 7837 5951 7871
rect 6101 7837 6135 7871
rect 7849 7837 7883 7871
rect 8033 7837 8067 7871
rect 9045 7837 9079 7871
rect 12173 7837 12207 7871
rect 14289 7837 14323 7871
rect 14473 7837 14507 7871
rect 15485 7837 15519 7871
rect 16865 7837 16899 7871
rect 6653 7769 6687 7803
rect 4169 7701 4203 7735
rect 7113 7701 7147 7735
rect 8493 7701 8527 7735
rect 11897 7701 11931 7735
rect 3157 7497 3191 7531
rect 4537 7497 4571 7531
rect 5273 7497 5307 7531
rect 5733 7497 5767 7531
rect 9045 7497 9079 7531
rect 17509 7497 17543 7531
rect 3801 7361 3835 7395
rect 6285 7361 6319 7395
rect 11621 7361 11655 7395
rect 1777 7293 1811 7327
rect 5457 7293 5491 7327
rect 7205 7293 7239 7327
rect 7665 7293 7699 7327
rect 7932 7293 7966 7327
rect 9321 7293 9355 7327
rect 9577 7293 9611 7327
rect 11989 7293 12023 7327
rect 14105 7293 14139 7327
rect 16129 7293 16163 7327
rect 2044 7225 2078 7259
rect 4997 7225 5031 7259
rect 6193 7225 6227 7259
rect 11437 7225 11471 7259
rect 14372 7225 14406 7259
rect 16396 7225 16430 7259
rect 3433 7157 3467 7191
rect 6101 7157 6135 7191
rect 7021 7157 7055 7191
rect 10701 7157 10735 7191
rect 10977 7157 11011 7191
rect 11345 7157 11379 7191
rect 12449 7157 12483 7191
rect 13001 7157 13035 7191
rect 13645 7157 13679 7191
rect 15485 7157 15519 7191
rect 5733 6953 5767 6987
rect 8861 6953 8895 6987
rect 11529 6953 11563 6987
rect 13645 6953 13679 6987
rect 2329 6885 2363 6919
rect 3341 6885 3375 6919
rect 10425 6885 10459 6919
rect 14565 6885 14599 6919
rect 3433 6817 3467 6851
rect 4344 6817 4378 6851
rect 6101 6817 6135 6851
rect 10885 6817 10919 6851
rect 11621 6817 11655 6851
rect 12725 6817 12759 6851
rect 13553 6817 13587 6851
rect 15301 6817 15335 6851
rect 16681 6817 16715 6851
rect 17325 6817 17359 6851
rect 2421 6749 2455 6783
rect 2605 6749 2639 6783
rect 3617 6749 3651 6783
rect 4077 6749 4111 6783
rect 11805 6749 11839 6783
rect 12265 6749 12299 6783
rect 13829 6749 13863 6783
rect 14657 6749 14691 6783
rect 14841 6749 14875 6783
rect 15485 6749 15519 6783
rect 16773 6749 16807 6783
rect 16957 6749 16991 6783
rect 1685 6681 1719 6715
rect 2973 6681 3007 6715
rect 11161 6681 11195 6715
rect 13185 6681 13219 6715
rect 17785 6681 17819 6715
rect 1961 6613 1995 6647
rect 5457 6613 5491 6647
rect 8493 6613 8527 6647
rect 10701 6613 10735 6647
rect 12541 6613 12575 6647
rect 14197 6613 14231 6647
rect 16313 6613 16347 6647
rect 2789 6409 2823 6443
rect 13829 6409 13863 6443
rect 15485 6409 15519 6443
rect 17417 6409 17451 6443
rect 9965 6341 9999 6375
rect 11897 6341 11931 6375
rect 3065 6273 3099 6307
rect 4261 6273 4295 6307
rect 4445 6273 4479 6307
rect 7481 6273 7515 6307
rect 18613 6273 18647 6307
rect 1409 6205 1443 6239
rect 1676 6205 1710 6239
rect 4629 6205 4663 6239
rect 6377 6205 6411 6239
rect 7297 6205 7331 6239
rect 8309 6205 8343 6239
rect 10517 6205 10551 6239
rect 12449 6205 12483 6239
rect 12705 6205 12739 6239
rect 14105 6205 14139 6239
rect 14361 6205 14395 6239
rect 16037 6205 16071 6239
rect 18429 6205 18463 6239
rect 4896 6137 4930 6171
rect 7205 6137 7239 6171
rect 7849 6137 7883 6171
rect 8554 6137 8588 6171
rect 10762 6137 10796 6171
rect 16304 6137 16338 6171
rect 3617 6069 3651 6103
rect 3985 6069 4019 6103
rect 4077 6069 4111 6103
rect 4445 6069 4479 6103
rect 6009 6069 6043 6103
rect 6837 6069 6871 6103
rect 9689 6069 9723 6103
rect 18061 6069 18095 6103
rect 18521 6069 18555 6103
rect 1961 5865 1995 5899
rect 2329 5865 2363 5899
rect 2421 5865 2455 5899
rect 2973 5865 3007 5899
rect 3433 5865 3467 5899
rect 11345 5865 11379 5899
rect 12817 5865 12851 5899
rect 15301 5865 15335 5899
rect 3341 5797 3375 5831
rect 3893 5797 3927 5831
rect 6276 5797 6310 5831
rect 9956 5797 9990 5831
rect 11713 5797 11747 5831
rect 11805 5797 11839 5831
rect 2513 5661 2547 5695
rect 3617 5661 3651 5695
rect 4445 5729 4479 5763
rect 6009 5729 6043 5763
rect 7481 5729 7515 5763
rect 7932 5729 7966 5763
rect 9689 5729 9723 5763
rect 12725 5729 12759 5763
rect 14289 5729 14323 5763
rect 15945 5729 15979 5763
rect 16856 5729 16890 5763
rect 4537 5661 4571 5695
rect 4721 5661 4755 5695
rect 7665 5661 7699 5695
rect 11897 5661 11931 5695
rect 13001 5661 13035 5695
rect 14473 5661 14507 5695
rect 16589 5661 16623 5695
rect 7389 5593 7423 5627
rect 7573 5593 7607 5627
rect 3893 5525 3927 5559
rect 4077 5525 4111 5559
rect 5089 5525 5123 5559
rect 9045 5525 9079 5559
rect 11069 5525 11103 5559
rect 12357 5525 12391 5559
rect 13369 5525 13403 5559
rect 15761 5525 15795 5559
rect 17969 5525 18003 5559
rect 3525 5321 3559 5355
rect 7849 5321 7883 5355
rect 11897 5321 11931 5355
rect 16497 5321 16531 5355
rect 16589 5321 16623 5355
rect 7021 5253 7055 5287
rect 6377 5185 6411 5219
rect 7573 5185 7607 5219
rect 3893 5117 3927 5151
rect 6101 5117 6135 5151
rect 6193 5049 6227 5083
rect 9321 5253 9355 5287
rect 8493 5185 8527 5219
rect 8677 5185 8711 5219
rect 9965 5185 9999 5219
rect 10793 5185 10827 5219
rect 10977 5185 11011 5219
rect 12449 5185 12483 5219
rect 13645 5185 13679 5219
rect 15485 5185 15519 5219
rect 16221 5185 16255 5219
rect 9689 5117 9723 5151
rect 14565 5117 14599 5151
rect 10701 5049 10735 5083
rect 11345 5049 11379 5083
rect 14841 5049 14875 5083
rect 15485 5049 15519 5083
rect 15945 5049 15979 5083
rect 17233 5185 17267 5219
rect 19993 5185 20027 5219
rect 16957 5117 16991 5151
rect 17601 5117 17635 5151
rect 20260 5117 20294 5151
rect 4261 4981 4295 5015
rect 5733 4981 5767 5015
rect 7389 4981 7423 5015
rect 7481 4981 7515 5015
rect 7849 4981 7883 5015
rect 8033 4981 8067 5015
rect 8401 4981 8435 5015
rect 9781 4981 9815 5015
rect 10333 4981 10367 5015
rect 13185 4981 13219 5015
rect 15577 4981 15611 5015
rect 16037 4981 16071 5015
rect 16497 4981 16531 5015
rect 17049 4981 17083 5015
rect 18061 4981 18095 5015
rect 21373 4981 21407 5015
rect 22017 4981 22051 5015
rect 1501 4777 1535 4811
rect 1869 4777 1903 4811
rect 3249 4777 3283 4811
rect 4537 4777 4571 4811
rect 6745 4777 6779 4811
rect 7113 4777 7147 4811
rect 14841 4777 14875 4811
rect 18061 4777 18095 4811
rect 21281 4777 21315 4811
rect 2329 4709 2363 4743
rect 7481 4709 7515 4743
rect 8585 4709 8619 4743
rect 10784 4709 10818 4743
rect 15485 4709 15519 4743
rect 2237 4641 2271 4675
rect 5641 4641 5675 4675
rect 8125 4641 8159 4675
rect 10149 4641 10183 4675
rect 13084 4641 13118 4675
rect 15945 4641 15979 4675
rect 16212 4641 16246 4675
rect 17969 4641 18003 4675
rect 2513 4573 2547 4607
rect 3341 4573 3375 4607
rect 3433 4573 3467 4607
rect 5733 4573 5767 4607
rect 5917 4573 5951 4607
rect 6377 4573 6411 4607
rect 7573 4573 7607 4607
rect 7665 4573 7699 4607
rect 9137 4573 9171 4607
rect 10517 4573 10551 4607
rect 12817 4573 12851 4607
rect 18153 4573 18187 4607
rect 17325 4505 17359 4539
rect 2881 4437 2915 4471
rect 4905 4437 4939 4471
rect 5273 4437 5307 4471
rect 9689 4437 9723 4471
rect 11897 4437 11931 4471
rect 14197 4437 14231 4471
rect 17601 4437 17635 4471
rect 3341 4233 3375 4267
rect 5273 4233 5307 4267
rect 8217 4233 8251 4267
rect 17141 4233 17175 4267
rect 4997 4165 5031 4199
rect 22017 4165 22051 4199
rect 1501 4097 1535 4131
rect 5733 4097 5767 4131
rect 5825 4097 5859 4131
rect 6285 4097 6319 4131
rect 6837 4097 6871 4131
rect 9505 4097 9539 4131
rect 10425 4097 10459 4131
rect 11437 4097 11471 4131
rect 11621 4097 11655 4131
rect 15761 4097 15795 4131
rect 17417 4097 17451 4131
rect 1961 4029 1995 4063
rect 3617 4029 3651 4063
rect 3873 4029 3907 4063
rect 5641 4029 5675 4063
rect 9229 4029 9263 4063
rect 12449 4029 12483 4063
rect 12705 4029 12739 4063
rect 14105 4029 14139 4063
rect 14361 4029 14395 4063
rect 2228 3961 2262 3995
rect 7082 3961 7116 3995
rect 9321 3961 9355 3995
rect 10333 3961 10367 3995
rect 16006 3961 16040 3995
rect 8493 3893 8527 3927
rect 8861 3893 8895 3927
rect 9873 3893 9907 3927
rect 10241 3893 10275 3927
rect 10977 3893 11011 3927
rect 11345 3893 11379 3927
rect 11989 3893 12023 3927
rect 13829 3893 13863 3927
rect 15485 3893 15519 3927
rect 21373 3893 21407 3927
rect 4077 3689 4111 3723
rect 6561 3689 6595 3723
rect 9505 3689 9539 3723
rect 10149 3689 10183 3723
rect 11069 3689 11103 3723
rect 11437 3689 11471 3723
rect 13185 3689 13219 3723
rect 14197 3689 14231 3723
rect 13277 3621 13311 3655
rect 1501 3553 1535 3587
rect 1768 3553 1802 3587
rect 3157 3553 3191 3587
rect 4445 3553 4479 3587
rect 5181 3553 5215 3587
rect 5448 3553 5482 3587
rect 7205 3553 7239 3587
rect 7297 3553 7331 3587
rect 7941 3553 7975 3587
rect 8208 3553 8242 3587
rect 9597 3553 9631 3587
rect 10057 3553 10091 3587
rect 11989 3553 12023 3587
rect 15301 3553 15335 3587
rect 15853 3553 15887 3587
rect 16773 3553 16807 3587
rect 17509 3553 17543 3587
rect 19717 3553 19751 3587
rect 20085 3553 20119 3587
rect 20913 3553 20947 3587
rect 3433 3485 3467 3519
rect 4537 3485 4571 3519
rect 4629 3485 4663 3519
rect 7481 3485 7515 3519
rect 10333 3485 10367 3519
rect 12265 3485 12299 3519
rect 13461 3485 13495 3519
rect 14289 3485 14323 3519
rect 14381 3485 14415 3519
rect 17049 3485 17083 3519
rect 2881 3417 2915 3451
rect 14841 3417 14875 3451
rect 6837 3349 6871 3383
rect 9321 3349 9355 3383
rect 9689 3349 9723 3383
rect 10701 3349 10735 3383
rect 12817 3349 12851 3383
rect 13829 3349 13863 3383
rect 15485 3349 15519 3383
rect 16037 3349 16071 3383
rect 17693 3349 17727 3383
rect 20269 3349 20303 3383
rect 21097 3349 21131 3383
rect 2329 3145 2363 3179
rect 10149 3145 10183 3179
rect 15209 3077 15243 3111
rect 2881 3009 2915 3043
rect 4997 3009 5031 3043
rect 7481 3009 7515 3043
rect 8769 3009 8803 3043
rect 10977 3009 11011 3043
rect 14749 3009 14783 3043
rect 15669 3009 15703 3043
rect 15853 3009 15887 3043
rect 20729 3009 20763 3043
rect 1961 2941 1995 2975
rect 2145 2941 2179 2975
rect 3341 2941 3375 2975
rect 3608 2941 3642 2975
rect 5264 2941 5298 2975
rect 8125 2941 8159 2975
rect 9036 2941 9070 2975
rect 11437 2941 11471 2975
rect 12449 2941 12483 2975
rect 13185 2941 13219 2975
rect 13921 2941 13955 2975
rect 14473 2941 14507 2975
rect 16221 2941 16255 2975
rect 16957 2941 16991 2975
rect 18061 2941 18095 2975
rect 18613 2941 18647 2975
rect 20545 2941 20579 2975
rect 2697 2873 2731 2907
rect 7297 2873 7331 2907
rect 7389 2873 7423 2907
rect 10793 2873 10827 2907
rect 11713 2873 11747 2907
rect 12725 2873 12759 2907
rect 13461 2873 13495 2907
rect 15577 2873 15611 2907
rect 16497 2873 16531 2907
rect 17233 2873 17267 2907
rect 1593 2805 1627 2839
rect 2145 2805 2179 2839
rect 2789 2805 2823 2839
rect 4721 2805 4755 2839
rect 6377 2805 6411 2839
rect 6929 2805 6963 2839
rect 7941 2805 7975 2839
rect 8125 2805 8159 2839
rect 8309 2805 8343 2839
rect 10425 2805 10459 2839
rect 10885 2805 10919 2839
rect 14105 2805 14139 2839
rect 18245 2805 18279 2839
rect 18797 2805 18831 2839
rect 2789 2601 2823 2635
rect 5825 2601 5859 2635
rect 6193 2601 6227 2635
rect 6285 2601 6319 2635
rect 6929 2601 6963 2635
rect 7297 2601 7331 2635
rect 8401 2601 8435 2635
rect 9137 2601 9171 2635
rect 9781 2601 9815 2635
rect 10241 2601 10275 2635
rect 16957 2601 16991 2635
rect 7389 2533 7423 2567
rect 9045 2533 9079 2567
rect 10149 2533 10183 2567
rect 3157 2465 3191 2499
rect 4077 2465 4111 2499
rect 11897 2465 11931 2499
rect 12633 2465 12667 2499
rect 13185 2465 13219 2499
rect 13737 2465 13771 2499
rect 14289 2465 14323 2499
rect 14841 2465 14875 2499
rect 15485 2465 15519 2499
rect 16405 2465 16439 2499
rect 17417 2465 17451 2499
rect 3249 2397 3283 2431
rect 3433 2397 3467 2431
rect 6469 2397 6503 2431
rect 7481 2397 7515 2431
rect 9321 2397 9355 2431
rect 10333 2397 10367 2431
rect 8677 2329 8711 2363
rect 2421 2261 2455 2295
rect 7941 2261 7975 2295
rect 11253 2261 11287 2295
rect 12081 2261 12115 2295
rect 12817 2261 12851 2295
rect 13369 2261 13403 2295
rect 13921 2261 13955 2295
rect 14473 2261 14507 2295
rect 15025 2261 15059 2295
rect 15669 2261 15703 2295
rect 16589 2261 16623 2295
rect 17601 2261 17635 2295
rect 21373 2261 21407 2295
<< metal1 >>
rect 3694 21768 3700 21820
rect 3752 21808 3758 21820
rect 10778 21808 10784 21820
rect 3752 21780 10784 21808
rect 3752 21768 3758 21780
rect 10778 21768 10784 21780
rect 10836 21768 10842 21820
rect 1104 20698 21896 20720
rect 1104 20646 4447 20698
rect 4499 20646 4511 20698
rect 4563 20646 4575 20698
rect 4627 20646 4639 20698
rect 4691 20646 11378 20698
rect 11430 20646 11442 20698
rect 11494 20646 11506 20698
rect 11558 20646 11570 20698
rect 11622 20646 18308 20698
rect 18360 20646 18372 20698
rect 18424 20646 18436 20698
rect 18488 20646 18500 20698
rect 18552 20646 21896 20698
rect 1104 20624 21896 20646
rect 1946 20584 1952 20596
rect 1907 20556 1952 20584
rect 1946 20544 1952 20556
rect 2004 20544 2010 20596
rect 2501 20587 2559 20593
rect 2501 20553 2513 20587
rect 2547 20584 2559 20587
rect 2774 20584 2780 20596
rect 2547 20556 2780 20584
rect 2547 20553 2559 20556
rect 2501 20547 2559 20553
rect 2774 20544 2780 20556
rect 2832 20544 2838 20596
rect 1765 20383 1823 20389
rect 1765 20349 1777 20383
rect 1811 20349 1823 20383
rect 1765 20343 1823 20349
rect 2317 20383 2375 20389
rect 2317 20349 2329 20383
rect 2363 20380 2375 20383
rect 2590 20380 2596 20392
rect 2363 20352 2596 20380
rect 2363 20349 2375 20352
rect 2317 20343 2375 20349
rect 1780 20312 1808 20343
rect 2590 20340 2596 20352
rect 2648 20340 2654 20392
rect 3234 20312 3240 20324
rect 1780 20284 3240 20312
rect 3234 20272 3240 20284
rect 3292 20272 3298 20324
rect 1104 20154 21896 20176
rect 1104 20102 7912 20154
rect 7964 20102 7976 20154
rect 8028 20102 8040 20154
rect 8092 20102 8104 20154
rect 8156 20102 14843 20154
rect 14895 20102 14907 20154
rect 14959 20102 14971 20154
rect 15023 20102 15035 20154
rect 15087 20102 21896 20154
rect 1104 20080 21896 20102
rect 2593 20043 2651 20049
rect 2593 20009 2605 20043
rect 2639 20040 2651 20043
rect 2774 20040 2780 20052
rect 2639 20012 2780 20040
rect 2639 20009 2651 20012
rect 2593 20003 2651 20009
rect 2774 20000 2780 20012
rect 2832 20000 2838 20052
rect 3142 20040 3148 20052
rect 3103 20012 3148 20040
rect 3142 20000 3148 20012
rect 3200 20000 3206 20052
rect 1857 19907 1915 19913
rect 1857 19873 1869 19907
rect 1903 19873 1915 19907
rect 1857 19867 1915 19873
rect 2409 19907 2467 19913
rect 2409 19873 2421 19907
rect 2455 19904 2467 19907
rect 2498 19904 2504 19916
rect 2455 19876 2504 19904
rect 2455 19873 2467 19876
rect 2409 19867 2467 19873
rect 1872 19836 1900 19867
rect 2498 19864 2504 19876
rect 2556 19864 2562 19916
rect 2958 19904 2964 19916
rect 2919 19876 2964 19904
rect 2958 19864 2964 19876
rect 3016 19864 3022 19916
rect 2774 19836 2780 19848
rect 1872 19808 2780 19836
rect 2774 19796 2780 19808
rect 2832 19796 2838 19848
rect 2038 19768 2044 19780
rect 1999 19740 2044 19768
rect 2038 19728 2044 19740
rect 2096 19728 2102 19780
rect 1104 19610 21896 19632
rect 1104 19558 4447 19610
rect 4499 19558 4511 19610
rect 4563 19558 4575 19610
rect 4627 19558 4639 19610
rect 4691 19558 11378 19610
rect 11430 19558 11442 19610
rect 11494 19558 11506 19610
rect 11558 19558 11570 19610
rect 11622 19558 18308 19610
rect 18360 19558 18372 19610
rect 18424 19558 18436 19610
rect 18488 19558 18500 19610
rect 18552 19558 21896 19610
rect 1104 19536 21896 19558
rect 1946 19428 1952 19440
rect 1907 19400 1952 19428
rect 1946 19388 1952 19400
rect 2004 19388 2010 19440
rect 2498 19360 2504 19372
rect 2459 19332 2504 19360
rect 2498 19320 2504 19332
rect 2556 19320 2562 19372
rect 3234 19360 3240 19372
rect 3195 19332 3240 19360
rect 3234 19320 3240 19332
rect 3292 19320 3298 19372
rect 1765 19295 1823 19301
rect 1765 19261 1777 19295
rect 1811 19261 1823 19295
rect 1765 19255 1823 19261
rect 2317 19295 2375 19301
rect 2317 19261 2329 19295
rect 2363 19292 2375 19295
rect 2961 19295 3019 19301
rect 2961 19292 2973 19295
rect 2363 19264 2973 19292
rect 2363 19261 2375 19264
rect 2317 19255 2375 19261
rect 2961 19261 2973 19264
rect 3007 19261 3019 19295
rect 2961 19255 3019 19261
rect 3053 19295 3111 19301
rect 3053 19261 3065 19295
rect 3099 19292 3111 19295
rect 8938 19292 8944 19304
rect 3099 19264 8944 19292
rect 3099 19261 3111 19264
rect 3053 19255 3111 19261
rect 1780 19224 1808 19255
rect 8938 19252 8944 19264
rect 8996 19252 9002 19304
rect 3234 19224 3240 19236
rect 1780 19196 3240 19224
rect 3234 19184 3240 19196
rect 3292 19184 3298 19236
rect 2961 19159 3019 19165
rect 2961 19125 2973 19159
rect 3007 19156 3019 19159
rect 10594 19156 10600 19168
rect 3007 19128 10600 19156
rect 3007 19125 3019 19128
rect 2961 19119 3019 19125
rect 10594 19116 10600 19128
rect 10652 19116 10658 19168
rect 1104 19066 21896 19088
rect 1104 19014 7912 19066
rect 7964 19014 7976 19066
rect 8028 19014 8040 19066
rect 8092 19014 8104 19066
rect 8156 19014 14843 19066
rect 14895 19014 14907 19066
rect 14959 19014 14971 19066
rect 15023 19014 15035 19066
rect 15087 19014 21896 19066
rect 1104 18992 21896 19014
rect 1946 18952 1952 18964
rect 1907 18924 1952 18952
rect 1946 18912 1952 18924
rect 2004 18912 2010 18964
rect 10778 18952 10784 18964
rect 10739 18924 10784 18952
rect 10778 18912 10784 18924
rect 10836 18912 10842 18964
rect 2590 18884 2596 18896
rect 2551 18856 2596 18884
rect 2590 18844 2596 18856
rect 2648 18844 2654 18896
rect 2958 18844 2964 18896
rect 3016 18884 3022 18896
rect 3329 18887 3387 18893
rect 3329 18884 3341 18887
rect 3016 18856 3341 18884
rect 3016 18844 3022 18856
rect 3329 18853 3341 18856
rect 3375 18853 3387 18887
rect 3329 18847 3387 18853
rect 1762 18816 1768 18828
rect 1723 18788 1768 18816
rect 1762 18776 1768 18788
rect 1820 18776 1826 18828
rect 2327 18819 2385 18825
rect 2327 18785 2339 18819
rect 2373 18785 2385 18819
rect 2327 18779 2385 18785
rect 3053 18819 3111 18825
rect 3053 18785 3065 18819
rect 3099 18816 3111 18819
rect 9674 18816 9680 18828
rect 3099 18788 9680 18816
rect 3099 18785 3111 18788
rect 3053 18779 3111 18785
rect 2332 18748 2360 18779
rect 9674 18776 9680 18788
rect 9732 18776 9738 18828
rect 10597 18819 10655 18825
rect 10597 18785 10609 18819
rect 10643 18816 10655 18819
rect 11054 18816 11060 18828
rect 10643 18788 11060 18816
rect 10643 18785 10655 18788
rect 10597 18779 10655 18785
rect 11054 18776 11060 18788
rect 11112 18776 11118 18828
rect 5626 18748 5632 18760
rect 2332 18720 5632 18748
rect 5626 18708 5632 18720
rect 5684 18708 5690 18760
rect 1104 18522 21896 18544
rect 1104 18470 4447 18522
rect 4499 18470 4511 18522
rect 4563 18470 4575 18522
rect 4627 18470 4639 18522
rect 4691 18470 11378 18522
rect 11430 18470 11442 18522
rect 11494 18470 11506 18522
rect 11558 18470 11570 18522
rect 11622 18470 18308 18522
rect 18360 18470 18372 18522
rect 18424 18470 18436 18522
rect 18488 18470 18500 18522
rect 18552 18470 21896 18522
rect 1104 18448 21896 18470
rect 2774 18232 2780 18284
rect 2832 18272 2838 18284
rect 11054 18272 11060 18284
rect 2832 18244 2877 18272
rect 11015 18244 11060 18272
rect 2832 18232 2838 18244
rect 11054 18232 11060 18244
rect 11112 18232 11118 18284
rect 1765 18207 1823 18213
rect 1765 18173 1777 18207
rect 1811 18173 1823 18207
rect 1765 18167 1823 18173
rect 2593 18207 2651 18213
rect 2593 18173 2605 18207
rect 2639 18204 2651 18207
rect 2682 18204 2688 18216
rect 2639 18176 2688 18204
rect 2639 18173 2651 18176
rect 2593 18167 2651 18173
rect 1780 18136 1808 18167
rect 2682 18164 2688 18176
rect 2740 18164 2746 18216
rect 10873 18207 10931 18213
rect 10873 18173 10885 18207
rect 10919 18204 10931 18207
rect 11422 18204 11428 18216
rect 10919 18176 11428 18204
rect 10919 18173 10931 18176
rect 10873 18167 10931 18173
rect 11422 18164 11428 18176
rect 11480 18164 11486 18216
rect 3326 18136 3332 18148
rect 1780 18108 3332 18136
rect 3326 18096 3332 18108
rect 3384 18096 3390 18148
rect 1946 18068 1952 18080
rect 1907 18040 1952 18068
rect 1946 18028 1952 18040
rect 2004 18028 2010 18080
rect 1104 17978 21896 18000
rect 1104 17926 7912 17978
rect 7964 17926 7976 17978
rect 8028 17926 8040 17978
rect 8092 17926 8104 17978
rect 8156 17926 14843 17978
rect 14895 17926 14907 17978
rect 14959 17926 14971 17978
rect 15023 17926 15035 17978
rect 15087 17926 21896 17978
rect 1104 17904 21896 17926
rect 1854 17864 1860 17876
rect 1815 17836 1860 17864
rect 1854 17824 1860 17836
rect 1912 17824 1918 17876
rect 5626 17824 5632 17876
rect 5684 17864 5690 17876
rect 8021 17867 8079 17873
rect 8021 17864 8033 17867
rect 5684 17836 8033 17864
rect 5684 17824 5690 17836
rect 8021 17833 8033 17836
rect 8067 17833 8079 17867
rect 9674 17864 9680 17876
rect 9635 17836 9680 17864
rect 8021 17827 8079 17833
rect 9674 17824 9680 17836
rect 9732 17824 9738 17876
rect 11422 17864 11428 17876
rect 11383 17836 11428 17864
rect 11422 17824 11428 17836
rect 11480 17824 11486 17876
rect 1762 17756 1768 17808
rect 1820 17796 1826 17808
rect 2501 17799 2559 17805
rect 2501 17796 2513 17799
rect 1820 17768 2513 17796
rect 1820 17756 1826 17768
rect 2501 17765 2513 17768
rect 2547 17765 2559 17799
rect 3234 17796 3240 17808
rect 3195 17768 3240 17796
rect 2501 17759 2559 17765
rect 3234 17756 3240 17768
rect 3292 17756 3298 17808
rect 5344 17799 5402 17805
rect 5344 17765 5356 17799
rect 5390 17796 5402 17799
rect 5534 17796 5540 17808
rect 5390 17768 5540 17796
rect 5390 17765 5402 17768
rect 5344 17759 5402 17765
rect 5534 17756 5540 17768
rect 5592 17756 5598 17808
rect 1670 17728 1676 17740
rect 1631 17700 1676 17728
rect 1670 17688 1676 17700
rect 1728 17688 1734 17740
rect 2214 17731 2272 17737
rect 2214 17697 2226 17731
rect 2260 17697 2272 17731
rect 2214 17691 2272 17697
rect 2961 17731 3019 17737
rect 2961 17697 2973 17731
rect 3007 17728 3019 17731
rect 7558 17728 7564 17740
rect 3007 17700 7564 17728
rect 3007 17697 3019 17700
rect 2961 17691 3019 17697
rect 2231 17524 2259 17691
rect 7558 17688 7564 17700
rect 7616 17688 7622 17740
rect 8202 17688 8208 17740
rect 8260 17728 8266 17740
rect 8389 17731 8447 17737
rect 8389 17728 8401 17731
rect 8260 17700 8401 17728
rect 8260 17688 8266 17700
rect 8389 17697 8401 17700
rect 8435 17697 8447 17731
rect 8389 17691 8447 17697
rect 10045 17731 10103 17737
rect 10045 17697 10057 17731
rect 10091 17728 10103 17731
rect 10689 17731 10747 17737
rect 10689 17728 10701 17731
rect 10091 17700 10701 17728
rect 10091 17697 10103 17700
rect 10045 17691 10103 17697
rect 10689 17697 10701 17700
rect 10735 17697 10747 17731
rect 10689 17691 10747 17697
rect 11793 17731 11851 17737
rect 11793 17697 11805 17731
rect 11839 17728 11851 17731
rect 12434 17728 12440 17740
rect 11839 17700 12440 17728
rect 11839 17697 11851 17700
rect 11793 17691 11851 17697
rect 12434 17688 12440 17700
rect 12492 17688 12498 17740
rect 4062 17620 4068 17672
rect 4120 17660 4126 17672
rect 5077 17663 5135 17669
rect 5077 17660 5089 17663
rect 4120 17632 5089 17660
rect 4120 17620 4126 17632
rect 5077 17629 5089 17632
rect 5123 17629 5135 17663
rect 8478 17660 8484 17672
rect 8439 17632 8484 17660
rect 5077 17623 5135 17629
rect 8478 17620 8484 17632
rect 8536 17620 8542 17672
rect 8665 17663 8723 17669
rect 8665 17629 8677 17663
rect 8711 17660 8723 17663
rect 9306 17660 9312 17672
rect 8711 17632 9312 17660
rect 8711 17629 8723 17632
rect 8665 17623 8723 17629
rect 9306 17620 9312 17632
rect 9364 17620 9370 17672
rect 9674 17620 9680 17672
rect 9732 17660 9738 17672
rect 10137 17663 10195 17669
rect 10137 17660 10149 17663
rect 9732 17632 10149 17660
rect 9732 17620 9738 17632
rect 10137 17629 10149 17632
rect 10183 17629 10195 17663
rect 10318 17660 10324 17672
rect 10279 17632 10324 17660
rect 10137 17623 10195 17629
rect 10318 17620 10324 17632
rect 10376 17620 10382 17672
rect 11882 17660 11888 17672
rect 11843 17632 11888 17660
rect 11882 17620 11888 17632
rect 11940 17620 11946 17672
rect 12069 17663 12127 17669
rect 12069 17629 12081 17663
rect 12115 17660 12127 17663
rect 13722 17660 13728 17672
rect 12115 17632 13728 17660
rect 12115 17629 12127 17632
rect 12069 17623 12127 17629
rect 13722 17620 13728 17632
rect 13780 17620 13786 17672
rect 8386 17592 8392 17604
rect 6012 17564 8392 17592
rect 6012 17524 6040 17564
rect 8386 17552 8392 17564
rect 8444 17552 8450 17604
rect 6454 17524 6460 17536
rect 2231 17496 6040 17524
rect 6415 17496 6460 17524
rect 6454 17484 6460 17496
rect 6512 17484 6518 17536
rect 1104 17434 21896 17456
rect 1104 17382 4447 17434
rect 4499 17382 4511 17434
rect 4563 17382 4575 17434
rect 4627 17382 4639 17434
rect 4691 17382 11378 17434
rect 11430 17382 11442 17434
rect 11494 17382 11506 17434
rect 11558 17382 11570 17434
rect 11622 17382 18308 17434
rect 18360 17382 18372 17434
rect 18424 17382 18436 17434
rect 18488 17382 18500 17434
rect 18552 17382 21896 17434
rect 1104 17360 21896 17382
rect 1946 17320 1952 17332
rect 1907 17292 1952 17320
rect 1946 17280 1952 17292
rect 2004 17280 2010 17332
rect 6825 17323 6883 17329
rect 6825 17320 6837 17323
rect 3160 17292 6837 17320
rect 2593 17187 2651 17193
rect 2593 17184 2605 17187
rect 1780 17156 2605 17184
rect 1780 17125 1808 17156
rect 2593 17153 2605 17156
rect 2639 17153 2651 17187
rect 2593 17147 2651 17153
rect 1765 17119 1823 17125
rect 1765 17085 1777 17119
rect 1811 17085 1823 17119
rect 1765 17079 1823 17085
rect 2409 17119 2467 17125
rect 2409 17085 2421 17119
rect 2455 17116 2467 17119
rect 2958 17116 2964 17128
rect 2455 17088 2964 17116
rect 2455 17085 2467 17088
rect 2409 17079 2467 17085
rect 2958 17076 2964 17088
rect 3016 17076 3022 17128
rect 3160 17125 3188 17292
rect 6825 17289 6837 17292
rect 6871 17289 6883 17323
rect 6825 17283 6883 17289
rect 3326 17184 3332 17196
rect 3287 17156 3332 17184
rect 3326 17144 3332 17156
rect 3384 17144 3390 17196
rect 6454 17144 6460 17196
rect 6512 17184 6518 17196
rect 7377 17187 7435 17193
rect 7377 17184 7389 17187
rect 6512 17156 7389 17184
rect 6512 17144 6518 17156
rect 7377 17153 7389 17156
rect 7423 17153 7435 17187
rect 8202 17184 8208 17196
rect 8163 17156 8208 17184
rect 7377 17147 7435 17153
rect 8202 17144 8208 17156
rect 8260 17144 8266 17196
rect 12434 17184 12440 17196
rect 12395 17156 12440 17184
rect 12434 17144 12440 17156
rect 12492 17144 12498 17196
rect 3145 17119 3203 17125
rect 3145 17085 3157 17119
rect 3191 17085 3203 17119
rect 3145 17079 3203 17085
rect 4062 17076 4068 17128
rect 4120 17116 4126 17128
rect 4157 17119 4215 17125
rect 4157 17116 4169 17119
rect 4120 17088 4169 17116
rect 4120 17076 4126 17088
rect 4157 17085 4169 17088
rect 4203 17116 4215 17119
rect 5718 17116 5724 17128
rect 4203 17088 5724 17116
rect 4203 17085 4215 17088
rect 4157 17079 4215 17085
rect 5718 17076 5724 17088
rect 5776 17076 5782 17128
rect 8665 17119 8723 17125
rect 8665 17085 8677 17119
rect 8711 17116 8723 17119
rect 8754 17116 8760 17128
rect 8711 17088 8760 17116
rect 8711 17085 8723 17088
rect 8665 17079 8723 17085
rect 8754 17076 8760 17088
rect 8812 17116 8818 17128
rect 10321 17119 10379 17125
rect 10321 17116 10333 17119
rect 8812 17088 10333 17116
rect 8812 17076 8818 17088
rect 10321 17085 10333 17088
rect 10367 17085 10379 17119
rect 10321 17079 10379 17085
rect 4424 17051 4482 17057
rect 4424 17048 4436 17051
rect 4172 17020 4436 17048
rect 4172 16992 4200 17020
rect 4424 17017 4436 17020
rect 4470 17048 4482 17051
rect 5442 17048 5448 17060
rect 4470 17020 5448 17048
rect 4470 17017 4482 17020
rect 4424 17011 4482 17017
rect 5442 17008 5448 17020
rect 5500 17008 5506 17060
rect 5813 17051 5871 17057
rect 5813 17017 5825 17051
rect 5859 17048 5871 17051
rect 7193 17051 7251 17057
rect 7193 17048 7205 17051
rect 5859 17020 7205 17048
rect 5859 17017 5871 17020
rect 5813 17011 5871 17017
rect 7193 17017 7205 17020
rect 7239 17017 7251 17051
rect 7193 17011 7251 17017
rect 8932 17051 8990 17057
rect 8932 17017 8944 17051
rect 8978 17048 8990 17051
rect 9306 17048 9312 17060
rect 8978 17020 9312 17048
rect 8978 17017 8990 17020
rect 8932 17011 8990 17017
rect 9306 17008 9312 17020
rect 9364 17008 9370 17060
rect 10226 17048 10232 17060
rect 10060 17020 10232 17048
rect 4154 16940 4160 16992
rect 4212 16940 4218 16992
rect 5534 16980 5540 16992
rect 5495 16952 5540 16980
rect 5534 16940 5540 16952
rect 5592 16940 5598 16992
rect 6270 16980 6276 16992
rect 6231 16952 6276 16980
rect 6270 16940 6276 16952
rect 6328 16940 6334 16992
rect 6914 16940 6920 16992
rect 6972 16980 6978 16992
rect 7285 16983 7343 16989
rect 7285 16980 7297 16983
rect 6972 16952 7297 16980
rect 6972 16940 6978 16952
rect 7285 16949 7297 16952
rect 7331 16949 7343 16983
rect 7285 16943 7343 16949
rect 7466 16940 7472 16992
rect 7524 16980 7530 16992
rect 10060 16989 10088 17020
rect 10226 17008 10232 17020
rect 10284 17048 10290 17060
rect 10566 17051 10624 17057
rect 10566 17048 10578 17051
rect 10284 17020 10578 17048
rect 10284 17008 10290 17020
rect 10566 17017 10578 17020
rect 10612 17017 10624 17051
rect 10566 17011 10624 17017
rect 7837 16983 7895 16989
rect 7837 16980 7849 16983
rect 7524 16952 7849 16980
rect 7524 16940 7530 16952
rect 7837 16949 7849 16952
rect 7883 16949 7895 16983
rect 7837 16943 7895 16949
rect 10045 16983 10103 16989
rect 10045 16949 10057 16983
rect 10091 16949 10103 16983
rect 10045 16943 10103 16949
rect 10318 16940 10324 16992
rect 10376 16980 10382 16992
rect 11701 16983 11759 16989
rect 11701 16980 11713 16983
rect 10376 16952 11713 16980
rect 10376 16940 10382 16952
rect 11701 16949 11713 16952
rect 11747 16949 11759 16983
rect 11701 16943 11759 16949
rect 1104 16890 21896 16912
rect 1104 16838 7912 16890
rect 7964 16838 7976 16890
rect 8028 16838 8040 16890
rect 8092 16838 8104 16890
rect 8156 16838 14843 16890
rect 14895 16838 14907 16890
rect 14959 16838 14971 16890
rect 15023 16838 15035 16890
rect 15087 16838 21896 16890
rect 1104 16816 21896 16838
rect 2958 16776 2964 16788
rect 2919 16748 2964 16776
rect 2958 16736 2964 16748
rect 3016 16736 3022 16788
rect 5442 16776 5448 16788
rect 3252 16748 4384 16776
rect 5403 16748 5448 16776
rect 1670 16668 1676 16720
rect 1728 16708 1734 16720
rect 2317 16711 2375 16717
rect 2317 16708 2329 16711
rect 1728 16680 2329 16708
rect 1728 16668 1734 16680
rect 2317 16677 2329 16680
rect 2363 16677 2375 16711
rect 2317 16671 2375 16677
rect 2041 16643 2099 16649
rect 2041 16609 2053 16643
rect 2087 16640 2099 16643
rect 3252 16640 3280 16748
rect 3329 16711 3387 16717
rect 3329 16677 3341 16711
rect 3375 16708 3387 16711
rect 4246 16708 4252 16720
rect 3375 16680 4252 16708
rect 3375 16677 3387 16680
rect 3329 16671 3387 16677
rect 4246 16668 4252 16680
rect 4304 16668 4310 16720
rect 4356 16708 4384 16748
rect 5442 16736 5448 16748
rect 5500 16736 5506 16788
rect 6270 16736 6276 16788
rect 6328 16776 6334 16788
rect 9306 16776 9312 16788
rect 6328 16748 8892 16776
rect 9267 16748 9312 16776
rect 6328 16736 6334 16748
rect 5902 16708 5908 16720
rect 4356 16680 5908 16708
rect 5902 16668 5908 16680
rect 5960 16668 5966 16720
rect 6172 16711 6230 16717
rect 6172 16677 6184 16711
rect 6218 16708 6230 16711
rect 6454 16708 6460 16720
rect 6218 16680 6460 16708
rect 6218 16677 6230 16680
rect 6172 16671 6230 16677
rect 6454 16668 6460 16680
rect 6512 16668 6518 16720
rect 8754 16708 8760 16720
rect 7944 16680 8760 16708
rect 4154 16640 4160 16652
rect 2087 16612 3280 16640
rect 3896 16612 4160 16640
rect 2087 16609 2099 16612
rect 2041 16603 2099 16609
rect 3418 16572 3424 16584
rect 3379 16544 3424 16572
rect 3418 16532 3424 16544
rect 3476 16532 3482 16584
rect 3605 16575 3663 16581
rect 3605 16541 3617 16575
rect 3651 16572 3663 16575
rect 3896 16572 3924 16612
rect 4154 16600 4160 16612
rect 4212 16600 4218 16652
rect 4338 16649 4344 16652
rect 4332 16603 4344 16649
rect 4396 16640 4402 16652
rect 4396 16612 4432 16640
rect 4338 16600 4344 16603
rect 4396 16600 4402 16612
rect 5718 16600 5724 16652
rect 5776 16640 5782 16652
rect 5776 16612 5948 16640
rect 5776 16600 5782 16612
rect 4062 16572 4068 16584
rect 3651 16544 3924 16572
rect 4023 16544 4068 16572
rect 3651 16541 3663 16544
rect 3605 16535 3663 16541
rect 4062 16532 4068 16544
rect 4120 16532 4126 16584
rect 5920 16581 5948 16612
rect 7006 16600 7012 16652
rect 7064 16640 7070 16652
rect 7944 16649 7972 16680
rect 8754 16668 8760 16680
rect 8812 16668 8818 16720
rect 8864 16708 8892 16748
rect 9306 16736 9312 16748
rect 9364 16736 9370 16788
rect 9674 16776 9680 16788
rect 9635 16748 9680 16776
rect 9674 16736 9680 16748
rect 9732 16736 9738 16788
rect 12069 16779 12127 16785
rect 12069 16745 12081 16779
rect 12115 16745 12127 16779
rect 13722 16776 13728 16788
rect 13635 16748 13728 16776
rect 12069 16739 12127 16745
rect 10042 16708 10048 16720
rect 8864 16680 10048 16708
rect 10042 16668 10048 16680
rect 10100 16668 10106 16720
rect 10318 16668 10324 16720
rect 10376 16708 10382 16720
rect 10934 16711 10992 16717
rect 10934 16708 10946 16711
rect 10376 16680 10946 16708
rect 10376 16668 10382 16680
rect 10934 16677 10946 16680
rect 10980 16677 10992 16711
rect 10934 16671 10992 16677
rect 11974 16668 11980 16720
rect 12032 16708 12038 16720
rect 12084 16708 12112 16739
rect 13722 16736 13728 16748
rect 13780 16776 13786 16788
rect 19242 16776 19248 16788
rect 13780 16748 19248 16776
rect 13780 16736 13786 16748
rect 19242 16736 19248 16748
rect 19300 16736 19306 16788
rect 12590 16711 12648 16717
rect 12590 16708 12602 16711
rect 12032 16680 12602 16708
rect 12032 16668 12038 16680
rect 12590 16677 12602 16680
rect 12636 16677 12648 16711
rect 12590 16671 12648 16677
rect 7561 16643 7619 16649
rect 7561 16640 7573 16643
rect 7064 16612 7573 16640
rect 7064 16600 7070 16612
rect 7561 16609 7573 16612
rect 7607 16609 7619 16643
rect 7561 16603 7619 16609
rect 7929 16643 7987 16649
rect 7929 16609 7941 16643
rect 7975 16609 7987 16643
rect 7929 16603 7987 16609
rect 8196 16643 8254 16649
rect 8196 16609 8208 16643
rect 8242 16640 8254 16643
rect 9030 16640 9036 16652
rect 8242 16612 9036 16640
rect 8242 16609 8254 16612
rect 8196 16603 8254 16609
rect 9030 16600 9036 16612
rect 9088 16600 9094 16652
rect 12342 16640 12348 16652
rect 12303 16612 12348 16640
rect 12342 16600 12348 16612
rect 12400 16600 12406 16652
rect 5905 16575 5963 16581
rect 5905 16541 5917 16575
rect 5951 16541 5963 16575
rect 10134 16572 10140 16584
rect 10095 16544 10140 16572
rect 5905 16535 5963 16541
rect 10134 16532 10140 16544
rect 10192 16532 10198 16584
rect 10226 16532 10232 16584
rect 10284 16572 10290 16584
rect 10686 16572 10692 16584
rect 10284 16544 10329 16572
rect 10647 16544 10692 16572
rect 10284 16532 10290 16544
rect 10686 16532 10692 16544
rect 10744 16532 10750 16584
rect 7282 16436 7288 16448
rect 7243 16408 7288 16436
rect 7282 16396 7288 16408
rect 7340 16396 7346 16448
rect 1104 16346 21896 16368
rect 1104 16294 4447 16346
rect 4499 16294 4511 16346
rect 4563 16294 4575 16346
rect 4627 16294 4639 16346
rect 4691 16294 11378 16346
rect 11430 16294 11442 16346
rect 11494 16294 11506 16346
rect 11558 16294 11570 16346
rect 11622 16294 18308 16346
rect 18360 16294 18372 16346
rect 18424 16294 18436 16346
rect 18488 16294 18500 16346
rect 18552 16294 21896 16346
rect 1104 16272 21896 16294
rect 1946 16232 1952 16244
rect 1907 16204 1952 16232
rect 1946 16192 1952 16204
rect 2004 16192 2010 16244
rect 2501 16235 2559 16241
rect 2501 16201 2513 16235
rect 2547 16232 2559 16235
rect 2774 16232 2780 16244
rect 2547 16204 2780 16232
rect 2547 16201 2559 16204
rect 2501 16195 2559 16201
rect 2774 16192 2780 16204
rect 2832 16192 2838 16244
rect 4338 16232 4344 16244
rect 4299 16204 4344 16232
rect 4338 16192 4344 16204
rect 4396 16192 4402 16244
rect 5721 16235 5779 16241
rect 5721 16201 5733 16235
rect 5767 16232 5779 16235
rect 6914 16232 6920 16244
rect 5767 16204 6920 16232
rect 5767 16201 5779 16204
rect 5721 16195 5779 16201
rect 6914 16192 6920 16204
rect 6972 16192 6978 16244
rect 9030 16192 9036 16244
rect 9088 16232 9094 16244
rect 10137 16235 10195 16241
rect 10137 16232 10149 16235
rect 9088 16204 10149 16232
rect 9088 16192 9094 16204
rect 10137 16201 10149 16204
rect 10183 16201 10195 16235
rect 10137 16195 10195 16201
rect 11333 16235 11391 16241
rect 11333 16201 11345 16235
rect 11379 16232 11391 16235
rect 11882 16232 11888 16244
rect 11379 16204 11888 16232
rect 11379 16201 11391 16204
rect 11333 16195 11391 16201
rect 11882 16192 11888 16204
rect 11940 16192 11946 16244
rect 4246 16056 4252 16108
rect 4304 16096 4310 16108
rect 4617 16099 4675 16105
rect 4617 16096 4629 16099
rect 4304 16068 4629 16096
rect 4304 16056 4310 16068
rect 4617 16065 4629 16068
rect 4663 16065 4675 16099
rect 4617 16059 4675 16065
rect 5534 16056 5540 16108
rect 5592 16096 5598 16108
rect 6273 16099 6331 16105
rect 6273 16096 6285 16099
rect 5592 16068 6285 16096
rect 5592 16056 5598 16068
rect 6273 16065 6285 16068
rect 6319 16065 6331 16099
rect 6273 16059 6331 16065
rect 7282 16056 7288 16108
rect 7340 16096 7346 16108
rect 7745 16099 7803 16105
rect 7745 16096 7757 16099
rect 7340 16068 7757 16096
rect 7340 16056 7346 16068
rect 7745 16065 7757 16068
rect 7791 16065 7803 16099
rect 8754 16096 8760 16108
rect 8715 16068 8760 16096
rect 7745 16059 7803 16065
rect 8754 16056 8760 16068
rect 8812 16056 8818 16108
rect 11974 16096 11980 16108
rect 11935 16068 11980 16096
rect 11974 16056 11980 16068
rect 12032 16056 12038 16108
rect 1762 16028 1768 16040
rect 1723 16000 1768 16028
rect 1762 15988 1768 16000
rect 1820 15988 1826 16040
rect 2314 16028 2320 16040
rect 2275 16000 2320 16028
rect 2314 15988 2320 16000
rect 2372 15988 2378 16040
rect 2961 16031 3019 16037
rect 2961 15997 2973 16031
rect 3007 16028 3019 16031
rect 4062 16028 4068 16040
rect 3007 16000 4068 16028
rect 3007 15997 3019 16000
rect 2961 15991 3019 15997
rect 4062 15988 4068 16000
rect 4120 15988 4126 16040
rect 11057 16031 11115 16037
rect 11057 16028 11069 16031
rect 7576 16000 11069 16028
rect 3228 15963 3286 15969
rect 3228 15929 3240 15963
rect 3274 15960 3286 15963
rect 3602 15960 3608 15972
rect 3274 15932 3608 15960
rect 3274 15929 3286 15932
rect 3228 15923 3286 15929
rect 3602 15920 3608 15932
rect 3660 15920 3666 15972
rect 6181 15963 6239 15969
rect 6181 15929 6193 15963
rect 6227 15960 6239 15963
rect 7006 15960 7012 15972
rect 6227 15932 7012 15960
rect 6227 15929 6239 15932
rect 6181 15923 6239 15929
rect 7006 15920 7012 15932
rect 7064 15920 7070 15972
rect 4982 15852 4988 15904
rect 5040 15892 5046 15904
rect 5077 15895 5135 15901
rect 5077 15892 5089 15895
rect 5040 15864 5089 15892
rect 5040 15852 5046 15864
rect 5077 15861 5089 15864
rect 5123 15861 5135 15895
rect 5077 15855 5135 15861
rect 6089 15895 6147 15901
rect 6089 15861 6101 15895
rect 6135 15892 6147 15895
rect 6270 15892 6276 15904
rect 6135 15864 6276 15892
rect 6135 15861 6147 15864
rect 6089 15855 6147 15861
rect 6270 15852 6276 15864
rect 6328 15852 6334 15904
rect 6546 15852 6552 15904
rect 6604 15892 6610 15904
rect 6825 15895 6883 15901
rect 6825 15892 6837 15895
rect 6604 15864 6837 15892
rect 6604 15852 6610 15864
rect 6825 15861 6837 15864
rect 6871 15861 6883 15895
rect 7190 15892 7196 15904
rect 7151 15864 7196 15892
rect 6825 15855 6883 15861
rect 7190 15852 7196 15864
rect 7248 15852 7254 15904
rect 7466 15852 7472 15904
rect 7524 15892 7530 15904
rect 7576 15901 7604 16000
rect 11057 15997 11069 16000
rect 11103 16028 11115 16031
rect 11701 16031 11759 16037
rect 11701 16028 11713 16031
rect 11103 16000 11713 16028
rect 11103 15997 11115 16000
rect 11057 15991 11115 15997
rect 11701 15997 11713 16000
rect 11747 15997 11759 16031
rect 11701 15991 11759 15997
rect 9024 15963 9082 15969
rect 9024 15929 9036 15963
rect 9070 15960 9082 15963
rect 9582 15960 9588 15972
rect 9070 15932 9588 15960
rect 9070 15929 9082 15932
rect 9024 15923 9082 15929
rect 9582 15920 9588 15932
rect 9640 15920 9646 15972
rect 10134 15920 10140 15972
rect 10192 15960 10198 15972
rect 10597 15963 10655 15969
rect 10597 15960 10609 15963
rect 10192 15932 10609 15960
rect 10192 15920 10198 15932
rect 10597 15929 10609 15932
rect 10643 15960 10655 15963
rect 11974 15960 11980 15972
rect 10643 15932 11980 15960
rect 10643 15929 10655 15932
rect 10597 15923 10655 15929
rect 11974 15920 11980 15932
rect 12032 15920 12038 15972
rect 7561 15895 7619 15901
rect 7561 15892 7573 15895
rect 7524 15864 7573 15892
rect 7524 15852 7530 15864
rect 7561 15861 7573 15864
rect 7607 15861 7619 15895
rect 7561 15855 7619 15861
rect 7650 15852 7656 15904
rect 7708 15892 7714 15904
rect 8205 15895 8263 15901
rect 8205 15892 8217 15895
rect 7708 15864 8217 15892
rect 7708 15852 7714 15864
rect 8205 15861 8217 15864
rect 8251 15861 8263 15895
rect 8205 15855 8263 15861
rect 11793 15895 11851 15901
rect 11793 15861 11805 15895
rect 11839 15892 11851 15895
rect 12434 15892 12440 15904
rect 11839 15864 12440 15892
rect 11839 15861 11851 15864
rect 11793 15855 11851 15861
rect 12434 15852 12440 15864
rect 12492 15852 12498 15904
rect 1104 15802 21896 15824
rect 1104 15750 7912 15802
rect 7964 15750 7976 15802
rect 8028 15750 8040 15802
rect 8092 15750 8104 15802
rect 8156 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 15035 15802
rect 15087 15750 21896 15802
rect 1104 15728 21896 15750
rect 1670 15688 1676 15700
rect 1631 15660 1676 15688
rect 1670 15648 1676 15660
rect 1728 15648 1734 15700
rect 3418 15648 3424 15700
rect 3476 15688 3482 15700
rect 4065 15691 4123 15697
rect 4065 15688 4077 15691
rect 3476 15660 4077 15688
rect 3476 15648 3482 15660
rect 4065 15657 4077 15660
rect 4111 15657 4123 15691
rect 8294 15688 8300 15700
rect 4065 15651 4123 15657
rect 4448 15660 8300 15688
rect 2314 15620 2320 15632
rect 2275 15592 2320 15620
rect 2314 15580 2320 15592
rect 2372 15580 2378 15632
rect 1489 15555 1547 15561
rect 1489 15521 1501 15555
rect 1535 15521 1547 15555
rect 1489 15515 1547 15521
rect 2041 15555 2099 15561
rect 2041 15521 2053 15555
rect 2087 15552 2099 15555
rect 2958 15552 2964 15564
rect 2087 15524 2964 15552
rect 2087 15521 2099 15524
rect 2041 15515 2099 15521
rect 1504 15484 1532 15515
rect 2958 15512 2964 15524
rect 3016 15512 3022 15564
rect 3694 15512 3700 15564
rect 3752 15552 3758 15564
rect 4448 15561 4476 15660
rect 8294 15648 8300 15660
rect 8352 15648 8358 15700
rect 8478 15688 8484 15700
rect 8439 15660 8484 15688
rect 8478 15648 8484 15660
rect 8536 15648 8542 15700
rect 10042 15688 10048 15700
rect 10003 15660 10048 15688
rect 10042 15648 10048 15660
rect 10100 15648 10106 15700
rect 4890 15580 4896 15632
rect 4948 15620 4954 15632
rect 5629 15623 5687 15629
rect 5629 15620 5641 15623
rect 4948 15592 5641 15620
rect 4948 15580 4954 15592
rect 5629 15589 5641 15592
rect 5675 15589 5687 15623
rect 5629 15583 5687 15589
rect 5721 15623 5779 15629
rect 5721 15589 5733 15623
rect 5767 15620 5779 15623
rect 6546 15620 6552 15632
rect 5767 15592 6552 15620
rect 5767 15589 5779 15592
rect 5721 15583 5779 15589
rect 4433 15555 4491 15561
rect 4433 15552 4445 15555
rect 3752 15524 4445 15552
rect 3752 15512 3758 15524
rect 4433 15521 4445 15524
rect 4479 15521 4491 15555
rect 4433 15515 4491 15521
rect 4525 15555 4583 15561
rect 4525 15521 4537 15555
rect 4571 15552 4583 15555
rect 5074 15552 5080 15564
rect 4571 15524 5080 15552
rect 4571 15521 4583 15524
rect 4525 15515 4583 15521
rect 5074 15512 5080 15524
rect 5132 15512 5138 15564
rect 5644 15552 5672 15583
rect 6546 15580 6552 15592
rect 6604 15580 6610 15632
rect 6816 15623 6874 15629
rect 6816 15589 6828 15623
rect 6862 15620 6874 15623
rect 7282 15620 7288 15632
rect 6862 15592 7288 15620
rect 6862 15589 6874 15592
rect 6816 15583 6874 15589
rect 7282 15580 7288 15592
rect 7340 15580 7346 15632
rect 8312 15620 8340 15648
rect 8849 15623 8907 15629
rect 8849 15620 8861 15623
rect 8312 15592 8861 15620
rect 8849 15589 8861 15592
rect 8895 15589 8907 15623
rect 8849 15583 8907 15589
rect 9122 15552 9128 15564
rect 5644 15524 9128 15552
rect 9122 15512 9128 15524
rect 9180 15512 9186 15564
rect 2590 15484 2596 15496
rect 1504 15456 2596 15484
rect 2590 15444 2596 15456
rect 2648 15444 2654 15496
rect 4617 15487 4675 15493
rect 4617 15453 4629 15487
rect 4663 15453 4675 15487
rect 4617 15447 4675 15453
rect 4338 15376 4344 15428
rect 4396 15416 4402 15428
rect 4632 15416 4660 15447
rect 5810 15444 5816 15496
rect 5868 15484 5874 15496
rect 6549 15487 6607 15493
rect 5868 15456 5913 15484
rect 5868 15444 5874 15456
rect 6549 15453 6561 15487
rect 6595 15453 6607 15487
rect 6549 15447 6607 15453
rect 8941 15487 8999 15493
rect 8941 15453 8953 15487
rect 8987 15453 8999 15487
rect 8941 15447 8999 15453
rect 4396 15388 4660 15416
rect 4396 15376 4402 15388
rect 3694 15348 3700 15360
rect 3655 15320 3700 15348
rect 3694 15308 3700 15320
rect 3752 15308 3758 15360
rect 4154 15308 4160 15360
rect 4212 15348 4218 15360
rect 5261 15351 5319 15357
rect 5261 15348 5273 15351
rect 4212 15320 5273 15348
rect 4212 15308 4218 15320
rect 5261 15317 5273 15320
rect 5307 15317 5319 15351
rect 6564 15348 6592 15447
rect 8956 15416 8984 15447
rect 9030 15444 9036 15496
rect 9088 15484 9094 15496
rect 9088 15456 9133 15484
rect 9088 15444 9094 15456
rect 9769 15419 9827 15425
rect 9769 15416 9781 15419
rect 8956 15388 9781 15416
rect 9769 15385 9781 15388
rect 9815 15416 9827 15419
rect 11146 15416 11152 15428
rect 9815 15388 11152 15416
rect 9815 15385 9827 15388
rect 9769 15379 9827 15385
rect 11146 15376 11152 15388
rect 11204 15376 11210 15428
rect 6914 15348 6920 15360
rect 6564 15320 6920 15348
rect 5261 15311 5319 15317
rect 6914 15308 6920 15320
rect 6972 15308 6978 15360
rect 7466 15308 7472 15360
rect 7524 15348 7530 15360
rect 7929 15351 7987 15357
rect 7929 15348 7941 15351
rect 7524 15320 7941 15348
rect 7524 15308 7530 15320
rect 7929 15317 7941 15320
rect 7975 15317 7987 15351
rect 7929 15311 7987 15317
rect 1104 15258 21896 15280
rect 1104 15206 4447 15258
rect 4499 15206 4511 15258
rect 4563 15206 4575 15258
rect 4627 15206 4639 15258
rect 4691 15206 11378 15258
rect 11430 15206 11442 15258
rect 11494 15206 11506 15258
rect 11558 15206 11570 15258
rect 11622 15206 18308 15258
rect 18360 15206 18372 15258
rect 18424 15206 18436 15258
rect 18488 15206 18500 15258
rect 18552 15206 21896 15258
rect 1104 15184 21896 15206
rect 1854 15144 1860 15156
rect 1815 15116 1860 15144
rect 1854 15104 1860 15116
rect 1912 15104 1918 15156
rect 2958 15144 2964 15156
rect 2919 15116 2964 15144
rect 2958 15104 2964 15116
rect 3016 15104 3022 15156
rect 6273 15147 6331 15153
rect 6273 15144 6285 15147
rect 4356 15116 6285 15144
rect 1762 14968 1768 15020
rect 1820 15008 1826 15020
rect 2409 15011 2467 15017
rect 2409 15008 2421 15011
rect 1820 14980 2421 15008
rect 1820 14968 1826 14980
rect 2409 14977 2421 14980
rect 2455 14977 2467 15011
rect 3602 15008 3608 15020
rect 3515 14980 3608 15008
rect 2409 14971 2467 14977
rect 3602 14968 3608 14980
rect 3660 15008 3666 15020
rect 4356 15008 4384 15116
rect 6273 15113 6285 15116
rect 6319 15113 6331 15147
rect 8294 15144 8300 15156
rect 8255 15116 8300 15144
rect 6273 15107 6331 15113
rect 8294 15104 8300 15116
rect 8352 15104 8358 15156
rect 8938 15104 8944 15156
rect 8996 15144 9002 15156
rect 9033 15147 9091 15153
rect 9033 15144 9045 15147
rect 8996 15116 9045 15144
rect 8996 15104 9002 15116
rect 9033 15113 9045 15116
rect 9079 15113 9091 15147
rect 9033 15107 9091 15113
rect 4617 15079 4675 15085
rect 4617 15045 4629 15079
rect 4663 15076 4675 15079
rect 4890 15076 4896 15088
rect 4663 15048 4896 15076
rect 4663 15045 4675 15048
rect 4617 15039 4675 15045
rect 4890 15036 4896 15048
rect 4948 15036 4954 15088
rect 5902 15036 5908 15088
rect 5960 15076 5966 15088
rect 6825 15079 6883 15085
rect 6825 15076 6837 15079
rect 5960 15048 6837 15076
rect 5960 15036 5966 15048
rect 6825 15045 6837 15048
rect 6871 15045 6883 15079
rect 6825 15039 6883 15045
rect 3660 14980 4384 15008
rect 3660 14968 3666 14980
rect 7190 14968 7196 15020
rect 7248 15008 7254 15020
rect 7285 15011 7343 15017
rect 7285 15008 7297 15011
rect 7248 14980 7297 15008
rect 7248 14968 7254 14980
rect 7285 14977 7297 14980
rect 7331 14977 7343 15011
rect 7466 15008 7472 15020
rect 7427 14980 7472 15008
rect 7285 14971 7343 14977
rect 7466 14968 7472 14980
rect 7524 14968 7530 15020
rect 9582 15008 9588 15020
rect 9543 14980 9588 15008
rect 9582 14968 9588 14980
rect 9640 14968 9646 15020
rect 1670 14940 1676 14952
rect 1631 14912 1676 14940
rect 1670 14900 1676 14912
rect 1728 14900 1734 14952
rect 2235 14943 2293 14949
rect 2235 14909 2247 14943
rect 2281 14909 2293 14943
rect 2235 14903 2293 14909
rect 3421 14943 3479 14949
rect 3421 14909 3433 14943
rect 3467 14940 3479 14943
rect 4154 14940 4160 14952
rect 3467 14912 4160 14940
rect 3467 14909 3479 14912
rect 3421 14903 3479 14909
rect 2240 14804 2268 14903
rect 4154 14900 4160 14912
rect 4212 14900 4218 14952
rect 4430 14900 4436 14952
rect 4488 14940 4494 14952
rect 4893 14943 4951 14949
rect 4893 14940 4905 14943
rect 4488 14912 4905 14940
rect 4488 14900 4494 14912
rect 4893 14909 4905 14912
rect 4939 14909 4951 14943
rect 4893 14903 4951 14909
rect 3329 14875 3387 14881
rect 3329 14841 3341 14875
rect 3375 14872 3387 14875
rect 3973 14875 4031 14881
rect 3973 14872 3985 14875
rect 3375 14844 3985 14872
rect 3375 14841 3387 14844
rect 3329 14835 3387 14841
rect 3973 14841 3985 14844
rect 4019 14841 4031 14875
rect 5160 14875 5218 14881
rect 3973 14835 4031 14841
rect 4172 14844 4660 14872
rect 4172 14804 4200 14844
rect 2240 14776 4200 14804
rect 4632 14804 4660 14844
rect 5160 14841 5172 14875
rect 5206 14872 5218 14875
rect 5810 14872 5816 14884
rect 5206 14844 5816 14872
rect 5206 14841 5218 14844
rect 5160 14835 5218 14841
rect 5810 14832 5816 14844
rect 5868 14832 5874 14884
rect 7193 14875 7251 14881
rect 7193 14841 7205 14875
rect 7239 14872 7251 14875
rect 7837 14875 7895 14881
rect 7837 14872 7849 14875
rect 7239 14844 7849 14872
rect 7239 14841 7251 14844
rect 7193 14835 7251 14841
rect 7837 14841 7849 14844
rect 7883 14841 7895 14875
rect 7837 14835 7895 14841
rect 9401 14875 9459 14881
rect 9401 14841 9413 14875
rect 9447 14872 9459 14875
rect 10045 14875 10103 14881
rect 10045 14872 10057 14875
rect 9447 14844 10057 14872
rect 9447 14841 9459 14844
rect 9401 14835 9459 14841
rect 10045 14841 10057 14844
rect 10091 14841 10103 14875
rect 10045 14835 10103 14841
rect 5626 14804 5632 14816
rect 4632 14776 5632 14804
rect 5626 14764 5632 14776
rect 5684 14764 5690 14816
rect 9493 14807 9551 14813
rect 9493 14773 9505 14807
rect 9539 14804 9551 14807
rect 11238 14804 11244 14816
rect 9539 14776 11244 14804
rect 9539 14773 9551 14776
rect 9493 14767 9551 14773
rect 11238 14764 11244 14776
rect 11296 14764 11302 14816
rect 1104 14714 21896 14736
rect 1104 14662 7912 14714
rect 7964 14662 7976 14714
rect 8028 14662 8040 14714
rect 8092 14662 8104 14714
rect 8156 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 15035 14714
rect 15087 14662 21896 14714
rect 1104 14640 21896 14662
rect 3234 14600 3240 14612
rect 3195 14572 3240 14600
rect 3234 14560 3240 14572
rect 3292 14560 3298 14612
rect 5810 14600 5816 14612
rect 5771 14572 5816 14600
rect 5810 14560 5816 14572
rect 5868 14560 5874 14612
rect 9582 14560 9588 14612
rect 9640 14600 9646 14612
rect 11425 14603 11483 14609
rect 11425 14600 11437 14603
rect 9640 14572 11437 14600
rect 9640 14560 9646 14572
rect 11425 14569 11437 14572
rect 11471 14569 11483 14603
rect 11425 14563 11483 14569
rect 7184 14535 7242 14541
rect 2332 14504 5856 14532
rect 1762 14464 1768 14476
rect 1723 14436 1768 14464
rect 1762 14424 1768 14436
rect 1820 14424 1826 14476
rect 2332 14473 2360 14504
rect 5828 14476 5856 14504
rect 7184 14501 7196 14535
rect 7230 14532 7242 14535
rect 7466 14532 7472 14544
rect 7230 14504 7472 14532
rect 7230 14501 7242 14504
rect 7184 14495 7242 14501
rect 7466 14492 7472 14504
rect 7524 14492 7530 14544
rect 2327 14467 2385 14473
rect 2327 14433 2339 14467
rect 2373 14433 2385 14467
rect 2327 14427 2385 14433
rect 2774 14424 2780 14476
rect 2832 14464 2838 14476
rect 3053 14467 3111 14473
rect 3053 14464 3065 14467
rect 2832 14436 3065 14464
rect 2832 14424 2838 14436
rect 3053 14433 3065 14436
rect 3099 14433 3111 14467
rect 3053 14427 3111 14433
rect 4700 14467 4758 14473
rect 4700 14433 4712 14467
rect 4746 14464 4758 14467
rect 5258 14464 5264 14476
rect 4746 14436 5264 14464
rect 4746 14433 4758 14436
rect 4700 14427 4758 14433
rect 5258 14424 5264 14436
rect 5316 14424 5322 14476
rect 5810 14424 5816 14476
rect 5868 14424 5874 14476
rect 6914 14464 6920 14476
rect 6827 14436 6920 14464
rect 6914 14424 6920 14436
rect 6972 14464 6978 14476
rect 8754 14464 8760 14476
rect 6972 14436 8760 14464
rect 6972 14424 6978 14436
rect 8754 14424 8760 14436
rect 8812 14464 8818 14476
rect 9582 14464 9588 14476
rect 8812 14436 9588 14464
rect 8812 14424 8818 14436
rect 9582 14424 9588 14436
rect 9640 14464 9646 14476
rect 10045 14467 10103 14473
rect 10045 14464 10057 14467
rect 9640 14436 10057 14464
rect 9640 14424 9646 14436
rect 10045 14433 10057 14436
rect 10091 14433 10103 14467
rect 10045 14427 10103 14433
rect 10312 14467 10370 14473
rect 10312 14433 10324 14467
rect 10358 14464 10370 14467
rect 10870 14464 10876 14476
rect 10358 14436 10876 14464
rect 10358 14433 10370 14436
rect 10312 14427 10370 14433
rect 10870 14424 10876 14436
rect 10928 14424 10934 14476
rect 1670 14356 1676 14408
rect 1728 14396 1734 14408
rect 2501 14399 2559 14405
rect 2501 14396 2513 14399
rect 1728 14368 2513 14396
rect 1728 14356 1734 14368
rect 2501 14365 2513 14368
rect 2547 14365 2559 14399
rect 2501 14359 2559 14365
rect 4154 14356 4160 14408
rect 4212 14396 4218 14408
rect 4430 14396 4436 14408
rect 4212 14368 4436 14396
rect 4212 14356 4218 14368
rect 4430 14356 4436 14368
rect 4488 14356 4494 14408
rect 1946 14260 1952 14272
rect 1907 14232 1952 14260
rect 1946 14220 1952 14232
rect 2004 14220 2010 14272
rect 8202 14220 8208 14272
rect 8260 14260 8266 14272
rect 8297 14263 8355 14269
rect 8297 14260 8309 14263
rect 8260 14232 8309 14260
rect 8260 14220 8266 14232
rect 8297 14229 8309 14232
rect 8343 14229 8355 14263
rect 11698 14260 11704 14272
rect 11659 14232 11704 14260
rect 8297 14223 8355 14229
rect 11698 14220 11704 14232
rect 11756 14220 11762 14272
rect 1104 14170 21896 14192
rect 1104 14118 4447 14170
rect 4499 14118 4511 14170
rect 4563 14118 4575 14170
rect 4627 14118 4639 14170
rect 4691 14118 11378 14170
rect 11430 14118 11442 14170
rect 11494 14118 11506 14170
rect 11558 14118 11570 14170
rect 11622 14118 18308 14170
rect 18360 14118 18372 14170
rect 18424 14118 18436 14170
rect 18488 14118 18500 14170
rect 18552 14118 21896 14170
rect 1104 14096 21896 14118
rect 2958 14016 2964 14068
rect 3016 14056 3022 14068
rect 3237 14059 3295 14065
rect 3237 14056 3249 14059
rect 3016 14028 3249 14056
rect 3016 14016 3022 14028
rect 3237 14025 3249 14028
rect 3283 14025 3295 14059
rect 3237 14019 3295 14025
rect 5258 14016 5264 14068
rect 5316 14056 5322 14068
rect 5353 14059 5411 14065
rect 5353 14056 5365 14059
rect 5316 14028 5365 14056
rect 5316 14016 5322 14028
rect 5353 14025 5365 14028
rect 5399 14025 5411 14059
rect 5626 14056 5632 14068
rect 5587 14028 5632 14056
rect 5353 14019 5411 14025
rect 1857 13923 1915 13929
rect 1857 13889 1869 13923
rect 1903 13920 1915 13923
rect 2774 13920 2780 13932
rect 1903 13892 2780 13920
rect 1903 13889 1915 13892
rect 1857 13883 1915 13889
rect 2774 13880 2780 13892
rect 2832 13880 2838 13932
rect 5368 13920 5396 14019
rect 5626 14016 5632 14028
rect 5684 14016 5690 14068
rect 7006 14016 7012 14068
rect 7064 14056 7070 14068
rect 9033 14059 9091 14065
rect 9033 14056 9045 14059
rect 7064 14028 9045 14056
rect 7064 14016 7070 14028
rect 9033 14025 9045 14028
rect 9079 14025 9091 14059
rect 9033 14019 9091 14025
rect 10870 14016 10876 14068
rect 10928 14056 10934 14068
rect 10965 14059 11023 14065
rect 10965 14056 10977 14059
rect 10928 14028 10977 14056
rect 10928 14016 10934 14028
rect 10965 14025 10977 14028
rect 11011 14025 11023 14059
rect 11238 14056 11244 14068
rect 11199 14028 11244 14056
rect 10965 14019 11023 14025
rect 7745 13991 7803 13997
rect 7745 13957 7757 13991
rect 7791 13988 7803 13991
rect 8938 13988 8944 14000
rect 7791 13960 8944 13988
rect 7791 13957 7803 13960
rect 7745 13951 7803 13957
rect 8938 13948 8944 13960
rect 8996 13948 9002 14000
rect 6181 13923 6239 13929
rect 6181 13920 6193 13923
rect 5368 13892 6193 13920
rect 6181 13889 6193 13892
rect 6227 13889 6239 13923
rect 6181 13883 6239 13889
rect 8202 13880 8208 13932
rect 8260 13920 8266 13932
rect 8297 13923 8355 13929
rect 8297 13920 8309 13923
rect 8260 13892 8309 13920
rect 8260 13880 8266 13892
rect 8297 13889 8309 13892
rect 8343 13889 8355 13923
rect 9217 13923 9275 13929
rect 9217 13920 9229 13923
rect 8297 13883 8355 13889
rect 8680 13892 9229 13920
rect 1578 13852 1584 13864
rect 1539 13824 1584 13852
rect 1578 13812 1584 13824
rect 1636 13812 1642 13864
rect 2327 13855 2385 13861
rect 2327 13821 2339 13855
rect 2373 13821 2385 13855
rect 3050 13852 3056 13864
rect 3011 13824 3056 13852
rect 2327 13815 2385 13821
rect 2332 13716 2360 13815
rect 3050 13812 3056 13824
rect 3108 13812 3114 13864
rect 3142 13812 3148 13864
rect 3200 13812 3206 13864
rect 3973 13855 4031 13861
rect 3973 13821 3985 13855
rect 4019 13852 4031 13855
rect 4062 13852 4068 13864
rect 4019 13824 4068 13852
rect 4019 13821 4031 13824
rect 3973 13815 4031 13821
rect 4062 13812 4068 13824
rect 4120 13812 4126 13864
rect 6822 13852 6828 13864
rect 5175 13824 6828 13852
rect 2590 13784 2596 13796
rect 2551 13756 2596 13784
rect 2590 13744 2596 13756
rect 2648 13744 2654 13796
rect 3160 13784 3188 13812
rect 2700 13756 3188 13784
rect 4240 13787 4298 13793
rect 2700 13716 2728 13756
rect 4240 13753 4252 13787
rect 4286 13784 4298 13787
rect 5074 13784 5080 13796
rect 4286 13756 5080 13784
rect 4286 13753 4298 13756
rect 4240 13747 4298 13753
rect 5074 13744 5080 13756
rect 5132 13744 5138 13796
rect 2332 13688 2728 13716
rect 2866 13676 2872 13728
rect 2924 13716 2930 13728
rect 5175 13716 5203 13824
rect 6822 13812 6828 13824
rect 6880 13852 6886 13864
rect 7377 13855 7435 13861
rect 7377 13852 7389 13855
rect 6880 13824 7389 13852
rect 6880 13812 6886 13824
rect 7377 13821 7389 13824
rect 7423 13852 7435 13855
rect 8113 13855 8171 13861
rect 8113 13852 8125 13855
rect 7423 13824 8125 13852
rect 7423 13821 7435 13824
rect 7377 13815 7435 13821
rect 8113 13821 8125 13824
rect 8159 13821 8171 13855
rect 8570 13852 8576 13864
rect 8113 13815 8171 13821
rect 8220 13824 8576 13852
rect 5534 13744 5540 13796
rect 5592 13784 5598 13796
rect 8220 13793 8248 13824
rect 8570 13812 8576 13824
rect 8628 13852 8634 13864
rect 8680 13852 8708 13892
rect 9217 13889 9229 13892
rect 9263 13889 9275 13923
rect 9582 13920 9588 13932
rect 9543 13892 9588 13920
rect 9217 13883 9275 13889
rect 9582 13880 9588 13892
rect 9640 13880 9646 13932
rect 10980 13920 11008 14019
rect 11238 14016 11244 14028
rect 11296 14016 11302 14068
rect 11793 13923 11851 13929
rect 11793 13920 11805 13923
rect 10980 13892 11805 13920
rect 11793 13889 11805 13892
rect 11839 13889 11851 13923
rect 11793 13883 11851 13889
rect 8628 13824 8708 13852
rect 8628 13812 8634 13824
rect 8754 13812 8760 13864
rect 8812 13812 8818 13864
rect 8941 13855 8999 13861
rect 8941 13821 8953 13855
rect 8987 13852 8999 13855
rect 9033 13855 9091 13861
rect 9033 13852 9045 13855
rect 8987 13824 9045 13852
rect 8987 13821 8999 13824
rect 8941 13815 8999 13821
rect 9033 13821 9045 13824
rect 9079 13821 9091 13855
rect 9033 13815 9091 13821
rect 9122 13812 9128 13864
rect 9180 13852 9186 13864
rect 9398 13852 9404 13864
rect 9180 13824 9404 13852
rect 9180 13812 9186 13824
rect 9398 13812 9404 13824
rect 9456 13852 9462 13864
rect 11609 13855 11667 13861
rect 11609 13852 11621 13855
rect 9456 13824 11621 13852
rect 9456 13812 9462 13824
rect 11609 13821 11621 13824
rect 11655 13852 11667 13855
rect 11698 13852 11704 13864
rect 11655 13824 11704 13852
rect 11655 13821 11667 13824
rect 11609 13815 11667 13821
rect 11698 13812 11704 13824
rect 11756 13812 11762 13864
rect 6089 13787 6147 13793
rect 6089 13784 6101 13787
rect 5592 13756 6101 13784
rect 5592 13744 5598 13756
rect 6089 13753 6101 13756
rect 6135 13753 6147 13787
rect 6089 13747 6147 13753
rect 8205 13787 8263 13793
rect 8205 13753 8217 13787
rect 8251 13753 8263 13787
rect 8205 13747 8263 13753
rect 5994 13716 6000 13728
rect 2924 13688 5203 13716
rect 5955 13688 6000 13716
rect 2924 13676 2930 13688
rect 5994 13676 6000 13688
rect 6052 13676 6058 13728
rect 8772 13725 8800 13812
rect 9852 13787 9910 13793
rect 9852 13753 9864 13787
rect 9898 13784 9910 13787
rect 10870 13784 10876 13796
rect 9898 13756 10876 13784
rect 9898 13753 9910 13756
rect 9852 13747 9910 13753
rect 10870 13744 10876 13756
rect 10928 13744 10934 13796
rect 8757 13719 8815 13725
rect 8757 13685 8769 13719
rect 8803 13685 8815 13719
rect 8757 13679 8815 13685
rect 11701 13719 11759 13725
rect 11701 13685 11713 13719
rect 11747 13716 11759 13719
rect 11882 13716 11888 13728
rect 11747 13688 11888 13716
rect 11747 13685 11759 13688
rect 11701 13679 11759 13685
rect 11882 13676 11888 13688
rect 11940 13676 11946 13728
rect 1104 13626 21896 13648
rect 1104 13574 7912 13626
rect 7964 13574 7976 13626
rect 8028 13574 8040 13626
rect 8092 13574 8104 13626
rect 8156 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 15035 13626
rect 15087 13574 21896 13626
rect 1104 13552 21896 13574
rect 3510 13512 3516 13524
rect 3471 13484 3516 13512
rect 3510 13472 3516 13484
rect 3568 13472 3574 13524
rect 4525 13515 4583 13521
rect 4525 13481 4537 13515
rect 4571 13512 4583 13515
rect 5994 13512 6000 13524
rect 4571 13484 6000 13512
rect 4571 13481 4583 13484
rect 4525 13475 4583 13481
rect 5994 13472 6000 13484
rect 6052 13472 6058 13524
rect 10870 13472 10876 13524
rect 10928 13512 10934 13524
rect 11333 13515 11391 13521
rect 11333 13512 11345 13515
rect 10928 13484 11345 13512
rect 10928 13472 10934 13484
rect 11333 13481 11345 13484
rect 11379 13481 11391 13515
rect 11333 13475 11391 13481
rect 1762 13404 1768 13456
rect 1820 13444 1826 13456
rect 2133 13447 2191 13453
rect 2133 13444 2145 13447
rect 1820 13416 2145 13444
rect 1820 13404 1826 13416
rect 2133 13413 2145 13416
rect 2179 13413 2191 13447
rect 2133 13407 2191 13413
rect 2869 13447 2927 13453
rect 2869 13413 2881 13447
rect 2915 13444 2927 13447
rect 3050 13444 3056 13456
rect 2915 13416 3056 13444
rect 2915 13413 2927 13416
rect 2869 13407 2927 13413
rect 3050 13404 3056 13416
rect 3108 13404 3114 13456
rect 5074 13404 5080 13456
rect 5132 13444 5138 13456
rect 7276 13447 7334 13453
rect 5132 13416 5672 13444
rect 5132 13404 5138 13416
rect 1857 13379 1915 13385
rect 1857 13345 1869 13379
rect 1903 13376 1915 13379
rect 1946 13376 1952 13388
rect 1903 13348 1952 13376
rect 1903 13345 1915 13348
rect 1857 13339 1915 13345
rect 1946 13336 1952 13348
rect 2004 13336 2010 13388
rect 2593 13379 2651 13385
rect 2593 13345 2605 13379
rect 2639 13376 2651 13379
rect 3234 13376 3240 13388
rect 2639 13348 3240 13376
rect 2639 13345 2651 13348
rect 2593 13339 2651 13345
rect 3234 13336 3240 13348
rect 3292 13336 3298 13388
rect 3329 13379 3387 13385
rect 3329 13345 3341 13379
rect 3375 13376 3387 13379
rect 3418 13376 3424 13388
rect 3375 13348 3424 13376
rect 3375 13345 3387 13348
rect 3329 13339 3387 13345
rect 3418 13336 3424 13348
rect 3476 13336 3482 13388
rect 4249 13379 4307 13385
rect 4249 13345 4261 13379
rect 4295 13376 4307 13379
rect 5258 13376 5264 13388
rect 4295 13348 5264 13376
rect 4295 13345 4307 13348
rect 4249 13339 4307 13345
rect 5258 13336 5264 13348
rect 5316 13376 5322 13388
rect 5445 13379 5503 13385
rect 5445 13376 5457 13379
rect 5316 13348 5457 13376
rect 5316 13336 5322 13348
rect 5445 13345 5457 13348
rect 5491 13345 5503 13379
rect 5445 13339 5503 13345
rect 5644 13317 5672 13416
rect 7276 13413 7288 13447
rect 7322 13444 7334 13447
rect 8202 13444 8208 13456
rect 7322 13416 8208 13444
rect 7322 13413 7334 13416
rect 7276 13407 7334 13413
rect 8202 13404 8208 13416
rect 8260 13404 8266 13456
rect 10042 13444 10048 13456
rect 9955 13416 10048 13444
rect 6914 13336 6920 13388
rect 6972 13376 6978 13388
rect 7009 13379 7067 13385
rect 7009 13376 7021 13379
rect 6972 13348 7021 13376
rect 6972 13336 6978 13348
rect 7009 13345 7021 13348
rect 7055 13376 7067 13379
rect 8110 13376 8116 13388
rect 7055 13348 8116 13376
rect 7055 13345 7067 13348
rect 7009 13339 7067 13345
rect 8110 13336 8116 13348
rect 8168 13336 8174 13388
rect 9968 13385 9996 13416
rect 10042 13404 10048 13416
rect 10100 13444 10106 13456
rect 10686 13444 10692 13456
rect 10100 13416 10692 13444
rect 10100 13404 10106 13416
rect 10686 13404 10692 13416
rect 10744 13404 10750 13456
rect 9953 13379 10011 13385
rect 9953 13345 9965 13379
rect 9999 13345 10011 13379
rect 9953 13339 10011 13345
rect 10220 13379 10278 13385
rect 10220 13345 10232 13379
rect 10266 13376 10278 13379
rect 11054 13376 11060 13388
rect 10266 13348 11060 13376
rect 10266 13345 10278 13348
rect 10220 13339 10278 13345
rect 11054 13336 11060 13348
rect 11112 13336 11118 13388
rect 5537 13311 5595 13317
rect 5537 13277 5549 13311
rect 5583 13277 5595 13311
rect 5537 13271 5595 13277
rect 5629 13311 5687 13317
rect 5629 13277 5641 13311
rect 5675 13277 5687 13311
rect 5629 13271 5687 13277
rect 5077 13243 5135 13249
rect 5077 13209 5089 13243
rect 5123 13240 5135 13243
rect 5442 13240 5448 13252
rect 5123 13212 5448 13240
rect 5123 13209 5135 13212
rect 5077 13203 5135 13209
rect 5442 13200 5448 13212
rect 5500 13200 5506 13252
rect 5552 13172 5580 13271
rect 8018 13268 8024 13320
rect 8076 13308 8082 13320
rect 8665 13311 8723 13317
rect 8665 13308 8677 13311
rect 8076 13280 8677 13308
rect 8076 13268 8082 13280
rect 8665 13277 8677 13280
rect 8711 13277 8723 13311
rect 8665 13271 8723 13277
rect 9125 13311 9183 13317
rect 9125 13277 9137 13311
rect 9171 13277 9183 13311
rect 9125 13271 9183 13277
rect 6086 13172 6092 13184
rect 5552 13144 6092 13172
rect 6086 13132 6092 13144
rect 6144 13132 6150 13184
rect 8386 13172 8392 13184
rect 8347 13144 8392 13172
rect 8386 13132 8392 13144
rect 8444 13132 8450 13184
rect 9140 13172 9168 13271
rect 10962 13172 10968 13184
rect 9140 13144 10968 13172
rect 10962 13132 10968 13144
rect 11020 13132 11026 13184
rect 11701 13175 11759 13181
rect 11701 13141 11713 13175
rect 11747 13172 11759 13175
rect 11882 13172 11888 13184
rect 11747 13144 11888 13172
rect 11747 13141 11759 13144
rect 11701 13135 11759 13141
rect 11882 13132 11888 13144
rect 11940 13132 11946 13184
rect 1104 13082 21896 13104
rect 1104 13030 4447 13082
rect 4499 13030 4511 13082
rect 4563 13030 4575 13082
rect 4627 13030 4639 13082
rect 4691 13030 11378 13082
rect 11430 13030 11442 13082
rect 11494 13030 11506 13082
rect 11558 13030 11570 13082
rect 11622 13030 18308 13082
rect 18360 13030 18372 13082
rect 18424 13030 18436 13082
rect 18488 13030 18500 13082
rect 18552 13030 21896 13082
rect 1104 13008 21896 13030
rect 1578 12928 1584 12980
rect 1636 12968 1642 12980
rect 2225 12971 2283 12977
rect 2225 12968 2237 12971
rect 1636 12940 2237 12968
rect 1636 12928 1642 12940
rect 2225 12937 2237 12940
rect 2271 12937 2283 12971
rect 2225 12931 2283 12937
rect 5074 12928 5080 12980
rect 5132 12968 5138 12980
rect 5537 12971 5595 12977
rect 5537 12968 5549 12971
rect 5132 12940 5549 12968
rect 5132 12928 5138 12940
rect 5537 12937 5549 12940
rect 5583 12937 5595 12971
rect 7006 12968 7012 12980
rect 6967 12940 7012 12968
rect 5537 12931 5595 12937
rect 7006 12928 7012 12940
rect 7064 12928 7070 12980
rect 7469 12971 7527 12977
rect 7469 12937 7481 12971
rect 7515 12968 7527 12971
rect 8297 12971 8355 12977
rect 8297 12968 8309 12971
rect 7515 12940 8309 12968
rect 7515 12937 7527 12940
rect 7469 12931 7527 12937
rect 8297 12937 8309 12940
rect 8343 12937 8355 12971
rect 8478 12968 8484 12980
rect 8439 12940 8484 12968
rect 8297 12931 8355 12937
rect 8478 12928 8484 12940
rect 8536 12928 8542 12980
rect 10594 12968 10600 12980
rect 10555 12940 10600 12968
rect 10594 12928 10600 12940
rect 10652 12928 10658 12980
rect 5258 12860 5264 12912
rect 5316 12900 5322 12912
rect 5442 12900 5448 12912
rect 5316 12872 5448 12900
rect 5316 12860 5322 12872
rect 5442 12860 5448 12872
rect 5500 12900 5506 12912
rect 8846 12900 8852 12912
rect 5500 12872 8852 12900
rect 5500 12860 5506 12872
rect 8846 12860 8852 12872
rect 8904 12860 8910 12912
rect 10870 12860 10876 12912
rect 10928 12900 10934 12912
rect 10928 12872 11192 12900
rect 10928 12860 10934 12872
rect 2866 12832 2872 12844
rect 2827 12804 2872 12832
rect 2866 12792 2872 12804
rect 2924 12792 2930 12844
rect 3418 12832 3424 12844
rect 3379 12804 3424 12832
rect 3418 12792 3424 12804
rect 3476 12792 3482 12844
rect 8113 12835 8171 12841
rect 8113 12801 8125 12835
rect 8159 12832 8171 12835
rect 8202 12832 8208 12844
rect 8159 12804 8208 12832
rect 8159 12801 8171 12804
rect 8113 12795 8171 12801
rect 8202 12792 8208 12804
rect 8260 12792 8266 12844
rect 8386 12792 8392 12844
rect 8444 12832 8450 12844
rect 9033 12835 9091 12841
rect 9033 12832 9045 12835
rect 8444 12804 9045 12832
rect 8444 12792 8450 12804
rect 9033 12801 9045 12804
rect 9079 12801 9091 12835
rect 9033 12795 9091 12801
rect 10229 12835 10287 12841
rect 10229 12801 10241 12835
rect 10275 12832 10287 12835
rect 11054 12832 11060 12844
rect 10275 12804 11060 12832
rect 10275 12801 10287 12804
rect 10229 12795 10287 12801
rect 11054 12792 11060 12804
rect 11112 12792 11118 12844
rect 11164 12841 11192 12872
rect 11149 12835 11207 12841
rect 11149 12801 11161 12835
rect 11195 12801 11207 12835
rect 11149 12795 11207 12801
rect 3237 12767 3295 12773
rect 3237 12733 3249 12767
rect 3283 12764 3295 12767
rect 4062 12764 4068 12776
rect 3283 12736 4068 12764
rect 3283 12733 3295 12736
rect 3237 12727 3295 12733
rect 4062 12724 4068 12736
rect 4120 12724 4126 12776
rect 4154 12724 4160 12776
rect 4212 12764 4218 12776
rect 5997 12767 6055 12773
rect 4212 12736 4257 12764
rect 4212 12724 4218 12736
rect 5997 12733 6009 12767
rect 6043 12764 6055 12767
rect 7006 12764 7012 12776
rect 6043 12736 7012 12764
rect 6043 12733 6055 12736
rect 5997 12727 6055 12733
rect 7006 12724 7012 12736
rect 7064 12724 7070 12776
rect 7193 12767 7251 12773
rect 7193 12733 7205 12767
rect 7239 12764 7251 12767
rect 7742 12764 7748 12776
rect 7239 12736 7748 12764
rect 7239 12733 7251 12736
rect 7193 12727 7251 12733
rect 7742 12724 7748 12736
rect 7800 12724 7806 12776
rect 8938 12764 8944 12776
rect 8899 12736 8944 12764
rect 8938 12724 8944 12736
rect 8996 12724 9002 12776
rect 9582 12724 9588 12776
rect 9640 12764 9646 12776
rect 9953 12767 10011 12773
rect 9953 12764 9965 12767
rect 9640 12736 9965 12764
rect 9640 12724 9646 12736
rect 9953 12733 9965 12736
rect 9999 12733 10011 12767
rect 9953 12727 10011 12733
rect 10045 12767 10103 12773
rect 10045 12733 10057 12767
rect 10091 12764 10103 12767
rect 10870 12764 10876 12776
rect 10091 12736 10876 12764
rect 10091 12733 10103 12736
rect 10045 12727 10103 12733
rect 10870 12724 10876 12736
rect 10928 12764 10934 12776
rect 11609 12767 11667 12773
rect 11609 12764 11621 12767
rect 10928 12736 11621 12764
rect 10928 12724 10934 12736
rect 11609 12733 11621 12736
rect 11655 12733 11667 12767
rect 11609 12727 11667 12733
rect 4424 12699 4482 12705
rect 4424 12665 4436 12699
rect 4470 12696 4482 12699
rect 4706 12696 4712 12708
rect 4470 12668 4712 12696
rect 4470 12665 4482 12668
rect 4424 12659 4482 12665
rect 4706 12656 4712 12668
rect 4764 12656 4770 12708
rect 7837 12699 7895 12705
rect 7837 12665 7849 12699
rect 7883 12696 7895 12699
rect 8018 12696 8024 12708
rect 7883 12668 8024 12696
rect 7883 12665 7895 12668
rect 7837 12659 7895 12665
rect 8018 12656 8024 12668
rect 8076 12656 8082 12708
rect 8297 12699 8355 12705
rect 8297 12665 8309 12699
rect 8343 12696 8355 12699
rect 8849 12699 8907 12705
rect 8849 12696 8861 12699
rect 8343 12668 8861 12696
rect 8343 12665 8355 12668
rect 8297 12659 8355 12665
rect 8849 12665 8861 12668
rect 8895 12665 8907 12699
rect 11057 12699 11115 12705
rect 11057 12696 11069 12699
rect 8849 12659 8907 12665
rect 9600 12668 11069 12696
rect 2590 12628 2596 12640
rect 2551 12600 2596 12628
rect 2590 12588 2596 12600
rect 2648 12588 2654 12640
rect 2685 12631 2743 12637
rect 2685 12597 2697 12631
rect 2731 12628 2743 12631
rect 2774 12628 2780 12640
rect 2731 12600 2780 12628
rect 2731 12597 2743 12600
rect 2685 12591 2743 12597
rect 2774 12588 2780 12600
rect 2832 12588 2838 12640
rect 5074 12588 5080 12640
rect 5132 12628 5138 12640
rect 5813 12631 5871 12637
rect 5813 12628 5825 12631
rect 5132 12600 5825 12628
rect 5132 12588 5138 12600
rect 5813 12597 5825 12600
rect 5859 12628 5871 12631
rect 6362 12628 6368 12640
rect 5859 12600 6368 12628
rect 5859 12597 5871 12600
rect 5813 12591 5871 12597
rect 6362 12588 6368 12600
rect 6420 12588 6426 12640
rect 6457 12631 6515 12637
rect 6457 12597 6469 12631
rect 6503 12628 6515 12631
rect 7929 12631 7987 12637
rect 7929 12628 7941 12631
rect 6503 12600 7941 12628
rect 6503 12597 6515 12600
rect 6457 12591 6515 12597
rect 7929 12597 7941 12600
rect 7975 12628 7987 12631
rect 8754 12628 8760 12640
rect 7975 12600 8760 12628
rect 7975 12597 7987 12600
rect 7929 12591 7987 12597
rect 8754 12588 8760 12600
rect 8812 12588 8818 12640
rect 9600 12637 9628 12668
rect 11057 12665 11069 12668
rect 11103 12665 11115 12699
rect 11057 12659 11115 12665
rect 9585 12631 9643 12637
rect 9585 12597 9597 12631
rect 9631 12597 9643 12631
rect 10962 12628 10968 12640
rect 10923 12600 10968 12628
rect 9585 12591 9643 12597
rect 10962 12588 10968 12600
rect 11020 12588 11026 12640
rect 1104 12538 21896 12560
rect 1104 12486 7912 12538
rect 7964 12486 7976 12538
rect 8028 12486 8040 12538
rect 8092 12486 8104 12538
rect 8156 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 15035 12538
rect 15087 12486 21896 12538
rect 1104 12464 21896 12486
rect 1486 12384 1492 12436
rect 1544 12424 1550 12436
rect 1581 12427 1639 12433
rect 1581 12424 1593 12427
rect 1544 12396 1593 12424
rect 1544 12384 1550 12396
rect 1581 12393 1593 12396
rect 1627 12393 1639 12427
rect 1581 12387 1639 12393
rect 3142 12384 3148 12436
rect 3200 12424 3206 12436
rect 4065 12427 4123 12433
rect 4065 12424 4077 12427
rect 3200 12396 4077 12424
rect 3200 12384 3206 12396
rect 4065 12393 4077 12396
rect 4111 12393 4123 12427
rect 8846 12424 8852 12436
rect 4065 12387 4123 12393
rect 4172 12396 8524 12424
rect 8807 12396 8852 12424
rect 2866 12316 2872 12368
rect 2924 12356 2930 12368
rect 3326 12356 3332 12368
rect 2924 12328 3332 12356
rect 2924 12316 2930 12328
rect 3326 12316 3332 12328
rect 3384 12316 3390 12368
rect 3970 12316 3976 12368
rect 4028 12356 4034 12368
rect 4172 12356 4200 12396
rect 4028 12328 4200 12356
rect 4525 12359 4583 12365
rect 4028 12316 4034 12328
rect 4525 12325 4537 12359
rect 4571 12356 4583 12359
rect 5626 12356 5632 12368
rect 4571 12328 5632 12356
rect 4571 12325 4583 12328
rect 4525 12319 4583 12325
rect 5626 12316 5632 12328
rect 5684 12316 5690 12368
rect 7092 12359 7150 12365
rect 7092 12325 7104 12359
rect 7138 12356 7150 12359
rect 8386 12356 8392 12368
rect 7138 12328 8392 12356
rect 7138 12325 7150 12328
rect 7092 12319 7150 12325
rect 8386 12316 8392 12328
rect 8444 12316 8450 12368
rect 8496 12356 8524 12396
rect 8846 12384 8852 12396
rect 8904 12424 8910 12436
rect 9582 12424 9588 12436
rect 8904 12396 9588 12424
rect 8904 12384 8910 12396
rect 9582 12384 9588 12396
rect 9640 12384 9646 12436
rect 11054 12384 11060 12436
rect 11112 12424 11118 12436
rect 11241 12427 11299 12433
rect 11241 12424 11253 12427
rect 11112 12396 11253 12424
rect 11112 12384 11118 12396
rect 11241 12393 11253 12396
rect 11287 12393 11299 12427
rect 11241 12387 11299 12393
rect 12158 12384 12164 12436
rect 12216 12424 12222 12436
rect 12434 12424 12440 12436
rect 12216 12396 12440 12424
rect 12216 12384 12222 12396
rect 12434 12384 12440 12396
rect 12492 12384 12498 12436
rect 19702 12384 19708 12436
rect 19760 12424 19766 12436
rect 20257 12427 20315 12433
rect 20257 12424 20269 12427
rect 19760 12396 20269 12424
rect 19760 12384 19766 12396
rect 20257 12393 20269 12396
rect 20303 12393 20315 12427
rect 20257 12387 20315 12393
rect 11698 12356 11704 12368
rect 8496 12328 11704 12356
rect 11698 12316 11704 12328
rect 11756 12316 11762 12368
rect 12360 12328 12480 12356
rect 1397 12291 1455 12297
rect 1397 12257 1409 12291
rect 1443 12257 1455 12291
rect 1397 12251 1455 12257
rect 1949 12291 2007 12297
rect 1949 12257 1961 12291
rect 1995 12288 2007 12291
rect 2038 12288 2044 12300
rect 1995 12260 2044 12288
rect 1995 12257 2007 12260
rect 1949 12251 2007 12257
rect 1412 12084 1440 12251
rect 2038 12248 2044 12260
rect 2096 12248 2102 12300
rect 2216 12291 2274 12297
rect 2216 12257 2228 12291
rect 2262 12288 2274 12291
rect 2958 12288 2964 12300
rect 2262 12260 2964 12288
rect 2262 12257 2274 12260
rect 2216 12251 2274 12257
rect 2958 12248 2964 12260
rect 3016 12248 3022 12300
rect 4433 12291 4491 12297
rect 4433 12257 4445 12291
rect 4479 12288 4491 12291
rect 4798 12288 4804 12300
rect 4479 12260 4804 12288
rect 4479 12257 4491 12260
rect 4433 12251 4491 12257
rect 4798 12248 4804 12260
rect 4856 12248 4862 12300
rect 4893 12291 4951 12297
rect 4893 12257 4905 12291
rect 4939 12288 4951 12291
rect 5074 12288 5080 12300
rect 4939 12260 5080 12288
rect 4939 12257 4951 12260
rect 4893 12251 4951 12257
rect 5074 12248 5080 12260
rect 5132 12248 5138 12300
rect 5344 12291 5402 12297
rect 5344 12257 5356 12291
rect 5390 12288 5402 12291
rect 5902 12288 5908 12300
rect 5390 12260 5908 12288
rect 5390 12257 5402 12260
rect 5344 12251 5402 12257
rect 5902 12248 5908 12260
rect 5960 12248 5966 12300
rect 9861 12291 9919 12297
rect 9861 12257 9873 12291
rect 9907 12288 9919 12291
rect 9950 12288 9956 12300
rect 9907 12260 9956 12288
rect 9907 12257 9919 12260
rect 9861 12251 9919 12257
rect 9950 12248 9956 12260
rect 10008 12248 10014 12300
rect 10128 12291 10186 12297
rect 10128 12257 10140 12291
rect 10174 12288 10186 12291
rect 11054 12288 11060 12300
rect 10174 12260 11060 12288
rect 10174 12257 10186 12260
rect 10128 12251 10186 12257
rect 11054 12248 11060 12260
rect 11112 12248 11118 12300
rect 4706 12220 4712 12232
rect 4619 12192 4712 12220
rect 4706 12180 4712 12192
rect 4764 12220 4770 12232
rect 4764 12192 5028 12220
rect 4764 12180 4770 12192
rect 4246 12152 4252 12164
rect 2884 12124 4252 12152
rect 2884 12084 2912 12124
rect 4246 12112 4252 12124
rect 4304 12112 4310 12164
rect 3326 12084 3332 12096
rect 1412 12056 2912 12084
rect 3287 12056 3332 12084
rect 3326 12044 3332 12056
rect 3384 12044 3390 12096
rect 4154 12044 4160 12096
rect 4212 12084 4218 12096
rect 4893 12087 4951 12093
rect 4893 12084 4905 12087
rect 4212 12056 4905 12084
rect 4212 12044 4218 12056
rect 4893 12053 4905 12056
rect 4939 12053 4951 12087
rect 5000 12084 5028 12192
rect 6362 12180 6368 12232
rect 6420 12220 6426 12232
rect 6822 12220 6828 12232
rect 6420 12192 6828 12220
rect 6420 12180 6426 12192
rect 6822 12180 6828 12192
rect 6880 12180 6886 12232
rect 9692 12192 9895 12220
rect 8294 12112 8300 12164
rect 8352 12152 8358 12164
rect 8352 12124 9619 12152
rect 8352 12112 8358 12124
rect 6457 12087 6515 12093
rect 6457 12084 6469 12087
rect 5000 12056 6469 12084
rect 4893 12047 4951 12053
rect 6457 12053 6469 12056
rect 6503 12053 6515 12087
rect 6457 12047 6515 12053
rect 8110 12044 8116 12096
rect 8168 12084 8174 12096
rect 8205 12087 8263 12093
rect 8205 12084 8217 12087
rect 8168 12056 8217 12084
rect 8168 12044 8174 12056
rect 8205 12053 8217 12056
rect 8251 12053 8263 12087
rect 9214 12084 9220 12096
rect 9175 12056 9220 12084
rect 8205 12047 8263 12053
rect 9214 12044 9220 12056
rect 9272 12044 9278 12096
rect 9591 12084 9619 12124
rect 9692 12084 9720 12192
rect 9591 12056 9720 12084
rect 9867 12084 9895 12192
rect 12360 12084 12388 12328
rect 12452 12288 12480 12328
rect 19702 12288 19708 12300
rect 12452 12260 19708 12288
rect 19702 12248 19708 12260
rect 19760 12248 19766 12300
rect 9867 12056 12388 12084
rect 19889 12087 19947 12093
rect 19889 12053 19901 12087
rect 19935 12084 19947 12087
rect 20530 12084 20536 12096
rect 19935 12056 20536 12084
rect 19935 12053 19947 12056
rect 19889 12047 19947 12053
rect 20530 12044 20536 12056
rect 20588 12044 20594 12096
rect 1104 11994 21896 12016
rect 1104 11942 4447 11994
rect 4499 11942 4511 11994
rect 4563 11942 4575 11994
rect 4627 11942 4639 11994
rect 4691 11942 11378 11994
rect 11430 11942 11442 11994
rect 11494 11942 11506 11994
rect 11558 11942 11570 11994
rect 11622 11942 18308 11994
rect 18360 11942 18372 11994
rect 18424 11942 18436 11994
rect 18488 11942 18500 11994
rect 18552 11942 21896 11994
rect 1104 11920 21896 11942
rect 2041 11883 2099 11889
rect 2041 11849 2053 11883
rect 2087 11880 2099 11883
rect 2590 11880 2596 11892
rect 2087 11852 2596 11880
rect 2087 11849 2099 11852
rect 2041 11843 2099 11849
rect 2590 11840 2596 11852
rect 2648 11840 2654 11892
rect 2682 11840 2688 11892
rect 2740 11880 2746 11892
rect 7009 11883 7067 11889
rect 2740 11852 6868 11880
rect 2740 11840 2746 11852
rect 6840 11812 6868 11852
rect 7009 11849 7021 11883
rect 7055 11880 7067 11883
rect 7558 11880 7564 11892
rect 7055 11852 7564 11880
rect 7055 11849 7067 11852
rect 7009 11843 7067 11849
rect 7558 11840 7564 11852
rect 7616 11840 7622 11892
rect 10965 11883 11023 11889
rect 10965 11880 10977 11883
rect 7668 11852 10977 11880
rect 7668 11812 7696 11852
rect 10965 11849 10977 11852
rect 11011 11849 11023 11883
rect 10965 11843 11023 11849
rect 6840 11784 7696 11812
rect 9585 11815 9643 11821
rect 9585 11781 9597 11815
rect 9631 11781 9643 11815
rect 9585 11775 9643 11781
rect 9953 11815 10011 11821
rect 9953 11781 9965 11815
rect 9999 11812 10011 11815
rect 9999 11784 11468 11812
rect 9999 11781 10011 11784
rect 9953 11775 10011 11781
rect 2685 11747 2743 11753
rect 2685 11713 2697 11747
rect 2731 11744 2743 11747
rect 2958 11744 2964 11756
rect 2731 11716 2964 11744
rect 2731 11713 2743 11716
rect 2685 11707 2743 11713
rect 2958 11704 2964 11716
rect 3016 11704 3022 11756
rect 4709 11747 4767 11753
rect 4709 11713 4721 11747
rect 4755 11744 4767 11747
rect 4798 11744 4804 11756
rect 4755 11716 4804 11744
rect 4755 11713 4767 11716
rect 4709 11707 4767 11713
rect 4798 11704 4804 11716
rect 4856 11704 4862 11756
rect 7653 11747 7711 11753
rect 7653 11713 7665 11747
rect 7699 11713 7711 11747
rect 8202 11744 8208 11756
rect 8163 11716 8208 11744
rect 7653 11707 7711 11713
rect 2038 11636 2044 11688
rect 2096 11676 2102 11688
rect 2406 11676 2412 11688
rect 2096 11648 2412 11676
rect 2096 11636 2102 11648
rect 2406 11636 2412 11648
rect 2464 11676 2470 11688
rect 3326 11685 3332 11688
rect 3053 11679 3111 11685
rect 3053 11676 3065 11679
rect 2464 11648 3065 11676
rect 2464 11636 2470 11648
rect 3053 11645 3065 11648
rect 3099 11645 3111 11679
rect 3320 11676 3332 11685
rect 3287 11648 3332 11676
rect 3053 11639 3111 11645
rect 3320 11639 3332 11648
rect 3326 11636 3332 11639
rect 3384 11636 3390 11688
rect 7668 11676 7696 11707
rect 8202 11704 8208 11716
rect 8260 11704 8266 11756
rect 9600 11744 9628 11775
rect 9858 11744 9864 11756
rect 9600 11716 9864 11744
rect 9858 11704 9864 11716
rect 9916 11744 9922 11756
rect 11440 11753 11468 11784
rect 10505 11747 10563 11753
rect 10505 11744 10517 11747
rect 9916 11716 10517 11744
rect 9916 11704 9922 11716
rect 10505 11713 10517 11716
rect 10551 11713 10563 11747
rect 10505 11707 10563 11713
rect 11425 11747 11483 11753
rect 11425 11713 11437 11747
rect 11471 11713 11483 11747
rect 11425 11707 11483 11713
rect 11517 11747 11575 11753
rect 11517 11713 11529 11747
rect 11563 11713 11575 11747
rect 11517 11707 11575 11713
rect 8478 11685 8484 11688
rect 8461 11679 8484 11685
rect 8461 11676 8473 11679
rect 7668 11648 8473 11676
rect 8461 11645 8473 11648
rect 8536 11676 8542 11688
rect 8536 11648 8609 11676
rect 8461 11639 8484 11645
rect 8478 11636 8484 11639
rect 8536 11636 8542 11648
rect 9398 11636 9404 11688
rect 9456 11676 9462 11688
rect 10413 11679 10471 11685
rect 10413 11676 10425 11679
rect 9456 11648 10425 11676
rect 9456 11636 9462 11648
rect 10413 11645 10425 11648
rect 10459 11645 10471 11679
rect 10413 11639 10471 11645
rect 11054 11636 11060 11688
rect 11112 11676 11118 11688
rect 11532 11676 11560 11707
rect 11112 11648 11560 11676
rect 11112 11636 11118 11648
rect 11698 11636 11704 11688
rect 11756 11676 11762 11688
rect 19245 11679 19303 11685
rect 19245 11676 19257 11679
rect 11756 11648 19257 11676
rect 11756 11636 11762 11648
rect 19245 11645 19257 11648
rect 19291 11676 19303 11679
rect 19797 11679 19855 11685
rect 19797 11676 19809 11679
rect 19291 11648 19809 11676
rect 19291 11645 19303 11648
rect 19245 11639 19303 11645
rect 19797 11645 19809 11648
rect 19843 11645 19855 11679
rect 19797 11639 19855 11645
rect 1765 11611 1823 11617
rect 1765 11577 1777 11611
rect 1811 11608 1823 11611
rect 1811 11580 2544 11608
rect 1811 11577 1823 11580
rect 1765 11571 1823 11577
rect 2314 11500 2320 11552
rect 2372 11540 2378 11552
rect 2516 11549 2544 11580
rect 3970 11568 3976 11620
rect 4028 11608 4034 11620
rect 10042 11608 10048 11620
rect 4028 11580 10048 11608
rect 4028 11568 4034 11580
rect 10042 11568 10048 11580
rect 10100 11568 10106 11620
rect 11333 11611 11391 11617
rect 11333 11577 11345 11611
rect 11379 11608 11391 11611
rect 12437 11611 12495 11617
rect 12437 11608 12449 11611
rect 11379 11580 12449 11608
rect 11379 11577 11391 11580
rect 11333 11571 11391 11577
rect 12437 11577 12449 11580
rect 12483 11577 12495 11611
rect 12437 11571 12495 11577
rect 2409 11543 2467 11549
rect 2409 11540 2421 11543
rect 2372 11512 2421 11540
rect 2372 11500 2378 11512
rect 2409 11509 2421 11512
rect 2455 11509 2467 11543
rect 2409 11503 2467 11509
rect 2501 11543 2559 11549
rect 2501 11509 2513 11543
rect 2547 11540 2559 11543
rect 3142 11540 3148 11552
rect 2547 11512 3148 11540
rect 2547 11509 2559 11512
rect 2501 11503 2559 11509
rect 3142 11500 3148 11512
rect 3200 11500 3206 11552
rect 4338 11500 4344 11552
rect 4396 11540 4402 11552
rect 4433 11543 4491 11549
rect 4433 11540 4445 11543
rect 4396 11512 4445 11540
rect 4396 11500 4402 11512
rect 4433 11509 4445 11512
rect 4479 11509 4491 11543
rect 7374 11540 7380 11552
rect 7335 11512 7380 11540
rect 4433 11503 4491 11509
rect 7374 11500 7380 11512
rect 7432 11500 7438 11552
rect 7466 11500 7472 11552
rect 7524 11540 7530 11552
rect 7524 11512 7569 11540
rect 7524 11500 7530 11512
rect 9214 11500 9220 11552
rect 9272 11540 9278 11552
rect 10321 11543 10379 11549
rect 10321 11540 10333 11543
rect 9272 11512 10333 11540
rect 9272 11500 9278 11512
rect 10321 11509 10333 11512
rect 10367 11509 10379 11543
rect 10321 11503 10379 11509
rect 19429 11543 19487 11549
rect 19429 11509 19441 11543
rect 19475 11540 19487 11543
rect 20070 11540 20076 11552
rect 19475 11512 20076 11540
rect 19475 11509 19487 11512
rect 19429 11503 19487 11509
rect 20070 11500 20076 11512
rect 20128 11500 20134 11552
rect 1104 11450 21896 11472
rect 1104 11398 7912 11450
rect 7964 11398 7976 11450
rect 8028 11398 8040 11450
rect 8092 11398 8104 11450
rect 8156 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 15035 11450
rect 15087 11398 21896 11450
rect 1104 11376 21896 11398
rect 2314 11336 2320 11348
rect 2275 11308 2320 11336
rect 2314 11296 2320 11308
rect 2372 11296 2378 11348
rect 2774 11296 2780 11348
rect 2832 11336 2838 11348
rect 2832 11308 2877 11336
rect 2832 11296 2838 11308
rect 3050 11296 3056 11348
rect 3108 11336 3114 11348
rect 3145 11339 3203 11345
rect 3145 11336 3157 11339
rect 3108 11308 3157 11336
rect 3108 11296 3114 11308
rect 3145 11305 3157 11308
rect 3191 11305 3203 11339
rect 3145 11299 3203 11305
rect 5902 11296 5908 11348
rect 5960 11336 5966 11348
rect 5997 11339 6055 11345
rect 5997 11336 6009 11339
rect 5960 11308 6009 11336
rect 5960 11296 5966 11308
rect 5997 11305 6009 11308
rect 6043 11336 6055 11339
rect 6086 11336 6092 11348
rect 6043 11308 6092 11336
rect 6043 11305 6055 11308
rect 5997 11299 6055 11305
rect 6086 11296 6092 11308
rect 6144 11296 6150 11348
rect 7374 11296 7380 11348
rect 7432 11336 7438 11348
rect 8757 11339 8815 11345
rect 8757 11336 8769 11339
rect 7432 11308 8769 11336
rect 7432 11296 7438 11308
rect 8757 11305 8769 11308
rect 8803 11305 8815 11339
rect 10134 11336 10140 11348
rect 8757 11299 8815 11305
rect 9692 11308 10140 11336
rect 2041 11271 2099 11277
rect 2041 11237 2053 11271
rect 2087 11268 2099 11271
rect 3068 11268 3096 11296
rect 2087 11240 3096 11268
rect 2087 11237 2099 11240
rect 2041 11231 2099 11237
rect 4246 11228 4252 11280
rect 4304 11268 4310 11280
rect 6641 11271 6699 11277
rect 6641 11268 6653 11271
rect 4304 11240 6653 11268
rect 4304 11228 4310 11240
rect 6641 11237 6653 11240
rect 6687 11237 6699 11271
rect 6641 11231 6699 11237
rect 9692 11212 9720 11308
rect 10134 11296 10140 11308
rect 10192 11296 10198 11348
rect 11054 11336 11060 11348
rect 11015 11308 11060 11336
rect 11054 11296 11060 11308
rect 11112 11296 11118 11348
rect 9858 11228 9864 11280
rect 9916 11277 9922 11280
rect 9916 11271 9980 11277
rect 9916 11237 9934 11271
rect 9968 11237 9980 11271
rect 9916 11231 9980 11237
rect 9916 11228 9922 11231
rect 10042 11228 10048 11280
rect 10100 11268 10106 11280
rect 10100 11240 18828 11268
rect 10100 11228 10106 11240
rect 2958 11160 2964 11212
rect 3016 11200 3022 11212
rect 4884 11203 4942 11209
rect 3016 11172 3372 11200
rect 3016 11160 3022 11172
rect 3344 11141 3372 11172
rect 4884 11169 4896 11203
rect 4930 11200 4942 11203
rect 5442 11200 5448 11212
rect 4930 11172 5448 11200
rect 4930 11169 4942 11172
rect 4884 11163 4942 11169
rect 5442 11160 5448 11172
rect 5500 11160 5506 11212
rect 6365 11203 6423 11209
rect 6365 11169 6377 11203
rect 6411 11200 6423 11203
rect 7190 11200 7196 11212
rect 6411 11172 7196 11200
rect 6411 11169 6423 11172
rect 6365 11163 6423 11169
rect 7190 11160 7196 11172
rect 7248 11160 7254 11212
rect 7368 11203 7426 11209
rect 7368 11169 7380 11203
rect 7414 11200 7426 11203
rect 8202 11200 8208 11212
rect 7414 11172 8208 11200
rect 7414 11169 7426 11172
rect 7368 11163 7426 11169
rect 8202 11160 8208 11172
rect 8260 11160 8266 11212
rect 9674 11160 9680 11212
rect 9732 11200 9738 11212
rect 9732 11172 10732 11200
rect 9732 11160 9738 11172
rect 3237 11135 3295 11141
rect 3237 11101 3249 11135
rect 3283 11101 3295 11135
rect 3237 11095 3295 11101
rect 3329 11135 3387 11141
rect 3329 11101 3341 11135
rect 3375 11101 3387 11135
rect 3329 11095 3387 11101
rect 3252 11064 3280 11095
rect 4154 11092 4160 11144
rect 4212 11132 4218 11144
rect 4617 11135 4675 11141
rect 4617 11132 4629 11135
rect 4212 11104 4629 11132
rect 4212 11092 4218 11104
rect 4617 11101 4629 11104
rect 4663 11101 4675 11135
rect 4617 11095 4675 11101
rect 6822 11092 6828 11144
rect 6880 11132 6886 11144
rect 7101 11135 7159 11141
rect 7101 11132 7113 11135
rect 6880 11104 7113 11132
rect 6880 11092 6886 11104
rect 7101 11101 7113 11104
rect 7147 11101 7159 11135
rect 7101 11095 7159 11101
rect 4065 11067 4123 11073
rect 4065 11064 4077 11067
rect 3252 11036 4077 11064
rect 4065 11033 4077 11036
rect 4111 11064 4123 11067
rect 4246 11064 4252 11076
rect 4111 11036 4252 11064
rect 4111 11033 4123 11036
rect 4065 11027 4123 11033
rect 4246 11024 4252 11036
rect 4304 11024 4310 11076
rect 8478 11064 8484 11076
rect 8439 11036 8484 11064
rect 8478 11024 8484 11036
rect 8536 11024 8542 11076
rect 9309 11067 9367 11073
rect 9309 11033 9321 11067
rect 9355 11064 9367 11067
rect 9398 11064 9404 11076
rect 9355 11036 9404 11064
rect 9355 11033 9367 11036
rect 9309 11027 9367 11033
rect 9398 11024 9404 11036
rect 9456 11024 9462 11076
rect 10704 11064 10732 11172
rect 11238 11160 11244 11212
rect 11296 11200 11302 11212
rect 18800 11209 18828 11240
rect 11517 11203 11575 11209
rect 11517 11200 11529 11203
rect 11296 11172 11529 11200
rect 11296 11160 11302 11172
rect 11517 11169 11529 11172
rect 11563 11169 11575 11203
rect 11517 11163 11575 11169
rect 18785 11203 18843 11209
rect 18785 11169 18797 11203
rect 18831 11200 18843 11203
rect 19337 11203 19395 11209
rect 19337 11200 19349 11203
rect 18831 11172 19349 11200
rect 18831 11169 18843 11172
rect 18785 11163 18843 11169
rect 19337 11169 19349 11172
rect 19383 11169 19395 11203
rect 19337 11163 19395 11169
rect 11333 11067 11391 11073
rect 11333 11064 11345 11067
rect 10704 11036 11345 11064
rect 11333 11033 11345 11036
rect 11379 11033 11391 11067
rect 11333 11027 11391 11033
rect 18969 11067 19027 11073
rect 18969 11033 18981 11067
rect 19015 11064 19027 11067
rect 19518 11064 19524 11076
rect 19015 11036 19524 11064
rect 19015 11033 19027 11036
rect 18969 11027 19027 11033
rect 19518 11024 19524 11036
rect 19576 11024 19582 11076
rect 3878 10956 3884 11008
rect 3936 10996 3942 11008
rect 11054 10996 11060 11008
rect 3936 10968 11060 10996
rect 3936 10956 3942 10968
rect 11054 10956 11060 10968
rect 11112 10956 11118 11008
rect 1104 10906 21896 10928
rect 1104 10854 4447 10906
rect 4499 10854 4511 10906
rect 4563 10854 4575 10906
rect 4627 10854 4639 10906
rect 4691 10854 11378 10906
rect 11430 10854 11442 10906
rect 11494 10854 11506 10906
rect 11558 10854 11570 10906
rect 11622 10854 18308 10906
rect 18360 10854 18372 10906
rect 18424 10854 18436 10906
rect 18488 10854 18500 10906
rect 18552 10854 21896 10906
rect 1104 10832 21896 10854
rect 2958 10752 2964 10804
rect 3016 10792 3022 10804
rect 3053 10795 3111 10801
rect 3053 10792 3065 10795
rect 3016 10764 3065 10792
rect 3016 10752 3022 10764
rect 3053 10761 3065 10764
rect 3099 10761 3111 10795
rect 5442 10792 5448 10804
rect 5403 10764 5448 10792
rect 3053 10755 3111 10761
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 5721 10795 5779 10801
rect 5721 10761 5733 10795
rect 5767 10792 5779 10795
rect 5810 10792 5816 10804
rect 5767 10764 5816 10792
rect 5767 10761 5779 10764
rect 5721 10755 5779 10761
rect 5810 10752 5816 10764
rect 5868 10752 5874 10804
rect 7377 10795 7435 10801
rect 7377 10761 7389 10795
rect 7423 10792 7435 10795
rect 7466 10792 7472 10804
rect 7423 10764 7472 10792
rect 7423 10761 7435 10764
rect 7377 10755 7435 10761
rect 7466 10752 7472 10764
rect 7524 10752 7530 10804
rect 7558 10752 7564 10804
rect 7616 10792 7622 10804
rect 7742 10792 7748 10804
rect 7616 10764 7748 10792
rect 7616 10752 7622 10764
rect 7742 10752 7748 10764
rect 7800 10792 7806 10804
rect 8389 10795 8447 10801
rect 8389 10792 8401 10795
rect 7800 10764 8401 10792
rect 7800 10752 7806 10764
rect 8389 10761 8401 10764
rect 8435 10761 8447 10795
rect 9122 10792 9128 10804
rect 8389 10755 8447 10761
rect 8496 10764 9128 10792
rect 8496 10724 8524 10764
rect 9122 10752 9128 10764
rect 9180 10792 9186 10804
rect 9953 10795 10011 10801
rect 9953 10792 9965 10795
rect 9180 10764 9965 10792
rect 9180 10752 9186 10764
rect 9953 10761 9965 10764
rect 9999 10761 10011 10795
rect 9953 10755 10011 10761
rect 12342 10752 12348 10804
rect 12400 10792 12406 10804
rect 12897 10795 12955 10801
rect 12897 10792 12909 10795
rect 12400 10764 12909 10792
rect 12400 10752 12406 10764
rect 12897 10761 12909 10764
rect 12943 10761 12955 10795
rect 12897 10755 12955 10761
rect 11609 10727 11667 10733
rect 11609 10724 11621 10727
rect 7852 10696 8524 10724
rect 8588 10696 11621 10724
rect 5442 10616 5448 10668
rect 5500 10656 5506 10668
rect 7852 10665 7880 10696
rect 6273 10659 6331 10665
rect 6273 10656 6285 10659
rect 5500 10628 6285 10656
rect 5500 10616 5506 10628
rect 6273 10625 6285 10628
rect 6319 10625 6331 10659
rect 6273 10619 6331 10625
rect 7837 10659 7895 10665
rect 7837 10625 7849 10659
rect 7883 10625 7895 10659
rect 7837 10619 7895 10625
rect 8021 10659 8079 10665
rect 8021 10625 8033 10659
rect 8067 10656 8079 10659
rect 8202 10656 8208 10668
rect 8067 10628 8208 10656
rect 8067 10625 8079 10628
rect 8021 10619 8079 10625
rect 8202 10616 8208 10628
rect 8260 10616 8266 10668
rect 1673 10591 1731 10597
rect 1673 10557 1685 10591
rect 1719 10588 1731 10591
rect 2406 10588 2412 10600
rect 1719 10560 2412 10588
rect 1719 10557 1731 10560
rect 1673 10551 1731 10557
rect 2406 10548 2412 10560
rect 2464 10588 2470 10600
rect 4065 10591 4123 10597
rect 4065 10588 4077 10591
rect 2464 10560 4077 10588
rect 2464 10548 2470 10560
rect 4065 10557 4077 10560
rect 4111 10588 4123 10591
rect 4154 10588 4160 10600
rect 4111 10560 4160 10588
rect 4111 10557 4123 10560
rect 4065 10551 4123 10557
rect 4154 10548 4160 10560
rect 4212 10548 4218 10600
rect 4338 10597 4344 10600
rect 4332 10588 4344 10597
rect 4299 10560 4344 10588
rect 4332 10551 4344 10560
rect 4338 10548 4344 10551
rect 4396 10548 4402 10600
rect 5810 10548 5816 10600
rect 5868 10588 5874 10600
rect 8588 10597 8616 10696
rect 11609 10693 11621 10696
rect 11655 10724 11667 10727
rect 11790 10724 11796 10736
rect 11655 10696 11796 10724
rect 11655 10693 11667 10696
rect 11609 10687 11667 10693
rect 11790 10684 11796 10696
rect 11848 10684 11854 10736
rect 18509 10727 18567 10733
rect 18509 10693 18521 10727
rect 18555 10724 18567 10727
rect 19150 10724 19156 10736
rect 18555 10696 19156 10724
rect 18555 10693 18567 10696
rect 18509 10687 18567 10693
rect 19150 10684 19156 10696
rect 19208 10684 19214 10736
rect 9490 10656 9496 10668
rect 9451 10628 9496 10656
rect 9490 10616 9496 10628
rect 9548 10616 9554 10668
rect 9600 10628 18368 10656
rect 7009 10591 7067 10597
rect 7009 10588 7021 10591
rect 5868 10560 7021 10588
rect 5868 10548 5874 10560
rect 7009 10557 7021 10560
rect 7055 10588 7067 10591
rect 7745 10591 7803 10597
rect 7745 10588 7757 10591
rect 7055 10560 7757 10588
rect 7055 10557 7067 10560
rect 7009 10551 7067 10557
rect 7745 10557 7757 10560
rect 7791 10557 7803 10591
rect 7745 10551 7803 10557
rect 8573 10591 8631 10597
rect 8573 10557 8585 10591
rect 8619 10557 8631 10591
rect 8573 10551 8631 10557
rect 1940 10523 1998 10529
rect 1940 10489 1952 10523
rect 1986 10520 1998 10523
rect 2958 10520 2964 10532
rect 1986 10492 2964 10520
rect 1986 10489 1998 10492
rect 1940 10483 1998 10489
rect 2958 10480 2964 10492
rect 3016 10480 3022 10532
rect 3970 10480 3976 10532
rect 4028 10520 4034 10532
rect 9600 10520 9628 10628
rect 11238 10548 11244 10600
rect 11296 10588 11302 10600
rect 18340 10597 18368 10628
rect 13081 10591 13139 10597
rect 13081 10588 13093 10591
rect 11296 10560 13093 10588
rect 11296 10548 11302 10560
rect 13081 10557 13093 10560
rect 13127 10557 13139 10591
rect 13081 10551 13139 10557
rect 18325 10591 18383 10597
rect 18325 10557 18337 10591
rect 18371 10588 18383 10591
rect 18877 10591 18935 10597
rect 18877 10588 18889 10591
rect 18371 10560 18889 10588
rect 18371 10557 18383 10560
rect 18325 10551 18383 10557
rect 18877 10557 18889 10560
rect 18923 10557 18935 10591
rect 18877 10551 18935 10557
rect 4028 10492 9628 10520
rect 10321 10523 10379 10529
rect 4028 10480 4034 10492
rect 10321 10489 10333 10523
rect 10367 10520 10379 10523
rect 10367 10492 12572 10520
rect 10367 10489 10379 10492
rect 10321 10483 10379 10489
rect 3789 10455 3847 10461
rect 3789 10421 3801 10455
rect 3835 10452 3847 10455
rect 3878 10452 3884 10464
rect 3835 10424 3884 10452
rect 3835 10421 3847 10424
rect 3789 10415 3847 10421
rect 3878 10412 3884 10424
rect 3936 10412 3942 10464
rect 4154 10412 4160 10464
rect 4212 10452 4218 10464
rect 6089 10455 6147 10461
rect 6089 10452 6101 10455
rect 4212 10424 6101 10452
rect 4212 10412 4218 10424
rect 6089 10421 6101 10424
rect 6135 10421 6147 10455
rect 6089 10415 6147 10421
rect 6178 10412 6184 10464
rect 6236 10452 6242 10464
rect 8938 10452 8944 10464
rect 6236 10424 6281 10452
rect 8899 10424 8944 10452
rect 6236 10412 6242 10424
rect 8938 10412 8944 10424
rect 8996 10412 9002 10464
rect 9306 10452 9312 10464
rect 9267 10424 9312 10452
rect 9306 10412 9312 10424
rect 9364 10412 9370 10464
rect 9401 10455 9459 10461
rect 9401 10421 9413 10455
rect 9447 10452 9459 10455
rect 9674 10452 9680 10464
rect 9447 10424 9680 10452
rect 9447 10421 9459 10424
rect 9401 10415 9459 10421
rect 9674 10412 9680 10424
rect 9732 10412 9738 10464
rect 12544 10461 12572 10492
rect 12529 10455 12587 10461
rect 12529 10421 12541 10455
rect 12575 10452 12587 10455
rect 20714 10452 20720 10464
rect 12575 10424 20720 10452
rect 12575 10421 12587 10424
rect 12529 10415 12587 10421
rect 20714 10412 20720 10424
rect 20772 10412 20778 10464
rect 1104 10362 21896 10384
rect 1104 10310 7912 10362
rect 7964 10310 7976 10362
rect 8028 10310 8040 10362
rect 8092 10310 8104 10362
rect 8156 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 15035 10362
rect 15087 10310 21896 10362
rect 1104 10288 21896 10310
rect 4154 10248 4160 10260
rect 4115 10220 4160 10248
rect 4154 10208 4160 10220
rect 4212 10208 4218 10260
rect 4617 10251 4675 10257
rect 4617 10217 4629 10251
rect 4663 10248 4675 10251
rect 6178 10248 6184 10260
rect 4663 10220 6184 10248
rect 4663 10217 4675 10220
rect 4617 10211 4675 10217
rect 6178 10208 6184 10220
rect 6236 10208 6242 10260
rect 7190 10208 7196 10260
rect 7248 10248 7254 10260
rect 7377 10251 7435 10257
rect 7377 10248 7389 10251
rect 7248 10220 7389 10248
rect 7248 10208 7254 10220
rect 7377 10217 7389 10220
rect 7423 10217 7435 10251
rect 7377 10211 7435 10217
rect 7837 10251 7895 10257
rect 7837 10217 7849 10251
rect 7883 10248 7895 10251
rect 8938 10248 8944 10260
rect 7883 10220 8944 10248
rect 7883 10217 7895 10220
rect 7837 10211 7895 10217
rect 8938 10208 8944 10220
rect 8996 10208 9002 10260
rect 9306 10208 9312 10260
rect 9364 10248 9370 10260
rect 9677 10251 9735 10257
rect 9677 10248 9689 10251
rect 9364 10220 9689 10248
rect 9364 10208 9370 10220
rect 9677 10217 9689 10220
rect 9723 10217 9735 10251
rect 9677 10211 9735 10217
rect 10689 10251 10747 10257
rect 10689 10217 10701 10251
rect 10735 10248 10747 10251
rect 11238 10248 11244 10260
rect 10735 10220 11244 10248
rect 10735 10217 10747 10220
rect 10689 10211 10747 10217
rect 11238 10208 11244 10220
rect 11296 10208 11302 10260
rect 2041 10183 2099 10189
rect 2041 10149 2053 10183
rect 2087 10180 2099 10183
rect 2777 10183 2835 10189
rect 2777 10180 2789 10183
rect 2087 10152 2789 10180
rect 2087 10149 2099 10152
rect 2041 10143 2099 10149
rect 2777 10149 2789 10152
rect 2823 10180 2835 10183
rect 5810 10180 5816 10192
rect 2823 10152 3832 10180
rect 2823 10149 2835 10152
rect 2777 10143 2835 10149
rect 2685 10115 2743 10121
rect 2685 10081 2697 10115
rect 2731 10112 2743 10115
rect 3329 10115 3387 10121
rect 3329 10112 3341 10115
rect 2731 10084 3341 10112
rect 2731 10081 2743 10084
rect 2685 10075 2743 10081
rect 3329 10081 3341 10084
rect 3375 10081 3387 10115
rect 3329 10075 3387 10081
rect 2869 10047 2927 10053
rect 2869 10013 2881 10047
rect 2915 10013 2927 10047
rect 3804 10044 3832 10152
rect 5000 10152 5816 10180
rect 3878 10072 3884 10124
rect 3936 10112 3942 10124
rect 5000 10121 5028 10152
rect 5810 10140 5816 10152
rect 5868 10140 5874 10192
rect 5902 10140 5908 10192
rect 5960 10180 5966 10192
rect 6089 10183 6147 10189
rect 6089 10180 6101 10183
rect 5960 10152 6101 10180
rect 5960 10140 5966 10152
rect 6089 10149 6101 10152
rect 6135 10180 6147 10183
rect 6641 10183 6699 10189
rect 6641 10180 6653 10183
rect 6135 10152 6653 10180
rect 6135 10149 6147 10152
rect 6089 10143 6147 10149
rect 6641 10149 6653 10152
rect 6687 10149 6699 10183
rect 8754 10180 8760 10192
rect 6641 10143 6699 10149
rect 6748 10152 8760 10180
rect 4985 10115 5043 10121
rect 4985 10112 4997 10115
rect 3936 10084 4997 10112
rect 3936 10072 3942 10084
rect 4985 10081 4997 10084
rect 5031 10081 5043 10115
rect 4985 10075 5043 10081
rect 5077 10115 5135 10121
rect 5077 10081 5089 10115
rect 5123 10112 5135 10115
rect 5350 10112 5356 10124
rect 5123 10084 5356 10112
rect 5123 10081 5135 10084
rect 5077 10075 5135 10081
rect 5350 10072 5356 10084
rect 5408 10072 5414 10124
rect 5718 10072 5724 10124
rect 5776 10112 5782 10124
rect 5997 10115 6055 10121
rect 5997 10112 6009 10115
rect 5776 10084 6009 10112
rect 5776 10072 5782 10084
rect 5997 10081 6009 10084
rect 6043 10081 6055 10115
rect 5997 10075 6055 10081
rect 4154 10044 4160 10056
rect 3804 10016 4160 10044
rect 2869 10007 2927 10013
rect 2682 9936 2688 9988
rect 2740 9976 2746 9988
rect 2884 9976 2912 10007
rect 4154 10004 4160 10016
rect 4212 10004 4218 10056
rect 4338 10004 4344 10056
rect 4396 10044 4402 10056
rect 5169 10047 5227 10053
rect 5169 10044 5181 10047
rect 4396 10016 5181 10044
rect 4396 10004 4402 10016
rect 5169 10013 5181 10016
rect 5215 10013 5227 10047
rect 6178 10044 6184 10056
rect 5169 10007 5227 10013
rect 5276 10016 5764 10044
rect 6139 10016 6184 10044
rect 2740 9948 2912 9976
rect 2740 9936 2746 9948
rect 3142 9936 3148 9988
rect 3200 9976 3206 9988
rect 5276 9976 5304 10016
rect 5626 9976 5632 9988
rect 3200 9948 5304 9976
rect 5587 9948 5632 9976
rect 3200 9936 3206 9948
rect 5626 9936 5632 9948
rect 5684 9936 5690 9988
rect 5736 9976 5764 10016
rect 6178 10004 6184 10016
rect 6236 10004 6242 10056
rect 6748 9976 6776 10152
rect 8754 10140 8760 10152
rect 8812 10140 8818 10192
rect 6914 10072 6920 10124
rect 6972 10112 6978 10124
rect 7009 10115 7067 10121
rect 7009 10112 7021 10115
rect 6972 10084 7021 10112
rect 6972 10072 6978 10084
rect 7009 10081 7021 10084
rect 7055 10081 7067 10115
rect 7742 10112 7748 10124
rect 7703 10084 7748 10112
rect 7009 10075 7067 10081
rect 7024 10044 7052 10075
rect 7742 10072 7748 10084
rect 7800 10072 7806 10124
rect 8849 10115 8907 10121
rect 8849 10112 8861 10115
rect 7852 10084 8861 10112
rect 7852 10044 7880 10084
rect 8849 10081 8861 10084
rect 8895 10081 8907 10115
rect 8849 10075 8907 10081
rect 9582 10072 9588 10124
rect 9640 10112 9646 10124
rect 10045 10115 10103 10121
rect 10045 10112 10057 10115
rect 9640 10084 10057 10112
rect 9640 10072 9646 10084
rect 10045 10081 10057 10084
rect 10091 10081 10103 10115
rect 10045 10075 10103 10081
rect 10873 10115 10931 10121
rect 10873 10081 10885 10115
rect 10919 10112 10931 10115
rect 11238 10112 11244 10124
rect 10919 10084 11244 10112
rect 10919 10081 10931 10084
rect 10873 10075 10931 10081
rect 11238 10072 11244 10084
rect 11296 10072 11302 10124
rect 11416 10115 11474 10121
rect 11416 10081 11428 10115
rect 11462 10112 11474 10115
rect 11698 10112 11704 10124
rect 11462 10084 11704 10112
rect 11462 10081 11474 10084
rect 11416 10075 11474 10081
rect 11698 10072 11704 10084
rect 11756 10072 11762 10124
rect 7024 10016 7880 10044
rect 8021 10047 8079 10053
rect 8021 10013 8033 10047
rect 8067 10044 8079 10047
rect 8202 10044 8208 10056
rect 8067 10016 8208 10044
rect 8067 10013 8079 10016
rect 8021 10007 8079 10013
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 9033 10047 9091 10053
rect 9033 10013 9045 10047
rect 9079 10013 9091 10047
rect 9033 10007 9091 10013
rect 7282 9976 7288 9988
rect 5736 9948 6776 9976
rect 6932 9948 7288 9976
rect 2317 9911 2375 9917
rect 2317 9877 2329 9911
rect 2363 9908 2375 9911
rect 3602 9908 3608 9920
rect 2363 9880 3608 9908
rect 2363 9877 2375 9880
rect 2317 9871 2375 9877
rect 3602 9868 3608 9880
rect 3660 9868 3666 9920
rect 4154 9868 4160 9920
rect 4212 9908 4218 9920
rect 6932 9908 6960 9948
rect 7282 9936 7288 9948
rect 7340 9936 7346 9988
rect 9048 9976 9076 10007
rect 9214 10004 9220 10056
rect 9272 10044 9278 10056
rect 10137 10047 10195 10053
rect 10137 10044 10149 10047
rect 9272 10016 10149 10044
rect 9272 10004 9278 10016
rect 10137 10013 10149 10016
rect 10183 10013 10195 10047
rect 10318 10044 10324 10056
rect 10279 10016 10324 10044
rect 10137 10007 10195 10013
rect 10318 10004 10324 10016
rect 10376 10004 10382 10056
rect 11149 10047 11207 10053
rect 11149 10013 11161 10047
rect 11195 10013 11207 10047
rect 11149 10007 11207 10013
rect 10336 9976 10364 10004
rect 9048 9948 10364 9976
rect 8386 9908 8392 9920
rect 4212 9880 6960 9908
rect 8347 9880 8392 9908
rect 4212 9868 4218 9880
rect 8386 9868 8392 9880
rect 8444 9868 8450 9920
rect 11164 9908 11192 10007
rect 12342 9908 12348 9920
rect 11164 9880 12348 9908
rect 12342 9868 12348 9880
rect 12400 9868 12406 9920
rect 12526 9908 12532 9920
rect 12487 9880 12532 9908
rect 12526 9868 12532 9880
rect 12584 9868 12590 9920
rect 1104 9818 21896 9840
rect 1104 9766 4447 9818
rect 4499 9766 4511 9818
rect 4563 9766 4575 9818
rect 4627 9766 4639 9818
rect 4691 9766 11378 9818
rect 11430 9766 11442 9818
rect 11494 9766 11506 9818
rect 11558 9766 11570 9818
rect 11622 9766 18308 9818
rect 18360 9766 18372 9818
rect 18424 9766 18436 9818
rect 18488 9766 18500 9818
rect 18552 9766 21896 9818
rect 1104 9744 21896 9766
rect 3970 9664 3976 9716
rect 4028 9704 4034 9716
rect 14182 9704 14188 9716
rect 4028 9676 14188 9704
rect 4028 9664 4034 9676
rect 14182 9664 14188 9676
rect 14240 9664 14246 9716
rect 2958 9636 2964 9648
rect 2919 9608 2964 9636
rect 2958 9596 2964 9608
rect 3016 9596 3022 9648
rect 3234 9636 3240 9648
rect 3195 9608 3240 9636
rect 3234 9596 3240 9608
rect 3292 9596 3298 9648
rect 3326 9596 3332 9648
rect 3384 9636 3390 9648
rect 3694 9636 3700 9648
rect 3384 9608 3700 9636
rect 3384 9596 3390 9608
rect 3694 9596 3700 9608
rect 3752 9596 3758 9648
rect 4062 9596 4068 9648
rect 4120 9636 4126 9648
rect 4525 9639 4583 9645
rect 4525 9636 4537 9639
rect 4120 9608 4537 9636
rect 4120 9596 4126 9608
rect 4525 9605 4537 9608
rect 4571 9605 4583 9639
rect 4525 9599 4583 9605
rect 12342 9596 12348 9648
rect 12400 9636 12406 9648
rect 15197 9639 15255 9645
rect 12400 9608 13860 9636
rect 12400 9596 12406 9608
rect 2976 9568 3004 9596
rect 3789 9571 3847 9577
rect 3789 9568 3801 9571
rect 2976 9540 3801 9568
rect 3789 9537 3801 9540
rect 3835 9537 3847 9571
rect 3789 9531 3847 9537
rect 5169 9571 5227 9577
rect 5169 9537 5181 9571
rect 5215 9568 5227 9571
rect 5442 9568 5448 9580
rect 5215 9540 5448 9568
rect 5215 9537 5227 9540
rect 5169 9531 5227 9537
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 11425 9571 11483 9577
rect 11425 9568 11437 9571
rect 10796 9540 11437 9568
rect 10796 9512 10824 9540
rect 11425 9537 11437 9540
rect 11471 9537 11483 9571
rect 11425 9531 11483 9537
rect 11609 9571 11667 9577
rect 11609 9537 11621 9571
rect 11655 9537 11667 9571
rect 11609 9531 11667 9537
rect 1581 9503 1639 9509
rect 1581 9469 1593 9503
rect 1627 9469 1639 9503
rect 1581 9463 1639 9469
rect 1848 9503 1906 9509
rect 1848 9469 1860 9503
rect 1894 9500 1906 9503
rect 2682 9500 2688 9512
rect 1894 9472 2688 9500
rect 1894 9469 1906 9472
rect 1848 9463 1906 9469
rect 1596 9364 1624 9463
rect 2682 9460 2688 9472
rect 2740 9460 2746 9512
rect 3602 9500 3608 9512
rect 3563 9472 3608 9500
rect 3602 9460 3608 9472
rect 3660 9460 3666 9512
rect 6638 9500 6644 9512
rect 3804 9472 6644 9500
rect 3804 9444 3832 9472
rect 6638 9460 6644 9472
rect 6696 9460 6702 9512
rect 6822 9500 6828 9512
rect 6783 9472 6828 9500
rect 6822 9460 6828 9472
rect 6880 9500 6886 9512
rect 9309 9503 9367 9509
rect 9309 9500 9321 9503
rect 6880 9472 9321 9500
rect 6880 9460 6886 9472
rect 9309 9469 9321 9472
rect 9355 9500 9367 9503
rect 9858 9500 9864 9512
rect 9355 9472 9864 9500
rect 9355 9469 9367 9472
rect 9309 9463 9367 9469
rect 9858 9460 9864 9472
rect 9916 9500 9922 9512
rect 10502 9500 10508 9512
rect 9916 9472 10508 9500
rect 9916 9460 9922 9472
rect 10502 9460 10508 9472
rect 10560 9460 10566 9512
rect 10778 9460 10784 9512
rect 10836 9460 10842 9512
rect 11054 9460 11060 9512
rect 11112 9500 11118 9512
rect 11333 9503 11391 9509
rect 11333 9500 11345 9503
rect 11112 9472 11345 9500
rect 11112 9460 11118 9472
rect 11333 9469 11345 9472
rect 11379 9469 11391 9503
rect 11624 9500 11652 9531
rect 12526 9528 12532 9580
rect 12584 9568 12590 9580
rect 13832 9577 13860 9608
rect 15197 9605 15209 9639
rect 15243 9605 15255 9639
rect 15197 9599 15255 9605
rect 12989 9571 13047 9577
rect 12989 9568 13001 9571
rect 12584 9540 13001 9568
rect 12584 9528 12590 9540
rect 12989 9537 13001 9540
rect 13035 9537 13047 9571
rect 12989 9531 13047 9537
rect 13817 9571 13875 9577
rect 13817 9537 13829 9571
rect 13863 9537 13875 9571
rect 13817 9531 13875 9537
rect 11698 9500 11704 9512
rect 11611 9472 11704 9500
rect 11333 9463 11391 9469
rect 11698 9460 11704 9472
rect 11756 9500 11762 9512
rect 15212 9500 15240 9599
rect 11756 9472 15240 9500
rect 11756 9460 11762 9472
rect 3786 9392 3792 9444
rect 3844 9392 3850 9444
rect 4798 9392 4804 9444
rect 4856 9432 4862 9444
rect 4985 9435 5043 9441
rect 4985 9432 4997 9435
rect 4856 9404 4997 9432
rect 4856 9392 4862 9404
rect 4985 9401 4997 9404
rect 5031 9401 5043 9435
rect 4985 9395 5043 9401
rect 7092 9435 7150 9441
rect 7092 9401 7104 9435
rect 7138 9432 7150 9435
rect 7190 9432 7196 9444
rect 7138 9404 7196 9432
rect 7138 9401 7150 9404
rect 7092 9395 7150 9401
rect 7190 9392 7196 9404
rect 7248 9392 7254 9444
rect 8941 9435 8999 9441
rect 8941 9432 8953 9435
rect 7291 9404 8953 9432
rect 1854 9364 1860 9376
rect 1596 9336 1860 9364
rect 1854 9324 1860 9336
rect 1912 9324 1918 9376
rect 3694 9364 3700 9376
rect 3655 9336 3700 9364
rect 3694 9324 3700 9336
rect 3752 9324 3758 9376
rect 4890 9364 4896 9376
rect 4851 9336 4896 9364
rect 4890 9324 4896 9336
rect 4948 9324 4954 9376
rect 5350 9324 5356 9376
rect 5408 9364 5414 9376
rect 5537 9367 5595 9373
rect 5537 9364 5549 9367
rect 5408 9336 5549 9364
rect 5408 9324 5414 9336
rect 5537 9333 5549 9336
rect 5583 9333 5595 9367
rect 5537 9327 5595 9333
rect 5718 9324 5724 9376
rect 5776 9364 5782 9376
rect 5905 9367 5963 9373
rect 5905 9364 5917 9367
rect 5776 9336 5917 9364
rect 5776 9324 5782 9336
rect 5905 9333 5917 9336
rect 5951 9364 5963 9367
rect 7291 9364 7319 9404
rect 8941 9401 8953 9404
rect 8987 9432 8999 9435
rect 9214 9432 9220 9444
rect 8987 9404 9220 9432
rect 8987 9401 8999 9404
rect 8941 9395 8999 9401
rect 9214 9392 9220 9404
rect 9272 9392 9278 9444
rect 9576 9435 9634 9441
rect 9576 9401 9588 9435
rect 9622 9432 9634 9435
rect 10318 9432 10324 9444
rect 9622 9404 10324 9432
rect 9622 9401 9634 9404
rect 9576 9395 9634 9401
rect 10318 9392 10324 9404
rect 10376 9392 10382 9444
rect 12897 9435 12955 9441
rect 12897 9432 12909 9435
rect 10980 9404 12909 9432
rect 8202 9364 8208 9376
rect 5951 9336 7319 9364
rect 8163 9336 8208 9364
rect 5951 9333 5963 9336
rect 5905 9327 5963 9333
rect 8202 9324 8208 9336
rect 8260 9324 8266 9376
rect 8478 9364 8484 9376
rect 8439 9336 8484 9364
rect 8478 9324 8484 9336
rect 8536 9324 8542 9376
rect 9490 9324 9496 9376
rect 9548 9364 9554 9376
rect 10980 9373 11008 9404
rect 12897 9401 12909 9404
rect 12943 9401 12955 9435
rect 12897 9395 12955 9401
rect 14084 9435 14142 9441
rect 14084 9401 14096 9435
rect 14130 9432 14142 9435
rect 14642 9432 14648 9444
rect 14130 9404 14648 9432
rect 14130 9401 14142 9404
rect 14084 9395 14142 9401
rect 14642 9392 14648 9404
rect 14700 9392 14706 9444
rect 10689 9367 10747 9373
rect 10689 9364 10701 9367
rect 9548 9336 10701 9364
rect 9548 9324 9554 9336
rect 10689 9333 10701 9336
rect 10735 9333 10747 9367
rect 10689 9327 10747 9333
rect 10965 9367 11023 9373
rect 10965 9333 10977 9367
rect 11011 9333 11023 9367
rect 10965 9327 11023 9333
rect 12437 9367 12495 9373
rect 12437 9333 12449 9367
rect 12483 9364 12495 9367
rect 12618 9364 12624 9376
rect 12483 9336 12624 9364
rect 12483 9333 12495 9336
rect 12437 9327 12495 9333
rect 12618 9324 12624 9336
rect 12676 9324 12682 9376
rect 12802 9364 12808 9376
rect 12763 9336 12808 9364
rect 12802 9324 12808 9336
rect 12860 9324 12866 9376
rect 1104 9274 21896 9296
rect 1104 9222 7912 9274
rect 7964 9222 7976 9274
rect 8028 9222 8040 9274
rect 8092 9222 8104 9274
rect 8156 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 15035 9274
rect 15087 9222 21896 9274
rect 1104 9200 21896 9222
rect 2409 9163 2467 9169
rect 2409 9129 2421 9163
rect 2455 9160 2467 9163
rect 3694 9160 3700 9172
rect 2455 9132 3700 9160
rect 2455 9129 2467 9132
rect 2409 9123 2467 9129
rect 3694 9120 3700 9132
rect 3752 9120 3758 9172
rect 4525 9163 4583 9169
rect 4525 9129 4537 9163
rect 4571 9160 4583 9163
rect 4890 9160 4896 9172
rect 4571 9132 4896 9160
rect 4571 9129 4583 9132
rect 4525 9123 4583 9129
rect 4890 9120 4896 9132
rect 4948 9120 4954 9172
rect 5074 9120 5080 9172
rect 5132 9160 5138 9172
rect 6730 9160 6736 9172
rect 5132 9132 6736 9160
rect 5132 9120 5138 9132
rect 6730 9120 6736 9132
rect 6788 9120 6794 9172
rect 7742 9160 7748 9172
rect 7703 9132 7748 9160
rect 7742 9120 7748 9132
rect 7800 9120 7806 9172
rect 8113 9163 8171 9169
rect 8113 9129 8125 9163
rect 8159 9160 8171 9163
rect 8478 9160 8484 9172
rect 8159 9132 8484 9160
rect 8159 9129 8171 9132
rect 8113 9123 8171 9129
rect 8478 9120 8484 9132
rect 8536 9120 8542 9172
rect 8754 9160 8760 9172
rect 8715 9132 8760 9160
rect 8754 9120 8760 9132
rect 8812 9120 8818 9172
rect 9674 9160 9680 9172
rect 9635 9132 9680 9160
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 11054 9120 11060 9172
rect 11112 9160 11118 9172
rect 11149 9163 11207 9169
rect 11149 9160 11161 9163
rect 11112 9132 11161 9160
rect 11112 9120 11118 9132
rect 11149 9129 11161 9132
rect 11195 9129 11207 9163
rect 11149 9123 11207 9129
rect 11698 9120 11704 9172
rect 11756 9160 11762 9172
rect 12342 9160 12348 9172
rect 11756 9132 12348 9160
rect 11756 9120 11762 9132
rect 12342 9120 12348 9132
rect 12400 9120 12406 9172
rect 2682 9052 2688 9104
rect 2740 9092 2746 9104
rect 2740 9064 3096 9092
rect 2740 9052 2746 9064
rect 2774 8984 2780 9036
rect 2832 9024 2838 9036
rect 2832 8996 2877 9024
rect 2832 8984 2838 8996
rect 3068 8968 3096 9064
rect 4062 9052 4068 9104
rect 4120 9092 4126 9104
rect 8205 9095 8263 9101
rect 4120 9064 7696 9092
rect 4120 9052 4126 9064
rect 4893 9027 4951 9033
rect 4893 8993 4905 9027
rect 4939 9024 4951 9027
rect 5626 9024 5632 9036
rect 4939 8996 5632 9024
rect 4939 8993 4951 8996
rect 4893 8987 4951 8993
rect 5626 8984 5632 8996
rect 5684 8984 5690 9036
rect 5804 9027 5862 9033
rect 5804 8993 5816 9027
rect 5850 9024 5862 9027
rect 6086 9024 6092 9036
rect 5850 8996 6092 9024
rect 5850 8993 5862 8996
rect 5804 8987 5862 8993
rect 6086 8984 6092 8996
rect 6144 8984 6150 9036
rect 7377 9027 7435 9033
rect 7377 8993 7389 9027
rect 7423 9024 7435 9027
rect 7558 9024 7564 9036
rect 7423 8996 7564 9024
rect 7423 8993 7435 8996
rect 7377 8987 7435 8993
rect 7558 8984 7564 8996
rect 7616 8984 7622 9036
rect 7668 9024 7696 9064
rect 8205 9061 8217 9095
rect 8251 9092 8263 9095
rect 8386 9092 8392 9104
rect 8251 9064 8392 9092
rect 8251 9061 8263 9064
rect 8205 9055 8263 9061
rect 8386 9052 8392 9064
rect 8444 9052 8450 9104
rect 11968 9095 12026 9101
rect 8496 9064 10180 9092
rect 8496 9024 8524 9064
rect 10042 9024 10048 9036
rect 7668 8996 8524 9024
rect 10003 8996 10048 9024
rect 10042 8984 10048 8996
rect 10100 8984 10106 9036
rect 10152 9024 10180 9064
rect 11968 9061 11980 9095
rect 12014 9092 12026 9095
rect 12526 9092 12532 9104
rect 12014 9064 12532 9092
rect 12014 9061 12026 9064
rect 11968 9055 12026 9061
rect 12526 9052 12532 9064
rect 12584 9052 12590 9104
rect 14366 9024 14372 9036
rect 10152 8996 14372 9024
rect 14366 8984 14372 8996
rect 14424 8984 14430 9036
rect 14461 9027 14519 9033
rect 14461 8993 14473 9027
rect 14507 9024 14519 9027
rect 15102 9024 15108 9036
rect 14507 8996 15108 9024
rect 14507 8993 14519 8996
rect 14461 8987 14519 8993
rect 15102 8984 15108 8996
rect 15160 8984 15166 9036
rect 2866 8956 2872 8968
rect 2827 8928 2872 8956
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 3050 8956 3056 8968
rect 3011 8928 3056 8956
rect 3050 8916 3056 8928
rect 3108 8916 3114 8968
rect 4985 8959 5043 8965
rect 4985 8925 4997 8959
rect 5031 8925 5043 8959
rect 4985 8919 5043 8925
rect 5169 8959 5227 8965
rect 5169 8925 5181 8959
rect 5215 8925 5227 8959
rect 5169 8919 5227 8925
rect 4154 8888 4160 8900
rect 4115 8860 4160 8888
rect 4154 8848 4160 8860
rect 4212 8888 4218 8900
rect 5000 8888 5028 8919
rect 4212 8860 5028 8888
rect 4212 8848 4218 8860
rect 4246 8780 4252 8832
rect 4304 8820 4310 8832
rect 4982 8820 4988 8832
rect 4304 8792 4988 8820
rect 4304 8780 4310 8792
rect 4982 8780 4988 8792
rect 5040 8780 5046 8832
rect 5074 8780 5080 8832
rect 5132 8820 5138 8832
rect 5184 8820 5212 8919
rect 5258 8916 5264 8968
rect 5316 8956 5322 8968
rect 5537 8959 5595 8965
rect 5537 8956 5549 8959
rect 5316 8928 5549 8956
rect 5316 8916 5322 8928
rect 5537 8925 5549 8928
rect 5583 8925 5595 8959
rect 5537 8919 5595 8925
rect 7190 8916 7196 8968
rect 7248 8956 7254 8968
rect 8389 8959 8447 8965
rect 8389 8956 8401 8959
rect 7248 8928 8401 8956
rect 7248 8916 7254 8928
rect 8389 8925 8401 8928
rect 8435 8956 8447 8959
rect 9490 8956 9496 8968
rect 8435 8928 9496 8956
rect 8435 8925 8447 8928
rect 8389 8919 8447 8925
rect 9490 8916 9496 8928
rect 9548 8916 9554 8968
rect 10137 8959 10195 8965
rect 10137 8925 10149 8959
rect 10183 8925 10195 8959
rect 10318 8956 10324 8968
rect 10231 8928 10324 8956
rect 10137 8919 10195 8925
rect 6638 8848 6644 8900
rect 6696 8888 6702 8900
rect 10152 8888 10180 8919
rect 10318 8916 10324 8928
rect 10376 8956 10382 8968
rect 11698 8956 11704 8968
rect 10376 8928 11284 8956
rect 11659 8928 11704 8956
rect 10376 8916 10382 8928
rect 10594 8888 10600 8900
rect 6696 8860 10088 8888
rect 10152 8860 10600 8888
rect 6696 8848 6702 8860
rect 6917 8823 6975 8829
rect 6917 8820 6929 8823
rect 5132 8792 6929 8820
rect 5132 8780 5138 8792
rect 6917 8789 6929 8792
rect 6963 8789 6975 8823
rect 7190 8820 7196 8832
rect 7151 8792 7196 8820
rect 6917 8783 6975 8789
rect 7190 8780 7196 8792
rect 7248 8780 7254 8832
rect 8938 8780 8944 8832
rect 8996 8820 9002 8832
rect 9217 8823 9275 8829
rect 9217 8820 9229 8823
rect 8996 8792 9229 8820
rect 8996 8780 9002 8792
rect 9217 8789 9229 8792
rect 9263 8820 9275 8823
rect 9582 8820 9588 8832
rect 9263 8792 9588 8820
rect 9263 8789 9275 8792
rect 9217 8783 9275 8789
rect 9582 8780 9588 8792
rect 9640 8780 9646 8832
rect 10060 8820 10088 8860
rect 10594 8848 10600 8860
rect 10652 8848 10658 8900
rect 11054 8888 11060 8900
rect 10704 8860 11060 8888
rect 10704 8820 10732 8860
rect 11054 8848 11060 8860
rect 11112 8848 11118 8900
rect 10060 8792 10732 8820
rect 10778 8780 10784 8832
rect 10836 8820 10842 8832
rect 11256 8820 11284 8928
rect 11698 8916 11704 8928
rect 11756 8916 11762 8968
rect 14550 8956 14556 8968
rect 14511 8928 14556 8956
rect 14550 8916 14556 8928
rect 14608 8916 14614 8968
rect 14642 8916 14648 8968
rect 14700 8956 14706 8968
rect 14700 8928 14745 8956
rect 14700 8916 14706 8928
rect 13081 8823 13139 8829
rect 13081 8820 13093 8823
rect 10836 8792 10881 8820
rect 11256 8792 13093 8820
rect 10836 8780 10842 8792
rect 13081 8789 13093 8792
rect 13127 8789 13139 8823
rect 13081 8783 13139 8789
rect 14093 8823 14151 8829
rect 14093 8789 14105 8823
rect 14139 8820 14151 8823
rect 16482 8820 16488 8832
rect 14139 8792 16488 8820
rect 14139 8789 14151 8792
rect 14093 8783 14151 8789
rect 16482 8780 16488 8792
rect 16540 8780 16546 8832
rect 1104 8730 21896 8752
rect 1104 8678 4447 8730
rect 4499 8678 4511 8730
rect 4563 8678 4575 8730
rect 4627 8678 4639 8730
rect 4691 8678 11378 8730
rect 11430 8678 11442 8730
rect 11494 8678 11506 8730
rect 11558 8678 11570 8730
rect 11622 8678 18308 8730
rect 18360 8678 18372 8730
rect 18424 8678 18436 8730
rect 18488 8678 18500 8730
rect 18552 8678 21896 8730
rect 1104 8656 21896 8678
rect 3050 8576 3056 8628
rect 3108 8616 3114 8628
rect 3329 8619 3387 8625
rect 3329 8616 3341 8619
rect 3108 8588 3341 8616
rect 3108 8576 3114 8588
rect 3329 8585 3341 8588
rect 3375 8585 3387 8619
rect 5258 8616 5264 8628
rect 3329 8579 3387 8585
rect 4264 8588 5264 8616
rect 4264 8489 4292 8588
rect 5258 8576 5264 8588
rect 5316 8576 5322 8628
rect 5442 8576 5448 8628
rect 5500 8616 5506 8628
rect 5629 8619 5687 8625
rect 5629 8616 5641 8619
rect 5500 8588 5641 8616
rect 5500 8576 5506 8588
rect 5629 8585 5641 8588
rect 5675 8585 5687 8619
rect 5629 8579 5687 8585
rect 6086 8576 6092 8628
rect 6144 8616 6150 8628
rect 8389 8619 8447 8625
rect 8389 8616 8401 8619
rect 6144 8588 8401 8616
rect 6144 8576 6150 8588
rect 8389 8585 8401 8588
rect 8435 8585 8447 8619
rect 8389 8579 8447 8585
rect 11238 8576 11244 8628
rect 11296 8616 11302 8628
rect 11609 8619 11667 8625
rect 11609 8616 11621 8619
rect 11296 8588 11621 8616
rect 11296 8576 11302 8588
rect 11609 8585 11621 8588
rect 11655 8616 11667 8619
rect 12158 8616 12164 8628
rect 11655 8588 12164 8616
rect 11655 8585 11667 8588
rect 11609 8579 11667 8585
rect 12158 8576 12164 8588
rect 12216 8576 12222 8628
rect 14642 8576 14648 8628
rect 14700 8616 14706 8628
rect 14829 8619 14887 8625
rect 14829 8616 14841 8619
rect 14700 8588 14841 8616
rect 14700 8576 14706 8588
rect 14829 8585 14841 8588
rect 14875 8585 14887 8619
rect 14829 8579 14887 8585
rect 12618 8508 12624 8560
rect 12676 8548 12682 8560
rect 12676 8520 13492 8548
rect 12676 8508 12682 8520
rect 4249 8483 4307 8489
rect 4249 8449 4261 8483
rect 4295 8449 4307 8483
rect 4249 8443 4307 8449
rect 5626 8440 5632 8492
rect 5684 8480 5690 8492
rect 5905 8483 5963 8489
rect 5905 8480 5917 8483
rect 5684 8452 5917 8480
rect 5684 8440 5690 8452
rect 5905 8449 5917 8452
rect 5951 8449 5963 8483
rect 5905 8443 5963 8449
rect 6822 8440 6828 8492
rect 6880 8480 6886 8492
rect 7009 8483 7067 8489
rect 7009 8480 7021 8483
rect 6880 8452 7021 8480
rect 6880 8440 6886 8452
rect 7009 8449 7021 8452
rect 7055 8449 7067 8483
rect 7009 8443 7067 8449
rect 8018 8440 8024 8492
rect 8076 8480 8082 8492
rect 9493 8483 9551 8489
rect 9493 8480 9505 8483
rect 8076 8452 9505 8480
rect 8076 8440 8082 8452
rect 9493 8449 9505 8452
rect 9539 8480 9551 8483
rect 10042 8480 10048 8492
rect 9539 8452 10048 8480
rect 9539 8449 9551 8452
rect 9493 8443 9551 8449
rect 10042 8440 10048 8452
rect 10100 8440 10106 8492
rect 12437 8483 12495 8489
rect 12437 8449 12449 8483
rect 12483 8480 12495 8483
rect 12802 8480 12808 8492
rect 12483 8452 12808 8480
rect 12483 8449 12495 8452
rect 12437 8443 12495 8449
rect 12802 8440 12808 8452
rect 12860 8440 12866 8492
rect 13464 8480 13492 8520
rect 15102 8480 15108 8492
rect 13464 8452 13584 8480
rect 15063 8452 15108 8480
rect 1854 8372 1860 8424
rect 1912 8412 1918 8424
rect 1949 8415 2007 8421
rect 1949 8412 1961 8415
rect 1912 8384 1961 8412
rect 1912 8372 1918 8384
rect 1949 8381 1961 8384
rect 1995 8381 2007 8415
rect 1949 8375 2007 8381
rect 4516 8415 4574 8421
rect 4516 8381 4528 8415
rect 4562 8412 4574 8415
rect 5074 8412 5080 8424
rect 4562 8384 5080 8412
rect 4562 8381 4574 8384
rect 4516 8375 4574 8381
rect 5074 8372 5080 8384
rect 5132 8372 5138 8424
rect 7276 8415 7334 8421
rect 7276 8381 7288 8415
rect 7322 8412 7334 8415
rect 8202 8412 8208 8424
rect 7322 8384 8208 8412
rect 7322 8381 7334 8384
rect 7276 8375 7334 8381
rect 8202 8372 8208 8384
rect 8260 8372 8266 8424
rect 10594 8412 10600 8424
rect 10555 8384 10600 8412
rect 10594 8372 10600 8384
rect 10652 8372 10658 8424
rect 11790 8412 11796 8424
rect 11751 8384 11796 8412
rect 11790 8372 11796 8384
rect 11848 8372 11854 8424
rect 11882 8372 11888 8424
rect 11940 8412 11946 8424
rect 12250 8412 12256 8424
rect 11940 8384 12256 8412
rect 11940 8372 11946 8384
rect 12250 8372 12256 8384
rect 12308 8372 12314 8424
rect 13449 8415 13507 8421
rect 13449 8381 13461 8415
rect 13495 8381 13507 8415
rect 13556 8412 13584 8452
rect 15102 8440 15108 8452
rect 15160 8440 15166 8492
rect 16853 8415 16911 8421
rect 16853 8412 16865 8415
rect 13556 8384 16865 8412
rect 13449 8375 13507 8381
rect 16853 8381 16865 8384
rect 16899 8381 16911 8415
rect 16853 8375 16911 8381
rect 2216 8347 2274 8353
rect 2216 8313 2228 8347
rect 2262 8344 2274 8347
rect 2498 8344 2504 8356
rect 2262 8316 2504 8344
rect 2262 8313 2274 8316
rect 2216 8307 2274 8313
rect 2498 8304 2504 8316
rect 2556 8304 2562 8356
rect 3326 8344 3332 8356
rect 3068 8316 3332 8344
rect 1578 8276 1584 8288
rect 1539 8248 1584 8276
rect 1578 8236 1584 8248
rect 1636 8276 1642 8288
rect 3068 8276 3096 8316
rect 3326 8304 3332 8316
rect 3384 8344 3390 8356
rect 3602 8344 3608 8356
rect 3384 8316 3608 8344
rect 3384 8304 3390 8316
rect 3602 8304 3608 8316
rect 3660 8304 3666 8356
rect 3970 8304 3976 8356
rect 4028 8344 4034 8356
rect 13354 8344 13360 8356
rect 4028 8316 13360 8344
rect 4028 8304 4034 8316
rect 13354 8304 13360 8316
rect 13412 8304 13418 8356
rect 1636 8248 3096 8276
rect 1636 8236 1642 8248
rect 3142 8236 3148 8288
rect 3200 8276 3206 8288
rect 5534 8276 5540 8288
rect 3200 8248 5540 8276
rect 3200 8236 3206 8248
rect 5534 8236 5540 8248
rect 5592 8236 5598 8288
rect 13464 8276 13492 8375
rect 13716 8347 13774 8353
rect 13716 8313 13728 8347
rect 13762 8344 13774 8347
rect 14458 8344 14464 8356
rect 13762 8316 14464 8344
rect 13762 8313 13774 8316
rect 13716 8307 13774 8313
rect 14458 8304 14464 8316
rect 14516 8304 14522 8356
rect 17129 8347 17187 8353
rect 17129 8313 17141 8347
rect 17175 8344 17187 8347
rect 18598 8344 18604 8356
rect 17175 8316 18604 8344
rect 17175 8313 17187 8316
rect 17129 8307 17187 8313
rect 18598 8304 18604 8316
rect 18656 8304 18662 8356
rect 14090 8276 14096 8288
rect 13464 8248 14096 8276
rect 14090 8236 14096 8248
rect 14148 8236 14154 8288
rect 1104 8186 21896 8208
rect 1104 8134 7912 8186
rect 7964 8134 7976 8186
rect 8028 8134 8040 8186
rect 8092 8134 8104 8186
rect 8156 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 15035 8186
rect 15087 8134 21896 8186
rect 1104 8112 21896 8134
rect 1949 8075 2007 8081
rect 1949 8041 1961 8075
rect 1995 8072 2007 8075
rect 2774 8072 2780 8084
rect 1995 8044 2780 8072
rect 1995 8041 2007 8044
rect 1949 8035 2007 8041
rect 2774 8032 2780 8044
rect 2832 8032 2838 8084
rect 2866 8032 2872 8084
rect 2924 8072 2930 8084
rect 2961 8075 3019 8081
rect 2961 8072 2973 8075
rect 2924 8044 2973 8072
rect 2924 8032 2930 8044
rect 2961 8041 2973 8044
rect 3007 8041 3019 8075
rect 2961 8035 3019 8041
rect 4433 8075 4491 8081
rect 4433 8041 4445 8075
rect 4479 8072 4491 8075
rect 4798 8072 4804 8084
rect 4479 8044 4804 8072
rect 4479 8041 4491 8044
rect 4433 8035 4491 8041
rect 4798 8032 4804 8044
rect 4856 8032 4862 8084
rect 4893 8075 4951 8081
rect 4893 8041 4905 8075
rect 4939 8072 4951 8075
rect 5445 8075 5503 8081
rect 5445 8072 5457 8075
rect 4939 8044 5457 8072
rect 4939 8041 4951 8044
rect 4893 8035 4951 8041
rect 5445 8041 5457 8044
rect 5491 8041 5503 8075
rect 5445 8035 5503 8041
rect 7377 8075 7435 8081
rect 7377 8041 7389 8075
rect 7423 8072 7435 8075
rect 8941 8075 8999 8081
rect 8941 8072 8953 8075
rect 7423 8044 8953 8072
rect 7423 8041 7435 8044
rect 7377 8035 7435 8041
rect 8941 8041 8953 8044
rect 8987 8041 8999 8075
rect 8941 8035 8999 8041
rect 13541 8075 13599 8081
rect 13541 8041 13553 8075
rect 13587 8041 13599 8075
rect 13541 8035 13599 8041
rect 13817 8075 13875 8081
rect 13817 8041 13829 8075
rect 13863 8072 13875 8075
rect 14550 8072 14556 8084
rect 13863 8044 14556 8072
rect 13863 8041 13875 8044
rect 13817 8035 13875 8041
rect 3878 8004 3884 8016
rect 2516 7976 2636 8004
rect 1578 7896 1584 7948
rect 1636 7936 1642 7948
rect 2317 7939 2375 7945
rect 2317 7936 2329 7939
rect 1636 7908 2329 7936
rect 1636 7896 1642 7908
rect 2317 7905 2329 7908
rect 2363 7905 2375 7939
rect 2516 7936 2544 7976
rect 2317 7899 2375 7905
rect 2424 7908 2544 7936
rect 2608 7936 2636 7976
rect 3344 7976 3884 8004
rect 3344 7948 3372 7976
rect 3878 7964 3884 7976
rect 3936 8004 3942 8016
rect 5813 8007 5871 8013
rect 5813 8004 5825 8007
rect 3936 7976 5825 8004
rect 3936 7964 3942 7976
rect 5813 7973 5825 7976
rect 5859 7973 5871 8007
rect 13556 8004 13584 8035
rect 14550 8032 14556 8044
rect 14608 8032 14614 8084
rect 14182 8004 14188 8016
rect 5813 7967 5871 7973
rect 8956 7976 13584 8004
rect 14143 7976 14188 8004
rect 3142 7936 3148 7948
rect 2608 7908 3148 7936
rect 2424 7877 2452 7908
rect 3142 7896 3148 7908
rect 3200 7896 3206 7948
rect 3326 7936 3332 7948
rect 3287 7908 3332 7936
rect 3326 7896 3332 7908
rect 3384 7896 3390 7948
rect 3421 7939 3479 7945
rect 3421 7905 3433 7939
rect 3467 7936 3479 7939
rect 4801 7939 4859 7945
rect 3467 7908 3924 7936
rect 3467 7905 3479 7908
rect 3421 7899 3479 7905
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7868 1731 7871
rect 2409 7871 2467 7877
rect 2409 7868 2421 7871
rect 1719 7840 2421 7868
rect 1719 7837 1731 7840
rect 1673 7831 1731 7837
rect 2409 7837 2421 7840
rect 2455 7837 2467 7871
rect 2409 7831 2467 7837
rect 2498 7828 2504 7880
rect 2556 7868 2562 7880
rect 3605 7871 3663 7877
rect 2556 7840 2601 7868
rect 2556 7828 2562 7840
rect 3605 7837 3617 7871
rect 3651 7837 3663 7871
rect 3605 7831 3663 7837
rect 3050 7760 3056 7812
rect 3108 7800 3114 7812
rect 3620 7800 3648 7831
rect 3108 7772 3648 7800
rect 3108 7760 3114 7772
rect 3896 7732 3924 7908
rect 4801 7905 4813 7939
rect 4847 7936 4859 7939
rect 5718 7936 5724 7948
rect 4847 7908 5724 7936
rect 4847 7905 4859 7908
rect 4801 7899 4859 7905
rect 5718 7896 5724 7908
rect 5776 7896 5782 7948
rect 7745 7939 7803 7945
rect 7745 7905 7757 7939
rect 7791 7905 7803 7939
rect 8846 7936 8852 7948
rect 8807 7908 8852 7936
rect 7745 7899 7803 7905
rect 5074 7868 5080 7880
rect 5035 7840 5080 7868
rect 5074 7828 5080 7840
rect 5132 7828 5138 7880
rect 5902 7868 5908 7880
rect 5863 7840 5908 7868
rect 5902 7828 5908 7840
rect 5960 7828 5966 7880
rect 6086 7868 6092 7880
rect 6047 7840 6092 7868
rect 6086 7828 6092 7840
rect 6144 7828 6150 7880
rect 3970 7760 3976 7812
rect 4028 7800 4034 7812
rect 6641 7803 6699 7809
rect 6641 7800 6653 7803
rect 4028 7772 6653 7800
rect 4028 7760 4034 7772
rect 6641 7769 6653 7772
rect 6687 7800 6699 7803
rect 7760 7800 7788 7899
rect 8846 7896 8852 7908
rect 8904 7896 8910 7948
rect 7837 7871 7895 7877
rect 7837 7837 7849 7871
rect 7883 7837 7895 7871
rect 7837 7831 7895 7837
rect 6687 7772 7788 7800
rect 6687 7769 6699 7772
rect 6641 7763 6699 7769
rect 4157 7735 4215 7741
rect 4157 7732 4169 7735
rect 3896 7704 4169 7732
rect 4157 7701 4169 7704
rect 4203 7732 4215 7735
rect 5074 7732 5080 7744
rect 4203 7704 5080 7732
rect 4203 7701 4215 7704
rect 4157 7695 4215 7701
rect 5074 7692 5080 7704
rect 5132 7692 5138 7744
rect 7101 7735 7159 7741
rect 7101 7701 7113 7735
rect 7147 7732 7159 7735
rect 7282 7732 7288 7744
rect 7147 7704 7288 7732
rect 7147 7701 7159 7704
rect 7101 7695 7159 7701
rect 7282 7692 7288 7704
rect 7340 7732 7346 7744
rect 7852 7732 7880 7831
rect 7926 7828 7932 7880
rect 7984 7868 7990 7880
rect 8021 7871 8079 7877
rect 8021 7868 8033 7871
rect 7984 7840 8033 7868
rect 7984 7828 7990 7840
rect 8021 7837 8033 7840
rect 8067 7868 8079 7871
rect 8956 7868 8984 7976
rect 14182 7964 14188 7976
rect 14240 8004 14246 8016
rect 14829 8007 14887 8013
rect 14829 8004 14841 8007
rect 14240 7976 14841 8004
rect 14240 7964 14246 7976
rect 14829 7973 14841 7976
rect 14875 7973 14887 8007
rect 14829 7967 14887 7973
rect 10502 7936 10508 7948
rect 10463 7908 10508 7936
rect 10502 7896 10508 7908
rect 10560 7896 10566 7948
rect 10772 7939 10830 7945
rect 10772 7905 10784 7939
rect 10818 7936 10830 7939
rect 11698 7936 11704 7948
rect 10818 7908 11704 7936
rect 10818 7905 10830 7908
rect 10772 7899 10830 7905
rect 11698 7896 11704 7908
rect 11756 7896 11762 7948
rect 11882 7896 11888 7948
rect 11940 7936 11946 7948
rect 12417 7939 12475 7945
rect 12417 7936 12429 7939
rect 11940 7908 12429 7936
rect 11940 7896 11946 7908
rect 12417 7905 12429 7908
rect 12463 7905 12475 7939
rect 12417 7899 12475 7905
rect 15289 7939 15347 7945
rect 15289 7905 15301 7939
rect 15335 7905 15347 7939
rect 15289 7899 15347 7905
rect 8067 7840 8984 7868
rect 8067 7837 8079 7840
rect 8021 7831 8079 7837
rect 9030 7828 9036 7880
rect 9088 7868 9094 7880
rect 9088 7840 9133 7868
rect 9088 7828 9094 7840
rect 11606 7828 11612 7880
rect 11664 7868 11670 7880
rect 12161 7871 12219 7877
rect 12161 7868 12173 7871
rect 11664 7840 12173 7868
rect 11664 7828 11670 7840
rect 12161 7837 12173 7840
rect 12207 7837 12219 7871
rect 12161 7831 12219 7837
rect 13630 7828 13636 7880
rect 13688 7868 13694 7880
rect 14277 7871 14335 7877
rect 14277 7868 14289 7871
rect 13688 7840 14289 7868
rect 13688 7828 13694 7840
rect 14277 7837 14289 7840
rect 14323 7837 14335 7871
rect 14458 7868 14464 7880
rect 14419 7840 14464 7868
rect 14277 7831 14335 7837
rect 14458 7828 14464 7840
rect 14516 7828 14522 7880
rect 15304 7800 15332 7899
rect 16482 7896 16488 7948
rect 16540 7936 16546 7948
rect 16577 7939 16635 7945
rect 16577 7936 16589 7939
rect 16540 7908 16589 7936
rect 16540 7896 16546 7908
rect 16577 7905 16589 7908
rect 16623 7905 16635 7939
rect 16577 7899 16635 7905
rect 15470 7868 15476 7880
rect 15431 7840 15476 7868
rect 15470 7828 15476 7840
rect 15528 7828 15534 7880
rect 16853 7871 16911 7877
rect 16853 7837 16865 7871
rect 16899 7868 16911 7871
rect 17494 7868 17500 7880
rect 16899 7840 17500 7868
rect 16899 7837 16911 7840
rect 16853 7831 16911 7837
rect 17494 7828 17500 7840
rect 17552 7828 17558 7880
rect 11716 7772 12020 7800
rect 7340 7704 7880 7732
rect 8481 7735 8539 7741
rect 7340 7692 7346 7704
rect 8481 7701 8493 7735
rect 8527 7732 8539 7735
rect 11716 7732 11744 7772
rect 11882 7732 11888 7744
rect 8527 7704 11744 7732
rect 11843 7704 11888 7732
rect 8527 7701 8539 7704
rect 8481 7695 8539 7701
rect 11882 7692 11888 7704
rect 11940 7692 11946 7744
rect 11992 7732 12020 7772
rect 13832 7772 15332 7800
rect 13832 7732 13860 7772
rect 11992 7704 13860 7732
rect 1104 7642 21896 7664
rect 1104 7590 4447 7642
rect 4499 7590 4511 7642
rect 4563 7590 4575 7642
rect 4627 7590 4639 7642
rect 4691 7590 11378 7642
rect 11430 7590 11442 7642
rect 11494 7590 11506 7642
rect 11558 7590 11570 7642
rect 11622 7590 18308 7642
rect 18360 7590 18372 7642
rect 18424 7590 18436 7642
rect 18488 7590 18500 7642
rect 18552 7590 21896 7642
rect 1104 7568 21896 7590
rect 2498 7488 2504 7540
rect 2556 7528 2562 7540
rect 3050 7528 3056 7540
rect 2556 7500 3056 7528
rect 2556 7488 2562 7500
rect 3050 7488 3056 7500
rect 3108 7528 3114 7540
rect 3145 7531 3203 7537
rect 3145 7528 3157 7531
rect 3108 7500 3157 7528
rect 3108 7488 3114 7500
rect 3145 7497 3157 7500
rect 3191 7497 3203 7531
rect 3145 7491 3203 7497
rect 3326 7488 3332 7540
rect 3384 7528 3390 7540
rect 4525 7531 4583 7537
rect 4525 7528 4537 7531
rect 3384 7500 4537 7528
rect 3384 7488 3390 7500
rect 4525 7497 4537 7500
rect 4571 7497 4583 7531
rect 4525 7491 4583 7497
rect 4890 7488 4896 7540
rect 4948 7528 4954 7540
rect 5258 7528 5264 7540
rect 4948 7500 5264 7528
rect 4948 7488 4954 7500
rect 5258 7488 5264 7500
rect 5316 7488 5322 7540
rect 5718 7528 5724 7540
rect 5679 7500 5724 7528
rect 5718 7488 5724 7500
rect 5776 7488 5782 7540
rect 9030 7528 9036 7540
rect 8991 7500 9036 7528
rect 9030 7488 9036 7500
rect 9088 7488 9094 7540
rect 14458 7488 14464 7540
rect 14516 7528 14522 7540
rect 17497 7531 17555 7537
rect 17497 7528 17509 7531
rect 14516 7500 17509 7528
rect 14516 7488 14522 7500
rect 17497 7497 17509 7500
rect 17543 7497 17555 7531
rect 17497 7491 17555 7497
rect 4062 7420 4068 7472
rect 4120 7460 4126 7472
rect 4120 7432 7604 7460
rect 4120 7420 4126 7432
rect 3234 7352 3240 7404
rect 3292 7392 3298 7404
rect 3789 7395 3847 7401
rect 3789 7392 3801 7395
rect 3292 7364 3801 7392
rect 3292 7352 3298 7364
rect 3789 7361 3801 7364
rect 3835 7361 3847 7395
rect 3789 7355 3847 7361
rect 6086 7352 6092 7404
rect 6144 7392 6150 7404
rect 6273 7395 6331 7401
rect 6273 7392 6285 7395
rect 6144 7364 6285 7392
rect 6144 7352 6150 7364
rect 6273 7361 6285 7364
rect 6319 7361 6331 7395
rect 6273 7355 6331 7361
rect 1765 7327 1823 7333
rect 1765 7293 1777 7327
rect 1811 7324 1823 7327
rect 1854 7324 1860 7336
rect 1811 7296 1860 7324
rect 1811 7293 1823 7296
rect 1765 7287 1823 7293
rect 1854 7284 1860 7296
rect 1912 7324 1918 7336
rect 4890 7324 4896 7336
rect 1912 7296 4896 7324
rect 1912 7284 1918 7296
rect 4890 7284 4896 7296
rect 4948 7284 4954 7336
rect 5445 7327 5503 7333
rect 5445 7293 5457 7327
rect 5491 7324 5503 7327
rect 7190 7324 7196 7336
rect 5491 7296 7196 7324
rect 5491 7293 5503 7296
rect 5445 7287 5503 7293
rect 7190 7284 7196 7296
rect 7248 7284 7254 7336
rect 2032 7259 2090 7265
rect 2032 7225 2044 7259
rect 2078 7256 2090 7259
rect 2406 7256 2412 7268
rect 2078 7228 2412 7256
rect 2078 7225 2090 7228
rect 2032 7219 2090 7225
rect 2406 7216 2412 7228
rect 2464 7216 2470 7268
rect 3694 7216 3700 7268
rect 3752 7256 3758 7268
rect 4985 7259 5043 7265
rect 4985 7256 4997 7259
rect 3752 7228 4997 7256
rect 3752 7216 3758 7228
rect 4985 7225 4997 7228
rect 5031 7256 5043 7259
rect 5902 7256 5908 7268
rect 5031 7228 5908 7256
rect 5031 7225 5043 7228
rect 4985 7219 5043 7225
rect 5902 7216 5908 7228
rect 5960 7216 5966 7268
rect 6181 7259 6239 7265
rect 6181 7256 6193 7259
rect 6012 7228 6193 7256
rect 2958 7148 2964 7200
rect 3016 7188 3022 7200
rect 3326 7188 3332 7200
rect 3016 7160 3332 7188
rect 3016 7148 3022 7160
rect 3326 7148 3332 7160
rect 3384 7188 3390 7200
rect 3421 7191 3479 7197
rect 3421 7188 3433 7191
rect 3384 7160 3433 7188
rect 3384 7148 3390 7160
rect 3421 7157 3433 7160
rect 3467 7157 3479 7191
rect 3421 7151 3479 7157
rect 5534 7148 5540 7200
rect 5592 7188 5598 7200
rect 6012 7188 6040 7228
rect 6181 7225 6193 7228
rect 6227 7225 6239 7259
rect 6181 7219 6239 7225
rect 5592 7160 6040 7188
rect 5592 7148 5598 7160
rect 6086 7148 6092 7200
rect 6144 7188 6150 7200
rect 7006 7188 7012 7200
rect 6144 7160 6189 7188
rect 6967 7160 7012 7188
rect 6144 7148 6150 7160
rect 7006 7148 7012 7160
rect 7064 7148 7070 7200
rect 7576 7188 7604 7432
rect 9048 7392 9076 7488
rect 11606 7392 11612 7404
rect 9048 7364 9444 7392
rect 11567 7364 11612 7392
rect 7926 7333 7932 7336
rect 7653 7327 7711 7333
rect 7653 7293 7665 7327
rect 7699 7293 7711 7327
rect 7920 7324 7932 7333
rect 7887 7296 7932 7324
rect 7653 7287 7711 7293
rect 7920 7287 7932 7296
rect 7668 7256 7696 7287
rect 7926 7284 7932 7287
rect 7984 7284 7990 7336
rect 9306 7324 9312 7336
rect 9267 7296 9312 7324
rect 9306 7284 9312 7296
rect 9364 7284 9370 7336
rect 9416 7324 9444 7364
rect 11606 7352 11612 7364
rect 11664 7352 11670 7404
rect 9565 7327 9623 7333
rect 9565 7324 9577 7327
rect 9416 7296 9577 7324
rect 9565 7293 9577 7296
rect 9611 7293 9623 7327
rect 11977 7327 12035 7333
rect 11977 7324 11989 7327
rect 9565 7287 9623 7293
rect 11440 7296 11989 7324
rect 9324 7256 9352 7284
rect 7668 7228 9352 7256
rect 10778 7216 10784 7268
rect 10836 7256 10842 7268
rect 11440 7265 11468 7296
rect 11977 7293 11989 7296
rect 12023 7293 12035 7327
rect 14090 7324 14096 7336
rect 14051 7296 14096 7324
rect 11977 7287 12035 7293
rect 14090 7284 14096 7296
rect 14148 7284 14154 7336
rect 16022 7284 16028 7336
rect 16080 7324 16086 7336
rect 16117 7327 16175 7333
rect 16117 7324 16129 7327
rect 16080 7296 16129 7324
rect 16080 7284 16086 7296
rect 16117 7293 16129 7296
rect 16163 7293 16175 7327
rect 16117 7287 16175 7293
rect 11425 7259 11483 7265
rect 11425 7256 11437 7259
rect 10836 7228 11437 7256
rect 10836 7216 10842 7228
rect 11425 7225 11437 7228
rect 11471 7225 11483 7259
rect 11425 7219 11483 7225
rect 11606 7216 11612 7268
rect 11664 7256 11670 7268
rect 14360 7259 14418 7265
rect 11664 7228 13759 7256
rect 11664 7216 11670 7228
rect 9950 7188 9956 7200
rect 7576 7160 9956 7188
rect 9950 7148 9956 7160
rect 10008 7148 10014 7200
rect 10686 7188 10692 7200
rect 10647 7160 10692 7188
rect 10686 7148 10692 7160
rect 10744 7148 10750 7200
rect 10965 7191 11023 7197
rect 10965 7157 10977 7191
rect 11011 7188 11023 7191
rect 11238 7188 11244 7200
rect 11011 7160 11244 7188
rect 11011 7157 11023 7160
rect 10965 7151 11023 7157
rect 11238 7148 11244 7160
rect 11296 7148 11302 7200
rect 11330 7148 11336 7200
rect 11388 7188 11394 7200
rect 11388 7160 11433 7188
rect 11388 7148 11394 7160
rect 12434 7148 12440 7200
rect 12492 7188 12498 7200
rect 12986 7188 12992 7200
rect 12492 7160 12537 7188
rect 12947 7160 12992 7188
rect 12492 7148 12498 7160
rect 12986 7148 12992 7160
rect 13044 7188 13050 7200
rect 13630 7188 13636 7200
rect 13044 7160 13636 7188
rect 13044 7148 13050 7160
rect 13630 7148 13636 7160
rect 13688 7148 13694 7200
rect 13731 7188 13759 7228
rect 14360 7225 14372 7259
rect 14406 7256 14418 7259
rect 14734 7256 14740 7268
rect 14406 7228 14740 7256
rect 14406 7225 14418 7228
rect 14360 7219 14418 7225
rect 14734 7216 14740 7228
rect 14792 7216 14798 7268
rect 16384 7259 16442 7265
rect 16384 7225 16396 7259
rect 16430 7256 16442 7259
rect 17402 7256 17408 7268
rect 16430 7228 17408 7256
rect 16430 7225 16442 7228
rect 16384 7219 16442 7225
rect 17402 7216 17408 7228
rect 17460 7216 17466 7268
rect 15473 7191 15531 7197
rect 15473 7188 15485 7191
rect 13731 7160 15485 7188
rect 15473 7157 15485 7160
rect 15519 7157 15531 7191
rect 15473 7151 15531 7157
rect 1104 7098 21896 7120
rect 1104 7046 7912 7098
rect 7964 7046 7976 7098
rect 8028 7046 8040 7098
rect 8092 7046 8104 7098
rect 8156 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 15035 7098
rect 15087 7046 21896 7098
rect 1104 7024 21896 7046
rect 5534 6944 5540 6996
rect 5592 6984 5598 6996
rect 5721 6987 5779 6993
rect 5721 6984 5733 6987
rect 5592 6956 5733 6984
rect 5592 6944 5598 6956
rect 5721 6953 5733 6956
rect 5767 6953 5779 6987
rect 8846 6984 8852 6996
rect 8807 6956 8852 6984
rect 5721 6947 5779 6953
rect 8846 6944 8852 6956
rect 8904 6944 8910 6996
rect 11517 6987 11575 6993
rect 11517 6953 11529 6987
rect 11563 6984 11575 6987
rect 12434 6984 12440 6996
rect 11563 6956 12440 6984
rect 11563 6953 11575 6956
rect 11517 6947 11575 6953
rect 12434 6944 12440 6956
rect 12492 6944 12498 6996
rect 13630 6984 13636 6996
rect 13591 6956 13636 6984
rect 13630 6944 13636 6956
rect 13688 6944 13694 6996
rect 2317 6919 2375 6925
rect 2317 6885 2329 6919
rect 2363 6916 2375 6919
rect 3050 6916 3056 6928
rect 2363 6888 3056 6916
rect 2363 6885 2375 6888
rect 2317 6879 2375 6885
rect 3050 6876 3056 6888
rect 3108 6876 3114 6928
rect 3234 6876 3240 6928
rect 3292 6916 3298 6928
rect 3329 6919 3387 6925
rect 3329 6916 3341 6919
rect 3292 6888 3341 6916
rect 3292 6876 3298 6888
rect 3329 6885 3341 6888
rect 3375 6885 3387 6919
rect 3329 6879 3387 6885
rect 3602 6876 3608 6928
rect 3660 6916 3666 6928
rect 3660 6888 4467 6916
rect 3660 6876 3666 6888
rect 2866 6808 2872 6860
rect 2924 6848 2930 6860
rect 3418 6848 3424 6860
rect 2924 6820 3424 6848
rect 2924 6808 2930 6820
rect 3418 6808 3424 6820
rect 3476 6808 3482 6860
rect 4338 6857 4344 6860
rect 4332 6848 4344 6857
rect 3620 6820 4344 6848
rect 3620 6789 3648 6820
rect 4332 6811 4344 6820
rect 4338 6808 4344 6811
rect 4396 6808 4402 6860
rect 4439 6848 4467 6888
rect 4614 6876 4620 6928
rect 4672 6916 4678 6928
rect 10413 6919 10471 6925
rect 10413 6916 10425 6919
rect 4672 6888 10425 6916
rect 4672 6876 4678 6888
rect 10413 6885 10425 6888
rect 10459 6916 10471 6919
rect 11330 6916 11336 6928
rect 10459 6888 11336 6916
rect 10459 6885 10471 6888
rect 10413 6879 10471 6885
rect 11330 6876 11336 6888
rect 11388 6876 11394 6928
rect 14553 6919 14611 6925
rect 14553 6885 14565 6919
rect 14599 6916 14611 6919
rect 15194 6916 15200 6928
rect 14599 6888 15200 6916
rect 14599 6885 14611 6888
rect 14553 6879 14611 6885
rect 15194 6876 15200 6888
rect 15252 6876 15258 6928
rect 6086 6848 6092 6860
rect 4439 6820 6092 6848
rect 6086 6808 6092 6820
rect 6144 6808 6150 6860
rect 10873 6851 10931 6857
rect 10873 6817 10885 6851
rect 10919 6817 10931 6851
rect 10873 6811 10931 6817
rect 2409 6783 2467 6789
rect 2409 6749 2421 6783
rect 2455 6780 2467 6783
rect 2593 6783 2651 6789
rect 2455 6752 2544 6780
rect 2455 6749 2467 6752
rect 2409 6743 2467 6749
rect 1673 6715 1731 6721
rect 1673 6681 1685 6715
rect 1719 6712 1731 6715
rect 2516 6712 2544 6752
rect 2593 6749 2605 6783
rect 2639 6780 2651 6783
rect 3605 6783 3663 6789
rect 2639 6752 3096 6780
rect 2639 6749 2651 6752
rect 2593 6743 2651 6749
rect 2961 6715 3019 6721
rect 2961 6712 2973 6715
rect 1719 6684 2452 6712
rect 2516 6684 2973 6712
rect 1719 6681 1731 6684
rect 1673 6675 1731 6681
rect 1949 6647 2007 6653
rect 1949 6613 1961 6647
rect 1995 6644 2007 6647
rect 2314 6644 2320 6656
rect 1995 6616 2320 6644
rect 1995 6613 2007 6616
rect 1949 6607 2007 6613
rect 2314 6604 2320 6616
rect 2372 6604 2378 6656
rect 2424 6644 2452 6684
rect 2961 6681 2973 6684
rect 3007 6681 3019 6715
rect 2961 6675 3019 6681
rect 2866 6644 2872 6656
rect 2424 6616 2872 6644
rect 2866 6604 2872 6616
rect 2924 6604 2930 6656
rect 3068 6644 3096 6752
rect 3605 6749 3617 6783
rect 3651 6749 3663 6783
rect 3605 6743 3663 6749
rect 3786 6740 3792 6792
rect 3844 6780 3850 6792
rect 4065 6783 4123 6789
rect 4065 6780 4077 6783
rect 3844 6752 4077 6780
rect 3844 6740 3850 6752
rect 4065 6749 4077 6752
rect 4111 6749 4123 6783
rect 4065 6743 4123 6749
rect 3602 6644 3608 6656
rect 3068 6616 3608 6644
rect 3602 6604 3608 6616
rect 3660 6644 3666 6656
rect 5445 6647 5503 6653
rect 5445 6644 5457 6647
rect 3660 6616 5457 6644
rect 3660 6604 3666 6616
rect 5445 6613 5457 6616
rect 5491 6613 5503 6647
rect 8478 6644 8484 6656
rect 8439 6616 8484 6644
rect 5445 6607 5503 6613
rect 8478 6604 8484 6616
rect 8536 6604 8542 6656
rect 9306 6604 9312 6656
rect 9364 6644 9370 6656
rect 10502 6644 10508 6656
rect 9364 6616 10508 6644
rect 9364 6604 9370 6616
rect 10502 6604 10508 6616
rect 10560 6644 10566 6656
rect 10689 6647 10747 6653
rect 10689 6644 10701 6647
rect 10560 6616 10701 6644
rect 10560 6604 10566 6616
rect 10689 6613 10701 6616
rect 10735 6613 10747 6647
rect 10888 6644 10916 6811
rect 11238 6808 11244 6860
rect 11296 6848 11302 6860
rect 11609 6851 11667 6857
rect 11609 6848 11621 6851
rect 11296 6820 11621 6848
rect 11296 6808 11302 6820
rect 11609 6817 11621 6820
rect 11655 6817 11667 6851
rect 11609 6811 11667 6817
rect 12158 6808 12164 6860
rect 12216 6848 12222 6860
rect 12713 6851 12771 6857
rect 12713 6848 12725 6851
rect 12216 6820 12725 6848
rect 12216 6808 12222 6820
rect 12713 6817 12725 6820
rect 12759 6817 12771 6851
rect 12713 6811 12771 6817
rect 13541 6851 13599 6857
rect 13541 6817 13553 6851
rect 13587 6817 13599 6851
rect 15289 6851 15347 6857
rect 15289 6848 15301 6851
rect 13541 6811 13599 6817
rect 14936 6820 15301 6848
rect 11793 6783 11851 6789
rect 11793 6749 11805 6783
rect 11839 6780 11851 6783
rect 11882 6780 11888 6792
rect 11839 6752 11888 6780
rect 11839 6749 11851 6752
rect 11793 6743 11851 6749
rect 11882 6740 11888 6752
rect 11940 6740 11946 6792
rect 12253 6783 12311 6789
rect 12253 6749 12265 6783
rect 12299 6780 12311 6783
rect 12434 6780 12440 6792
rect 12299 6752 12440 6780
rect 12299 6749 12311 6752
rect 12253 6743 12311 6749
rect 12434 6740 12440 6752
rect 12492 6780 12498 6792
rect 13556 6780 13584 6811
rect 13814 6780 13820 6792
rect 12492 6752 13584 6780
rect 13775 6752 13820 6780
rect 12492 6740 12498 6752
rect 13814 6740 13820 6752
rect 13872 6740 13878 6792
rect 14645 6783 14703 6789
rect 14645 6780 14657 6783
rect 13924 6752 14657 6780
rect 11149 6715 11207 6721
rect 11149 6681 11161 6715
rect 11195 6712 11207 6715
rect 13173 6715 13231 6721
rect 11195 6684 13124 6712
rect 11195 6681 11207 6684
rect 11149 6675 11207 6681
rect 12526 6644 12532 6656
rect 10888 6616 12532 6644
rect 10689 6607 10747 6613
rect 12526 6604 12532 6616
rect 12584 6604 12590 6656
rect 13096 6644 13124 6684
rect 13173 6681 13185 6715
rect 13219 6712 13231 6715
rect 13924 6712 13952 6752
rect 14645 6749 14657 6752
rect 14691 6749 14703 6783
rect 14826 6780 14832 6792
rect 14787 6752 14832 6780
rect 14645 6743 14703 6749
rect 14826 6740 14832 6752
rect 14884 6740 14890 6792
rect 14936 6712 14964 6820
rect 15289 6817 15301 6820
rect 15335 6817 15347 6851
rect 15289 6811 15347 6817
rect 16669 6851 16727 6857
rect 16669 6817 16681 6851
rect 16715 6848 16727 6851
rect 17313 6851 17371 6857
rect 17313 6848 17325 6851
rect 16715 6820 17325 6848
rect 16715 6817 16727 6820
rect 16669 6811 16727 6817
rect 17313 6817 17325 6820
rect 17359 6817 17371 6851
rect 17313 6811 17371 6817
rect 15473 6783 15531 6789
rect 15473 6780 15485 6783
rect 15304 6752 15485 6780
rect 15304 6724 15332 6752
rect 15473 6749 15485 6752
rect 15519 6749 15531 6783
rect 15473 6743 15531 6749
rect 16482 6740 16488 6792
rect 16540 6780 16546 6792
rect 16761 6783 16819 6789
rect 16761 6780 16773 6783
rect 16540 6752 16773 6780
rect 16540 6740 16546 6752
rect 16761 6749 16773 6752
rect 16807 6749 16819 6783
rect 16761 6743 16819 6749
rect 16945 6783 17003 6789
rect 16945 6749 16957 6783
rect 16991 6780 17003 6783
rect 17218 6780 17224 6792
rect 16991 6752 17224 6780
rect 16991 6749 17003 6752
rect 16945 6743 17003 6749
rect 13219 6684 13952 6712
rect 14108 6684 14964 6712
rect 13219 6681 13231 6684
rect 13173 6675 13231 6681
rect 14108 6644 14136 6684
rect 15286 6672 15292 6724
rect 15344 6672 15350 6724
rect 16776 6712 16804 6743
rect 17218 6740 17224 6752
rect 17276 6740 17282 6792
rect 17773 6715 17831 6721
rect 17773 6712 17785 6715
rect 16776 6684 17785 6712
rect 17773 6681 17785 6684
rect 17819 6681 17831 6715
rect 17773 6675 17831 6681
rect 13096 6616 14136 6644
rect 14185 6647 14243 6653
rect 14185 6613 14197 6647
rect 14231 6644 14243 6647
rect 14274 6644 14280 6656
rect 14231 6616 14280 6644
rect 14231 6613 14243 6616
rect 14185 6607 14243 6613
rect 14274 6604 14280 6616
rect 14332 6604 14338 6656
rect 16301 6647 16359 6653
rect 16301 6613 16313 6647
rect 16347 6644 16359 6647
rect 17678 6644 17684 6656
rect 16347 6616 17684 6644
rect 16347 6613 16359 6616
rect 16301 6607 16359 6613
rect 17678 6604 17684 6616
rect 17736 6604 17742 6656
rect 1104 6554 21896 6576
rect 1104 6502 4447 6554
rect 4499 6502 4511 6554
rect 4563 6502 4575 6554
rect 4627 6502 4639 6554
rect 4691 6502 11378 6554
rect 11430 6502 11442 6554
rect 11494 6502 11506 6554
rect 11558 6502 11570 6554
rect 11622 6502 18308 6554
rect 18360 6502 18372 6554
rect 18424 6502 18436 6554
rect 18488 6502 18500 6554
rect 18552 6502 21896 6554
rect 1104 6480 21896 6502
rect 2406 6400 2412 6452
rect 2464 6440 2470 6452
rect 2777 6443 2835 6449
rect 2777 6440 2789 6443
rect 2464 6412 2789 6440
rect 2464 6400 2470 6412
rect 2777 6409 2789 6412
rect 2823 6409 2835 6443
rect 2777 6403 2835 6409
rect 4062 6400 4068 6452
rect 4120 6440 4126 6452
rect 12434 6440 12440 6452
rect 4120 6412 12440 6440
rect 4120 6400 4126 6412
rect 12434 6400 12440 6412
rect 12492 6400 12498 6452
rect 13814 6440 13820 6452
rect 13775 6412 13820 6440
rect 13814 6400 13820 6412
rect 13872 6400 13878 6452
rect 14826 6400 14832 6452
rect 14884 6440 14890 6452
rect 15473 6443 15531 6449
rect 15473 6440 15485 6443
rect 14884 6412 15485 6440
rect 14884 6400 14890 6412
rect 15473 6409 15485 6412
rect 15519 6409 15531 6443
rect 17402 6440 17408 6452
rect 17363 6412 17408 6440
rect 15473 6403 15531 6409
rect 17402 6400 17408 6412
rect 17460 6400 17466 6452
rect 9950 6372 9956 6384
rect 9911 6344 9956 6372
rect 9950 6332 9956 6344
rect 10008 6332 10014 6384
rect 11885 6375 11943 6381
rect 11885 6341 11897 6375
rect 11931 6341 11943 6375
rect 11885 6335 11943 6341
rect 3050 6304 3056 6316
rect 3011 6276 3056 6304
rect 3050 6264 3056 6276
rect 3108 6264 3114 6316
rect 4249 6307 4307 6313
rect 4249 6273 4261 6307
rect 4295 6304 4307 6307
rect 4338 6304 4344 6316
rect 4295 6276 4344 6304
rect 4295 6273 4307 6276
rect 4249 6267 4307 6273
rect 4338 6264 4344 6276
rect 4396 6304 4402 6316
rect 4433 6307 4491 6313
rect 4433 6304 4445 6307
rect 4396 6276 4445 6304
rect 4396 6264 4402 6276
rect 4433 6273 4445 6276
rect 4479 6273 4491 6307
rect 7466 6304 7472 6316
rect 7427 6276 7472 6304
rect 4433 6267 4491 6273
rect 7466 6264 7472 6276
rect 7524 6264 7530 6316
rect 11900 6304 11928 6335
rect 13832 6304 13860 6400
rect 17420 6304 17448 6400
rect 18601 6307 18659 6313
rect 18601 6304 18613 6307
rect 11900 6276 12572 6304
rect 13832 6276 14228 6304
rect 17420 6276 18613 6304
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6205 1455 6239
rect 1397 6199 1455 6205
rect 1664 6239 1722 6245
rect 1664 6205 1676 6239
rect 1710 6236 1722 6239
rect 3602 6236 3608 6248
rect 1710 6208 3608 6236
rect 1710 6205 1722 6208
rect 1664 6199 1722 6205
rect 1412 6168 1440 6199
rect 3602 6196 3608 6208
rect 3660 6196 3666 6248
rect 4617 6239 4675 6245
rect 4617 6205 4629 6239
rect 4663 6236 4675 6239
rect 4706 6236 4712 6248
rect 4663 6208 4712 6236
rect 4663 6205 4675 6208
rect 4617 6199 4675 6205
rect 4706 6196 4712 6208
rect 4764 6196 4770 6248
rect 6365 6239 6423 6245
rect 6365 6236 6377 6239
rect 4816 6208 6377 6236
rect 2682 6168 2688 6180
rect 1412 6140 2688 6168
rect 2682 6128 2688 6140
rect 2740 6168 2746 6180
rect 3786 6168 3792 6180
rect 2740 6140 3792 6168
rect 2740 6128 2746 6140
rect 3786 6128 3792 6140
rect 3844 6128 3850 6180
rect 3878 6128 3884 6180
rect 3936 6168 3942 6180
rect 4816 6168 4844 6208
rect 6365 6205 6377 6208
rect 6411 6236 6423 6239
rect 7285 6239 7343 6245
rect 7285 6236 7297 6239
rect 6411 6208 7297 6236
rect 6411 6205 6423 6208
rect 6365 6199 6423 6205
rect 7285 6205 7297 6208
rect 7331 6205 7343 6239
rect 7285 6199 7343 6205
rect 8297 6239 8355 6245
rect 8297 6205 8309 6239
rect 8343 6236 8355 6239
rect 9306 6236 9312 6248
rect 8343 6208 9312 6236
rect 8343 6205 8355 6208
rect 8297 6199 8355 6205
rect 9306 6196 9312 6208
rect 9364 6196 9370 6248
rect 10502 6236 10508 6248
rect 10415 6208 10508 6236
rect 10502 6196 10508 6208
rect 10560 6236 10566 6248
rect 12342 6236 12348 6248
rect 10560 6208 12348 6236
rect 10560 6196 10566 6208
rect 12342 6196 12348 6208
rect 12400 6236 12406 6248
rect 12437 6239 12495 6245
rect 12437 6236 12449 6239
rect 12400 6208 12449 6236
rect 12400 6196 12406 6208
rect 12437 6205 12449 6208
rect 12483 6205 12495 6239
rect 12544 6236 12572 6276
rect 12693 6239 12751 6245
rect 12693 6236 12705 6239
rect 12544 6208 12705 6236
rect 12437 6199 12495 6205
rect 12693 6205 12705 6208
rect 12739 6236 12751 6239
rect 13078 6236 13084 6248
rect 12739 6208 13084 6236
rect 12739 6205 12751 6208
rect 12693 6199 12751 6205
rect 13078 6196 13084 6208
rect 13136 6196 13142 6248
rect 14090 6236 14096 6248
rect 14003 6208 14096 6236
rect 14090 6196 14096 6208
rect 14148 6196 14154 6248
rect 14200 6236 14228 6276
rect 18601 6273 18613 6276
rect 18647 6273 18659 6307
rect 18601 6267 18659 6273
rect 14349 6239 14407 6245
rect 14349 6236 14361 6239
rect 14200 6208 14361 6236
rect 14349 6205 14361 6208
rect 14395 6205 14407 6239
rect 16022 6236 16028 6248
rect 15983 6208 16028 6236
rect 14349 6199 14407 6205
rect 16022 6196 16028 6208
rect 16080 6196 16086 6248
rect 17678 6196 17684 6248
rect 17736 6236 17742 6248
rect 18417 6239 18475 6245
rect 18417 6236 18429 6239
rect 17736 6208 18429 6236
rect 17736 6196 17742 6208
rect 18417 6205 18429 6208
rect 18463 6205 18475 6239
rect 18417 6199 18475 6205
rect 3936 6140 4844 6168
rect 4884 6171 4942 6177
rect 3936 6128 3942 6140
rect 4884 6137 4896 6171
rect 4930 6168 4942 6171
rect 5442 6168 5448 6180
rect 4930 6140 5448 6168
rect 4930 6137 4942 6140
rect 4884 6131 4942 6137
rect 5442 6128 5448 6140
rect 5500 6128 5506 6180
rect 7193 6171 7251 6177
rect 7193 6137 7205 6171
rect 7239 6168 7251 6171
rect 7837 6171 7895 6177
rect 7837 6168 7849 6171
rect 7239 6140 7849 6168
rect 7239 6137 7251 6140
rect 7193 6131 7251 6137
rect 7837 6137 7849 6140
rect 7883 6137 7895 6171
rect 7837 6131 7895 6137
rect 8202 6128 8208 6180
rect 8260 6168 8266 6180
rect 8542 6171 8600 6177
rect 8542 6168 8554 6171
rect 8260 6140 8554 6168
rect 8260 6128 8266 6140
rect 8542 6137 8554 6140
rect 8588 6137 8600 6171
rect 10750 6171 10808 6177
rect 10750 6168 10762 6171
rect 8542 6131 8600 6137
rect 9692 6140 10762 6168
rect 2866 6060 2872 6112
rect 2924 6100 2930 6112
rect 3050 6100 3056 6112
rect 2924 6072 3056 6100
rect 2924 6060 2930 6072
rect 3050 6060 3056 6072
rect 3108 6060 3114 6112
rect 3418 6060 3424 6112
rect 3476 6100 3482 6112
rect 3605 6103 3663 6109
rect 3605 6100 3617 6103
rect 3476 6072 3617 6100
rect 3476 6060 3482 6072
rect 3605 6069 3617 6072
rect 3651 6069 3663 6103
rect 3970 6100 3976 6112
rect 3931 6072 3976 6100
rect 3605 6063 3663 6069
rect 3970 6060 3976 6072
rect 4028 6060 4034 6112
rect 4065 6103 4123 6109
rect 4065 6069 4077 6103
rect 4111 6100 4123 6103
rect 4246 6100 4252 6112
rect 4111 6072 4252 6100
rect 4111 6069 4123 6072
rect 4065 6063 4123 6069
rect 4246 6060 4252 6072
rect 4304 6060 4310 6112
rect 4433 6103 4491 6109
rect 4433 6069 4445 6103
rect 4479 6100 4491 6103
rect 4706 6100 4712 6112
rect 4479 6072 4712 6100
rect 4479 6069 4491 6072
rect 4433 6063 4491 6069
rect 4706 6060 4712 6072
rect 4764 6100 4770 6112
rect 5997 6103 6055 6109
rect 5997 6100 6009 6103
rect 4764 6072 6009 6100
rect 4764 6060 4770 6072
rect 5997 6069 6009 6072
rect 6043 6069 6055 6103
rect 6822 6100 6828 6112
rect 6783 6072 6828 6100
rect 5997 6063 6055 6069
rect 6822 6060 6828 6072
rect 6880 6060 6886 6112
rect 9692 6109 9720 6140
rect 10750 6137 10762 6140
rect 10796 6168 10808 6171
rect 11790 6168 11796 6180
rect 10796 6140 11796 6168
rect 10796 6137 10808 6140
rect 10750 6131 10808 6137
rect 11790 6128 11796 6140
rect 11848 6128 11854 6180
rect 14108 6168 14136 6196
rect 16040 6168 16068 6196
rect 14108 6140 16068 6168
rect 16292 6171 16350 6177
rect 16292 6137 16304 6171
rect 16338 6168 16350 6171
rect 17218 6168 17224 6180
rect 16338 6140 17224 6168
rect 16338 6137 16350 6140
rect 16292 6131 16350 6137
rect 17218 6128 17224 6140
rect 17276 6128 17282 6180
rect 9677 6103 9735 6109
rect 9677 6069 9689 6103
rect 9723 6069 9735 6103
rect 9677 6063 9735 6069
rect 16942 6060 16948 6112
rect 17000 6100 17006 6112
rect 18049 6103 18107 6109
rect 18049 6100 18061 6103
rect 17000 6072 18061 6100
rect 17000 6060 17006 6072
rect 18049 6069 18061 6072
rect 18095 6069 18107 6103
rect 18049 6063 18107 6069
rect 18138 6060 18144 6112
rect 18196 6100 18202 6112
rect 18509 6103 18567 6109
rect 18509 6100 18521 6103
rect 18196 6072 18521 6100
rect 18196 6060 18202 6072
rect 18509 6069 18521 6072
rect 18555 6069 18567 6103
rect 18509 6063 18567 6069
rect 1104 6010 21896 6032
rect 1104 5958 7912 6010
rect 7964 5958 7976 6010
rect 8028 5958 8040 6010
rect 8092 5958 8104 6010
rect 8156 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 15035 6010
rect 15087 5958 21896 6010
rect 1104 5936 21896 5958
rect 1946 5896 1952 5908
rect 1907 5868 1952 5896
rect 1946 5856 1952 5868
rect 2004 5856 2010 5908
rect 2314 5896 2320 5908
rect 2275 5868 2320 5896
rect 2314 5856 2320 5868
rect 2372 5856 2378 5908
rect 2409 5899 2467 5905
rect 2409 5865 2421 5899
rect 2455 5896 2467 5899
rect 2961 5899 3019 5905
rect 2961 5896 2973 5899
rect 2455 5868 2973 5896
rect 2455 5865 2467 5868
rect 2409 5859 2467 5865
rect 2961 5865 2973 5868
rect 3007 5865 3019 5899
rect 3418 5896 3424 5908
rect 3379 5868 3424 5896
rect 2961 5859 3019 5865
rect 3418 5856 3424 5868
rect 3476 5856 3482 5908
rect 3510 5856 3516 5908
rect 3568 5896 3574 5908
rect 11333 5899 11391 5905
rect 3568 5868 10824 5896
rect 3568 5856 3574 5868
rect 3329 5831 3387 5837
rect 3329 5797 3341 5831
rect 3375 5828 3387 5831
rect 3881 5831 3939 5837
rect 3881 5828 3893 5831
rect 3375 5800 3893 5828
rect 3375 5797 3387 5800
rect 3329 5791 3387 5797
rect 3881 5797 3893 5800
rect 3927 5797 3939 5831
rect 6264 5831 6322 5837
rect 3881 5791 3939 5797
rect 4356 5800 6040 5828
rect 3786 5720 3792 5772
rect 3844 5760 3850 5772
rect 4356 5760 4384 5800
rect 3844 5732 4384 5760
rect 4433 5763 4491 5769
rect 3844 5720 3850 5732
rect 4433 5729 4445 5763
rect 4479 5760 4491 5763
rect 4890 5760 4896 5772
rect 4479 5732 4896 5760
rect 4479 5729 4491 5732
rect 4433 5723 4491 5729
rect 4890 5720 4896 5732
rect 4948 5720 4954 5772
rect 6012 5769 6040 5800
rect 6264 5797 6276 5831
rect 6310 5828 6322 5831
rect 7558 5828 7564 5840
rect 6310 5800 7564 5828
rect 6310 5797 6322 5800
rect 6264 5791 6322 5797
rect 7558 5788 7564 5800
rect 7616 5788 7622 5840
rect 9950 5837 9956 5840
rect 9944 5828 9956 5837
rect 9863 5800 9956 5828
rect 9944 5791 9956 5800
rect 10008 5828 10014 5840
rect 10686 5828 10692 5840
rect 10008 5800 10692 5828
rect 9950 5788 9956 5791
rect 10008 5788 10014 5800
rect 10686 5788 10692 5800
rect 10744 5788 10750 5840
rect 10796 5828 10824 5868
rect 11333 5865 11345 5899
rect 11379 5896 11391 5899
rect 12805 5899 12863 5905
rect 12805 5896 12817 5899
rect 11379 5868 12817 5896
rect 11379 5865 11391 5868
rect 11333 5859 11391 5865
rect 12805 5865 12817 5868
rect 12851 5865 12863 5899
rect 12805 5859 12863 5865
rect 15194 5856 15200 5908
rect 15252 5896 15258 5908
rect 15289 5899 15347 5905
rect 15289 5896 15301 5899
rect 15252 5868 15301 5896
rect 15252 5856 15258 5868
rect 15289 5865 15301 5868
rect 15335 5865 15347 5899
rect 15289 5859 15347 5865
rect 11701 5831 11759 5837
rect 11701 5828 11713 5831
rect 10796 5800 11713 5828
rect 11701 5797 11713 5800
rect 11747 5797 11759 5831
rect 11701 5791 11759 5797
rect 11793 5831 11851 5837
rect 11793 5797 11805 5831
rect 11839 5828 11851 5831
rect 12158 5828 12164 5840
rect 11839 5800 12164 5828
rect 11839 5797 11851 5800
rect 11793 5791 11851 5797
rect 5997 5763 6055 5769
rect 5997 5729 6009 5763
rect 6043 5760 6055 5763
rect 7006 5760 7012 5772
rect 6043 5732 7012 5760
rect 6043 5729 6055 5732
rect 5997 5723 6055 5729
rect 7006 5720 7012 5732
rect 7064 5720 7070 5772
rect 7466 5760 7472 5772
rect 7379 5732 7472 5760
rect 7466 5720 7472 5732
rect 7524 5760 7530 5772
rect 7920 5763 7978 5769
rect 7920 5760 7932 5763
rect 7524 5732 7932 5760
rect 7524 5720 7530 5732
rect 7920 5729 7932 5732
rect 7966 5760 7978 5763
rect 8662 5760 8668 5772
rect 7966 5732 8668 5760
rect 7966 5729 7978 5732
rect 7920 5723 7978 5729
rect 8662 5720 8668 5732
rect 8720 5720 8726 5772
rect 9677 5763 9735 5769
rect 9677 5729 9689 5763
rect 9723 5760 9735 5763
rect 10502 5760 10508 5772
rect 9723 5732 10508 5760
rect 9723 5729 9735 5732
rect 9677 5723 9735 5729
rect 10502 5720 10508 5732
rect 10560 5720 10566 5772
rect 11716 5760 11744 5791
rect 12158 5788 12164 5800
rect 12216 5788 12222 5840
rect 12526 5788 12532 5840
rect 12584 5828 12590 5840
rect 12584 5800 15976 5828
rect 12584 5788 12590 5800
rect 11974 5760 11980 5772
rect 11716 5732 11980 5760
rect 11974 5720 11980 5732
rect 12032 5720 12038 5772
rect 12710 5760 12716 5772
rect 12671 5732 12716 5760
rect 12710 5720 12716 5732
rect 12768 5720 12774 5772
rect 14274 5760 14280 5772
rect 14235 5732 14280 5760
rect 14274 5720 14280 5732
rect 14332 5720 14338 5772
rect 15948 5769 15976 5800
rect 15933 5763 15991 5769
rect 15933 5729 15945 5763
rect 15979 5729 15991 5763
rect 15933 5723 15991 5729
rect 16844 5763 16902 5769
rect 16844 5729 16856 5763
rect 16890 5760 16902 5763
rect 17310 5760 17316 5772
rect 16890 5732 17316 5760
rect 16890 5729 16902 5732
rect 16844 5723 16902 5729
rect 17310 5720 17316 5732
rect 17368 5720 17374 5772
rect 2406 5652 2412 5704
rect 2464 5692 2470 5704
rect 2501 5695 2559 5701
rect 2501 5692 2513 5695
rect 2464 5664 2513 5692
rect 2464 5652 2470 5664
rect 2501 5661 2513 5664
rect 2547 5661 2559 5695
rect 3602 5692 3608 5704
rect 3563 5664 3608 5692
rect 2501 5655 2559 5661
rect 3602 5652 3608 5664
rect 3660 5652 3666 5704
rect 3878 5652 3884 5704
rect 3936 5692 3942 5704
rect 4525 5695 4583 5701
rect 4525 5692 4537 5695
rect 3936 5664 4537 5692
rect 3936 5652 3942 5664
rect 4525 5661 4537 5664
rect 4571 5661 4583 5695
rect 4706 5692 4712 5704
rect 4667 5664 4712 5692
rect 4525 5655 4583 5661
rect 4540 5624 4568 5655
rect 4706 5652 4712 5664
rect 4764 5652 4770 5704
rect 4798 5652 4804 5704
rect 4856 5692 4862 5704
rect 5074 5692 5080 5704
rect 4856 5664 5080 5692
rect 4856 5652 4862 5664
rect 5074 5652 5080 5664
rect 5132 5652 5138 5704
rect 7024 5692 7052 5720
rect 7653 5695 7711 5701
rect 7653 5692 7665 5695
rect 7024 5664 7665 5692
rect 7653 5661 7665 5664
rect 7699 5661 7711 5695
rect 7653 5655 7711 5661
rect 11790 5652 11796 5704
rect 11848 5692 11854 5704
rect 11885 5695 11943 5701
rect 11885 5692 11897 5695
rect 11848 5664 11897 5692
rect 11848 5652 11854 5664
rect 11885 5661 11897 5664
rect 11931 5661 11943 5695
rect 11885 5655 11943 5661
rect 12989 5695 13047 5701
rect 12989 5661 13001 5695
rect 13035 5692 13047 5695
rect 13078 5692 13084 5704
rect 13035 5664 13084 5692
rect 13035 5661 13047 5664
rect 12989 5655 13047 5661
rect 13078 5652 13084 5664
rect 13136 5652 13142 5704
rect 14458 5692 14464 5704
rect 14419 5664 14464 5692
rect 14458 5652 14464 5664
rect 14516 5652 14522 5704
rect 16390 5652 16396 5704
rect 16448 5692 16454 5704
rect 16577 5695 16635 5701
rect 16577 5692 16589 5695
rect 16448 5664 16589 5692
rect 16448 5652 16454 5664
rect 16577 5661 16589 5664
rect 16623 5661 16635 5695
rect 16577 5655 16635 5661
rect 5626 5624 5632 5636
rect 4540 5596 5632 5624
rect 5626 5584 5632 5596
rect 5684 5584 5690 5636
rect 7377 5627 7435 5633
rect 7377 5593 7389 5627
rect 7423 5624 7435 5627
rect 7561 5627 7619 5633
rect 7561 5624 7573 5627
rect 7423 5596 7573 5624
rect 7423 5593 7435 5596
rect 7377 5587 7435 5593
rect 7561 5593 7573 5596
rect 7607 5593 7619 5627
rect 16482 5624 16488 5636
rect 7561 5587 7619 5593
rect 10612 5596 16488 5624
rect 3142 5516 3148 5568
rect 3200 5556 3206 5568
rect 3786 5556 3792 5568
rect 3200 5528 3792 5556
rect 3200 5516 3206 5528
rect 3786 5516 3792 5528
rect 3844 5516 3850 5568
rect 3881 5559 3939 5565
rect 3881 5525 3893 5559
rect 3927 5556 3939 5559
rect 4065 5559 4123 5565
rect 4065 5556 4077 5559
rect 3927 5528 4077 5556
rect 3927 5525 3939 5528
rect 3881 5519 3939 5525
rect 4065 5525 4077 5528
rect 4111 5525 4123 5559
rect 4065 5519 4123 5525
rect 4246 5516 4252 5568
rect 4304 5556 4310 5568
rect 5077 5559 5135 5565
rect 5077 5556 5089 5559
rect 4304 5528 5089 5556
rect 4304 5516 4310 5528
rect 5077 5525 5089 5528
rect 5123 5525 5135 5559
rect 5077 5519 5135 5525
rect 7466 5516 7472 5568
rect 7524 5556 7530 5568
rect 8018 5556 8024 5568
rect 7524 5528 8024 5556
rect 7524 5516 7530 5528
rect 8018 5516 8024 5528
rect 8076 5556 8082 5568
rect 9033 5559 9091 5565
rect 9033 5556 9045 5559
rect 8076 5528 9045 5556
rect 8076 5516 8082 5528
rect 9033 5525 9045 5528
rect 9079 5525 9091 5559
rect 9033 5519 9091 5525
rect 9214 5516 9220 5568
rect 9272 5556 9278 5568
rect 10612 5556 10640 5596
rect 16482 5584 16488 5596
rect 16540 5584 16546 5636
rect 11054 5556 11060 5568
rect 9272 5528 10640 5556
rect 11015 5528 11060 5556
rect 9272 5516 9278 5528
rect 11054 5516 11060 5528
rect 11112 5516 11118 5568
rect 12345 5559 12403 5565
rect 12345 5525 12357 5559
rect 12391 5556 12403 5559
rect 12802 5556 12808 5568
rect 12391 5528 12808 5556
rect 12391 5525 12403 5528
rect 12345 5519 12403 5525
rect 12802 5516 12808 5528
rect 12860 5516 12866 5568
rect 13262 5516 13268 5568
rect 13320 5556 13326 5568
rect 13357 5559 13415 5565
rect 13357 5556 13369 5559
rect 13320 5528 13369 5556
rect 13320 5516 13326 5528
rect 13357 5525 13369 5528
rect 13403 5525 13415 5559
rect 13357 5519 13415 5525
rect 15749 5559 15807 5565
rect 15749 5525 15761 5559
rect 15795 5556 15807 5559
rect 16022 5556 16028 5568
rect 15795 5528 16028 5556
rect 15795 5525 15807 5528
rect 15749 5519 15807 5525
rect 16022 5516 16028 5528
rect 16080 5556 16086 5568
rect 16390 5556 16396 5568
rect 16080 5528 16396 5556
rect 16080 5516 16086 5528
rect 16390 5516 16396 5528
rect 16448 5516 16454 5568
rect 17218 5516 17224 5568
rect 17276 5556 17282 5568
rect 17957 5559 18015 5565
rect 17957 5556 17969 5559
rect 17276 5528 17969 5556
rect 17276 5516 17282 5528
rect 17957 5525 17969 5528
rect 18003 5525 18015 5559
rect 17957 5519 18015 5525
rect 1104 5466 21896 5488
rect 1104 5414 4447 5466
rect 4499 5414 4511 5466
rect 4563 5414 4575 5466
rect 4627 5414 4639 5466
rect 4691 5414 11378 5466
rect 11430 5414 11442 5466
rect 11494 5414 11506 5466
rect 11558 5414 11570 5466
rect 11622 5414 18308 5466
rect 18360 5414 18372 5466
rect 18424 5414 18436 5466
rect 18488 5414 18500 5466
rect 18552 5414 21896 5466
rect 1104 5392 21896 5414
rect 3513 5355 3571 5361
rect 3513 5321 3525 5355
rect 3559 5352 3571 5355
rect 3970 5352 3976 5364
rect 3559 5324 3976 5352
rect 3559 5321 3571 5324
rect 3513 5315 3571 5321
rect 3970 5312 3976 5324
rect 4028 5312 4034 5364
rect 6730 5312 6736 5364
rect 6788 5352 6794 5364
rect 7837 5355 7895 5361
rect 7837 5352 7849 5355
rect 6788 5324 7849 5352
rect 6788 5312 6794 5324
rect 7837 5321 7849 5324
rect 7883 5352 7895 5355
rect 11885 5355 11943 5361
rect 7883 5324 10916 5352
rect 7883 5321 7895 5324
rect 7837 5315 7895 5321
rect 7009 5287 7067 5293
rect 7009 5253 7021 5287
rect 7055 5284 7067 5287
rect 9309 5287 9367 5293
rect 7055 5256 8524 5284
rect 7055 5253 7067 5256
rect 7009 5247 7067 5253
rect 6365 5219 6423 5225
rect 6365 5185 6377 5219
rect 6411 5216 6423 5219
rect 7466 5216 7472 5228
rect 6411 5188 7472 5216
rect 6411 5185 6423 5188
rect 6365 5179 6423 5185
rect 7466 5176 7472 5188
rect 7524 5176 7530 5228
rect 7558 5176 7564 5228
rect 7616 5216 7622 5228
rect 8496 5225 8524 5256
rect 9309 5253 9321 5287
rect 9355 5284 9367 5287
rect 10888 5284 10916 5324
rect 11885 5321 11897 5355
rect 11931 5352 11943 5355
rect 11974 5352 11980 5364
rect 11931 5324 11980 5352
rect 11931 5321 11943 5324
rect 11885 5315 11943 5321
rect 11974 5312 11980 5324
rect 12032 5312 12038 5364
rect 12158 5312 12164 5364
rect 12216 5352 12222 5364
rect 13262 5352 13268 5364
rect 12216 5324 13268 5352
rect 12216 5312 12222 5324
rect 13262 5312 13268 5324
rect 13320 5352 13326 5364
rect 16485 5355 16543 5361
rect 16485 5352 16497 5355
rect 13320 5324 16497 5352
rect 13320 5312 13326 5324
rect 16485 5321 16497 5324
rect 16531 5321 16543 5355
rect 16485 5315 16543 5321
rect 16577 5355 16635 5361
rect 16577 5321 16589 5355
rect 16623 5352 16635 5355
rect 18138 5352 18144 5364
rect 16623 5324 18144 5352
rect 16623 5321 16635 5324
rect 16577 5315 16635 5321
rect 18138 5312 18144 5324
rect 18196 5312 18202 5364
rect 12986 5284 12992 5296
rect 9355 5256 10824 5284
rect 10888 5256 12992 5284
rect 9355 5253 9367 5256
rect 9309 5247 9367 5253
rect 8481 5219 8539 5225
rect 7616 5188 7661 5216
rect 7616 5176 7622 5188
rect 8481 5185 8493 5219
rect 8527 5185 8539 5219
rect 8662 5216 8668 5228
rect 8623 5188 8668 5216
rect 8481 5179 8539 5185
rect 8662 5176 8668 5188
rect 8720 5176 8726 5228
rect 9950 5216 9956 5228
rect 9911 5188 9956 5216
rect 9950 5176 9956 5188
rect 10008 5176 10014 5228
rect 10796 5225 10824 5256
rect 12986 5244 12992 5256
rect 13044 5244 13050 5296
rect 16390 5244 16396 5296
rect 16448 5284 16454 5296
rect 16448 5256 20024 5284
rect 16448 5244 16454 5256
rect 10781 5219 10839 5225
rect 10781 5185 10793 5219
rect 10827 5185 10839 5219
rect 10781 5179 10839 5185
rect 10965 5219 11023 5225
rect 10965 5185 10977 5219
rect 11011 5216 11023 5219
rect 11054 5216 11060 5228
rect 11011 5188 11060 5216
rect 11011 5185 11023 5188
rect 10965 5179 11023 5185
rect 11054 5176 11060 5188
rect 11112 5176 11118 5228
rect 12437 5219 12495 5225
rect 12437 5185 12449 5219
rect 12483 5216 12495 5219
rect 12710 5216 12716 5228
rect 12483 5188 12716 5216
rect 12483 5185 12495 5188
rect 12437 5179 12495 5185
rect 12710 5176 12716 5188
rect 12768 5176 12774 5228
rect 13354 5176 13360 5228
rect 13412 5216 13418 5228
rect 13633 5219 13691 5225
rect 13633 5216 13645 5219
rect 13412 5188 13645 5216
rect 13412 5176 13418 5188
rect 13633 5185 13645 5188
rect 13679 5216 13691 5219
rect 14090 5216 14096 5228
rect 13679 5188 14096 5216
rect 13679 5185 13691 5188
rect 13633 5179 13691 5185
rect 14090 5176 14096 5188
rect 14148 5176 14154 5228
rect 14366 5176 14372 5228
rect 14424 5216 14430 5228
rect 15473 5219 15531 5225
rect 15473 5216 15485 5219
rect 14424 5188 15485 5216
rect 14424 5176 14430 5188
rect 15473 5185 15485 5188
rect 15519 5185 15531 5219
rect 15473 5179 15531 5185
rect 16209 5219 16267 5225
rect 16209 5185 16221 5219
rect 16255 5216 16267 5219
rect 16574 5216 16580 5228
rect 16255 5188 16580 5216
rect 16255 5185 16267 5188
rect 16209 5179 16267 5185
rect 16574 5176 16580 5188
rect 16632 5176 16638 5228
rect 17218 5216 17224 5228
rect 17179 5188 17224 5216
rect 17218 5176 17224 5188
rect 17276 5176 17282 5228
rect 19996 5225 20024 5256
rect 19981 5219 20039 5225
rect 19981 5185 19993 5219
rect 20027 5185 20039 5219
rect 19981 5179 20039 5185
rect 3510 5108 3516 5160
rect 3568 5148 3574 5160
rect 3878 5148 3884 5160
rect 3568 5120 3884 5148
rect 3568 5108 3574 5120
rect 3878 5108 3884 5120
rect 3936 5108 3942 5160
rect 6089 5151 6147 5157
rect 6089 5117 6101 5151
rect 6135 5148 6147 5151
rect 6822 5148 6828 5160
rect 6135 5120 6828 5148
rect 6135 5117 6147 5120
rect 6089 5111 6147 5117
rect 6822 5108 6828 5120
rect 6880 5108 6886 5160
rect 9677 5151 9735 5157
rect 9677 5117 9689 5151
rect 9723 5148 9735 5151
rect 9858 5148 9864 5160
rect 9723 5120 9864 5148
rect 9723 5117 9735 5120
rect 9677 5111 9735 5117
rect 9858 5108 9864 5120
rect 9916 5108 9922 5160
rect 14553 5151 14611 5157
rect 14553 5148 14565 5151
rect 10336 5120 14565 5148
rect 6181 5083 6239 5089
rect 6181 5049 6193 5083
rect 6227 5080 6239 5083
rect 6227 5052 8064 5080
rect 6227 5049 6239 5052
rect 6181 5043 6239 5049
rect 3878 4972 3884 5024
rect 3936 5012 3942 5024
rect 4249 5015 4307 5021
rect 4249 5012 4261 5015
rect 3936 4984 4261 5012
rect 3936 4972 3942 4984
rect 4249 4981 4261 4984
rect 4295 5012 4307 5015
rect 4890 5012 4896 5024
rect 4295 4984 4896 5012
rect 4295 4981 4307 4984
rect 4249 4975 4307 4981
rect 4890 4972 4896 4984
rect 4948 4972 4954 5024
rect 5721 5015 5779 5021
rect 5721 4981 5733 5015
rect 5767 5012 5779 5015
rect 7006 5012 7012 5024
rect 5767 4984 7012 5012
rect 5767 4981 5779 4984
rect 5721 4975 5779 4981
rect 7006 4972 7012 4984
rect 7064 4972 7070 5024
rect 7282 4972 7288 5024
rect 7340 5012 7346 5024
rect 8036 5021 8064 5052
rect 7377 5015 7435 5021
rect 7377 5012 7389 5015
rect 7340 4984 7389 5012
rect 7340 4972 7346 4984
rect 7377 4981 7389 4984
rect 7423 4981 7435 5015
rect 7377 4975 7435 4981
rect 7469 5015 7527 5021
rect 7469 4981 7481 5015
rect 7515 5012 7527 5015
rect 7837 5015 7895 5021
rect 7837 5012 7849 5015
rect 7515 4984 7849 5012
rect 7515 4981 7527 4984
rect 7469 4975 7527 4981
rect 7837 4981 7849 4984
rect 7883 4981 7895 5015
rect 7837 4975 7895 4981
rect 8021 5015 8079 5021
rect 8021 4981 8033 5015
rect 8067 4981 8079 5015
rect 8021 4975 8079 4981
rect 8202 4972 8208 5024
rect 8260 5012 8266 5024
rect 8389 5015 8447 5021
rect 8389 5012 8401 5015
rect 8260 4984 8401 5012
rect 8260 4972 8266 4984
rect 8389 4981 8401 4984
rect 8435 4981 8447 5015
rect 9766 5012 9772 5024
rect 9727 4984 9772 5012
rect 8389 4975 8447 4981
rect 9766 4972 9772 4984
rect 9824 4972 9830 5024
rect 10336 5021 10364 5120
rect 14553 5117 14565 5120
rect 14599 5117 14611 5151
rect 14553 5111 14611 5117
rect 16114 5108 16120 5160
rect 16172 5148 16178 5160
rect 16945 5151 17003 5157
rect 16945 5148 16957 5151
rect 16172 5120 16957 5148
rect 16172 5108 16178 5120
rect 16945 5117 16957 5120
rect 16991 5148 17003 5151
rect 17589 5151 17647 5157
rect 17589 5148 17601 5151
rect 16991 5120 17601 5148
rect 16991 5117 17003 5120
rect 16945 5111 17003 5117
rect 17589 5117 17601 5120
rect 17635 5117 17647 5151
rect 17589 5111 17647 5117
rect 20248 5151 20306 5157
rect 20248 5117 20260 5151
rect 20294 5148 20306 5151
rect 20622 5148 20628 5160
rect 20294 5120 20628 5148
rect 20294 5117 20306 5120
rect 20248 5111 20306 5117
rect 20622 5108 20628 5120
rect 20680 5108 20686 5160
rect 10689 5083 10747 5089
rect 10689 5049 10701 5083
rect 10735 5080 10747 5083
rect 11333 5083 11391 5089
rect 11333 5080 11345 5083
rect 10735 5052 11345 5080
rect 10735 5049 10747 5052
rect 10689 5043 10747 5049
rect 11333 5049 11345 5052
rect 11379 5049 11391 5083
rect 11333 5043 11391 5049
rect 14829 5083 14887 5089
rect 14829 5049 14841 5083
rect 14875 5080 14887 5083
rect 15378 5080 15384 5092
rect 14875 5052 15384 5080
rect 14875 5049 14887 5052
rect 14829 5043 14887 5049
rect 15378 5040 15384 5052
rect 15436 5040 15442 5092
rect 15473 5083 15531 5089
rect 15473 5049 15485 5083
rect 15519 5080 15531 5083
rect 15933 5083 15991 5089
rect 15933 5080 15945 5083
rect 15519 5052 15945 5080
rect 15519 5049 15531 5052
rect 15473 5043 15531 5049
rect 15933 5049 15945 5052
rect 15979 5049 15991 5083
rect 15933 5043 15991 5049
rect 10321 5015 10379 5021
rect 10321 4981 10333 5015
rect 10367 4981 10379 5015
rect 10321 4975 10379 4981
rect 11790 4972 11796 5024
rect 11848 5012 11854 5024
rect 12434 5012 12440 5024
rect 11848 4984 12440 5012
rect 11848 4972 11854 4984
rect 12434 4972 12440 4984
rect 12492 4972 12498 5024
rect 13170 5012 13176 5024
rect 13131 4984 13176 5012
rect 13170 4972 13176 4984
rect 13228 4972 13234 5024
rect 15562 5012 15568 5024
rect 15523 4984 15568 5012
rect 15562 4972 15568 4984
rect 15620 4972 15626 5024
rect 16022 5012 16028 5024
rect 15983 4984 16028 5012
rect 16022 4972 16028 4984
rect 16080 4972 16086 5024
rect 16485 5015 16543 5021
rect 16485 4981 16497 5015
rect 16531 5012 16543 5015
rect 17037 5015 17095 5021
rect 17037 5012 17049 5015
rect 16531 4984 17049 5012
rect 16531 4981 16543 4984
rect 16485 4975 16543 4981
rect 17037 4981 17049 4984
rect 17083 5012 17095 5015
rect 18049 5015 18107 5021
rect 18049 5012 18061 5015
rect 17083 4984 18061 5012
rect 17083 4981 17095 4984
rect 17037 4975 17095 4981
rect 18049 4981 18061 4984
rect 18095 5012 18107 5015
rect 21266 5012 21272 5024
rect 18095 4984 21272 5012
rect 18095 4981 18107 4984
rect 18049 4975 18107 4981
rect 21266 4972 21272 4984
rect 21324 4972 21330 5024
rect 21361 5015 21419 5021
rect 21361 4981 21373 5015
rect 21407 5012 21419 5015
rect 22005 5015 22063 5021
rect 22005 5012 22017 5015
rect 21407 4984 22017 5012
rect 21407 4981 21419 4984
rect 21361 4975 21419 4981
rect 22005 4981 22017 4984
rect 22051 4981 22063 5015
rect 22005 4975 22063 4981
rect 1104 4922 21896 4944
rect 1104 4870 7912 4922
rect 7964 4870 7976 4922
rect 8028 4870 8040 4922
rect 8092 4870 8104 4922
rect 8156 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 15035 4922
rect 15087 4870 21896 4922
rect 1104 4848 21896 4870
rect 1486 4808 1492 4820
rect 1447 4780 1492 4808
rect 1486 4768 1492 4780
rect 1544 4768 1550 4820
rect 1857 4811 1915 4817
rect 1857 4777 1869 4811
rect 1903 4808 1915 4811
rect 3237 4811 3295 4817
rect 3237 4808 3249 4811
rect 1903 4780 3249 4808
rect 1903 4777 1915 4780
rect 1857 4771 1915 4777
rect 3237 4777 3249 4780
rect 3283 4777 3295 4811
rect 3237 4771 3295 4777
rect 4062 4768 4068 4820
rect 4120 4808 4126 4820
rect 4525 4811 4583 4817
rect 4525 4808 4537 4811
rect 4120 4780 4537 4808
rect 4120 4768 4126 4780
rect 4525 4777 4537 4780
rect 4571 4808 4583 4811
rect 5626 4808 5632 4820
rect 4571 4780 5632 4808
rect 4571 4777 4583 4780
rect 4525 4771 4583 4777
rect 5626 4768 5632 4780
rect 5684 4768 5690 4820
rect 5718 4768 5724 4820
rect 5776 4808 5782 4820
rect 6730 4808 6736 4820
rect 5776 4780 6736 4808
rect 5776 4768 5782 4780
rect 6730 4768 6736 4780
rect 6788 4768 6794 4820
rect 7101 4811 7159 4817
rect 7101 4777 7113 4811
rect 7147 4808 7159 4811
rect 8202 4808 8208 4820
rect 7147 4780 8208 4808
rect 7147 4777 7159 4780
rect 7101 4771 7159 4777
rect 8202 4768 8208 4780
rect 8260 4768 8266 4820
rect 9950 4768 9956 4820
rect 10008 4808 10014 4820
rect 10870 4808 10876 4820
rect 10008 4780 10876 4808
rect 10008 4768 10014 4780
rect 10870 4768 10876 4780
rect 10928 4768 10934 4820
rect 14366 4768 14372 4820
rect 14424 4808 14430 4820
rect 14829 4811 14887 4817
rect 14829 4808 14841 4811
rect 14424 4780 14841 4808
rect 14424 4768 14430 4780
rect 14829 4777 14841 4780
rect 14875 4777 14887 4811
rect 14829 4771 14887 4777
rect 15562 4768 15568 4820
rect 15620 4808 15626 4820
rect 18049 4811 18107 4817
rect 18049 4808 18061 4811
rect 15620 4780 18061 4808
rect 15620 4768 15626 4780
rect 18049 4777 18061 4780
rect 18095 4777 18107 4811
rect 18049 4771 18107 4777
rect 20622 4768 20628 4820
rect 20680 4808 20686 4820
rect 21269 4811 21327 4817
rect 21269 4808 21281 4811
rect 20680 4780 21281 4808
rect 20680 4768 20686 4780
rect 21269 4777 21281 4780
rect 21315 4777 21327 4811
rect 21269 4771 21327 4777
rect 1504 4740 1532 4768
rect 2317 4743 2375 4749
rect 2317 4740 2329 4743
rect 1504 4712 2329 4740
rect 2317 4709 2329 4712
rect 2363 4709 2375 4743
rect 2317 4703 2375 4709
rect 3970 4700 3976 4752
rect 4028 4740 4034 4752
rect 7374 4740 7380 4752
rect 4028 4712 7380 4740
rect 4028 4700 4034 4712
rect 7374 4700 7380 4712
rect 7432 4740 7438 4752
rect 7466 4740 7472 4752
rect 7432 4712 7472 4740
rect 7432 4700 7438 4712
rect 7466 4700 7472 4712
rect 7524 4740 7530 4752
rect 8573 4743 8631 4749
rect 8573 4740 8585 4743
rect 7524 4712 8585 4740
rect 7524 4700 7530 4712
rect 8573 4709 8585 4712
rect 8619 4740 8631 4743
rect 10772 4743 10830 4749
rect 8619 4712 10732 4740
rect 8619 4709 8631 4712
rect 8573 4703 8631 4709
rect 1486 4632 1492 4684
rect 1544 4672 1550 4684
rect 2225 4675 2283 4681
rect 2225 4672 2237 4675
rect 1544 4644 2237 4672
rect 1544 4632 1550 4644
rect 2225 4641 2237 4644
rect 2271 4641 2283 4675
rect 2225 4635 2283 4641
rect 5629 4675 5687 4681
rect 5629 4641 5641 4675
rect 5675 4672 5687 4675
rect 6270 4672 6276 4684
rect 5675 4644 6276 4672
rect 5675 4641 5687 4644
rect 5629 4635 5687 4641
rect 6270 4632 6276 4644
rect 6328 4632 6334 4684
rect 7282 4672 7288 4684
rect 6380 4644 7288 4672
rect 2498 4604 2504 4616
rect 2459 4576 2504 4604
rect 2498 4564 2504 4576
rect 2556 4564 2562 4616
rect 3326 4604 3332 4616
rect 3287 4576 3332 4604
rect 3326 4564 3332 4576
rect 3384 4564 3390 4616
rect 3418 4564 3424 4616
rect 3476 4604 3482 4616
rect 3476 4576 3521 4604
rect 3476 4564 3482 4576
rect 5258 4564 5264 4616
rect 5316 4604 5322 4616
rect 5721 4607 5779 4613
rect 5721 4604 5733 4607
rect 5316 4576 5733 4604
rect 5316 4564 5322 4576
rect 5721 4573 5733 4576
rect 5767 4573 5779 4607
rect 5902 4604 5908 4616
rect 5863 4576 5908 4604
rect 5721 4567 5779 4573
rect 5902 4564 5908 4576
rect 5960 4564 5966 4616
rect 6086 4564 6092 4616
rect 6144 4604 6150 4616
rect 6380 4613 6408 4644
rect 7282 4632 7288 4644
rect 7340 4632 7346 4684
rect 8110 4672 8116 4684
rect 7576 4644 8116 4672
rect 6365 4607 6423 4613
rect 6365 4604 6377 4607
rect 6144 4576 6377 4604
rect 6144 4564 6150 4576
rect 6365 4573 6377 4576
rect 6411 4573 6423 4607
rect 6365 4567 6423 4573
rect 6914 4564 6920 4616
rect 6972 4604 6978 4616
rect 7576 4613 7604 4644
rect 8110 4632 8116 4644
rect 8168 4632 8174 4684
rect 10134 4672 10140 4684
rect 10095 4644 10140 4672
rect 10134 4632 10140 4644
rect 10192 4632 10198 4684
rect 10704 4672 10732 4712
rect 10772 4709 10784 4743
rect 10818 4740 10830 4743
rect 11054 4740 11060 4752
rect 10818 4712 11060 4740
rect 10818 4709 10830 4712
rect 10772 4703 10830 4709
rect 11054 4700 11060 4712
rect 11112 4700 11118 4752
rect 15473 4743 15531 4749
rect 15473 4740 15485 4743
rect 11256 4712 15485 4740
rect 11256 4672 11284 4712
rect 15473 4709 15485 4712
rect 15519 4740 15531 4743
rect 16022 4740 16028 4752
rect 15519 4712 16028 4740
rect 15519 4709 15531 4712
rect 15473 4703 15531 4709
rect 16022 4700 16028 4712
rect 16080 4700 16086 4752
rect 16390 4740 16396 4752
rect 16132 4712 16396 4740
rect 10704 4644 11284 4672
rect 13072 4675 13130 4681
rect 13072 4641 13084 4675
rect 13118 4672 13130 4675
rect 13630 4672 13636 4684
rect 13118 4644 13636 4672
rect 13118 4641 13130 4644
rect 13072 4635 13130 4641
rect 13630 4632 13636 4644
rect 13688 4632 13694 4684
rect 15746 4632 15752 4684
rect 15804 4672 15810 4684
rect 15933 4675 15991 4681
rect 15933 4672 15945 4675
rect 15804 4644 15945 4672
rect 15804 4632 15810 4644
rect 15933 4641 15945 4644
rect 15979 4672 15991 4675
rect 16132 4672 16160 4712
rect 16390 4700 16396 4712
rect 16448 4700 16454 4752
rect 15979 4644 16160 4672
rect 16200 4675 16258 4681
rect 15979 4641 15991 4644
rect 15933 4635 15991 4641
rect 16200 4641 16212 4675
rect 16246 4672 16258 4675
rect 16574 4672 16580 4684
rect 16246 4644 16580 4672
rect 16246 4641 16258 4644
rect 16200 4635 16258 4641
rect 16574 4632 16580 4644
rect 16632 4672 16638 4684
rect 17126 4672 17132 4684
rect 16632 4644 17132 4672
rect 16632 4632 16638 4644
rect 17126 4632 17132 4644
rect 17184 4632 17190 4684
rect 17954 4672 17960 4684
rect 17915 4644 17960 4672
rect 17954 4632 17960 4644
rect 18012 4632 18018 4684
rect 7561 4607 7619 4613
rect 7561 4604 7573 4607
rect 6972 4576 7573 4604
rect 6972 4564 6978 4576
rect 7561 4573 7573 4576
rect 7607 4573 7619 4607
rect 7561 4567 7619 4573
rect 7650 4564 7656 4616
rect 7708 4604 7714 4616
rect 7708 4576 7753 4604
rect 7708 4564 7714 4576
rect 8202 4564 8208 4616
rect 8260 4604 8266 4616
rect 9125 4607 9183 4613
rect 9125 4604 9137 4607
rect 8260 4576 9137 4604
rect 8260 4564 8266 4576
rect 9125 4573 9137 4576
rect 9171 4573 9183 4607
rect 9125 4567 9183 4573
rect 4062 4496 4068 4548
rect 4120 4536 4126 4548
rect 9140 4536 9168 4567
rect 9306 4564 9312 4616
rect 9364 4604 9370 4616
rect 10152 4604 10180 4632
rect 10502 4604 10508 4616
rect 9364 4576 10180 4604
rect 10463 4576 10508 4604
rect 9364 4564 9370 4576
rect 10502 4564 10508 4576
rect 10560 4564 10566 4616
rect 12805 4607 12863 4613
rect 12805 4573 12817 4607
rect 12851 4573 12863 4607
rect 12805 4567 12863 4573
rect 18141 4607 18199 4613
rect 18141 4573 18153 4607
rect 18187 4573 18199 4607
rect 18141 4567 18199 4573
rect 9766 4536 9772 4548
rect 4120 4508 8248 4536
rect 9140 4508 9772 4536
rect 4120 4496 4126 4508
rect 2869 4471 2927 4477
rect 2869 4437 2881 4471
rect 2915 4468 2927 4471
rect 3142 4468 3148 4480
rect 2915 4440 3148 4468
rect 2915 4437 2927 4440
rect 2869 4431 2927 4437
rect 3142 4428 3148 4440
rect 3200 4428 3206 4480
rect 4890 4468 4896 4480
rect 4851 4440 4896 4468
rect 4890 4428 4896 4440
rect 4948 4428 4954 4480
rect 5261 4471 5319 4477
rect 5261 4437 5273 4471
rect 5307 4468 5319 4471
rect 6178 4468 6184 4480
rect 5307 4440 6184 4468
rect 5307 4437 5319 4440
rect 5261 4431 5319 4437
rect 6178 4428 6184 4440
rect 6236 4428 6242 4480
rect 8220 4468 8248 4508
rect 9766 4496 9772 4508
rect 9824 4536 9830 4548
rect 10134 4536 10140 4548
rect 9824 4508 10140 4536
rect 9824 4496 9830 4508
rect 10134 4496 10140 4508
rect 10192 4496 10198 4548
rect 8386 4468 8392 4480
rect 8220 4440 8392 4468
rect 8386 4428 8392 4440
rect 8444 4428 8450 4480
rect 9674 4468 9680 4480
rect 9635 4440 9680 4468
rect 9674 4428 9680 4440
rect 9732 4428 9738 4480
rect 11885 4471 11943 4477
rect 11885 4437 11897 4471
rect 11931 4468 11943 4471
rect 12434 4468 12440 4480
rect 11931 4440 12440 4468
rect 11931 4437 11943 4440
rect 11885 4431 11943 4437
rect 12434 4428 12440 4440
rect 12492 4428 12498 4480
rect 12820 4468 12848 4567
rect 17310 4536 17316 4548
rect 17271 4508 17316 4536
rect 17310 4496 17316 4508
rect 17368 4536 17374 4548
rect 18156 4536 18184 4567
rect 17368 4508 18184 4536
rect 17368 4496 17374 4508
rect 13814 4468 13820 4480
rect 12820 4440 13820 4468
rect 13814 4428 13820 4440
rect 13872 4428 13878 4480
rect 14182 4468 14188 4480
rect 14143 4440 14188 4468
rect 14182 4428 14188 4440
rect 14240 4428 14246 4480
rect 16850 4428 16856 4480
rect 16908 4468 16914 4480
rect 17589 4471 17647 4477
rect 17589 4468 17601 4471
rect 16908 4440 17601 4468
rect 16908 4428 16914 4440
rect 17589 4437 17601 4440
rect 17635 4437 17647 4471
rect 17589 4431 17647 4437
rect 1104 4378 21896 4400
rect 1104 4326 4447 4378
rect 4499 4326 4511 4378
rect 4563 4326 4575 4378
rect 4627 4326 4639 4378
rect 4691 4326 11378 4378
rect 11430 4326 11442 4378
rect 11494 4326 11506 4378
rect 11558 4326 11570 4378
rect 11622 4326 18308 4378
rect 18360 4326 18372 4378
rect 18424 4326 18436 4378
rect 18488 4326 18500 4378
rect 18552 4326 21896 4378
rect 1104 4304 21896 4326
rect 3329 4267 3387 4273
rect 3329 4233 3341 4267
rect 3375 4264 3387 4267
rect 3418 4264 3424 4276
rect 3375 4236 3424 4264
rect 3375 4233 3387 4236
rect 3329 4227 3387 4233
rect 3418 4224 3424 4236
rect 3476 4224 3482 4276
rect 4890 4224 4896 4276
rect 4948 4264 4954 4276
rect 5258 4264 5264 4276
rect 4948 4236 5120 4264
rect 5219 4236 5264 4264
rect 4948 4224 4954 4236
rect 1486 4128 1492 4140
rect 1447 4100 1492 4128
rect 1486 4088 1492 4100
rect 1544 4088 1550 4140
rect 3436 4128 3464 4224
rect 4985 4199 5043 4205
rect 4985 4165 4997 4199
rect 5031 4165 5043 4199
rect 5092 4196 5120 4236
rect 5258 4224 5264 4236
rect 5316 4224 5322 4276
rect 5534 4224 5540 4276
rect 5592 4264 5598 4276
rect 6454 4264 6460 4276
rect 5592 4236 6460 4264
rect 5592 4224 5598 4236
rect 5092 4168 5672 4196
rect 4985 4159 5043 4165
rect 5000 4128 5028 4159
rect 5534 4128 5540 4140
rect 3436 4100 3740 4128
rect 5000 4100 5540 4128
rect 1946 4060 1952 4072
rect 1907 4032 1952 4060
rect 1946 4020 1952 4032
rect 2004 4020 2010 4072
rect 2682 4060 2688 4072
rect 2056 4032 2688 4060
rect 1486 3952 1492 4004
rect 1544 3992 1550 4004
rect 2056 3992 2084 4032
rect 2682 4020 2688 4032
rect 2740 4060 2746 4072
rect 3605 4063 3663 4069
rect 3605 4060 3617 4063
rect 2740 4032 3617 4060
rect 2740 4020 2746 4032
rect 3605 4029 3617 4032
rect 3651 4029 3663 4063
rect 3712 4060 3740 4100
rect 5534 4088 5540 4100
rect 5592 4088 5598 4140
rect 5644 4128 5672 4168
rect 5828 4137 5856 4236
rect 6454 4224 6460 4236
rect 6512 4224 6518 4276
rect 7558 4224 7564 4276
rect 7616 4264 7622 4276
rect 8205 4267 8263 4273
rect 8205 4264 8217 4267
rect 7616 4236 8217 4264
rect 7616 4224 7622 4236
rect 8205 4233 8217 4236
rect 8251 4233 8263 4267
rect 8205 4227 8263 4233
rect 10870 4224 10876 4276
rect 10928 4264 10934 4276
rect 17126 4264 17132 4276
rect 10928 4236 16896 4264
rect 17087 4236 17132 4264
rect 10928 4224 10934 4236
rect 10888 4196 10916 4224
rect 12434 4196 12440 4208
rect 9508 4168 10916 4196
rect 11624 4168 12440 4196
rect 5721 4131 5779 4137
rect 5721 4128 5733 4131
rect 5644 4100 5733 4128
rect 5721 4097 5733 4100
rect 5767 4097 5779 4131
rect 5721 4091 5779 4097
rect 5813 4131 5871 4137
rect 5813 4097 5825 4131
rect 5859 4097 5871 4131
rect 6270 4128 6276 4140
rect 6231 4100 6276 4128
rect 5813 4091 5871 4097
rect 3861 4063 3919 4069
rect 3861 4060 3873 4063
rect 3712 4032 3873 4060
rect 3605 4023 3663 4029
rect 3861 4029 3873 4032
rect 3907 4029 3919 4063
rect 5626 4060 5632 4072
rect 5587 4032 5632 4060
rect 3861 4023 3919 4029
rect 1544 3964 2084 3992
rect 2216 3995 2274 4001
rect 1544 3952 1550 3964
rect 2216 3961 2228 3995
rect 2262 3992 2274 3995
rect 2498 3992 2504 4004
rect 2262 3964 2504 3992
rect 2262 3961 2274 3964
rect 2216 3955 2274 3961
rect 2498 3952 2504 3964
rect 2556 3952 2562 4004
rect 3620 3992 3648 4023
rect 5626 4020 5632 4032
rect 5684 4020 5690 4072
rect 5166 3992 5172 4004
rect 3620 3964 5172 3992
rect 5166 3952 5172 3964
rect 5224 3952 5230 4004
rect 1302 3884 1308 3936
rect 1360 3924 1366 3936
rect 5626 3924 5632 3936
rect 1360 3896 5632 3924
rect 1360 3884 1366 3896
rect 5626 3884 5632 3896
rect 5684 3884 5690 3936
rect 5736 3924 5764 4091
rect 6270 4088 6276 4100
rect 6328 4088 6334 4140
rect 6822 4128 6828 4140
rect 6783 4100 6828 4128
rect 6822 4088 6828 4100
rect 6880 4088 6886 4140
rect 8110 4088 8116 4140
rect 8168 4128 8174 4140
rect 9508 4137 9536 4168
rect 9493 4131 9551 4137
rect 8168 4100 9352 4128
rect 8168 4088 8174 4100
rect 6840 4060 6868 4088
rect 6840 4032 7328 4060
rect 6638 3952 6644 4004
rect 6696 3992 6702 4004
rect 7070 3995 7128 4001
rect 7070 3992 7082 3995
rect 6696 3964 7082 3992
rect 6696 3952 6702 3964
rect 7070 3961 7082 3964
rect 7116 3961 7128 3995
rect 7300 3992 7328 4032
rect 7374 4020 7380 4072
rect 7432 4060 7438 4072
rect 8202 4060 8208 4072
rect 7432 4032 8208 4060
rect 7432 4020 7438 4032
rect 8202 4020 8208 4032
rect 8260 4020 8266 4072
rect 8386 4020 8392 4072
rect 8444 4060 8450 4072
rect 9217 4063 9275 4069
rect 9217 4060 9229 4063
rect 8444 4032 9229 4060
rect 8444 4020 8450 4032
rect 9217 4029 9229 4032
rect 9263 4029 9275 4063
rect 9324 4060 9352 4100
rect 9493 4097 9505 4131
rect 9539 4097 9551 4131
rect 10410 4128 10416 4140
rect 10371 4100 10416 4128
rect 9493 4091 9551 4097
rect 10410 4088 10416 4100
rect 10468 4088 10474 4140
rect 11422 4128 11428 4140
rect 10520 4100 11428 4128
rect 10520 4060 10548 4100
rect 11422 4088 11428 4100
rect 11480 4088 11486 4140
rect 11624 4137 11652 4168
rect 11609 4131 11667 4137
rect 11609 4097 11621 4131
rect 11655 4097 11667 4131
rect 12360 4128 12388 4168
rect 12434 4156 12440 4168
rect 12492 4156 12498 4208
rect 16868 4196 16896 4236
rect 17126 4224 17132 4236
rect 17184 4224 17190 4276
rect 22005 4199 22063 4205
rect 22005 4196 22017 4199
rect 16868 4168 22017 4196
rect 22005 4165 22017 4168
rect 22051 4165 22063 4199
rect 22005 4159 22063 4165
rect 15746 4128 15752 4140
rect 12360 4100 12572 4128
rect 15707 4100 15752 4128
rect 11609 4091 11667 4097
rect 9324 4032 10548 4060
rect 9217 4023 9275 4029
rect 10594 4020 10600 4072
rect 10652 4060 10658 4072
rect 12066 4060 12072 4072
rect 10652 4032 12072 4060
rect 10652 4020 10658 4032
rect 12066 4020 12072 4032
rect 12124 4020 12130 4072
rect 12342 4020 12348 4072
rect 12400 4060 12406 4072
rect 12437 4063 12495 4069
rect 12437 4060 12449 4063
rect 12400 4032 12449 4060
rect 12400 4020 12406 4032
rect 12437 4029 12449 4032
rect 12483 4029 12495 4063
rect 12544 4060 12572 4100
rect 15746 4088 15752 4100
rect 15804 4088 15810 4140
rect 17405 4131 17463 4137
rect 17405 4097 17417 4131
rect 17451 4128 17463 4131
rect 17954 4128 17960 4140
rect 17451 4100 17960 4128
rect 17451 4097 17463 4100
rect 17405 4091 17463 4097
rect 17954 4088 17960 4100
rect 18012 4088 18018 4140
rect 12693 4063 12751 4069
rect 12693 4060 12705 4063
rect 12544 4032 12705 4060
rect 12437 4023 12495 4029
rect 12693 4029 12705 4032
rect 12739 4029 12751 4063
rect 12693 4023 12751 4029
rect 13814 4020 13820 4072
rect 13872 4060 13878 4072
rect 14093 4063 14151 4069
rect 14093 4060 14105 4063
rect 13872 4032 14105 4060
rect 13872 4020 13878 4032
rect 14093 4029 14105 4032
rect 14139 4029 14151 4063
rect 14093 4023 14151 4029
rect 7558 3992 7564 4004
rect 7300 3964 7564 3992
rect 7070 3955 7128 3961
rect 7558 3952 7564 3964
rect 7616 3952 7622 4004
rect 9306 3992 9312 4004
rect 7668 3964 9312 3992
rect 7668 3924 7696 3964
rect 9306 3952 9312 3964
rect 9364 3952 9370 4004
rect 9766 3952 9772 4004
rect 9824 3992 9830 4004
rect 10321 3995 10379 4001
rect 10321 3992 10333 3995
rect 9824 3964 10333 3992
rect 9824 3952 9830 3964
rect 10321 3961 10333 3964
rect 10367 3961 10379 3995
rect 10321 3955 10379 3961
rect 10502 3952 10508 4004
rect 10560 3992 10566 4004
rect 12360 3992 12388 4020
rect 10560 3964 12388 3992
rect 14108 3992 14136 4023
rect 14182 4020 14188 4072
rect 14240 4060 14246 4072
rect 14366 4069 14372 4072
rect 14349 4063 14372 4069
rect 14349 4060 14361 4063
rect 14240 4032 14361 4060
rect 14240 4020 14246 4032
rect 14349 4029 14361 4032
rect 14424 4060 14430 4072
rect 15764 4060 15792 4088
rect 14424 4032 14497 4060
rect 14568 4032 15792 4060
rect 14349 4023 14372 4029
rect 14366 4020 14372 4023
rect 14424 4020 14430 4032
rect 14568 3992 14596 4032
rect 15838 3992 15844 4004
rect 14108 3964 14596 3992
rect 15488 3964 15844 3992
rect 10560 3952 10566 3964
rect 8478 3924 8484 3936
rect 5736 3896 7696 3924
rect 8439 3896 8484 3924
rect 8478 3884 8484 3896
rect 8536 3884 8542 3936
rect 8849 3927 8907 3933
rect 8849 3893 8861 3927
rect 8895 3924 8907 3927
rect 9122 3924 9128 3936
rect 8895 3896 9128 3924
rect 8895 3893 8907 3896
rect 8849 3887 8907 3893
rect 9122 3884 9128 3896
rect 9180 3884 9186 3936
rect 9858 3924 9864 3936
rect 9819 3896 9864 3924
rect 9858 3884 9864 3896
rect 9916 3884 9922 3936
rect 10226 3924 10232 3936
rect 10187 3896 10232 3924
rect 10226 3884 10232 3896
rect 10284 3884 10290 3936
rect 10962 3924 10968 3936
rect 10923 3896 10968 3924
rect 10962 3884 10968 3896
rect 11020 3884 11026 3936
rect 11238 3884 11244 3936
rect 11296 3924 11302 3936
rect 11333 3927 11391 3933
rect 11333 3924 11345 3927
rect 11296 3896 11345 3924
rect 11296 3884 11302 3896
rect 11333 3893 11345 3896
rect 11379 3924 11391 3927
rect 11977 3927 12035 3933
rect 11977 3924 11989 3927
rect 11379 3896 11989 3924
rect 11379 3893 11391 3896
rect 11333 3887 11391 3893
rect 11977 3893 11989 3896
rect 12023 3893 12035 3927
rect 11977 3887 12035 3893
rect 13630 3884 13636 3936
rect 13688 3924 13694 3936
rect 15488 3933 15516 3964
rect 15838 3952 15844 3964
rect 15896 3992 15902 4004
rect 15994 3995 16052 4001
rect 15994 3992 16006 3995
rect 15896 3964 16006 3992
rect 15896 3952 15902 3964
rect 15994 3961 16006 3964
rect 16040 3961 16052 3995
rect 15994 3955 16052 3961
rect 13817 3927 13875 3933
rect 13817 3924 13829 3927
rect 13688 3896 13829 3924
rect 13688 3884 13694 3896
rect 13817 3893 13829 3896
rect 13863 3893 13875 3927
rect 13817 3887 13875 3893
rect 15473 3927 15531 3933
rect 15473 3893 15485 3927
rect 15519 3893 15531 3927
rect 15473 3887 15531 3893
rect 21361 3927 21419 3933
rect 21361 3893 21373 3927
rect 21407 3924 21419 3927
rect 21818 3924 21824 3936
rect 21407 3896 21824 3924
rect 21407 3893 21419 3896
rect 21361 3887 21419 3893
rect 21818 3884 21824 3896
rect 21876 3884 21882 3936
rect 1104 3834 21896 3856
rect 1104 3782 7912 3834
rect 7964 3782 7976 3834
rect 8028 3782 8040 3834
rect 8092 3782 8104 3834
rect 8156 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 15035 3834
rect 15087 3782 21896 3834
rect 1104 3760 21896 3782
rect 3326 3680 3332 3732
rect 3384 3720 3390 3732
rect 4065 3723 4123 3729
rect 4065 3720 4077 3723
rect 3384 3692 4077 3720
rect 3384 3680 3390 3692
rect 4065 3689 4077 3692
rect 4111 3689 4123 3723
rect 4065 3683 4123 3689
rect 6549 3723 6607 3729
rect 6549 3689 6561 3723
rect 6595 3720 6607 3723
rect 6638 3720 6644 3732
rect 6595 3692 6644 3720
rect 6595 3689 6607 3692
rect 6549 3683 6607 3689
rect 6638 3680 6644 3692
rect 6696 3680 6702 3732
rect 8478 3720 8484 3732
rect 6932 3692 8484 3720
rect 2406 3612 2412 3664
rect 2464 3652 2470 3664
rect 6932 3652 6960 3692
rect 8478 3680 8484 3692
rect 8536 3720 8542 3732
rect 9493 3723 9551 3729
rect 9493 3720 9505 3723
rect 8536 3692 9505 3720
rect 8536 3680 8542 3692
rect 9493 3689 9505 3692
rect 9539 3689 9551 3723
rect 10134 3720 10140 3732
rect 10095 3692 10140 3720
rect 9493 3683 9551 3689
rect 10134 3680 10140 3692
rect 10192 3720 10198 3732
rect 11057 3723 11115 3729
rect 11057 3720 11069 3723
rect 10192 3692 11069 3720
rect 10192 3680 10198 3692
rect 11057 3689 11069 3692
rect 11103 3689 11115 3723
rect 11422 3720 11428 3732
rect 11383 3692 11428 3720
rect 11057 3683 11115 3689
rect 11422 3680 11428 3692
rect 11480 3680 11486 3732
rect 13170 3720 13176 3732
rect 13131 3692 13176 3720
rect 13170 3680 13176 3692
rect 13228 3680 13234 3732
rect 14090 3680 14096 3732
rect 14148 3720 14154 3732
rect 14185 3723 14243 3729
rect 14185 3720 14197 3723
rect 14148 3692 14197 3720
rect 14148 3680 14154 3692
rect 14185 3689 14197 3692
rect 14231 3689 14243 3723
rect 14185 3683 14243 3689
rect 2464 3624 4108 3652
rect 2464 3612 2470 3624
rect 1486 3584 1492 3596
rect 1447 3556 1492 3584
rect 1486 3544 1492 3556
rect 1544 3544 1550 3596
rect 1756 3587 1814 3593
rect 1756 3553 1768 3587
rect 1802 3584 1814 3587
rect 2866 3584 2872 3596
rect 1802 3556 2872 3584
rect 1802 3553 1814 3556
rect 1756 3547 1814 3553
rect 2866 3544 2872 3556
rect 2924 3544 2930 3596
rect 3142 3584 3148 3596
rect 3103 3556 3148 3584
rect 3142 3544 3148 3556
rect 3200 3544 3206 3596
rect 4080 3584 4108 3624
rect 4264 3624 6960 3652
rect 4264 3584 4292 3624
rect 4080 3556 4292 3584
rect 4338 3544 4344 3596
rect 4396 3584 4402 3596
rect 4433 3587 4491 3593
rect 4433 3584 4445 3587
rect 4396 3556 4445 3584
rect 4396 3544 4402 3556
rect 4433 3553 4445 3556
rect 4479 3553 4491 3587
rect 5166 3584 5172 3596
rect 5127 3556 5172 3584
rect 4433 3547 4491 3553
rect 5166 3544 5172 3556
rect 5224 3544 5230 3596
rect 5436 3587 5494 3593
rect 5436 3553 5448 3587
rect 5482 3584 5494 3587
rect 5902 3584 5908 3596
rect 5482 3556 5908 3584
rect 5482 3553 5494 3556
rect 5436 3547 5494 3553
rect 5902 3544 5908 3556
rect 5960 3584 5966 3596
rect 6362 3584 6368 3596
rect 5960 3556 6368 3584
rect 5960 3544 5966 3556
rect 6362 3544 6368 3556
rect 6420 3544 6426 3596
rect 6932 3584 6960 3624
rect 7006 3612 7012 3664
rect 7064 3652 7070 3664
rect 7064 3624 10180 3652
rect 7064 3612 7070 3624
rect 7193 3587 7251 3593
rect 7193 3584 7205 3587
rect 6932 3556 7205 3584
rect 7193 3553 7205 3556
rect 7239 3553 7251 3587
rect 7193 3547 7251 3553
rect 7285 3587 7343 3593
rect 7285 3553 7297 3587
rect 7331 3584 7343 3587
rect 7374 3584 7380 3596
rect 7331 3556 7380 3584
rect 7331 3553 7343 3556
rect 7285 3547 7343 3553
rect 7374 3544 7380 3556
rect 7432 3544 7438 3596
rect 7558 3544 7564 3596
rect 7616 3584 7622 3596
rect 7929 3587 7987 3593
rect 7929 3584 7941 3587
rect 7616 3556 7941 3584
rect 7616 3544 7622 3556
rect 7929 3553 7941 3556
rect 7975 3553 7987 3587
rect 7929 3547 7987 3553
rect 8196 3587 8254 3593
rect 8196 3553 8208 3587
rect 8242 3584 8254 3587
rect 9214 3584 9220 3596
rect 8242 3556 9220 3584
rect 8242 3553 8254 3556
rect 8196 3547 8254 3553
rect 9214 3544 9220 3556
rect 9272 3584 9278 3596
rect 9490 3584 9496 3596
rect 9272 3556 9496 3584
rect 9272 3544 9278 3556
rect 9490 3544 9496 3556
rect 9548 3544 9554 3596
rect 9585 3587 9643 3593
rect 9585 3553 9597 3587
rect 9631 3584 9643 3587
rect 9674 3584 9680 3596
rect 9631 3556 9680 3584
rect 9631 3553 9643 3556
rect 9585 3547 9643 3553
rect 9674 3544 9680 3556
rect 9732 3584 9738 3596
rect 10042 3584 10048 3596
rect 9732 3556 10048 3584
rect 9732 3544 9738 3556
rect 10042 3544 10048 3556
rect 10100 3544 10106 3596
rect 10152 3584 10180 3624
rect 10962 3612 10968 3664
rect 11020 3652 11026 3664
rect 13265 3655 13323 3661
rect 13265 3652 13277 3655
rect 11020 3624 13277 3652
rect 11020 3612 11026 3624
rect 13265 3621 13277 3624
rect 13311 3621 13323 3655
rect 13265 3615 13323 3621
rect 11977 3587 12035 3593
rect 11977 3584 11989 3587
rect 10152 3556 11989 3584
rect 11977 3553 11989 3556
rect 12023 3553 12035 3587
rect 11977 3547 12035 3553
rect 15289 3587 15347 3593
rect 15289 3553 15301 3587
rect 15335 3584 15347 3587
rect 15470 3584 15476 3596
rect 15335 3556 15476 3584
rect 15335 3553 15347 3556
rect 15289 3547 15347 3553
rect 15470 3544 15476 3556
rect 15528 3544 15534 3596
rect 15841 3587 15899 3593
rect 15841 3553 15853 3587
rect 15887 3553 15899 3587
rect 15841 3547 15899 3553
rect 16761 3587 16819 3593
rect 16761 3553 16773 3587
rect 16807 3584 16819 3587
rect 16850 3584 16856 3596
rect 16807 3556 16856 3584
rect 16807 3553 16819 3556
rect 16761 3547 16819 3553
rect 3418 3516 3424 3528
rect 3379 3488 3424 3516
rect 3418 3476 3424 3488
rect 3476 3476 3482 3528
rect 3602 3476 3608 3528
rect 3660 3516 3666 3528
rect 4525 3519 4583 3525
rect 4525 3516 4537 3519
rect 3660 3488 4537 3516
rect 3660 3476 3666 3488
rect 4525 3485 4537 3488
rect 4571 3485 4583 3519
rect 4525 3479 4583 3485
rect 4617 3519 4675 3525
rect 4617 3485 4629 3519
rect 4663 3485 4675 3519
rect 4617 3479 4675 3485
rect 2498 3408 2504 3460
rect 2556 3448 2562 3460
rect 2869 3451 2927 3457
rect 2869 3448 2881 3451
rect 2556 3420 2881 3448
rect 2556 3408 2562 3420
rect 2869 3417 2881 3420
rect 2915 3448 2927 3451
rect 4632 3448 4660 3479
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 7466 3516 7472 3528
rect 6512 3488 7472 3516
rect 6512 3476 6518 3488
rect 7466 3476 7472 3488
rect 7524 3476 7530 3528
rect 10321 3519 10379 3525
rect 10321 3485 10333 3519
rect 10367 3516 10379 3519
rect 10870 3516 10876 3528
rect 10367 3488 10876 3516
rect 10367 3485 10379 3488
rect 10321 3479 10379 3485
rect 10870 3476 10876 3488
rect 10928 3476 10934 3528
rect 12253 3519 12311 3525
rect 12253 3485 12265 3519
rect 12299 3516 12311 3519
rect 13262 3516 13268 3528
rect 12299 3488 13268 3516
rect 12299 3485 12311 3488
rect 12253 3479 12311 3485
rect 13262 3476 13268 3488
rect 13320 3476 13326 3528
rect 13449 3519 13507 3525
rect 13449 3485 13461 3519
rect 13495 3516 13507 3519
rect 13630 3516 13636 3528
rect 13495 3488 13636 3516
rect 13495 3485 13507 3488
rect 13449 3479 13507 3485
rect 13630 3476 13636 3488
rect 13688 3476 13694 3528
rect 14277 3519 14335 3525
rect 14277 3485 14289 3519
rect 14323 3485 14335 3519
rect 14277 3479 14335 3485
rect 10410 3448 10416 3460
rect 2915 3420 4660 3448
rect 6748 3420 7788 3448
rect 2915 3417 2927 3420
rect 2869 3411 2927 3417
rect 3234 3340 3240 3392
rect 3292 3380 3298 3392
rect 4890 3380 4896 3392
rect 3292 3352 4896 3380
rect 3292 3340 3298 3352
rect 4890 3340 4896 3352
rect 4948 3340 4954 3392
rect 5074 3340 5080 3392
rect 5132 3380 5138 3392
rect 6748 3380 6776 3420
rect 5132 3352 6776 3380
rect 6825 3383 6883 3389
rect 5132 3340 5138 3352
rect 6825 3349 6837 3383
rect 6871 3380 6883 3383
rect 7282 3380 7288 3392
rect 6871 3352 7288 3380
rect 6871 3349 6883 3352
rect 6825 3343 6883 3349
rect 7282 3340 7288 3352
rect 7340 3340 7346 3392
rect 7760 3380 7788 3420
rect 9324 3420 10416 3448
rect 9324 3389 9352 3420
rect 10410 3408 10416 3420
rect 10468 3408 10474 3460
rect 14292 3448 14320 3479
rect 14366 3476 14372 3528
rect 14424 3516 14430 3528
rect 14424 3488 14469 3516
rect 14424 3476 14430 3488
rect 14734 3476 14740 3528
rect 14792 3516 14798 3528
rect 15856 3516 15884 3547
rect 16850 3544 16856 3556
rect 16908 3544 16914 3596
rect 17494 3584 17500 3596
rect 17455 3556 17500 3584
rect 17494 3544 17500 3556
rect 17552 3544 17558 3596
rect 19702 3584 19708 3596
rect 19663 3556 19708 3584
rect 19702 3544 19708 3556
rect 19760 3584 19766 3596
rect 20073 3587 20131 3593
rect 20073 3584 20085 3587
rect 19760 3556 20085 3584
rect 19760 3544 19766 3556
rect 20073 3553 20085 3556
rect 20119 3553 20131 3587
rect 20073 3547 20131 3553
rect 20901 3587 20959 3593
rect 20901 3553 20913 3587
rect 20947 3584 20959 3587
rect 21818 3584 21824 3596
rect 20947 3556 21824 3584
rect 20947 3553 20959 3556
rect 20901 3547 20959 3553
rect 21818 3544 21824 3556
rect 21876 3544 21882 3596
rect 14792 3488 15884 3516
rect 17037 3519 17095 3525
rect 14792 3476 14798 3488
rect 17037 3485 17049 3519
rect 17083 3516 17095 3519
rect 18046 3516 18052 3528
rect 17083 3488 18052 3516
rect 17083 3485 17095 3488
rect 17037 3479 17095 3485
rect 18046 3476 18052 3488
rect 18104 3476 18110 3528
rect 14829 3451 14887 3457
rect 14829 3448 14841 3451
rect 10520 3420 14841 3448
rect 9309 3383 9367 3389
rect 9309 3380 9321 3383
rect 7760 3352 9321 3380
rect 9309 3349 9321 3352
rect 9355 3349 9367 3383
rect 9674 3380 9680 3392
rect 9635 3352 9680 3380
rect 9309 3343 9367 3349
rect 9674 3340 9680 3352
rect 9732 3340 9738 3392
rect 10042 3340 10048 3392
rect 10100 3380 10106 3392
rect 10520 3380 10548 3420
rect 14829 3417 14841 3420
rect 14875 3417 14887 3451
rect 14829 3411 14887 3417
rect 10686 3380 10692 3392
rect 10100 3352 10548 3380
rect 10647 3352 10692 3380
rect 10100 3340 10106 3352
rect 10686 3340 10692 3352
rect 10744 3340 10750 3392
rect 12805 3383 12863 3389
rect 12805 3349 12817 3383
rect 12851 3380 12863 3383
rect 13722 3380 13728 3392
rect 12851 3352 13728 3380
rect 12851 3349 12863 3352
rect 12805 3343 12863 3349
rect 13722 3340 13728 3352
rect 13780 3340 13786 3392
rect 13814 3340 13820 3392
rect 13872 3380 13878 3392
rect 15473 3383 15531 3389
rect 13872 3352 13917 3380
rect 13872 3340 13878 3352
rect 15473 3349 15485 3383
rect 15519 3380 15531 3383
rect 15654 3380 15660 3392
rect 15519 3352 15660 3380
rect 15519 3349 15531 3352
rect 15473 3343 15531 3349
rect 15654 3340 15660 3352
rect 15712 3340 15718 3392
rect 16025 3383 16083 3389
rect 16025 3349 16037 3383
rect 16071 3380 16083 3383
rect 16482 3380 16488 3392
rect 16071 3352 16488 3380
rect 16071 3349 16083 3352
rect 16025 3343 16083 3349
rect 16482 3340 16488 3352
rect 16540 3340 16546 3392
rect 17681 3383 17739 3389
rect 17681 3349 17693 3383
rect 17727 3380 17739 3383
rect 18138 3380 18144 3392
rect 17727 3352 18144 3380
rect 17727 3349 17739 3352
rect 17681 3343 17739 3349
rect 18138 3340 18144 3352
rect 18196 3340 18202 3392
rect 20257 3383 20315 3389
rect 20257 3349 20269 3383
rect 20303 3380 20315 3383
rect 20898 3380 20904 3392
rect 20303 3352 20904 3380
rect 20303 3349 20315 3352
rect 20257 3343 20315 3349
rect 20898 3340 20904 3352
rect 20956 3340 20962 3392
rect 21085 3383 21143 3389
rect 21085 3349 21097 3383
rect 21131 3380 21143 3383
rect 22278 3380 22284 3392
rect 21131 3352 22284 3380
rect 21131 3349 21143 3352
rect 21085 3343 21143 3349
rect 22278 3340 22284 3352
rect 22336 3340 22342 3392
rect 1104 3290 21896 3312
rect 1104 3238 4447 3290
rect 4499 3238 4511 3290
rect 4563 3238 4575 3290
rect 4627 3238 4639 3290
rect 4691 3238 11378 3290
rect 11430 3238 11442 3290
rect 11494 3238 11506 3290
rect 11558 3238 11570 3290
rect 11622 3238 18308 3290
rect 18360 3238 18372 3290
rect 18424 3238 18436 3290
rect 18488 3238 18500 3290
rect 18552 3238 21896 3290
rect 1104 3216 21896 3238
rect 2317 3179 2375 3185
rect 2317 3145 2329 3179
rect 2363 3176 2375 3179
rect 3602 3176 3608 3188
rect 2363 3148 3608 3176
rect 2363 3145 2375 3148
rect 2317 3139 2375 3145
rect 3602 3136 3608 3148
rect 3660 3136 3666 3188
rect 5166 3176 5172 3188
rect 5000 3148 5172 3176
rect 1946 3068 1952 3120
rect 2004 3108 2010 3120
rect 2004 3080 2268 3108
rect 2004 3068 2010 3080
rect 198 2932 204 2984
rect 256 2972 262 2984
rect 1302 2972 1308 2984
rect 256 2944 1308 2972
rect 256 2932 262 2944
rect 1302 2932 1308 2944
rect 1360 2972 1366 2984
rect 1949 2975 2007 2981
rect 1949 2972 1961 2975
rect 1360 2944 1961 2972
rect 1360 2932 1366 2944
rect 1949 2941 1961 2944
rect 1995 2972 2007 2975
rect 2133 2975 2191 2981
rect 2133 2972 2145 2975
rect 1995 2944 2145 2972
rect 1995 2941 2007 2944
rect 1949 2935 2007 2941
rect 2133 2941 2145 2944
rect 2179 2941 2191 2975
rect 2240 2972 2268 3080
rect 2866 3040 2872 3052
rect 2827 3012 2872 3040
rect 2866 3000 2872 3012
rect 2924 3000 2930 3052
rect 5000 3049 5028 3148
rect 5166 3136 5172 3148
rect 5224 3136 5230 3188
rect 9490 3136 9496 3188
rect 9548 3176 9554 3188
rect 10137 3179 10195 3185
rect 10137 3176 10149 3179
rect 9548 3148 10149 3176
rect 9548 3136 9554 3148
rect 10137 3145 10149 3148
rect 10183 3145 10195 3179
rect 10137 3139 10195 3145
rect 10318 3136 10324 3188
rect 10376 3176 10382 3188
rect 12250 3176 12256 3188
rect 10376 3148 12256 3176
rect 10376 3136 10382 3148
rect 12250 3136 12256 3148
rect 12308 3136 12314 3188
rect 13814 3136 13820 3188
rect 13872 3176 13878 3188
rect 13872 3148 15700 3176
rect 13872 3136 13878 3148
rect 15197 3111 15255 3117
rect 15197 3077 15209 3111
rect 15243 3077 15255 3111
rect 15197 3071 15255 3077
rect 4985 3043 5043 3049
rect 4985 3009 4997 3043
rect 5031 3009 5043 3043
rect 7466 3040 7472 3052
rect 7427 3012 7472 3040
rect 4985 3003 5043 3009
rect 7466 3000 7472 3012
rect 7524 3000 7530 3052
rect 7558 3000 7564 3052
rect 7616 3040 7622 3052
rect 8757 3043 8815 3049
rect 8757 3040 8769 3043
rect 7616 3012 8769 3040
rect 7616 3000 7622 3012
rect 8757 3009 8769 3012
rect 8803 3009 8815 3043
rect 10870 3040 10876 3052
rect 8757 3003 8815 3009
rect 9784 3012 10876 3040
rect 3329 2975 3387 2981
rect 3329 2972 3341 2975
rect 2240 2944 3341 2972
rect 2133 2935 2191 2941
rect 3329 2941 3341 2944
rect 3375 2941 3387 2975
rect 3329 2935 3387 2941
rect 3596 2975 3654 2981
rect 3596 2941 3608 2975
rect 3642 2972 3654 2975
rect 5074 2972 5080 2984
rect 3642 2944 5080 2972
rect 3642 2941 3654 2944
rect 3596 2935 3654 2941
rect 5074 2932 5080 2944
rect 5132 2932 5138 2984
rect 5252 2975 5310 2981
rect 5252 2941 5264 2975
rect 5298 2972 5310 2975
rect 5534 2972 5540 2984
rect 5298 2944 5540 2972
rect 5298 2941 5310 2944
rect 5252 2935 5310 2941
rect 5534 2932 5540 2944
rect 5592 2932 5598 2984
rect 8113 2975 8171 2981
rect 8113 2941 8125 2975
rect 8159 2972 8171 2975
rect 9024 2975 9082 2981
rect 8159 2944 8524 2972
rect 8159 2941 8171 2944
rect 8113 2935 8171 2941
rect 2685 2907 2743 2913
rect 2685 2904 2697 2907
rect 1596 2876 2697 2904
rect 1026 2796 1032 2848
rect 1084 2836 1090 2848
rect 1596 2845 1624 2876
rect 2685 2873 2697 2876
rect 2731 2904 2743 2907
rect 6086 2904 6092 2916
rect 2731 2876 6092 2904
rect 2731 2873 2743 2876
rect 2685 2867 2743 2873
rect 6086 2864 6092 2876
rect 6144 2864 6150 2916
rect 7006 2864 7012 2916
rect 7064 2904 7070 2916
rect 7285 2907 7343 2913
rect 7285 2904 7297 2907
rect 7064 2876 7297 2904
rect 7064 2864 7070 2876
rect 7285 2873 7297 2876
rect 7331 2873 7343 2907
rect 7285 2867 7343 2873
rect 7377 2907 7435 2913
rect 7377 2873 7389 2907
rect 7423 2904 7435 2907
rect 8386 2904 8392 2916
rect 7423 2876 8392 2904
rect 7423 2873 7435 2876
rect 7377 2867 7435 2873
rect 1581 2839 1639 2845
rect 1581 2836 1593 2839
rect 1084 2808 1593 2836
rect 1084 2796 1090 2808
rect 1581 2805 1593 2808
rect 1627 2805 1639 2839
rect 1581 2799 1639 2805
rect 2133 2839 2191 2845
rect 2133 2805 2145 2839
rect 2179 2836 2191 2839
rect 2777 2839 2835 2845
rect 2777 2836 2789 2839
rect 2179 2808 2789 2836
rect 2179 2805 2191 2808
rect 2133 2799 2191 2805
rect 2777 2805 2789 2808
rect 2823 2805 2835 2839
rect 2777 2799 2835 2805
rect 2866 2796 2872 2848
rect 2924 2836 2930 2848
rect 4709 2839 4767 2845
rect 4709 2836 4721 2839
rect 2924 2808 4721 2836
rect 2924 2796 2930 2808
rect 4709 2805 4721 2808
rect 4755 2805 4767 2839
rect 6362 2836 6368 2848
rect 6275 2808 6368 2836
rect 4709 2799 4767 2805
rect 6362 2796 6368 2808
rect 6420 2836 6426 2848
rect 6822 2836 6828 2848
rect 6420 2808 6828 2836
rect 6420 2796 6426 2808
rect 6822 2796 6828 2808
rect 6880 2796 6886 2848
rect 6917 2839 6975 2845
rect 6917 2805 6929 2839
rect 6963 2836 6975 2839
rect 7190 2836 7196 2848
rect 6963 2808 7196 2836
rect 6963 2805 6975 2808
rect 6917 2799 6975 2805
rect 7190 2796 7196 2808
rect 7248 2796 7254 2848
rect 7300 2836 7328 2867
rect 8386 2864 8392 2876
rect 8444 2864 8450 2916
rect 8496 2904 8524 2944
rect 9024 2941 9036 2975
rect 9070 2972 9082 2975
rect 9784 2972 9812 3012
rect 10870 3000 10876 3012
rect 10928 3040 10934 3052
rect 10965 3043 11023 3049
rect 10965 3040 10977 3043
rect 10928 3012 10977 3040
rect 10928 3000 10934 3012
rect 10965 3009 10977 3012
rect 11011 3009 11023 3043
rect 10965 3003 11023 3009
rect 13722 3000 13728 3052
rect 13780 3040 13786 3052
rect 14734 3040 14740 3052
rect 13780 3012 14504 3040
rect 14695 3012 14740 3040
rect 13780 3000 13786 3012
rect 9070 2944 9812 2972
rect 9070 2941 9082 2944
rect 9024 2935 9082 2941
rect 9858 2932 9864 2984
rect 9916 2972 9922 2984
rect 11425 2975 11483 2981
rect 11425 2972 11437 2975
rect 9916 2944 11437 2972
rect 9916 2932 9922 2944
rect 11425 2941 11437 2944
rect 11471 2941 11483 2975
rect 11425 2935 11483 2941
rect 12434 2932 12440 2984
rect 12492 2972 12498 2984
rect 12492 2944 12537 2972
rect 12492 2932 12498 2944
rect 12802 2932 12808 2984
rect 12860 2972 12866 2984
rect 13173 2975 13231 2981
rect 13173 2972 13185 2975
rect 12860 2944 13185 2972
rect 12860 2932 12866 2944
rect 13173 2941 13185 2944
rect 13219 2941 13231 2975
rect 13173 2935 13231 2941
rect 13262 2932 13268 2984
rect 13320 2972 13326 2984
rect 14476 2981 14504 3012
rect 14734 3000 14740 3012
rect 14792 3000 14798 3052
rect 13909 2975 13967 2981
rect 13909 2972 13921 2975
rect 13320 2944 13921 2972
rect 13320 2932 13326 2944
rect 13909 2941 13921 2944
rect 13955 2941 13967 2975
rect 13909 2935 13967 2941
rect 14461 2975 14519 2981
rect 14461 2941 14473 2975
rect 14507 2941 14519 2975
rect 15212 2972 15240 3071
rect 15672 3049 15700 3148
rect 15657 3043 15715 3049
rect 15657 3009 15669 3043
rect 15703 3009 15715 3043
rect 15838 3040 15844 3052
rect 15799 3012 15844 3040
rect 15657 3003 15715 3009
rect 15838 3000 15844 3012
rect 15896 3000 15902 3052
rect 20714 3040 20720 3052
rect 20675 3012 20720 3040
rect 20714 3000 20720 3012
rect 20772 3000 20778 3052
rect 16209 2975 16267 2981
rect 16209 2972 16221 2975
rect 15212 2944 16221 2972
rect 14461 2935 14519 2941
rect 16209 2941 16221 2944
rect 16255 2941 16267 2975
rect 16942 2972 16948 2984
rect 16903 2944 16948 2972
rect 16209 2935 16267 2941
rect 16942 2932 16948 2944
rect 17000 2932 17006 2984
rect 18046 2972 18052 2984
rect 18007 2944 18052 2972
rect 18046 2932 18052 2944
rect 18104 2932 18110 2984
rect 18598 2972 18604 2984
rect 18559 2944 18604 2972
rect 18598 2932 18604 2944
rect 18656 2932 18662 2984
rect 20533 2975 20591 2981
rect 20533 2941 20545 2975
rect 20579 2972 20591 2975
rect 21358 2972 21364 2984
rect 20579 2944 21364 2972
rect 20579 2941 20591 2944
rect 20533 2935 20591 2941
rect 21358 2932 21364 2944
rect 21416 2932 21422 2984
rect 10686 2904 10692 2916
rect 8496 2876 10692 2904
rect 10686 2864 10692 2876
rect 10744 2904 10750 2916
rect 10781 2907 10839 2913
rect 10781 2904 10793 2907
rect 10744 2876 10793 2904
rect 10744 2864 10750 2876
rect 10781 2873 10793 2876
rect 10827 2873 10839 2907
rect 10781 2867 10839 2873
rect 11701 2907 11759 2913
rect 11701 2873 11713 2907
rect 11747 2904 11759 2907
rect 11882 2904 11888 2916
rect 11747 2876 11888 2904
rect 11747 2873 11759 2876
rect 11701 2867 11759 2873
rect 11882 2864 11888 2876
rect 11940 2864 11946 2916
rect 12710 2904 12716 2916
rect 12671 2876 12716 2904
rect 12710 2864 12716 2876
rect 12768 2864 12774 2916
rect 13449 2907 13507 2913
rect 13449 2873 13461 2907
rect 13495 2904 13507 2907
rect 13722 2904 13728 2916
rect 13495 2876 13728 2904
rect 13495 2873 13507 2876
rect 13449 2867 13507 2873
rect 13722 2864 13728 2876
rect 13780 2864 13786 2916
rect 15565 2907 15623 2913
rect 15565 2873 15577 2907
rect 15611 2904 15623 2907
rect 15611 2876 16344 2904
rect 15611 2873 15623 2876
rect 15565 2867 15623 2873
rect 7929 2839 7987 2845
rect 7929 2836 7941 2839
rect 7300 2808 7941 2836
rect 7929 2805 7941 2808
rect 7975 2836 7987 2839
rect 8113 2839 8171 2845
rect 8113 2836 8125 2839
rect 7975 2808 8125 2836
rect 7975 2805 7987 2808
rect 7929 2799 7987 2805
rect 8113 2805 8125 2808
rect 8159 2805 8171 2839
rect 8294 2836 8300 2848
rect 8255 2808 8300 2836
rect 8113 2799 8171 2805
rect 8294 2796 8300 2808
rect 8352 2796 8358 2848
rect 10410 2836 10416 2848
rect 10371 2808 10416 2836
rect 10410 2796 10416 2808
rect 10468 2796 10474 2848
rect 10870 2836 10876 2848
rect 10831 2808 10876 2836
rect 10870 2796 10876 2808
rect 10928 2836 10934 2848
rect 12158 2836 12164 2848
rect 10928 2808 12164 2836
rect 10928 2796 10934 2808
rect 12158 2796 12164 2808
rect 12216 2796 12222 2848
rect 13906 2796 13912 2848
rect 13964 2836 13970 2848
rect 14093 2839 14151 2845
rect 14093 2836 14105 2839
rect 13964 2808 14105 2836
rect 13964 2796 13970 2808
rect 14093 2805 14105 2808
rect 14139 2805 14151 2839
rect 16316 2836 16344 2876
rect 16390 2864 16396 2916
rect 16448 2904 16454 2916
rect 16485 2907 16543 2913
rect 16485 2904 16497 2907
rect 16448 2876 16497 2904
rect 16448 2864 16454 2876
rect 16485 2873 16497 2876
rect 16531 2873 16543 2907
rect 16485 2867 16543 2873
rect 17221 2907 17279 2913
rect 17221 2873 17233 2907
rect 17267 2904 17279 2907
rect 17402 2904 17408 2916
rect 17267 2876 17408 2904
rect 17267 2873 17279 2876
rect 17221 2867 17279 2873
rect 17402 2864 17408 2876
rect 17460 2864 17466 2916
rect 16942 2836 16948 2848
rect 16316 2808 16948 2836
rect 14093 2799 14151 2805
rect 16942 2796 16948 2808
rect 17000 2796 17006 2848
rect 17494 2796 17500 2848
rect 17552 2836 17558 2848
rect 18233 2839 18291 2845
rect 18233 2836 18245 2839
rect 17552 2808 18245 2836
rect 17552 2796 17558 2808
rect 18233 2805 18245 2808
rect 18279 2805 18291 2839
rect 18233 2799 18291 2805
rect 18690 2796 18696 2848
rect 18748 2836 18754 2848
rect 18785 2839 18843 2845
rect 18785 2836 18797 2839
rect 18748 2808 18797 2836
rect 18748 2796 18754 2808
rect 18785 2805 18797 2808
rect 18831 2805 18843 2839
rect 18785 2799 18843 2805
rect 1104 2746 21896 2768
rect 1104 2694 7912 2746
rect 7964 2694 7976 2746
rect 8028 2694 8040 2746
rect 8092 2694 8104 2746
rect 8156 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 15035 2746
rect 15087 2694 21896 2746
rect 1104 2672 21896 2694
rect 2777 2635 2835 2641
rect 2777 2601 2789 2635
rect 2823 2632 2835 2635
rect 4338 2632 4344 2644
rect 2823 2604 4344 2632
rect 2823 2601 2835 2604
rect 2777 2595 2835 2601
rect 4338 2592 4344 2604
rect 4396 2592 4402 2644
rect 5813 2635 5871 2641
rect 5813 2601 5825 2635
rect 5859 2601 5871 2635
rect 6178 2632 6184 2644
rect 6139 2604 6184 2632
rect 5813 2595 5871 2601
rect 2774 2456 2780 2508
rect 2832 2496 2838 2508
rect 3145 2499 3203 2505
rect 3145 2496 3157 2499
rect 2832 2468 3157 2496
rect 2832 2456 2838 2468
rect 3145 2465 3157 2468
rect 3191 2496 3203 2499
rect 3970 2496 3976 2508
rect 3191 2468 3976 2496
rect 3191 2465 3203 2468
rect 3145 2459 3203 2465
rect 3970 2456 3976 2468
rect 4028 2496 4034 2508
rect 4065 2499 4123 2505
rect 4065 2496 4077 2499
rect 4028 2468 4077 2496
rect 4028 2456 4034 2468
rect 4065 2465 4077 2468
rect 4111 2465 4123 2499
rect 5828 2496 5856 2595
rect 6178 2592 6184 2604
rect 6236 2592 6242 2644
rect 6273 2635 6331 2641
rect 6273 2601 6285 2635
rect 6319 2632 6331 2635
rect 6917 2635 6975 2641
rect 6917 2632 6929 2635
rect 6319 2604 6929 2632
rect 6319 2601 6331 2604
rect 6273 2595 6331 2601
rect 6917 2601 6929 2604
rect 6963 2601 6975 2635
rect 7282 2632 7288 2644
rect 7243 2604 7288 2632
rect 6917 2595 6975 2601
rect 7282 2592 7288 2604
rect 7340 2592 7346 2644
rect 8386 2632 8392 2644
rect 8347 2604 8392 2632
rect 8386 2592 8392 2604
rect 8444 2592 8450 2644
rect 9122 2632 9128 2644
rect 9083 2604 9128 2632
rect 9122 2592 9128 2604
rect 9180 2592 9186 2644
rect 9766 2632 9772 2644
rect 9727 2604 9772 2632
rect 9766 2592 9772 2604
rect 9824 2592 9830 2644
rect 10229 2635 10287 2641
rect 10229 2601 10241 2635
rect 10275 2632 10287 2635
rect 10410 2632 10416 2644
rect 10275 2604 10416 2632
rect 10275 2601 10287 2604
rect 10229 2595 10287 2601
rect 10410 2592 10416 2604
rect 10468 2592 10474 2644
rect 16942 2632 16948 2644
rect 16903 2604 16948 2632
rect 16942 2592 16948 2604
rect 17000 2592 17006 2644
rect 7190 2524 7196 2576
rect 7248 2564 7254 2576
rect 7377 2567 7435 2573
rect 7377 2564 7389 2567
rect 7248 2536 7389 2564
rect 7248 2524 7254 2536
rect 7377 2533 7389 2536
rect 7423 2533 7435 2567
rect 7377 2527 7435 2533
rect 8294 2524 8300 2576
rect 8352 2564 8358 2576
rect 9033 2567 9091 2573
rect 9033 2564 9045 2567
rect 8352 2536 9045 2564
rect 8352 2524 8358 2536
rect 9033 2533 9045 2536
rect 9079 2533 9091 2567
rect 9033 2527 9091 2533
rect 9674 2524 9680 2576
rect 9732 2564 9738 2576
rect 10137 2567 10195 2573
rect 10137 2564 10149 2567
rect 9732 2536 10149 2564
rect 9732 2524 9738 2536
rect 10137 2533 10149 2536
rect 10183 2533 10195 2567
rect 12434 2564 12440 2576
rect 10137 2527 10195 2533
rect 10244 2536 12440 2564
rect 10244 2496 10272 2536
rect 12434 2524 12440 2536
rect 12492 2524 12498 2576
rect 11882 2496 11888 2508
rect 5828 2468 10272 2496
rect 11843 2468 11888 2496
rect 4065 2459 4123 2465
rect 11882 2456 11888 2468
rect 11940 2456 11946 2508
rect 12618 2496 12624 2508
rect 12579 2468 12624 2496
rect 12618 2456 12624 2468
rect 12676 2456 12682 2508
rect 12710 2456 12716 2508
rect 12768 2496 12774 2508
rect 13173 2499 13231 2505
rect 13173 2496 13185 2499
rect 12768 2468 13185 2496
rect 12768 2456 12774 2468
rect 13173 2465 13185 2468
rect 13219 2465 13231 2499
rect 13722 2496 13728 2508
rect 13683 2468 13728 2496
rect 13173 2459 13231 2465
rect 13722 2456 13728 2468
rect 13780 2456 13786 2508
rect 14277 2499 14335 2505
rect 14277 2465 14289 2499
rect 14323 2496 14335 2499
rect 14458 2496 14464 2508
rect 14323 2468 14464 2496
rect 14323 2465 14335 2468
rect 14277 2459 14335 2465
rect 14458 2456 14464 2468
rect 14516 2456 14522 2508
rect 14829 2499 14887 2505
rect 14829 2465 14841 2499
rect 14875 2496 14887 2499
rect 15286 2496 15292 2508
rect 14875 2468 15292 2496
rect 14875 2465 14887 2468
rect 14829 2459 14887 2465
rect 15286 2456 15292 2468
rect 15344 2456 15350 2508
rect 15378 2456 15384 2508
rect 15436 2496 15442 2508
rect 15473 2499 15531 2505
rect 15473 2496 15485 2499
rect 15436 2468 15485 2496
rect 15436 2456 15442 2468
rect 15473 2465 15485 2468
rect 15519 2465 15531 2499
rect 16390 2496 16396 2508
rect 16351 2468 16396 2496
rect 15473 2459 15531 2465
rect 16390 2456 16396 2468
rect 16448 2456 16454 2508
rect 17402 2496 17408 2508
rect 17363 2468 17408 2496
rect 17402 2456 17408 2468
rect 17460 2456 17466 2508
rect 3237 2431 3295 2437
rect 3237 2428 3249 2431
rect 3068 2400 3249 2428
rect 3068 2360 3096 2400
rect 3237 2397 3249 2400
rect 3283 2397 3295 2431
rect 3418 2428 3424 2440
rect 3379 2400 3424 2428
rect 3237 2391 3295 2397
rect 2424 2332 3096 2360
rect 3252 2360 3280 2391
rect 3418 2388 3424 2400
rect 3476 2388 3482 2440
rect 6457 2431 6515 2437
rect 6457 2397 6469 2431
rect 6503 2428 6515 2431
rect 6638 2428 6644 2440
rect 6503 2400 6644 2428
rect 6503 2397 6515 2400
rect 6457 2391 6515 2397
rect 6638 2388 6644 2400
rect 6696 2388 6702 2440
rect 6822 2388 6828 2440
rect 6880 2428 6886 2440
rect 7469 2431 7527 2437
rect 7469 2428 7481 2431
rect 6880 2400 7481 2428
rect 6880 2388 6886 2400
rect 7469 2397 7481 2400
rect 7515 2397 7527 2431
rect 7469 2391 7527 2397
rect 9214 2388 9220 2440
rect 9272 2428 9278 2440
rect 9309 2431 9367 2437
rect 9309 2428 9321 2431
rect 9272 2400 9321 2428
rect 9272 2388 9278 2400
rect 9309 2397 9321 2400
rect 9355 2428 9367 2431
rect 10321 2431 10379 2437
rect 10321 2428 10333 2431
rect 9355 2400 10333 2428
rect 9355 2397 9367 2400
rect 9309 2391 9367 2397
rect 10321 2397 10333 2400
rect 10367 2397 10379 2431
rect 10321 2391 10379 2397
rect 6914 2360 6920 2372
rect 3252 2332 6920 2360
rect 1946 2252 1952 2304
rect 2004 2292 2010 2304
rect 2424 2301 2452 2332
rect 6914 2320 6920 2332
rect 6972 2320 6978 2372
rect 8665 2363 8723 2369
rect 8665 2329 8677 2363
rect 8711 2360 8723 2363
rect 10226 2360 10232 2372
rect 8711 2332 10232 2360
rect 8711 2329 8723 2332
rect 8665 2323 8723 2329
rect 10226 2320 10232 2332
rect 10284 2320 10290 2372
rect 2409 2295 2467 2301
rect 2409 2292 2421 2295
rect 2004 2264 2421 2292
rect 2004 2252 2010 2264
rect 2409 2261 2421 2264
rect 2455 2261 2467 2295
rect 2409 2255 2467 2261
rect 6730 2252 6736 2304
rect 6788 2292 6794 2304
rect 7190 2292 7196 2304
rect 6788 2264 7196 2292
rect 6788 2252 6794 2264
rect 7190 2252 7196 2264
rect 7248 2252 7254 2304
rect 7926 2292 7932 2304
rect 7887 2264 7932 2292
rect 7926 2252 7932 2264
rect 7984 2252 7990 2304
rect 8386 2252 8392 2304
rect 8444 2292 8450 2304
rect 10870 2292 10876 2304
rect 8444 2264 10876 2292
rect 8444 2252 8450 2264
rect 10870 2252 10876 2264
rect 10928 2292 10934 2304
rect 11241 2295 11299 2301
rect 11241 2292 11253 2295
rect 10928 2264 11253 2292
rect 10928 2252 10934 2264
rect 11241 2261 11253 2264
rect 11287 2261 11299 2295
rect 11241 2255 11299 2261
rect 12069 2295 12127 2301
rect 12069 2261 12081 2295
rect 12115 2292 12127 2295
rect 12526 2292 12532 2304
rect 12115 2264 12532 2292
rect 12115 2261 12127 2264
rect 12069 2255 12127 2261
rect 12526 2252 12532 2264
rect 12584 2252 12590 2304
rect 12805 2295 12863 2301
rect 12805 2261 12817 2295
rect 12851 2292 12863 2295
rect 12986 2292 12992 2304
rect 12851 2264 12992 2292
rect 12851 2261 12863 2264
rect 12805 2255 12863 2261
rect 12986 2252 12992 2264
rect 13044 2252 13050 2304
rect 13357 2295 13415 2301
rect 13357 2261 13369 2295
rect 13403 2292 13415 2295
rect 13446 2292 13452 2304
rect 13403 2264 13452 2292
rect 13403 2261 13415 2264
rect 13357 2255 13415 2261
rect 13446 2252 13452 2264
rect 13504 2252 13510 2304
rect 13909 2295 13967 2301
rect 13909 2261 13921 2295
rect 13955 2292 13967 2295
rect 14274 2292 14280 2304
rect 13955 2264 14280 2292
rect 13955 2261 13967 2264
rect 13909 2255 13967 2261
rect 14274 2252 14280 2264
rect 14332 2252 14338 2304
rect 14461 2295 14519 2301
rect 14461 2261 14473 2295
rect 14507 2292 14519 2295
rect 14734 2292 14740 2304
rect 14507 2264 14740 2292
rect 14507 2261 14519 2264
rect 14461 2255 14519 2261
rect 14734 2252 14740 2264
rect 14792 2252 14798 2304
rect 15013 2295 15071 2301
rect 15013 2261 15025 2295
rect 15059 2292 15071 2295
rect 15194 2292 15200 2304
rect 15059 2264 15200 2292
rect 15059 2261 15071 2264
rect 15013 2255 15071 2261
rect 15194 2252 15200 2264
rect 15252 2252 15258 2304
rect 15657 2295 15715 2301
rect 15657 2261 15669 2295
rect 15703 2292 15715 2295
rect 16114 2292 16120 2304
rect 15703 2264 16120 2292
rect 15703 2261 15715 2264
rect 15657 2255 15715 2261
rect 16114 2252 16120 2264
rect 16172 2252 16178 2304
rect 16577 2295 16635 2301
rect 16577 2261 16589 2295
rect 16623 2292 16635 2295
rect 16942 2292 16948 2304
rect 16623 2264 16948 2292
rect 16623 2261 16635 2264
rect 16577 2255 16635 2261
rect 16942 2252 16948 2264
rect 17000 2252 17006 2304
rect 17589 2295 17647 2301
rect 17589 2261 17601 2295
rect 17635 2292 17647 2295
rect 17862 2292 17868 2304
rect 17635 2264 17868 2292
rect 17635 2261 17647 2264
rect 17589 2255 17647 2261
rect 17862 2252 17868 2264
rect 17920 2252 17926 2304
rect 21358 2292 21364 2304
rect 21271 2264 21364 2292
rect 21358 2252 21364 2264
rect 21416 2292 21422 2304
rect 22738 2292 22744 2304
rect 21416 2264 22744 2292
rect 21416 2252 21422 2264
rect 22738 2252 22744 2264
rect 22796 2252 22802 2304
rect 1104 2202 21896 2224
rect 1104 2150 4447 2202
rect 4499 2150 4511 2202
rect 4563 2150 4575 2202
rect 4627 2150 4639 2202
rect 4691 2150 11378 2202
rect 11430 2150 11442 2202
rect 11494 2150 11506 2202
rect 11558 2150 11570 2202
rect 11622 2150 18308 2202
rect 18360 2150 18372 2202
rect 18424 2150 18436 2202
rect 18488 2150 18500 2202
rect 18552 2150 21896 2202
rect 1104 2128 21896 2150
rect 1486 2048 1492 2100
rect 1544 2088 1550 2100
rect 7374 2088 7380 2100
rect 1544 2060 7380 2088
rect 1544 2048 1550 2060
rect 7374 2048 7380 2060
rect 7432 2088 7438 2100
rect 7926 2088 7932 2100
rect 7432 2060 7932 2088
rect 7432 2048 7438 2060
rect 7926 2048 7932 2060
rect 7984 2048 7990 2100
rect 566 1980 572 2032
rect 624 2020 630 2032
rect 7006 2020 7012 2032
rect 624 1992 7012 2020
rect 624 1980 630 1992
rect 7006 1980 7012 1992
rect 7064 1980 7070 2032
<< via1 >>
rect 3700 21768 3752 21820
rect 10784 21768 10836 21820
rect 4447 20646 4499 20698
rect 4511 20646 4563 20698
rect 4575 20646 4627 20698
rect 4639 20646 4691 20698
rect 11378 20646 11430 20698
rect 11442 20646 11494 20698
rect 11506 20646 11558 20698
rect 11570 20646 11622 20698
rect 18308 20646 18360 20698
rect 18372 20646 18424 20698
rect 18436 20646 18488 20698
rect 18500 20646 18552 20698
rect 1952 20587 2004 20596
rect 1952 20553 1961 20587
rect 1961 20553 1995 20587
rect 1995 20553 2004 20587
rect 1952 20544 2004 20553
rect 2780 20544 2832 20596
rect 2596 20340 2648 20392
rect 3240 20272 3292 20324
rect 7912 20102 7964 20154
rect 7976 20102 8028 20154
rect 8040 20102 8092 20154
rect 8104 20102 8156 20154
rect 14843 20102 14895 20154
rect 14907 20102 14959 20154
rect 14971 20102 15023 20154
rect 15035 20102 15087 20154
rect 2780 20000 2832 20052
rect 3148 20043 3200 20052
rect 3148 20009 3157 20043
rect 3157 20009 3191 20043
rect 3191 20009 3200 20043
rect 3148 20000 3200 20009
rect 2504 19864 2556 19916
rect 2964 19907 3016 19916
rect 2964 19873 2973 19907
rect 2973 19873 3007 19907
rect 3007 19873 3016 19907
rect 2964 19864 3016 19873
rect 2780 19796 2832 19848
rect 2044 19771 2096 19780
rect 2044 19737 2053 19771
rect 2053 19737 2087 19771
rect 2087 19737 2096 19771
rect 2044 19728 2096 19737
rect 4447 19558 4499 19610
rect 4511 19558 4563 19610
rect 4575 19558 4627 19610
rect 4639 19558 4691 19610
rect 11378 19558 11430 19610
rect 11442 19558 11494 19610
rect 11506 19558 11558 19610
rect 11570 19558 11622 19610
rect 18308 19558 18360 19610
rect 18372 19558 18424 19610
rect 18436 19558 18488 19610
rect 18500 19558 18552 19610
rect 1952 19431 2004 19440
rect 1952 19397 1961 19431
rect 1961 19397 1995 19431
rect 1995 19397 2004 19431
rect 1952 19388 2004 19397
rect 2504 19363 2556 19372
rect 2504 19329 2513 19363
rect 2513 19329 2547 19363
rect 2547 19329 2556 19363
rect 2504 19320 2556 19329
rect 3240 19363 3292 19372
rect 3240 19329 3249 19363
rect 3249 19329 3283 19363
rect 3283 19329 3292 19363
rect 3240 19320 3292 19329
rect 8944 19252 8996 19304
rect 3240 19184 3292 19236
rect 10600 19116 10652 19168
rect 7912 19014 7964 19066
rect 7976 19014 8028 19066
rect 8040 19014 8092 19066
rect 8104 19014 8156 19066
rect 14843 19014 14895 19066
rect 14907 19014 14959 19066
rect 14971 19014 15023 19066
rect 15035 19014 15087 19066
rect 1952 18955 2004 18964
rect 1952 18921 1961 18955
rect 1961 18921 1995 18955
rect 1995 18921 2004 18955
rect 1952 18912 2004 18921
rect 10784 18955 10836 18964
rect 10784 18921 10793 18955
rect 10793 18921 10827 18955
rect 10827 18921 10836 18955
rect 10784 18912 10836 18921
rect 2596 18887 2648 18896
rect 2596 18853 2605 18887
rect 2605 18853 2639 18887
rect 2639 18853 2648 18887
rect 2596 18844 2648 18853
rect 2964 18844 3016 18896
rect 1768 18819 1820 18828
rect 1768 18785 1777 18819
rect 1777 18785 1811 18819
rect 1811 18785 1820 18819
rect 1768 18776 1820 18785
rect 9680 18776 9732 18828
rect 11060 18776 11112 18828
rect 5632 18708 5684 18760
rect 4447 18470 4499 18522
rect 4511 18470 4563 18522
rect 4575 18470 4627 18522
rect 4639 18470 4691 18522
rect 11378 18470 11430 18522
rect 11442 18470 11494 18522
rect 11506 18470 11558 18522
rect 11570 18470 11622 18522
rect 18308 18470 18360 18522
rect 18372 18470 18424 18522
rect 18436 18470 18488 18522
rect 18500 18470 18552 18522
rect 2780 18275 2832 18284
rect 2780 18241 2789 18275
rect 2789 18241 2823 18275
rect 2823 18241 2832 18275
rect 11060 18275 11112 18284
rect 2780 18232 2832 18241
rect 11060 18241 11069 18275
rect 11069 18241 11103 18275
rect 11103 18241 11112 18275
rect 11060 18232 11112 18241
rect 2688 18164 2740 18216
rect 11428 18164 11480 18216
rect 3332 18096 3384 18148
rect 1952 18071 2004 18080
rect 1952 18037 1961 18071
rect 1961 18037 1995 18071
rect 1995 18037 2004 18071
rect 1952 18028 2004 18037
rect 7912 17926 7964 17978
rect 7976 17926 8028 17978
rect 8040 17926 8092 17978
rect 8104 17926 8156 17978
rect 14843 17926 14895 17978
rect 14907 17926 14959 17978
rect 14971 17926 15023 17978
rect 15035 17926 15087 17978
rect 1860 17867 1912 17876
rect 1860 17833 1869 17867
rect 1869 17833 1903 17867
rect 1903 17833 1912 17867
rect 1860 17824 1912 17833
rect 5632 17824 5684 17876
rect 9680 17867 9732 17876
rect 9680 17833 9689 17867
rect 9689 17833 9723 17867
rect 9723 17833 9732 17867
rect 9680 17824 9732 17833
rect 11428 17867 11480 17876
rect 11428 17833 11437 17867
rect 11437 17833 11471 17867
rect 11471 17833 11480 17867
rect 11428 17824 11480 17833
rect 1768 17756 1820 17808
rect 3240 17799 3292 17808
rect 3240 17765 3249 17799
rect 3249 17765 3283 17799
rect 3283 17765 3292 17799
rect 3240 17756 3292 17765
rect 5540 17756 5592 17808
rect 1676 17731 1728 17740
rect 1676 17697 1685 17731
rect 1685 17697 1719 17731
rect 1719 17697 1728 17731
rect 1676 17688 1728 17697
rect 7564 17688 7616 17740
rect 8208 17688 8260 17740
rect 12440 17688 12492 17740
rect 4068 17620 4120 17672
rect 8484 17663 8536 17672
rect 8484 17629 8493 17663
rect 8493 17629 8527 17663
rect 8527 17629 8536 17663
rect 8484 17620 8536 17629
rect 9312 17620 9364 17672
rect 9680 17620 9732 17672
rect 10324 17663 10376 17672
rect 10324 17629 10333 17663
rect 10333 17629 10367 17663
rect 10367 17629 10376 17663
rect 10324 17620 10376 17629
rect 11888 17663 11940 17672
rect 11888 17629 11897 17663
rect 11897 17629 11931 17663
rect 11931 17629 11940 17663
rect 11888 17620 11940 17629
rect 13728 17620 13780 17672
rect 8392 17552 8444 17604
rect 6460 17527 6512 17536
rect 6460 17493 6469 17527
rect 6469 17493 6503 17527
rect 6503 17493 6512 17527
rect 6460 17484 6512 17493
rect 4447 17382 4499 17434
rect 4511 17382 4563 17434
rect 4575 17382 4627 17434
rect 4639 17382 4691 17434
rect 11378 17382 11430 17434
rect 11442 17382 11494 17434
rect 11506 17382 11558 17434
rect 11570 17382 11622 17434
rect 18308 17382 18360 17434
rect 18372 17382 18424 17434
rect 18436 17382 18488 17434
rect 18500 17382 18552 17434
rect 1952 17323 2004 17332
rect 1952 17289 1961 17323
rect 1961 17289 1995 17323
rect 1995 17289 2004 17323
rect 1952 17280 2004 17289
rect 2964 17076 3016 17128
rect 3332 17187 3384 17196
rect 3332 17153 3341 17187
rect 3341 17153 3375 17187
rect 3375 17153 3384 17187
rect 3332 17144 3384 17153
rect 6460 17144 6512 17196
rect 8208 17187 8260 17196
rect 8208 17153 8217 17187
rect 8217 17153 8251 17187
rect 8251 17153 8260 17187
rect 8208 17144 8260 17153
rect 12440 17187 12492 17196
rect 12440 17153 12449 17187
rect 12449 17153 12483 17187
rect 12483 17153 12492 17187
rect 12440 17144 12492 17153
rect 4068 17076 4120 17128
rect 5724 17076 5776 17128
rect 8760 17076 8812 17128
rect 5448 17008 5500 17060
rect 9312 17008 9364 17060
rect 4160 16940 4212 16992
rect 5540 16983 5592 16992
rect 5540 16949 5549 16983
rect 5549 16949 5583 16983
rect 5583 16949 5592 16983
rect 5540 16940 5592 16949
rect 6276 16983 6328 16992
rect 6276 16949 6285 16983
rect 6285 16949 6319 16983
rect 6319 16949 6328 16983
rect 6276 16940 6328 16949
rect 6920 16940 6972 16992
rect 7472 16940 7524 16992
rect 10232 17008 10284 17060
rect 10324 16940 10376 16992
rect 7912 16838 7964 16890
rect 7976 16838 8028 16890
rect 8040 16838 8092 16890
rect 8104 16838 8156 16890
rect 14843 16838 14895 16890
rect 14907 16838 14959 16890
rect 14971 16838 15023 16890
rect 15035 16838 15087 16890
rect 2964 16779 3016 16788
rect 2964 16745 2973 16779
rect 2973 16745 3007 16779
rect 3007 16745 3016 16779
rect 2964 16736 3016 16745
rect 5448 16779 5500 16788
rect 1676 16668 1728 16720
rect 4252 16668 4304 16720
rect 5448 16745 5457 16779
rect 5457 16745 5491 16779
rect 5491 16745 5500 16779
rect 5448 16736 5500 16745
rect 6276 16736 6328 16788
rect 9312 16779 9364 16788
rect 5908 16668 5960 16720
rect 6460 16668 6512 16720
rect 3424 16575 3476 16584
rect 3424 16541 3433 16575
rect 3433 16541 3467 16575
rect 3467 16541 3476 16575
rect 3424 16532 3476 16541
rect 4160 16600 4212 16652
rect 4344 16643 4396 16652
rect 4344 16609 4378 16643
rect 4378 16609 4396 16643
rect 4344 16600 4396 16609
rect 5724 16600 5776 16652
rect 4068 16575 4120 16584
rect 4068 16541 4077 16575
rect 4077 16541 4111 16575
rect 4111 16541 4120 16575
rect 4068 16532 4120 16541
rect 7012 16600 7064 16652
rect 8760 16668 8812 16720
rect 9312 16745 9321 16779
rect 9321 16745 9355 16779
rect 9355 16745 9364 16779
rect 9312 16736 9364 16745
rect 9680 16779 9732 16788
rect 9680 16745 9689 16779
rect 9689 16745 9723 16779
rect 9723 16745 9732 16779
rect 9680 16736 9732 16745
rect 13728 16779 13780 16788
rect 10048 16711 10100 16720
rect 10048 16677 10057 16711
rect 10057 16677 10091 16711
rect 10091 16677 10100 16711
rect 10048 16668 10100 16677
rect 10324 16668 10376 16720
rect 11980 16668 12032 16720
rect 13728 16745 13737 16779
rect 13737 16745 13771 16779
rect 13771 16745 13780 16779
rect 13728 16736 13780 16745
rect 19248 16736 19300 16788
rect 9036 16600 9088 16652
rect 12348 16643 12400 16652
rect 12348 16609 12357 16643
rect 12357 16609 12391 16643
rect 12391 16609 12400 16643
rect 12348 16600 12400 16609
rect 10140 16575 10192 16584
rect 10140 16541 10149 16575
rect 10149 16541 10183 16575
rect 10183 16541 10192 16575
rect 10140 16532 10192 16541
rect 10232 16575 10284 16584
rect 10232 16541 10241 16575
rect 10241 16541 10275 16575
rect 10275 16541 10284 16575
rect 10692 16575 10744 16584
rect 10232 16532 10284 16541
rect 10692 16541 10701 16575
rect 10701 16541 10735 16575
rect 10735 16541 10744 16575
rect 10692 16532 10744 16541
rect 7288 16439 7340 16448
rect 7288 16405 7297 16439
rect 7297 16405 7331 16439
rect 7331 16405 7340 16439
rect 7288 16396 7340 16405
rect 4447 16294 4499 16346
rect 4511 16294 4563 16346
rect 4575 16294 4627 16346
rect 4639 16294 4691 16346
rect 11378 16294 11430 16346
rect 11442 16294 11494 16346
rect 11506 16294 11558 16346
rect 11570 16294 11622 16346
rect 18308 16294 18360 16346
rect 18372 16294 18424 16346
rect 18436 16294 18488 16346
rect 18500 16294 18552 16346
rect 1952 16235 2004 16244
rect 1952 16201 1961 16235
rect 1961 16201 1995 16235
rect 1995 16201 2004 16235
rect 1952 16192 2004 16201
rect 2780 16192 2832 16244
rect 4344 16235 4396 16244
rect 4344 16201 4353 16235
rect 4353 16201 4387 16235
rect 4387 16201 4396 16235
rect 4344 16192 4396 16201
rect 6920 16192 6972 16244
rect 9036 16192 9088 16244
rect 11888 16192 11940 16244
rect 4252 16056 4304 16108
rect 5540 16056 5592 16108
rect 7288 16056 7340 16108
rect 8760 16099 8812 16108
rect 8760 16065 8769 16099
rect 8769 16065 8803 16099
rect 8803 16065 8812 16099
rect 8760 16056 8812 16065
rect 11980 16099 12032 16108
rect 11980 16065 11989 16099
rect 11989 16065 12023 16099
rect 12023 16065 12032 16099
rect 11980 16056 12032 16065
rect 1768 16031 1820 16040
rect 1768 15997 1777 16031
rect 1777 15997 1811 16031
rect 1811 15997 1820 16031
rect 1768 15988 1820 15997
rect 2320 16031 2372 16040
rect 2320 15997 2329 16031
rect 2329 15997 2363 16031
rect 2363 15997 2372 16031
rect 2320 15988 2372 15997
rect 4068 15988 4120 16040
rect 3608 15920 3660 15972
rect 7012 15920 7064 15972
rect 4988 15852 5040 15904
rect 6276 15852 6328 15904
rect 6552 15852 6604 15904
rect 7196 15895 7248 15904
rect 7196 15861 7205 15895
rect 7205 15861 7239 15895
rect 7239 15861 7248 15895
rect 7196 15852 7248 15861
rect 7472 15852 7524 15904
rect 9588 15920 9640 15972
rect 10140 15920 10192 15972
rect 11980 15920 12032 15972
rect 7656 15895 7708 15904
rect 7656 15861 7665 15895
rect 7665 15861 7699 15895
rect 7699 15861 7708 15895
rect 7656 15852 7708 15861
rect 12440 15895 12492 15904
rect 12440 15861 12449 15895
rect 12449 15861 12483 15895
rect 12483 15861 12492 15895
rect 12440 15852 12492 15861
rect 7912 15750 7964 15802
rect 7976 15750 8028 15802
rect 8040 15750 8092 15802
rect 8104 15750 8156 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 15035 15750 15087 15802
rect 1676 15691 1728 15700
rect 1676 15657 1685 15691
rect 1685 15657 1719 15691
rect 1719 15657 1728 15691
rect 1676 15648 1728 15657
rect 3424 15648 3476 15700
rect 2320 15623 2372 15632
rect 2320 15589 2329 15623
rect 2329 15589 2363 15623
rect 2363 15589 2372 15623
rect 2320 15580 2372 15589
rect 2964 15512 3016 15564
rect 3700 15512 3752 15564
rect 8300 15648 8352 15700
rect 8484 15691 8536 15700
rect 8484 15657 8493 15691
rect 8493 15657 8527 15691
rect 8527 15657 8536 15691
rect 8484 15648 8536 15657
rect 10048 15691 10100 15700
rect 10048 15657 10057 15691
rect 10057 15657 10091 15691
rect 10091 15657 10100 15691
rect 10048 15648 10100 15657
rect 4896 15580 4948 15632
rect 5080 15512 5132 15564
rect 6552 15580 6604 15632
rect 7288 15580 7340 15632
rect 9128 15512 9180 15564
rect 2596 15444 2648 15496
rect 4344 15376 4396 15428
rect 5816 15487 5868 15496
rect 5816 15453 5825 15487
rect 5825 15453 5859 15487
rect 5859 15453 5868 15487
rect 5816 15444 5868 15453
rect 3700 15351 3752 15360
rect 3700 15317 3709 15351
rect 3709 15317 3743 15351
rect 3743 15317 3752 15351
rect 3700 15308 3752 15317
rect 4160 15308 4212 15360
rect 9036 15487 9088 15496
rect 9036 15453 9045 15487
rect 9045 15453 9079 15487
rect 9079 15453 9088 15487
rect 9036 15444 9088 15453
rect 11152 15376 11204 15428
rect 6920 15308 6972 15360
rect 7472 15308 7524 15360
rect 4447 15206 4499 15258
rect 4511 15206 4563 15258
rect 4575 15206 4627 15258
rect 4639 15206 4691 15258
rect 11378 15206 11430 15258
rect 11442 15206 11494 15258
rect 11506 15206 11558 15258
rect 11570 15206 11622 15258
rect 18308 15206 18360 15258
rect 18372 15206 18424 15258
rect 18436 15206 18488 15258
rect 18500 15206 18552 15258
rect 1860 15147 1912 15156
rect 1860 15113 1869 15147
rect 1869 15113 1903 15147
rect 1903 15113 1912 15147
rect 1860 15104 1912 15113
rect 2964 15147 3016 15156
rect 2964 15113 2973 15147
rect 2973 15113 3007 15147
rect 3007 15113 3016 15147
rect 2964 15104 3016 15113
rect 1768 14968 1820 15020
rect 3608 15011 3660 15020
rect 3608 14977 3617 15011
rect 3617 14977 3651 15011
rect 3651 14977 3660 15011
rect 8300 15147 8352 15156
rect 8300 15113 8309 15147
rect 8309 15113 8343 15147
rect 8343 15113 8352 15147
rect 8300 15104 8352 15113
rect 8944 15104 8996 15156
rect 4896 15036 4948 15088
rect 5908 15036 5960 15088
rect 3608 14968 3660 14977
rect 7196 14968 7248 15020
rect 7472 15011 7524 15020
rect 7472 14977 7481 15011
rect 7481 14977 7515 15011
rect 7515 14977 7524 15011
rect 7472 14968 7524 14977
rect 9588 15011 9640 15020
rect 9588 14977 9597 15011
rect 9597 14977 9631 15011
rect 9631 14977 9640 15011
rect 9588 14968 9640 14977
rect 1676 14943 1728 14952
rect 1676 14909 1685 14943
rect 1685 14909 1719 14943
rect 1719 14909 1728 14943
rect 1676 14900 1728 14909
rect 4160 14900 4212 14952
rect 4436 14900 4488 14952
rect 5816 14832 5868 14884
rect 5632 14764 5684 14816
rect 11244 14764 11296 14816
rect 7912 14662 7964 14714
rect 7976 14662 8028 14714
rect 8040 14662 8092 14714
rect 8104 14662 8156 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 15035 14662 15087 14714
rect 3240 14603 3292 14612
rect 3240 14569 3249 14603
rect 3249 14569 3283 14603
rect 3283 14569 3292 14603
rect 3240 14560 3292 14569
rect 5816 14603 5868 14612
rect 5816 14569 5825 14603
rect 5825 14569 5859 14603
rect 5859 14569 5868 14603
rect 5816 14560 5868 14569
rect 9588 14560 9640 14612
rect 1768 14467 1820 14476
rect 1768 14433 1777 14467
rect 1777 14433 1811 14467
rect 1811 14433 1820 14467
rect 1768 14424 1820 14433
rect 7472 14492 7524 14544
rect 2780 14424 2832 14476
rect 5264 14424 5316 14476
rect 5816 14424 5868 14476
rect 6920 14467 6972 14476
rect 6920 14433 6929 14467
rect 6929 14433 6963 14467
rect 6963 14433 6972 14467
rect 6920 14424 6972 14433
rect 8760 14424 8812 14476
rect 9588 14424 9640 14476
rect 10876 14424 10928 14476
rect 1676 14356 1728 14408
rect 4160 14356 4212 14408
rect 4436 14399 4488 14408
rect 4436 14365 4445 14399
rect 4445 14365 4479 14399
rect 4479 14365 4488 14399
rect 4436 14356 4488 14365
rect 1952 14263 2004 14272
rect 1952 14229 1961 14263
rect 1961 14229 1995 14263
rect 1995 14229 2004 14263
rect 1952 14220 2004 14229
rect 8208 14220 8260 14272
rect 11704 14263 11756 14272
rect 11704 14229 11713 14263
rect 11713 14229 11747 14263
rect 11747 14229 11756 14263
rect 11704 14220 11756 14229
rect 4447 14118 4499 14170
rect 4511 14118 4563 14170
rect 4575 14118 4627 14170
rect 4639 14118 4691 14170
rect 11378 14118 11430 14170
rect 11442 14118 11494 14170
rect 11506 14118 11558 14170
rect 11570 14118 11622 14170
rect 18308 14118 18360 14170
rect 18372 14118 18424 14170
rect 18436 14118 18488 14170
rect 18500 14118 18552 14170
rect 2964 14016 3016 14068
rect 5264 14016 5316 14068
rect 5632 14059 5684 14068
rect 2780 13880 2832 13932
rect 5632 14025 5641 14059
rect 5641 14025 5675 14059
rect 5675 14025 5684 14059
rect 5632 14016 5684 14025
rect 7012 14016 7064 14068
rect 10876 14016 10928 14068
rect 11244 14059 11296 14068
rect 8944 13948 8996 14000
rect 8208 13880 8260 13932
rect 1584 13855 1636 13864
rect 1584 13821 1593 13855
rect 1593 13821 1627 13855
rect 1627 13821 1636 13855
rect 1584 13812 1636 13821
rect 3056 13855 3108 13864
rect 3056 13821 3065 13855
rect 3065 13821 3099 13855
rect 3099 13821 3108 13855
rect 3056 13812 3108 13821
rect 3148 13812 3200 13864
rect 4068 13812 4120 13864
rect 2596 13787 2648 13796
rect 2596 13753 2605 13787
rect 2605 13753 2639 13787
rect 2639 13753 2648 13787
rect 2596 13744 2648 13753
rect 5080 13744 5132 13796
rect 2872 13676 2924 13728
rect 6828 13812 6880 13864
rect 5540 13744 5592 13796
rect 8576 13812 8628 13864
rect 9588 13923 9640 13932
rect 9588 13889 9597 13923
rect 9597 13889 9631 13923
rect 9631 13889 9640 13923
rect 9588 13880 9640 13889
rect 11244 14025 11253 14059
rect 11253 14025 11287 14059
rect 11287 14025 11296 14059
rect 11244 14016 11296 14025
rect 8760 13812 8812 13864
rect 9128 13812 9180 13864
rect 9404 13812 9456 13864
rect 11704 13812 11756 13864
rect 6000 13719 6052 13728
rect 6000 13685 6009 13719
rect 6009 13685 6043 13719
rect 6043 13685 6052 13719
rect 6000 13676 6052 13685
rect 10876 13744 10928 13796
rect 11888 13676 11940 13728
rect 7912 13574 7964 13626
rect 7976 13574 8028 13626
rect 8040 13574 8092 13626
rect 8104 13574 8156 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 15035 13574 15087 13626
rect 3516 13515 3568 13524
rect 3516 13481 3525 13515
rect 3525 13481 3559 13515
rect 3559 13481 3568 13515
rect 3516 13472 3568 13481
rect 6000 13472 6052 13524
rect 10876 13472 10928 13524
rect 1768 13404 1820 13456
rect 3056 13404 3108 13456
rect 5080 13404 5132 13456
rect 1952 13336 2004 13388
rect 3240 13336 3292 13388
rect 3424 13336 3476 13388
rect 5264 13336 5316 13388
rect 8208 13404 8260 13456
rect 6920 13336 6972 13388
rect 8116 13336 8168 13388
rect 10048 13404 10100 13456
rect 10692 13404 10744 13456
rect 11060 13336 11112 13388
rect 5448 13200 5500 13252
rect 8024 13268 8076 13320
rect 6092 13175 6144 13184
rect 6092 13141 6101 13175
rect 6101 13141 6135 13175
rect 6135 13141 6144 13175
rect 6092 13132 6144 13141
rect 8392 13175 8444 13184
rect 8392 13141 8401 13175
rect 8401 13141 8435 13175
rect 8435 13141 8444 13175
rect 8392 13132 8444 13141
rect 10968 13132 11020 13184
rect 11888 13132 11940 13184
rect 4447 13030 4499 13082
rect 4511 13030 4563 13082
rect 4575 13030 4627 13082
rect 4639 13030 4691 13082
rect 11378 13030 11430 13082
rect 11442 13030 11494 13082
rect 11506 13030 11558 13082
rect 11570 13030 11622 13082
rect 18308 13030 18360 13082
rect 18372 13030 18424 13082
rect 18436 13030 18488 13082
rect 18500 13030 18552 13082
rect 1584 12928 1636 12980
rect 5080 12928 5132 12980
rect 7012 12971 7064 12980
rect 7012 12937 7021 12971
rect 7021 12937 7055 12971
rect 7055 12937 7064 12971
rect 7012 12928 7064 12937
rect 8484 12971 8536 12980
rect 8484 12937 8493 12971
rect 8493 12937 8527 12971
rect 8527 12937 8536 12971
rect 8484 12928 8536 12937
rect 10600 12971 10652 12980
rect 10600 12937 10609 12971
rect 10609 12937 10643 12971
rect 10643 12937 10652 12971
rect 10600 12928 10652 12937
rect 5264 12860 5316 12912
rect 5448 12860 5500 12912
rect 8852 12860 8904 12912
rect 10876 12860 10928 12912
rect 2872 12835 2924 12844
rect 2872 12801 2881 12835
rect 2881 12801 2915 12835
rect 2915 12801 2924 12835
rect 2872 12792 2924 12801
rect 3424 12835 3476 12844
rect 3424 12801 3433 12835
rect 3433 12801 3467 12835
rect 3467 12801 3476 12835
rect 3424 12792 3476 12801
rect 8208 12792 8260 12844
rect 8392 12792 8444 12844
rect 11060 12792 11112 12844
rect 4068 12724 4120 12776
rect 4160 12767 4212 12776
rect 4160 12733 4169 12767
rect 4169 12733 4203 12767
rect 4203 12733 4212 12767
rect 4160 12724 4212 12733
rect 7012 12724 7064 12776
rect 7748 12724 7800 12776
rect 8944 12767 8996 12776
rect 8944 12733 8953 12767
rect 8953 12733 8987 12767
rect 8987 12733 8996 12767
rect 8944 12724 8996 12733
rect 9588 12724 9640 12776
rect 10876 12724 10928 12776
rect 4712 12656 4764 12708
rect 8024 12656 8076 12708
rect 2596 12631 2648 12640
rect 2596 12597 2605 12631
rect 2605 12597 2639 12631
rect 2639 12597 2648 12631
rect 2596 12588 2648 12597
rect 2780 12588 2832 12640
rect 5080 12588 5132 12640
rect 6368 12588 6420 12640
rect 8760 12588 8812 12640
rect 10968 12631 11020 12640
rect 10968 12597 10977 12631
rect 10977 12597 11011 12631
rect 11011 12597 11020 12631
rect 10968 12588 11020 12597
rect 7912 12486 7964 12538
rect 7976 12486 8028 12538
rect 8040 12486 8092 12538
rect 8104 12486 8156 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 15035 12486 15087 12538
rect 1492 12384 1544 12436
rect 3148 12384 3200 12436
rect 8852 12427 8904 12436
rect 2872 12316 2924 12368
rect 3332 12316 3384 12368
rect 3976 12316 4028 12368
rect 5632 12316 5684 12368
rect 8392 12316 8444 12368
rect 8852 12393 8861 12427
rect 8861 12393 8895 12427
rect 8895 12393 8904 12427
rect 8852 12384 8904 12393
rect 9588 12384 9640 12436
rect 11060 12384 11112 12436
rect 12164 12384 12216 12436
rect 12440 12384 12492 12436
rect 19708 12384 19760 12436
rect 11704 12316 11756 12368
rect 2044 12248 2096 12300
rect 2964 12248 3016 12300
rect 4804 12248 4856 12300
rect 5080 12291 5132 12300
rect 5080 12257 5089 12291
rect 5089 12257 5123 12291
rect 5123 12257 5132 12291
rect 5080 12248 5132 12257
rect 5908 12248 5960 12300
rect 9956 12248 10008 12300
rect 11060 12248 11112 12300
rect 4712 12223 4764 12232
rect 4712 12189 4721 12223
rect 4721 12189 4755 12223
rect 4755 12189 4764 12223
rect 4712 12180 4764 12189
rect 4252 12112 4304 12164
rect 3332 12087 3384 12096
rect 3332 12053 3341 12087
rect 3341 12053 3375 12087
rect 3375 12053 3384 12087
rect 3332 12044 3384 12053
rect 4160 12044 4212 12096
rect 6368 12180 6420 12232
rect 6828 12223 6880 12232
rect 6828 12189 6837 12223
rect 6837 12189 6871 12223
rect 6871 12189 6880 12223
rect 6828 12180 6880 12189
rect 8300 12112 8352 12164
rect 8116 12044 8168 12096
rect 9220 12087 9272 12096
rect 9220 12053 9229 12087
rect 9229 12053 9263 12087
rect 9263 12053 9272 12087
rect 9220 12044 9272 12053
rect 19708 12291 19760 12300
rect 19708 12257 19717 12291
rect 19717 12257 19751 12291
rect 19751 12257 19760 12291
rect 19708 12248 19760 12257
rect 20536 12044 20588 12096
rect 4447 11942 4499 11994
rect 4511 11942 4563 11994
rect 4575 11942 4627 11994
rect 4639 11942 4691 11994
rect 11378 11942 11430 11994
rect 11442 11942 11494 11994
rect 11506 11942 11558 11994
rect 11570 11942 11622 11994
rect 18308 11942 18360 11994
rect 18372 11942 18424 11994
rect 18436 11942 18488 11994
rect 18500 11942 18552 11994
rect 2596 11840 2648 11892
rect 2688 11840 2740 11892
rect 7564 11840 7616 11892
rect 2964 11704 3016 11756
rect 4804 11704 4856 11756
rect 8208 11747 8260 11756
rect 2044 11636 2096 11688
rect 2412 11636 2464 11688
rect 3332 11679 3384 11688
rect 3332 11645 3366 11679
rect 3366 11645 3384 11679
rect 3332 11636 3384 11645
rect 8208 11713 8217 11747
rect 8217 11713 8251 11747
rect 8251 11713 8260 11747
rect 8208 11704 8260 11713
rect 9864 11704 9916 11756
rect 8484 11679 8536 11688
rect 8484 11645 8507 11679
rect 8507 11645 8536 11679
rect 8484 11636 8536 11645
rect 9404 11636 9456 11688
rect 11060 11636 11112 11688
rect 11704 11636 11756 11688
rect 2320 11500 2372 11552
rect 3976 11568 4028 11620
rect 10048 11568 10100 11620
rect 3148 11500 3200 11552
rect 4344 11500 4396 11552
rect 7380 11543 7432 11552
rect 7380 11509 7389 11543
rect 7389 11509 7423 11543
rect 7423 11509 7432 11543
rect 7380 11500 7432 11509
rect 7472 11543 7524 11552
rect 7472 11509 7481 11543
rect 7481 11509 7515 11543
rect 7515 11509 7524 11543
rect 7472 11500 7524 11509
rect 9220 11500 9272 11552
rect 20076 11500 20128 11552
rect 7912 11398 7964 11450
rect 7976 11398 8028 11450
rect 8040 11398 8092 11450
rect 8104 11398 8156 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 15035 11398 15087 11450
rect 2320 11339 2372 11348
rect 2320 11305 2329 11339
rect 2329 11305 2363 11339
rect 2363 11305 2372 11339
rect 2320 11296 2372 11305
rect 2780 11339 2832 11348
rect 2780 11305 2789 11339
rect 2789 11305 2823 11339
rect 2823 11305 2832 11339
rect 2780 11296 2832 11305
rect 3056 11296 3108 11348
rect 5908 11296 5960 11348
rect 6092 11296 6144 11348
rect 7380 11296 7432 11348
rect 4252 11228 4304 11280
rect 10140 11296 10192 11348
rect 11060 11339 11112 11348
rect 11060 11305 11069 11339
rect 11069 11305 11103 11339
rect 11103 11305 11112 11339
rect 11060 11296 11112 11305
rect 9864 11228 9916 11280
rect 10048 11228 10100 11280
rect 2964 11160 3016 11212
rect 5448 11160 5500 11212
rect 7196 11160 7248 11212
rect 8208 11160 8260 11212
rect 9680 11203 9732 11212
rect 9680 11169 9689 11203
rect 9689 11169 9723 11203
rect 9723 11169 9732 11203
rect 9680 11160 9732 11169
rect 4160 11092 4212 11144
rect 6828 11092 6880 11144
rect 4252 11024 4304 11076
rect 8484 11067 8536 11076
rect 8484 11033 8493 11067
rect 8493 11033 8527 11067
rect 8527 11033 8536 11067
rect 8484 11024 8536 11033
rect 9404 11024 9456 11076
rect 11244 11160 11296 11212
rect 19524 11024 19576 11076
rect 3884 10956 3936 11008
rect 11060 10956 11112 11008
rect 4447 10854 4499 10906
rect 4511 10854 4563 10906
rect 4575 10854 4627 10906
rect 4639 10854 4691 10906
rect 11378 10854 11430 10906
rect 11442 10854 11494 10906
rect 11506 10854 11558 10906
rect 11570 10854 11622 10906
rect 18308 10854 18360 10906
rect 18372 10854 18424 10906
rect 18436 10854 18488 10906
rect 18500 10854 18552 10906
rect 2964 10752 3016 10804
rect 5448 10795 5500 10804
rect 5448 10761 5457 10795
rect 5457 10761 5491 10795
rect 5491 10761 5500 10795
rect 5448 10752 5500 10761
rect 5816 10752 5868 10804
rect 7472 10752 7524 10804
rect 7564 10752 7616 10804
rect 7748 10752 7800 10804
rect 9128 10752 9180 10804
rect 12348 10752 12400 10804
rect 5448 10616 5500 10668
rect 8208 10616 8260 10668
rect 2412 10548 2464 10600
rect 4160 10548 4212 10600
rect 4344 10591 4396 10600
rect 4344 10557 4378 10591
rect 4378 10557 4396 10591
rect 4344 10548 4396 10557
rect 5816 10548 5868 10600
rect 11796 10684 11848 10736
rect 19156 10684 19208 10736
rect 9496 10659 9548 10668
rect 9496 10625 9505 10659
rect 9505 10625 9539 10659
rect 9539 10625 9548 10659
rect 9496 10616 9548 10625
rect 2964 10480 3016 10532
rect 3976 10480 4028 10532
rect 11244 10548 11296 10600
rect 3884 10412 3936 10464
rect 4160 10412 4212 10464
rect 6184 10455 6236 10464
rect 6184 10421 6193 10455
rect 6193 10421 6227 10455
rect 6227 10421 6236 10455
rect 8944 10455 8996 10464
rect 6184 10412 6236 10421
rect 8944 10421 8953 10455
rect 8953 10421 8987 10455
rect 8987 10421 8996 10455
rect 8944 10412 8996 10421
rect 9312 10455 9364 10464
rect 9312 10421 9321 10455
rect 9321 10421 9355 10455
rect 9355 10421 9364 10455
rect 9312 10412 9364 10421
rect 9680 10412 9732 10464
rect 20720 10412 20772 10464
rect 7912 10310 7964 10362
rect 7976 10310 8028 10362
rect 8040 10310 8092 10362
rect 8104 10310 8156 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 15035 10310 15087 10362
rect 4160 10251 4212 10260
rect 4160 10217 4169 10251
rect 4169 10217 4203 10251
rect 4203 10217 4212 10251
rect 4160 10208 4212 10217
rect 6184 10208 6236 10260
rect 7196 10208 7248 10260
rect 8944 10208 8996 10260
rect 9312 10208 9364 10260
rect 11244 10208 11296 10260
rect 3884 10072 3936 10124
rect 5816 10140 5868 10192
rect 5908 10140 5960 10192
rect 8760 10183 8812 10192
rect 5356 10072 5408 10124
rect 5724 10072 5776 10124
rect 2688 9936 2740 9988
rect 4160 10004 4212 10056
rect 4344 10004 4396 10056
rect 6184 10047 6236 10056
rect 3148 9936 3200 9988
rect 5632 9979 5684 9988
rect 5632 9945 5641 9979
rect 5641 9945 5675 9979
rect 5675 9945 5684 9979
rect 5632 9936 5684 9945
rect 6184 10013 6193 10047
rect 6193 10013 6227 10047
rect 6227 10013 6236 10047
rect 6184 10004 6236 10013
rect 8760 10149 8769 10183
rect 8769 10149 8803 10183
rect 8803 10149 8812 10183
rect 8760 10140 8812 10149
rect 6920 10072 6972 10124
rect 7748 10115 7800 10124
rect 7748 10081 7757 10115
rect 7757 10081 7791 10115
rect 7791 10081 7800 10115
rect 7748 10072 7800 10081
rect 9588 10072 9640 10124
rect 11244 10072 11296 10124
rect 11704 10072 11756 10124
rect 8208 10004 8260 10056
rect 3608 9868 3660 9920
rect 4160 9868 4212 9920
rect 7288 9936 7340 9988
rect 9220 10004 9272 10056
rect 10324 10047 10376 10056
rect 10324 10013 10333 10047
rect 10333 10013 10367 10047
rect 10367 10013 10376 10047
rect 10324 10004 10376 10013
rect 8392 9911 8444 9920
rect 8392 9877 8401 9911
rect 8401 9877 8435 9911
rect 8435 9877 8444 9911
rect 8392 9868 8444 9877
rect 12348 9868 12400 9920
rect 12532 9911 12584 9920
rect 12532 9877 12541 9911
rect 12541 9877 12575 9911
rect 12575 9877 12584 9911
rect 12532 9868 12584 9877
rect 4447 9766 4499 9818
rect 4511 9766 4563 9818
rect 4575 9766 4627 9818
rect 4639 9766 4691 9818
rect 11378 9766 11430 9818
rect 11442 9766 11494 9818
rect 11506 9766 11558 9818
rect 11570 9766 11622 9818
rect 18308 9766 18360 9818
rect 18372 9766 18424 9818
rect 18436 9766 18488 9818
rect 18500 9766 18552 9818
rect 3976 9664 4028 9716
rect 14188 9664 14240 9716
rect 2964 9639 3016 9648
rect 2964 9605 2973 9639
rect 2973 9605 3007 9639
rect 3007 9605 3016 9639
rect 2964 9596 3016 9605
rect 3240 9639 3292 9648
rect 3240 9605 3249 9639
rect 3249 9605 3283 9639
rect 3283 9605 3292 9639
rect 3240 9596 3292 9605
rect 3332 9596 3384 9648
rect 3700 9596 3752 9648
rect 4068 9596 4120 9648
rect 12348 9596 12400 9648
rect 5448 9528 5500 9580
rect 2688 9460 2740 9512
rect 3608 9503 3660 9512
rect 3608 9469 3617 9503
rect 3617 9469 3651 9503
rect 3651 9469 3660 9503
rect 3608 9460 3660 9469
rect 6644 9460 6696 9512
rect 6828 9503 6880 9512
rect 6828 9469 6837 9503
rect 6837 9469 6871 9503
rect 6871 9469 6880 9503
rect 6828 9460 6880 9469
rect 9864 9460 9916 9512
rect 10508 9460 10560 9512
rect 10784 9460 10836 9512
rect 11060 9460 11112 9512
rect 12532 9528 12584 9580
rect 11704 9460 11756 9512
rect 3792 9392 3844 9444
rect 4804 9392 4856 9444
rect 7196 9392 7248 9444
rect 1860 9324 1912 9376
rect 3700 9367 3752 9376
rect 3700 9333 3709 9367
rect 3709 9333 3743 9367
rect 3743 9333 3752 9367
rect 3700 9324 3752 9333
rect 4896 9367 4948 9376
rect 4896 9333 4905 9367
rect 4905 9333 4939 9367
rect 4939 9333 4948 9367
rect 4896 9324 4948 9333
rect 5356 9324 5408 9376
rect 5724 9324 5776 9376
rect 9220 9392 9272 9444
rect 10324 9392 10376 9444
rect 8208 9367 8260 9376
rect 8208 9333 8217 9367
rect 8217 9333 8251 9367
rect 8251 9333 8260 9367
rect 8208 9324 8260 9333
rect 8484 9367 8536 9376
rect 8484 9333 8493 9367
rect 8493 9333 8527 9367
rect 8527 9333 8536 9367
rect 8484 9324 8536 9333
rect 9496 9324 9548 9376
rect 14648 9392 14700 9444
rect 12624 9324 12676 9376
rect 12808 9367 12860 9376
rect 12808 9333 12817 9367
rect 12817 9333 12851 9367
rect 12851 9333 12860 9367
rect 12808 9324 12860 9333
rect 7912 9222 7964 9274
rect 7976 9222 8028 9274
rect 8040 9222 8092 9274
rect 8104 9222 8156 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 15035 9222 15087 9274
rect 3700 9120 3752 9172
rect 4896 9120 4948 9172
rect 5080 9120 5132 9172
rect 6736 9120 6788 9172
rect 7748 9163 7800 9172
rect 7748 9129 7757 9163
rect 7757 9129 7791 9163
rect 7791 9129 7800 9163
rect 7748 9120 7800 9129
rect 8484 9120 8536 9172
rect 8760 9163 8812 9172
rect 8760 9129 8769 9163
rect 8769 9129 8803 9163
rect 8803 9129 8812 9163
rect 8760 9120 8812 9129
rect 9680 9163 9732 9172
rect 9680 9129 9689 9163
rect 9689 9129 9723 9163
rect 9723 9129 9732 9163
rect 9680 9120 9732 9129
rect 11060 9120 11112 9172
rect 11704 9120 11756 9172
rect 12348 9120 12400 9172
rect 2688 9052 2740 9104
rect 2780 9027 2832 9036
rect 2780 8993 2789 9027
rect 2789 8993 2823 9027
rect 2823 8993 2832 9027
rect 2780 8984 2832 8993
rect 4068 9052 4120 9104
rect 5632 8984 5684 9036
rect 6092 8984 6144 9036
rect 7564 8984 7616 9036
rect 8392 9052 8444 9104
rect 10048 9027 10100 9036
rect 10048 8993 10057 9027
rect 10057 8993 10091 9027
rect 10091 8993 10100 9027
rect 10048 8984 10100 8993
rect 12532 9052 12584 9104
rect 14372 8984 14424 9036
rect 15108 8984 15160 9036
rect 2872 8959 2924 8968
rect 2872 8925 2881 8959
rect 2881 8925 2915 8959
rect 2915 8925 2924 8959
rect 2872 8916 2924 8925
rect 3056 8959 3108 8968
rect 3056 8925 3065 8959
rect 3065 8925 3099 8959
rect 3099 8925 3108 8959
rect 3056 8916 3108 8925
rect 4160 8891 4212 8900
rect 4160 8857 4169 8891
rect 4169 8857 4203 8891
rect 4203 8857 4212 8891
rect 4160 8848 4212 8857
rect 4252 8780 4304 8832
rect 4988 8780 5040 8832
rect 5080 8780 5132 8832
rect 5264 8916 5316 8968
rect 7196 8916 7248 8968
rect 9496 8916 9548 8968
rect 10324 8959 10376 8968
rect 6644 8848 6696 8900
rect 10324 8925 10333 8959
rect 10333 8925 10367 8959
rect 10367 8925 10376 8959
rect 11704 8959 11756 8968
rect 10324 8916 10376 8925
rect 7196 8823 7248 8832
rect 7196 8789 7205 8823
rect 7205 8789 7239 8823
rect 7239 8789 7248 8823
rect 7196 8780 7248 8789
rect 8944 8780 8996 8832
rect 9588 8780 9640 8832
rect 10600 8848 10652 8900
rect 11060 8848 11112 8900
rect 10784 8823 10836 8832
rect 10784 8789 10793 8823
rect 10793 8789 10827 8823
rect 10827 8789 10836 8823
rect 11704 8925 11713 8959
rect 11713 8925 11747 8959
rect 11747 8925 11756 8959
rect 11704 8916 11756 8925
rect 14556 8959 14608 8968
rect 14556 8925 14565 8959
rect 14565 8925 14599 8959
rect 14599 8925 14608 8959
rect 14556 8916 14608 8925
rect 14648 8959 14700 8968
rect 14648 8925 14657 8959
rect 14657 8925 14691 8959
rect 14691 8925 14700 8959
rect 14648 8916 14700 8925
rect 10784 8780 10836 8789
rect 16488 8780 16540 8832
rect 4447 8678 4499 8730
rect 4511 8678 4563 8730
rect 4575 8678 4627 8730
rect 4639 8678 4691 8730
rect 11378 8678 11430 8730
rect 11442 8678 11494 8730
rect 11506 8678 11558 8730
rect 11570 8678 11622 8730
rect 18308 8678 18360 8730
rect 18372 8678 18424 8730
rect 18436 8678 18488 8730
rect 18500 8678 18552 8730
rect 3056 8576 3108 8628
rect 5264 8576 5316 8628
rect 5448 8576 5500 8628
rect 6092 8576 6144 8628
rect 11244 8576 11296 8628
rect 12164 8576 12216 8628
rect 14648 8576 14700 8628
rect 12624 8508 12676 8560
rect 5632 8440 5684 8492
rect 6828 8440 6880 8492
rect 8024 8440 8076 8492
rect 10048 8440 10100 8492
rect 12808 8440 12860 8492
rect 15108 8483 15160 8492
rect 1860 8372 1912 8424
rect 5080 8372 5132 8424
rect 8208 8372 8260 8424
rect 10600 8415 10652 8424
rect 10600 8381 10609 8415
rect 10609 8381 10643 8415
rect 10643 8381 10652 8415
rect 10600 8372 10652 8381
rect 11796 8415 11848 8424
rect 11796 8381 11805 8415
rect 11805 8381 11839 8415
rect 11839 8381 11848 8415
rect 11796 8372 11848 8381
rect 11888 8372 11940 8424
rect 12256 8372 12308 8424
rect 15108 8449 15117 8483
rect 15117 8449 15151 8483
rect 15151 8449 15160 8483
rect 15108 8440 15160 8449
rect 2504 8304 2556 8356
rect 1584 8279 1636 8288
rect 1584 8245 1593 8279
rect 1593 8245 1627 8279
rect 1627 8245 1636 8279
rect 3332 8304 3384 8356
rect 3608 8304 3660 8356
rect 3976 8304 4028 8356
rect 13360 8304 13412 8356
rect 1584 8236 1636 8245
rect 3148 8236 3200 8288
rect 5540 8236 5592 8288
rect 14464 8304 14516 8356
rect 18604 8304 18656 8356
rect 14096 8236 14148 8288
rect 7912 8134 7964 8186
rect 7976 8134 8028 8186
rect 8040 8134 8092 8186
rect 8104 8134 8156 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 15035 8134 15087 8186
rect 2780 8032 2832 8084
rect 2872 8032 2924 8084
rect 4804 8032 4856 8084
rect 1584 7896 1636 7948
rect 3884 7964 3936 8016
rect 14556 8032 14608 8084
rect 14188 8007 14240 8016
rect 3148 7896 3200 7948
rect 3332 7939 3384 7948
rect 3332 7905 3341 7939
rect 3341 7905 3375 7939
rect 3375 7905 3384 7939
rect 3332 7896 3384 7905
rect 2504 7871 2556 7880
rect 2504 7837 2513 7871
rect 2513 7837 2547 7871
rect 2547 7837 2556 7871
rect 2504 7828 2556 7837
rect 3056 7760 3108 7812
rect 5724 7896 5776 7948
rect 8852 7939 8904 7948
rect 5080 7871 5132 7880
rect 5080 7837 5089 7871
rect 5089 7837 5123 7871
rect 5123 7837 5132 7871
rect 5080 7828 5132 7837
rect 5908 7871 5960 7880
rect 5908 7837 5917 7871
rect 5917 7837 5951 7871
rect 5951 7837 5960 7871
rect 5908 7828 5960 7837
rect 6092 7871 6144 7880
rect 6092 7837 6101 7871
rect 6101 7837 6135 7871
rect 6135 7837 6144 7871
rect 6092 7828 6144 7837
rect 3976 7760 4028 7812
rect 8852 7905 8861 7939
rect 8861 7905 8895 7939
rect 8895 7905 8904 7939
rect 8852 7896 8904 7905
rect 5080 7692 5132 7744
rect 7288 7692 7340 7744
rect 7932 7828 7984 7880
rect 14188 7973 14197 8007
rect 14197 7973 14231 8007
rect 14231 7973 14240 8007
rect 14188 7964 14240 7973
rect 10508 7939 10560 7948
rect 10508 7905 10517 7939
rect 10517 7905 10551 7939
rect 10551 7905 10560 7939
rect 10508 7896 10560 7905
rect 11704 7896 11756 7948
rect 11888 7896 11940 7948
rect 9036 7871 9088 7880
rect 9036 7837 9045 7871
rect 9045 7837 9079 7871
rect 9079 7837 9088 7871
rect 9036 7828 9088 7837
rect 11612 7828 11664 7880
rect 13636 7828 13688 7880
rect 14464 7871 14516 7880
rect 14464 7837 14473 7871
rect 14473 7837 14507 7871
rect 14507 7837 14516 7871
rect 14464 7828 14516 7837
rect 16488 7896 16540 7948
rect 15476 7871 15528 7880
rect 15476 7837 15485 7871
rect 15485 7837 15519 7871
rect 15519 7837 15528 7871
rect 15476 7828 15528 7837
rect 17500 7828 17552 7880
rect 11888 7735 11940 7744
rect 11888 7701 11897 7735
rect 11897 7701 11931 7735
rect 11931 7701 11940 7735
rect 11888 7692 11940 7701
rect 4447 7590 4499 7642
rect 4511 7590 4563 7642
rect 4575 7590 4627 7642
rect 4639 7590 4691 7642
rect 11378 7590 11430 7642
rect 11442 7590 11494 7642
rect 11506 7590 11558 7642
rect 11570 7590 11622 7642
rect 18308 7590 18360 7642
rect 18372 7590 18424 7642
rect 18436 7590 18488 7642
rect 18500 7590 18552 7642
rect 2504 7488 2556 7540
rect 3056 7488 3108 7540
rect 3332 7488 3384 7540
rect 4896 7488 4948 7540
rect 5264 7531 5316 7540
rect 5264 7497 5273 7531
rect 5273 7497 5307 7531
rect 5307 7497 5316 7531
rect 5264 7488 5316 7497
rect 5724 7531 5776 7540
rect 5724 7497 5733 7531
rect 5733 7497 5767 7531
rect 5767 7497 5776 7531
rect 5724 7488 5776 7497
rect 9036 7531 9088 7540
rect 9036 7497 9045 7531
rect 9045 7497 9079 7531
rect 9079 7497 9088 7531
rect 9036 7488 9088 7497
rect 14464 7488 14516 7540
rect 4068 7420 4120 7472
rect 3240 7352 3292 7404
rect 6092 7352 6144 7404
rect 1860 7284 1912 7336
rect 4896 7284 4948 7336
rect 7196 7327 7248 7336
rect 7196 7293 7205 7327
rect 7205 7293 7239 7327
rect 7239 7293 7248 7327
rect 7196 7284 7248 7293
rect 2412 7216 2464 7268
rect 3700 7216 3752 7268
rect 5908 7216 5960 7268
rect 2964 7148 3016 7200
rect 3332 7148 3384 7200
rect 5540 7148 5592 7200
rect 6092 7191 6144 7200
rect 6092 7157 6101 7191
rect 6101 7157 6135 7191
rect 6135 7157 6144 7191
rect 7012 7191 7064 7200
rect 6092 7148 6144 7157
rect 7012 7157 7021 7191
rect 7021 7157 7055 7191
rect 7055 7157 7064 7191
rect 7012 7148 7064 7157
rect 11612 7395 11664 7404
rect 7932 7327 7984 7336
rect 7932 7293 7966 7327
rect 7966 7293 7984 7327
rect 7932 7284 7984 7293
rect 9312 7327 9364 7336
rect 9312 7293 9321 7327
rect 9321 7293 9355 7327
rect 9355 7293 9364 7327
rect 9312 7284 9364 7293
rect 11612 7361 11621 7395
rect 11621 7361 11655 7395
rect 11655 7361 11664 7395
rect 11612 7352 11664 7361
rect 10784 7216 10836 7268
rect 14096 7327 14148 7336
rect 14096 7293 14105 7327
rect 14105 7293 14139 7327
rect 14139 7293 14148 7327
rect 14096 7284 14148 7293
rect 16028 7284 16080 7336
rect 11612 7216 11664 7268
rect 9956 7148 10008 7200
rect 10692 7191 10744 7200
rect 10692 7157 10701 7191
rect 10701 7157 10735 7191
rect 10735 7157 10744 7191
rect 10692 7148 10744 7157
rect 11244 7148 11296 7200
rect 11336 7191 11388 7200
rect 11336 7157 11345 7191
rect 11345 7157 11379 7191
rect 11379 7157 11388 7191
rect 11336 7148 11388 7157
rect 12440 7191 12492 7200
rect 12440 7157 12449 7191
rect 12449 7157 12483 7191
rect 12483 7157 12492 7191
rect 12992 7191 13044 7200
rect 12440 7148 12492 7157
rect 12992 7157 13001 7191
rect 13001 7157 13035 7191
rect 13035 7157 13044 7191
rect 13636 7191 13688 7200
rect 12992 7148 13044 7157
rect 13636 7157 13645 7191
rect 13645 7157 13679 7191
rect 13679 7157 13688 7191
rect 13636 7148 13688 7157
rect 14740 7216 14792 7268
rect 17408 7216 17460 7268
rect 7912 7046 7964 7098
rect 7976 7046 8028 7098
rect 8040 7046 8092 7098
rect 8104 7046 8156 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 15035 7046 15087 7098
rect 5540 6944 5592 6996
rect 8852 6987 8904 6996
rect 8852 6953 8861 6987
rect 8861 6953 8895 6987
rect 8895 6953 8904 6987
rect 8852 6944 8904 6953
rect 12440 6944 12492 6996
rect 13636 6987 13688 6996
rect 13636 6953 13645 6987
rect 13645 6953 13679 6987
rect 13679 6953 13688 6987
rect 13636 6944 13688 6953
rect 3056 6876 3108 6928
rect 3240 6876 3292 6928
rect 3608 6876 3660 6928
rect 2872 6808 2924 6860
rect 3424 6851 3476 6860
rect 3424 6817 3433 6851
rect 3433 6817 3467 6851
rect 3467 6817 3476 6851
rect 3424 6808 3476 6817
rect 4344 6851 4396 6860
rect 4344 6817 4378 6851
rect 4378 6817 4396 6851
rect 4344 6808 4396 6817
rect 4620 6876 4672 6928
rect 11336 6876 11388 6928
rect 15200 6876 15252 6928
rect 6092 6851 6144 6860
rect 6092 6817 6101 6851
rect 6101 6817 6135 6851
rect 6135 6817 6144 6851
rect 6092 6808 6144 6817
rect 2320 6604 2372 6656
rect 2872 6604 2924 6656
rect 3792 6740 3844 6792
rect 3608 6604 3660 6656
rect 8484 6647 8536 6656
rect 8484 6613 8493 6647
rect 8493 6613 8527 6647
rect 8527 6613 8536 6647
rect 8484 6604 8536 6613
rect 9312 6604 9364 6656
rect 10508 6604 10560 6656
rect 11244 6808 11296 6860
rect 12164 6808 12216 6860
rect 11888 6740 11940 6792
rect 12440 6740 12492 6792
rect 13820 6783 13872 6792
rect 13820 6749 13829 6783
rect 13829 6749 13863 6783
rect 13863 6749 13872 6783
rect 13820 6740 13872 6749
rect 12532 6647 12584 6656
rect 12532 6613 12541 6647
rect 12541 6613 12575 6647
rect 12575 6613 12584 6647
rect 12532 6604 12584 6613
rect 14832 6783 14884 6792
rect 14832 6749 14841 6783
rect 14841 6749 14875 6783
rect 14875 6749 14884 6783
rect 14832 6740 14884 6749
rect 16488 6740 16540 6792
rect 15292 6672 15344 6724
rect 17224 6740 17276 6792
rect 14280 6604 14332 6656
rect 17684 6604 17736 6656
rect 4447 6502 4499 6554
rect 4511 6502 4563 6554
rect 4575 6502 4627 6554
rect 4639 6502 4691 6554
rect 11378 6502 11430 6554
rect 11442 6502 11494 6554
rect 11506 6502 11558 6554
rect 11570 6502 11622 6554
rect 18308 6502 18360 6554
rect 18372 6502 18424 6554
rect 18436 6502 18488 6554
rect 18500 6502 18552 6554
rect 2412 6400 2464 6452
rect 4068 6400 4120 6452
rect 12440 6400 12492 6452
rect 13820 6443 13872 6452
rect 13820 6409 13829 6443
rect 13829 6409 13863 6443
rect 13863 6409 13872 6443
rect 13820 6400 13872 6409
rect 14832 6400 14884 6452
rect 17408 6443 17460 6452
rect 17408 6409 17417 6443
rect 17417 6409 17451 6443
rect 17451 6409 17460 6443
rect 17408 6400 17460 6409
rect 9956 6375 10008 6384
rect 9956 6341 9965 6375
rect 9965 6341 9999 6375
rect 9999 6341 10008 6375
rect 9956 6332 10008 6341
rect 3056 6307 3108 6316
rect 3056 6273 3065 6307
rect 3065 6273 3099 6307
rect 3099 6273 3108 6307
rect 3056 6264 3108 6273
rect 4344 6264 4396 6316
rect 7472 6307 7524 6316
rect 7472 6273 7481 6307
rect 7481 6273 7515 6307
rect 7515 6273 7524 6307
rect 7472 6264 7524 6273
rect 3608 6196 3660 6248
rect 4712 6196 4764 6248
rect 2688 6128 2740 6180
rect 3792 6128 3844 6180
rect 3884 6128 3936 6180
rect 9312 6196 9364 6248
rect 10508 6239 10560 6248
rect 10508 6205 10517 6239
rect 10517 6205 10551 6239
rect 10551 6205 10560 6239
rect 10508 6196 10560 6205
rect 12348 6196 12400 6248
rect 13084 6196 13136 6248
rect 14096 6239 14148 6248
rect 14096 6205 14105 6239
rect 14105 6205 14139 6239
rect 14139 6205 14148 6239
rect 14096 6196 14148 6205
rect 16028 6239 16080 6248
rect 16028 6205 16037 6239
rect 16037 6205 16071 6239
rect 16071 6205 16080 6239
rect 16028 6196 16080 6205
rect 17684 6196 17736 6248
rect 5448 6128 5500 6180
rect 8208 6128 8260 6180
rect 2872 6060 2924 6112
rect 3056 6060 3108 6112
rect 3424 6060 3476 6112
rect 3976 6103 4028 6112
rect 3976 6069 3985 6103
rect 3985 6069 4019 6103
rect 4019 6069 4028 6103
rect 3976 6060 4028 6069
rect 4252 6060 4304 6112
rect 4712 6060 4764 6112
rect 6828 6103 6880 6112
rect 6828 6069 6837 6103
rect 6837 6069 6871 6103
rect 6871 6069 6880 6103
rect 6828 6060 6880 6069
rect 11796 6128 11848 6180
rect 17224 6128 17276 6180
rect 16948 6060 17000 6112
rect 18144 6060 18196 6112
rect 7912 5958 7964 6010
rect 7976 5958 8028 6010
rect 8040 5958 8092 6010
rect 8104 5958 8156 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 15035 5958 15087 6010
rect 1952 5899 2004 5908
rect 1952 5865 1961 5899
rect 1961 5865 1995 5899
rect 1995 5865 2004 5899
rect 1952 5856 2004 5865
rect 2320 5899 2372 5908
rect 2320 5865 2329 5899
rect 2329 5865 2363 5899
rect 2363 5865 2372 5899
rect 2320 5856 2372 5865
rect 3424 5899 3476 5908
rect 3424 5865 3433 5899
rect 3433 5865 3467 5899
rect 3467 5865 3476 5899
rect 3424 5856 3476 5865
rect 3516 5856 3568 5908
rect 3792 5720 3844 5772
rect 4896 5720 4948 5772
rect 7564 5788 7616 5840
rect 9956 5831 10008 5840
rect 9956 5797 9990 5831
rect 9990 5797 10008 5831
rect 9956 5788 10008 5797
rect 10692 5788 10744 5840
rect 15200 5856 15252 5908
rect 7012 5720 7064 5772
rect 7472 5763 7524 5772
rect 7472 5729 7481 5763
rect 7481 5729 7515 5763
rect 7515 5729 7524 5763
rect 7472 5720 7524 5729
rect 8668 5720 8720 5772
rect 10508 5720 10560 5772
rect 12164 5788 12216 5840
rect 12532 5788 12584 5840
rect 11980 5720 12032 5772
rect 12716 5763 12768 5772
rect 12716 5729 12725 5763
rect 12725 5729 12759 5763
rect 12759 5729 12768 5763
rect 12716 5720 12768 5729
rect 14280 5763 14332 5772
rect 14280 5729 14289 5763
rect 14289 5729 14323 5763
rect 14323 5729 14332 5763
rect 14280 5720 14332 5729
rect 17316 5720 17368 5772
rect 2412 5652 2464 5704
rect 3608 5695 3660 5704
rect 3608 5661 3617 5695
rect 3617 5661 3651 5695
rect 3651 5661 3660 5695
rect 3608 5652 3660 5661
rect 3884 5652 3936 5704
rect 4712 5695 4764 5704
rect 4712 5661 4721 5695
rect 4721 5661 4755 5695
rect 4755 5661 4764 5695
rect 4712 5652 4764 5661
rect 4804 5652 4856 5704
rect 5080 5652 5132 5704
rect 11796 5652 11848 5704
rect 13084 5652 13136 5704
rect 14464 5695 14516 5704
rect 14464 5661 14473 5695
rect 14473 5661 14507 5695
rect 14507 5661 14516 5695
rect 14464 5652 14516 5661
rect 16396 5652 16448 5704
rect 5632 5584 5684 5636
rect 3148 5516 3200 5568
rect 3792 5516 3844 5568
rect 4252 5516 4304 5568
rect 7472 5516 7524 5568
rect 8024 5516 8076 5568
rect 9220 5516 9272 5568
rect 16488 5584 16540 5636
rect 11060 5559 11112 5568
rect 11060 5525 11069 5559
rect 11069 5525 11103 5559
rect 11103 5525 11112 5559
rect 11060 5516 11112 5525
rect 12808 5516 12860 5568
rect 13268 5516 13320 5568
rect 16028 5516 16080 5568
rect 16396 5516 16448 5568
rect 17224 5516 17276 5568
rect 4447 5414 4499 5466
rect 4511 5414 4563 5466
rect 4575 5414 4627 5466
rect 4639 5414 4691 5466
rect 11378 5414 11430 5466
rect 11442 5414 11494 5466
rect 11506 5414 11558 5466
rect 11570 5414 11622 5466
rect 18308 5414 18360 5466
rect 18372 5414 18424 5466
rect 18436 5414 18488 5466
rect 18500 5414 18552 5466
rect 3976 5312 4028 5364
rect 6736 5312 6788 5364
rect 7472 5176 7524 5228
rect 7564 5219 7616 5228
rect 7564 5185 7573 5219
rect 7573 5185 7607 5219
rect 7607 5185 7616 5219
rect 11980 5312 12032 5364
rect 12164 5312 12216 5364
rect 13268 5312 13320 5364
rect 18144 5312 18196 5364
rect 7564 5176 7616 5185
rect 8668 5219 8720 5228
rect 8668 5185 8677 5219
rect 8677 5185 8711 5219
rect 8711 5185 8720 5219
rect 8668 5176 8720 5185
rect 9956 5219 10008 5228
rect 9956 5185 9965 5219
rect 9965 5185 9999 5219
rect 9999 5185 10008 5219
rect 9956 5176 10008 5185
rect 12992 5244 13044 5296
rect 16396 5244 16448 5296
rect 11060 5176 11112 5228
rect 12716 5176 12768 5228
rect 13360 5176 13412 5228
rect 14096 5176 14148 5228
rect 14372 5176 14424 5228
rect 16580 5176 16632 5228
rect 17224 5219 17276 5228
rect 17224 5185 17233 5219
rect 17233 5185 17267 5219
rect 17267 5185 17276 5219
rect 17224 5176 17276 5185
rect 3516 5108 3568 5160
rect 3884 5151 3936 5160
rect 3884 5117 3893 5151
rect 3893 5117 3927 5151
rect 3927 5117 3936 5151
rect 3884 5108 3936 5117
rect 6828 5108 6880 5160
rect 9864 5108 9916 5160
rect 3884 4972 3936 5024
rect 4896 4972 4948 5024
rect 7012 4972 7064 5024
rect 7288 4972 7340 5024
rect 8208 4972 8260 5024
rect 9772 5015 9824 5024
rect 9772 4981 9781 5015
rect 9781 4981 9815 5015
rect 9815 4981 9824 5015
rect 9772 4972 9824 4981
rect 16120 5108 16172 5160
rect 20628 5108 20680 5160
rect 15384 5040 15436 5092
rect 11796 4972 11848 5024
rect 12440 4972 12492 5024
rect 13176 5015 13228 5024
rect 13176 4981 13185 5015
rect 13185 4981 13219 5015
rect 13219 4981 13228 5015
rect 13176 4972 13228 4981
rect 15568 5015 15620 5024
rect 15568 4981 15577 5015
rect 15577 4981 15611 5015
rect 15611 4981 15620 5015
rect 15568 4972 15620 4981
rect 16028 5015 16080 5024
rect 16028 4981 16037 5015
rect 16037 4981 16071 5015
rect 16071 4981 16080 5015
rect 16028 4972 16080 4981
rect 21272 4972 21324 5024
rect 7912 4870 7964 4922
rect 7976 4870 8028 4922
rect 8040 4870 8092 4922
rect 8104 4870 8156 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 15035 4870 15087 4922
rect 1492 4811 1544 4820
rect 1492 4777 1501 4811
rect 1501 4777 1535 4811
rect 1535 4777 1544 4811
rect 1492 4768 1544 4777
rect 4068 4768 4120 4820
rect 5632 4768 5684 4820
rect 5724 4768 5776 4820
rect 6736 4811 6788 4820
rect 6736 4777 6745 4811
rect 6745 4777 6779 4811
rect 6779 4777 6788 4811
rect 6736 4768 6788 4777
rect 8208 4768 8260 4820
rect 9956 4768 10008 4820
rect 10876 4768 10928 4820
rect 14372 4768 14424 4820
rect 15568 4768 15620 4820
rect 20628 4768 20680 4820
rect 3976 4700 4028 4752
rect 7380 4700 7432 4752
rect 7472 4743 7524 4752
rect 7472 4709 7481 4743
rect 7481 4709 7515 4743
rect 7515 4709 7524 4743
rect 7472 4700 7524 4709
rect 1492 4632 1544 4684
rect 6276 4632 6328 4684
rect 2504 4607 2556 4616
rect 2504 4573 2513 4607
rect 2513 4573 2547 4607
rect 2547 4573 2556 4607
rect 2504 4564 2556 4573
rect 3332 4607 3384 4616
rect 3332 4573 3341 4607
rect 3341 4573 3375 4607
rect 3375 4573 3384 4607
rect 3332 4564 3384 4573
rect 3424 4607 3476 4616
rect 3424 4573 3433 4607
rect 3433 4573 3467 4607
rect 3467 4573 3476 4607
rect 3424 4564 3476 4573
rect 5264 4564 5316 4616
rect 5908 4607 5960 4616
rect 5908 4573 5917 4607
rect 5917 4573 5951 4607
rect 5951 4573 5960 4607
rect 5908 4564 5960 4573
rect 6092 4564 6144 4616
rect 7288 4632 7340 4684
rect 8116 4675 8168 4684
rect 6920 4564 6972 4616
rect 8116 4641 8125 4675
rect 8125 4641 8159 4675
rect 8159 4641 8168 4675
rect 8116 4632 8168 4641
rect 10140 4675 10192 4684
rect 10140 4641 10149 4675
rect 10149 4641 10183 4675
rect 10183 4641 10192 4675
rect 10140 4632 10192 4641
rect 11060 4700 11112 4752
rect 16028 4700 16080 4752
rect 13636 4632 13688 4684
rect 15752 4632 15804 4684
rect 16396 4700 16448 4752
rect 16580 4632 16632 4684
rect 17132 4632 17184 4684
rect 17960 4675 18012 4684
rect 17960 4641 17969 4675
rect 17969 4641 18003 4675
rect 18003 4641 18012 4675
rect 17960 4632 18012 4641
rect 7656 4607 7708 4616
rect 7656 4573 7665 4607
rect 7665 4573 7699 4607
rect 7699 4573 7708 4607
rect 7656 4564 7708 4573
rect 8208 4564 8260 4616
rect 4068 4496 4120 4548
rect 9312 4564 9364 4616
rect 10508 4607 10560 4616
rect 10508 4573 10517 4607
rect 10517 4573 10551 4607
rect 10551 4573 10560 4607
rect 10508 4564 10560 4573
rect 3148 4428 3200 4480
rect 4896 4471 4948 4480
rect 4896 4437 4905 4471
rect 4905 4437 4939 4471
rect 4939 4437 4948 4471
rect 4896 4428 4948 4437
rect 6184 4428 6236 4480
rect 9772 4496 9824 4548
rect 10140 4496 10192 4548
rect 8392 4428 8444 4480
rect 9680 4471 9732 4480
rect 9680 4437 9689 4471
rect 9689 4437 9723 4471
rect 9723 4437 9732 4471
rect 9680 4428 9732 4437
rect 12440 4428 12492 4480
rect 17316 4539 17368 4548
rect 17316 4505 17325 4539
rect 17325 4505 17359 4539
rect 17359 4505 17368 4539
rect 17316 4496 17368 4505
rect 13820 4428 13872 4480
rect 14188 4471 14240 4480
rect 14188 4437 14197 4471
rect 14197 4437 14231 4471
rect 14231 4437 14240 4471
rect 14188 4428 14240 4437
rect 16856 4428 16908 4480
rect 4447 4326 4499 4378
rect 4511 4326 4563 4378
rect 4575 4326 4627 4378
rect 4639 4326 4691 4378
rect 11378 4326 11430 4378
rect 11442 4326 11494 4378
rect 11506 4326 11558 4378
rect 11570 4326 11622 4378
rect 18308 4326 18360 4378
rect 18372 4326 18424 4378
rect 18436 4326 18488 4378
rect 18500 4326 18552 4378
rect 3424 4224 3476 4276
rect 4896 4224 4948 4276
rect 5264 4267 5316 4276
rect 1492 4131 1544 4140
rect 1492 4097 1501 4131
rect 1501 4097 1535 4131
rect 1535 4097 1544 4131
rect 1492 4088 1544 4097
rect 5264 4233 5273 4267
rect 5273 4233 5307 4267
rect 5307 4233 5316 4267
rect 5264 4224 5316 4233
rect 5540 4224 5592 4276
rect 1952 4063 2004 4072
rect 1952 4029 1961 4063
rect 1961 4029 1995 4063
rect 1995 4029 2004 4063
rect 1952 4020 2004 4029
rect 1492 3952 1544 4004
rect 2688 4020 2740 4072
rect 5540 4088 5592 4140
rect 6460 4224 6512 4276
rect 7564 4224 7616 4276
rect 10876 4224 10928 4276
rect 17132 4267 17184 4276
rect 6276 4131 6328 4140
rect 5632 4063 5684 4072
rect 2504 3952 2556 4004
rect 5632 4029 5641 4063
rect 5641 4029 5675 4063
rect 5675 4029 5684 4063
rect 5632 4020 5684 4029
rect 5172 3952 5224 4004
rect 1308 3884 1360 3936
rect 5632 3884 5684 3936
rect 6276 4097 6285 4131
rect 6285 4097 6319 4131
rect 6319 4097 6328 4131
rect 6276 4088 6328 4097
rect 6828 4131 6880 4140
rect 6828 4097 6837 4131
rect 6837 4097 6871 4131
rect 6871 4097 6880 4131
rect 6828 4088 6880 4097
rect 8116 4088 8168 4140
rect 6644 3952 6696 4004
rect 7380 4020 7432 4072
rect 8208 4020 8260 4072
rect 8392 4020 8444 4072
rect 10416 4131 10468 4140
rect 10416 4097 10425 4131
rect 10425 4097 10459 4131
rect 10459 4097 10468 4131
rect 10416 4088 10468 4097
rect 11428 4131 11480 4140
rect 11428 4097 11437 4131
rect 11437 4097 11471 4131
rect 11471 4097 11480 4131
rect 11428 4088 11480 4097
rect 12440 4156 12492 4208
rect 17132 4233 17141 4267
rect 17141 4233 17175 4267
rect 17175 4233 17184 4267
rect 17132 4224 17184 4233
rect 15752 4131 15804 4140
rect 10600 4020 10652 4072
rect 12072 4020 12124 4072
rect 12348 4020 12400 4072
rect 15752 4097 15761 4131
rect 15761 4097 15795 4131
rect 15795 4097 15804 4131
rect 15752 4088 15804 4097
rect 17960 4088 18012 4140
rect 13820 4020 13872 4072
rect 7564 3952 7616 4004
rect 9312 3995 9364 4004
rect 9312 3961 9321 3995
rect 9321 3961 9355 3995
rect 9355 3961 9364 3995
rect 9312 3952 9364 3961
rect 9772 3952 9824 4004
rect 10508 3952 10560 4004
rect 14188 4020 14240 4072
rect 14372 4063 14424 4072
rect 14372 4029 14395 4063
rect 14395 4029 14424 4063
rect 14372 4020 14424 4029
rect 8484 3927 8536 3936
rect 8484 3893 8493 3927
rect 8493 3893 8527 3927
rect 8527 3893 8536 3927
rect 8484 3884 8536 3893
rect 9128 3884 9180 3936
rect 9864 3927 9916 3936
rect 9864 3893 9873 3927
rect 9873 3893 9907 3927
rect 9907 3893 9916 3927
rect 9864 3884 9916 3893
rect 10232 3927 10284 3936
rect 10232 3893 10241 3927
rect 10241 3893 10275 3927
rect 10275 3893 10284 3927
rect 10232 3884 10284 3893
rect 10968 3927 11020 3936
rect 10968 3893 10977 3927
rect 10977 3893 11011 3927
rect 11011 3893 11020 3927
rect 10968 3884 11020 3893
rect 11244 3884 11296 3936
rect 13636 3884 13688 3936
rect 15844 3952 15896 4004
rect 21824 3884 21876 3936
rect 7912 3782 7964 3834
rect 7976 3782 8028 3834
rect 8040 3782 8092 3834
rect 8104 3782 8156 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 15035 3782 15087 3834
rect 3332 3680 3384 3732
rect 6644 3680 6696 3732
rect 2412 3612 2464 3664
rect 8484 3680 8536 3732
rect 10140 3723 10192 3732
rect 10140 3689 10149 3723
rect 10149 3689 10183 3723
rect 10183 3689 10192 3723
rect 10140 3680 10192 3689
rect 11428 3723 11480 3732
rect 11428 3689 11437 3723
rect 11437 3689 11471 3723
rect 11471 3689 11480 3723
rect 11428 3680 11480 3689
rect 13176 3723 13228 3732
rect 13176 3689 13185 3723
rect 13185 3689 13219 3723
rect 13219 3689 13228 3723
rect 13176 3680 13228 3689
rect 14096 3680 14148 3732
rect 1492 3587 1544 3596
rect 1492 3553 1501 3587
rect 1501 3553 1535 3587
rect 1535 3553 1544 3587
rect 1492 3544 1544 3553
rect 2872 3544 2924 3596
rect 3148 3587 3200 3596
rect 3148 3553 3157 3587
rect 3157 3553 3191 3587
rect 3191 3553 3200 3587
rect 3148 3544 3200 3553
rect 4344 3544 4396 3596
rect 5172 3587 5224 3596
rect 5172 3553 5181 3587
rect 5181 3553 5215 3587
rect 5215 3553 5224 3587
rect 5172 3544 5224 3553
rect 5908 3544 5960 3596
rect 6368 3544 6420 3596
rect 7012 3612 7064 3664
rect 7380 3544 7432 3596
rect 7564 3544 7616 3596
rect 9220 3544 9272 3596
rect 9496 3544 9548 3596
rect 9680 3544 9732 3596
rect 10048 3587 10100 3596
rect 10048 3553 10057 3587
rect 10057 3553 10091 3587
rect 10091 3553 10100 3587
rect 10048 3544 10100 3553
rect 10968 3612 11020 3664
rect 15476 3544 15528 3596
rect 3424 3519 3476 3528
rect 3424 3485 3433 3519
rect 3433 3485 3467 3519
rect 3467 3485 3476 3519
rect 3424 3476 3476 3485
rect 3608 3476 3660 3528
rect 2504 3408 2556 3460
rect 6460 3476 6512 3528
rect 7472 3519 7524 3528
rect 7472 3485 7481 3519
rect 7481 3485 7515 3519
rect 7515 3485 7524 3519
rect 7472 3476 7524 3485
rect 10876 3476 10928 3528
rect 13268 3476 13320 3528
rect 13636 3476 13688 3528
rect 3240 3340 3292 3392
rect 4896 3340 4948 3392
rect 5080 3340 5132 3392
rect 7288 3340 7340 3392
rect 10416 3408 10468 3460
rect 14372 3519 14424 3528
rect 14372 3485 14381 3519
rect 14381 3485 14415 3519
rect 14415 3485 14424 3519
rect 14372 3476 14424 3485
rect 14740 3476 14792 3528
rect 16856 3544 16908 3596
rect 17500 3587 17552 3596
rect 17500 3553 17509 3587
rect 17509 3553 17543 3587
rect 17543 3553 17552 3587
rect 17500 3544 17552 3553
rect 19708 3587 19760 3596
rect 19708 3553 19717 3587
rect 19717 3553 19751 3587
rect 19751 3553 19760 3587
rect 19708 3544 19760 3553
rect 21824 3544 21876 3596
rect 18052 3476 18104 3528
rect 9680 3383 9732 3392
rect 9680 3349 9689 3383
rect 9689 3349 9723 3383
rect 9723 3349 9732 3383
rect 9680 3340 9732 3349
rect 10048 3340 10100 3392
rect 10692 3383 10744 3392
rect 10692 3349 10701 3383
rect 10701 3349 10735 3383
rect 10735 3349 10744 3383
rect 10692 3340 10744 3349
rect 13728 3340 13780 3392
rect 13820 3383 13872 3392
rect 13820 3349 13829 3383
rect 13829 3349 13863 3383
rect 13863 3349 13872 3383
rect 13820 3340 13872 3349
rect 15660 3340 15712 3392
rect 16488 3340 16540 3392
rect 18144 3340 18196 3392
rect 20904 3340 20956 3392
rect 22284 3340 22336 3392
rect 4447 3238 4499 3290
rect 4511 3238 4563 3290
rect 4575 3238 4627 3290
rect 4639 3238 4691 3290
rect 11378 3238 11430 3290
rect 11442 3238 11494 3290
rect 11506 3238 11558 3290
rect 11570 3238 11622 3290
rect 18308 3238 18360 3290
rect 18372 3238 18424 3290
rect 18436 3238 18488 3290
rect 18500 3238 18552 3290
rect 3608 3136 3660 3188
rect 1952 3068 2004 3120
rect 204 2932 256 2984
rect 1308 2932 1360 2984
rect 2872 3043 2924 3052
rect 2872 3009 2881 3043
rect 2881 3009 2915 3043
rect 2915 3009 2924 3043
rect 2872 3000 2924 3009
rect 5172 3136 5224 3188
rect 9496 3136 9548 3188
rect 10324 3136 10376 3188
rect 12256 3136 12308 3188
rect 13820 3136 13872 3188
rect 7472 3043 7524 3052
rect 7472 3009 7481 3043
rect 7481 3009 7515 3043
rect 7515 3009 7524 3043
rect 7472 3000 7524 3009
rect 7564 3000 7616 3052
rect 5080 2932 5132 2984
rect 5540 2932 5592 2984
rect 1032 2796 1084 2848
rect 6092 2864 6144 2916
rect 7012 2864 7064 2916
rect 2872 2796 2924 2848
rect 6368 2839 6420 2848
rect 6368 2805 6377 2839
rect 6377 2805 6411 2839
rect 6411 2805 6420 2839
rect 6368 2796 6420 2805
rect 6828 2796 6880 2848
rect 7196 2796 7248 2848
rect 8392 2864 8444 2916
rect 10876 3000 10928 3052
rect 13728 3000 13780 3052
rect 14740 3043 14792 3052
rect 9864 2932 9916 2984
rect 12440 2975 12492 2984
rect 12440 2941 12449 2975
rect 12449 2941 12483 2975
rect 12483 2941 12492 2975
rect 12440 2932 12492 2941
rect 12808 2932 12860 2984
rect 13268 2932 13320 2984
rect 14740 3009 14749 3043
rect 14749 3009 14783 3043
rect 14783 3009 14792 3043
rect 14740 3000 14792 3009
rect 15844 3043 15896 3052
rect 15844 3009 15853 3043
rect 15853 3009 15887 3043
rect 15887 3009 15896 3043
rect 15844 3000 15896 3009
rect 20720 3043 20772 3052
rect 20720 3009 20729 3043
rect 20729 3009 20763 3043
rect 20763 3009 20772 3043
rect 20720 3000 20772 3009
rect 16948 2975 17000 2984
rect 16948 2941 16957 2975
rect 16957 2941 16991 2975
rect 16991 2941 17000 2975
rect 16948 2932 17000 2941
rect 18052 2975 18104 2984
rect 18052 2941 18061 2975
rect 18061 2941 18095 2975
rect 18095 2941 18104 2975
rect 18052 2932 18104 2941
rect 18604 2975 18656 2984
rect 18604 2941 18613 2975
rect 18613 2941 18647 2975
rect 18647 2941 18656 2975
rect 18604 2932 18656 2941
rect 21364 2932 21416 2984
rect 10692 2864 10744 2916
rect 11888 2864 11940 2916
rect 12716 2907 12768 2916
rect 12716 2873 12725 2907
rect 12725 2873 12759 2907
rect 12759 2873 12768 2907
rect 12716 2864 12768 2873
rect 13728 2864 13780 2916
rect 8300 2839 8352 2848
rect 8300 2805 8309 2839
rect 8309 2805 8343 2839
rect 8343 2805 8352 2839
rect 8300 2796 8352 2805
rect 10416 2839 10468 2848
rect 10416 2805 10425 2839
rect 10425 2805 10459 2839
rect 10459 2805 10468 2839
rect 10416 2796 10468 2805
rect 10876 2839 10928 2848
rect 10876 2805 10885 2839
rect 10885 2805 10919 2839
rect 10919 2805 10928 2839
rect 10876 2796 10928 2805
rect 12164 2796 12216 2848
rect 13912 2796 13964 2848
rect 16396 2864 16448 2916
rect 17408 2864 17460 2916
rect 16948 2796 17000 2848
rect 17500 2796 17552 2848
rect 18696 2796 18748 2848
rect 7912 2694 7964 2746
rect 7976 2694 8028 2746
rect 8040 2694 8092 2746
rect 8104 2694 8156 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 15035 2694 15087 2746
rect 4344 2592 4396 2644
rect 6184 2635 6236 2644
rect 2780 2456 2832 2508
rect 3976 2456 4028 2508
rect 6184 2601 6193 2635
rect 6193 2601 6227 2635
rect 6227 2601 6236 2635
rect 6184 2592 6236 2601
rect 7288 2635 7340 2644
rect 7288 2601 7297 2635
rect 7297 2601 7331 2635
rect 7331 2601 7340 2635
rect 7288 2592 7340 2601
rect 8392 2635 8444 2644
rect 8392 2601 8401 2635
rect 8401 2601 8435 2635
rect 8435 2601 8444 2635
rect 8392 2592 8444 2601
rect 9128 2635 9180 2644
rect 9128 2601 9137 2635
rect 9137 2601 9171 2635
rect 9171 2601 9180 2635
rect 9128 2592 9180 2601
rect 9772 2635 9824 2644
rect 9772 2601 9781 2635
rect 9781 2601 9815 2635
rect 9815 2601 9824 2635
rect 9772 2592 9824 2601
rect 10416 2592 10468 2644
rect 16948 2635 17000 2644
rect 16948 2601 16957 2635
rect 16957 2601 16991 2635
rect 16991 2601 17000 2635
rect 16948 2592 17000 2601
rect 7196 2524 7248 2576
rect 8300 2524 8352 2576
rect 9680 2524 9732 2576
rect 12440 2524 12492 2576
rect 11888 2499 11940 2508
rect 11888 2465 11897 2499
rect 11897 2465 11931 2499
rect 11931 2465 11940 2499
rect 11888 2456 11940 2465
rect 12624 2499 12676 2508
rect 12624 2465 12633 2499
rect 12633 2465 12667 2499
rect 12667 2465 12676 2499
rect 12624 2456 12676 2465
rect 12716 2456 12768 2508
rect 13728 2499 13780 2508
rect 13728 2465 13737 2499
rect 13737 2465 13771 2499
rect 13771 2465 13780 2499
rect 13728 2456 13780 2465
rect 14464 2456 14516 2508
rect 15292 2456 15344 2508
rect 15384 2456 15436 2508
rect 16396 2499 16448 2508
rect 16396 2465 16405 2499
rect 16405 2465 16439 2499
rect 16439 2465 16448 2499
rect 16396 2456 16448 2465
rect 17408 2499 17460 2508
rect 17408 2465 17417 2499
rect 17417 2465 17451 2499
rect 17451 2465 17460 2499
rect 17408 2456 17460 2465
rect 3424 2431 3476 2440
rect 3424 2397 3433 2431
rect 3433 2397 3467 2431
rect 3467 2397 3476 2431
rect 3424 2388 3476 2397
rect 6644 2388 6696 2440
rect 6828 2388 6880 2440
rect 9220 2388 9272 2440
rect 1952 2252 2004 2304
rect 6920 2320 6972 2372
rect 10232 2320 10284 2372
rect 6736 2252 6788 2304
rect 7196 2252 7248 2304
rect 7932 2295 7984 2304
rect 7932 2261 7941 2295
rect 7941 2261 7975 2295
rect 7975 2261 7984 2295
rect 7932 2252 7984 2261
rect 8392 2252 8444 2304
rect 10876 2252 10928 2304
rect 12532 2252 12584 2304
rect 12992 2252 13044 2304
rect 13452 2252 13504 2304
rect 14280 2252 14332 2304
rect 14740 2252 14792 2304
rect 15200 2252 15252 2304
rect 16120 2252 16172 2304
rect 16948 2252 17000 2304
rect 17868 2252 17920 2304
rect 21364 2295 21416 2304
rect 21364 2261 21373 2295
rect 21373 2261 21407 2295
rect 21407 2261 21416 2295
rect 21364 2252 21416 2261
rect 22744 2252 22796 2304
rect 4447 2150 4499 2202
rect 4511 2150 4563 2202
rect 4575 2150 4627 2202
rect 4639 2150 4691 2202
rect 11378 2150 11430 2202
rect 11442 2150 11494 2202
rect 11506 2150 11558 2202
rect 11570 2150 11622 2202
rect 18308 2150 18360 2202
rect 18372 2150 18424 2202
rect 18436 2150 18488 2202
rect 18500 2150 18552 2202
rect 1492 2048 1544 2100
rect 7380 2048 7432 2100
rect 7932 2048 7984 2100
rect 572 1980 624 2032
rect 7012 1980 7064 2032
<< metal2 >>
rect 2870 22672 2926 22681
rect 2870 22607 2926 22616
rect 2778 21312 2834 21321
rect 2778 21247 2834 21256
rect 1950 20768 2006 20777
rect 1950 20703 2006 20712
rect 1964 20602 1992 20703
rect 2792 20602 2820 21247
rect 1952 20596 2004 20602
rect 1952 20538 2004 20544
rect 2780 20596 2832 20602
rect 2780 20538 2832 20544
rect 2596 20392 2648 20398
rect 2596 20334 2648 20340
rect 2778 20360 2834 20369
rect 2504 19916 2556 19922
rect 2504 19858 2556 19864
rect 2042 19816 2098 19825
rect 2042 19751 2044 19760
rect 2096 19751 2098 19760
rect 2044 19722 2096 19728
rect 1952 19440 2004 19446
rect 1950 19408 1952 19417
rect 2004 19408 2006 19417
rect 2516 19378 2544 19858
rect 1950 19343 2006 19352
rect 2504 19372 2556 19378
rect 2504 19314 2556 19320
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 1964 18873 1992 18906
rect 2608 18902 2636 20334
rect 2778 20295 2834 20304
rect 2792 20058 2820 20295
rect 2780 20052 2832 20058
rect 2780 19994 2832 20000
rect 2780 19848 2832 19854
rect 2780 19790 2832 19796
rect 2596 18896 2648 18902
rect 1950 18864 2006 18873
rect 1768 18828 1820 18834
rect 2596 18838 2648 18844
rect 1950 18799 2006 18808
rect 1768 18770 1820 18776
rect 1780 17814 1808 18770
rect 1858 18456 1914 18465
rect 1858 18391 1914 18400
rect 1872 17882 1900 18391
rect 2792 18290 2820 19790
rect 2780 18284 2832 18290
rect 2780 18226 2832 18232
rect 2688 18216 2740 18222
rect 2688 18158 2740 18164
rect 1952 18080 2004 18086
rect 1950 18048 1952 18057
rect 2004 18048 2006 18057
rect 1950 17983 2006 17992
rect 1860 17876 1912 17882
rect 1860 17818 1912 17824
rect 1768 17808 1820 17814
rect 1768 17750 1820 17756
rect 1676 17740 1728 17746
rect 1676 17682 1728 17688
rect 1688 16726 1716 17682
rect 1950 17504 2006 17513
rect 1950 17439 2006 17448
rect 1964 17338 1992 17439
rect 1952 17332 2004 17338
rect 1952 17274 2004 17280
rect 1676 16720 1728 16726
rect 1676 16662 1728 16668
rect 1950 16552 2006 16561
rect 1950 16487 2006 16496
rect 1964 16250 1992 16487
rect 1952 16244 2004 16250
rect 1952 16186 2004 16192
rect 1674 16144 1730 16153
rect 1674 16079 1730 16088
rect 1688 15706 1716 16079
rect 1768 16040 1820 16046
rect 1768 15982 1820 15988
rect 2320 16040 2372 16046
rect 2320 15982 2372 15988
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 1780 15026 1808 15982
rect 2332 15638 2360 15982
rect 2320 15632 2372 15638
rect 1858 15600 1914 15609
rect 2320 15574 2372 15580
rect 1858 15535 1914 15544
rect 1872 15162 1900 15535
rect 2596 15496 2648 15502
rect 2596 15438 2648 15444
rect 1860 15156 1912 15162
rect 1860 15098 1912 15104
rect 1768 15020 1820 15026
rect 1768 14962 1820 14968
rect 1676 14952 1728 14958
rect 1676 14894 1728 14900
rect 1688 14414 1716 14894
rect 1768 14476 1820 14482
rect 1768 14418 1820 14424
rect 1676 14408 1728 14414
rect 1676 14350 1728 14356
rect 1584 13864 1636 13870
rect 1584 13806 1636 13812
rect 1490 13288 1546 13297
rect 1490 13223 1546 13232
rect 1504 12442 1532 13223
rect 1596 12986 1624 13806
rect 1780 13462 1808 14418
rect 1952 14272 2004 14278
rect 1950 14240 1952 14249
rect 2004 14240 2006 14249
rect 1950 14175 2006 14184
rect 2608 13802 2636 15438
rect 2596 13796 2648 13802
rect 2596 13738 2648 13744
rect 1768 13456 1820 13462
rect 1768 13398 1820 13404
rect 1952 13388 2004 13394
rect 1952 13330 2004 13336
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 1492 12436 1544 12442
rect 1492 12378 1544 12384
rect 1860 9376 1912 9382
rect 1860 9318 1912 9324
rect 1872 8430 1900 9318
rect 1860 8424 1912 8430
rect 1860 8366 1912 8372
rect 1584 8288 1636 8294
rect 1584 8230 1636 8236
rect 1596 7954 1624 8230
rect 1584 7948 1636 7954
rect 1584 7890 1636 7896
rect 1490 4856 1546 4865
rect 1490 4791 1492 4800
rect 1544 4791 1546 4800
rect 1492 4762 1544 4768
rect 1492 4684 1544 4690
rect 1492 4626 1544 4632
rect 1504 4146 1532 4626
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 1492 4004 1544 4010
rect 1492 3946 1544 3952
rect 1308 3936 1360 3942
rect 1308 3878 1360 3884
rect 1320 2990 1348 3878
rect 1504 3602 1532 3946
rect 1492 3596 1544 3602
rect 1492 3538 1544 3544
rect 204 2984 256 2990
rect 204 2926 256 2932
rect 1308 2984 1360 2990
rect 1308 2926 1360 2932
rect 216 800 244 2926
rect 1032 2848 1084 2854
rect 1032 2790 1084 2796
rect 572 2032 624 2038
rect 572 1974 624 1980
rect 584 800 612 1974
rect 1044 800 1072 2790
rect 1492 2100 1544 2106
rect 1492 2042 1544 2048
rect 1504 800 1532 2042
rect 1596 2009 1624 7890
rect 1872 7342 1900 8366
rect 1860 7336 1912 7342
rect 1860 7278 1912 7284
rect 1872 5794 1900 7278
rect 1964 5914 1992 13330
rect 2596 12640 2648 12646
rect 2596 12582 2648 12588
rect 2044 12300 2096 12306
rect 2044 12242 2096 12248
rect 2056 11694 2084 12242
rect 2608 11898 2636 12582
rect 2700 11898 2728 18158
rect 2778 17096 2834 17105
rect 2778 17031 2834 17040
rect 2792 16250 2820 17031
rect 2780 16244 2832 16250
rect 2780 16186 2832 16192
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 2792 13938 2820 14418
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 2884 13734 2912 22607
rect 3698 22264 3754 22273
rect 3698 22199 3754 22208
rect 3712 21826 3740 22199
rect 3700 21820 3752 21826
rect 3700 21762 3752 21768
rect 10784 21820 10836 21826
rect 10784 21762 10836 21768
rect 3146 21720 3202 21729
rect 3146 21655 3202 21664
rect 3160 20058 3188 21655
rect 4421 20700 4717 20720
rect 4477 20698 4501 20700
rect 4557 20698 4581 20700
rect 4637 20698 4661 20700
rect 4499 20646 4501 20698
rect 4563 20646 4575 20698
rect 4637 20646 4639 20698
rect 4477 20644 4501 20646
rect 4557 20644 4581 20646
rect 4637 20644 4661 20646
rect 4421 20624 4717 20644
rect 3240 20324 3292 20330
rect 3240 20266 3292 20272
rect 3148 20052 3200 20058
rect 3148 19994 3200 20000
rect 2964 19916 3016 19922
rect 2964 19858 3016 19864
rect 2976 18902 3004 19858
rect 3252 19378 3280 20266
rect 7886 20156 8182 20176
rect 7942 20154 7966 20156
rect 8022 20154 8046 20156
rect 8102 20154 8126 20156
rect 7964 20102 7966 20154
rect 8028 20102 8040 20154
rect 8102 20102 8104 20154
rect 7942 20100 7966 20102
rect 8022 20100 8046 20102
rect 8102 20100 8126 20102
rect 7886 20080 8182 20100
rect 4421 19612 4717 19632
rect 4477 19610 4501 19612
rect 4557 19610 4581 19612
rect 4637 19610 4661 19612
rect 4499 19558 4501 19610
rect 4563 19558 4575 19610
rect 4637 19558 4639 19610
rect 4477 19556 4501 19558
rect 4557 19556 4581 19558
rect 4637 19556 4661 19558
rect 4421 19536 4717 19556
rect 3240 19372 3292 19378
rect 3240 19314 3292 19320
rect 8944 19304 8996 19310
rect 8944 19246 8996 19252
rect 3240 19236 3292 19242
rect 3240 19178 3292 19184
rect 2964 18896 3016 18902
rect 2964 18838 3016 18844
rect 3252 17814 3280 19178
rect 7886 19068 8182 19088
rect 7942 19066 7966 19068
rect 8022 19066 8046 19068
rect 8102 19066 8126 19068
rect 7964 19014 7966 19066
rect 8028 19014 8040 19066
rect 8102 19014 8104 19066
rect 7942 19012 7966 19014
rect 8022 19012 8046 19014
rect 8102 19012 8126 19014
rect 7886 18992 8182 19012
rect 5632 18760 5684 18766
rect 5632 18702 5684 18708
rect 4421 18524 4717 18544
rect 4477 18522 4501 18524
rect 4557 18522 4581 18524
rect 4637 18522 4661 18524
rect 4499 18470 4501 18522
rect 4563 18470 4575 18522
rect 4637 18470 4639 18522
rect 4477 18468 4501 18470
rect 4557 18468 4581 18470
rect 4637 18468 4661 18470
rect 4421 18448 4717 18468
rect 3332 18148 3384 18154
rect 3332 18090 3384 18096
rect 3240 17808 3292 17814
rect 3240 17750 3292 17756
rect 3344 17202 3372 18090
rect 5644 17882 5672 18702
rect 7886 17980 8182 18000
rect 7942 17978 7966 17980
rect 8022 17978 8046 17980
rect 8102 17978 8126 17980
rect 7964 17926 7966 17978
rect 8028 17926 8040 17978
rect 8102 17926 8104 17978
rect 7942 17924 7966 17926
rect 8022 17924 8046 17926
rect 8102 17924 8126 17926
rect 7886 17904 8182 17924
rect 5632 17876 5684 17882
rect 5632 17818 5684 17824
rect 5540 17808 5592 17814
rect 5540 17750 5592 17756
rect 4068 17672 4120 17678
rect 4068 17614 4120 17620
rect 3332 17196 3384 17202
rect 3332 17138 3384 17144
rect 4080 17134 4108 17614
rect 4421 17436 4717 17456
rect 4477 17434 4501 17436
rect 4557 17434 4581 17436
rect 4637 17434 4661 17436
rect 4499 17382 4501 17434
rect 4563 17382 4575 17434
rect 4637 17382 4639 17434
rect 4477 17380 4501 17382
rect 4557 17380 4581 17382
rect 4637 17380 4661 17382
rect 4421 17360 4717 17380
rect 2964 17128 3016 17134
rect 2964 17070 3016 17076
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 2976 16794 3004 17070
rect 2964 16788 3016 16794
rect 2964 16730 3016 16736
rect 4080 16590 4108 17070
rect 5448 17060 5500 17066
rect 5448 17002 5500 17008
rect 4160 16992 4212 16998
rect 4160 16934 4212 16940
rect 4172 16658 4200 16934
rect 5460 16794 5488 17002
rect 5552 16998 5580 17750
rect 7564 17740 7616 17746
rect 7564 17682 7616 17688
rect 8208 17740 8260 17746
rect 8208 17682 8260 17688
rect 6460 17536 6512 17542
rect 6460 17478 6512 17484
rect 6472 17202 6500 17478
rect 6460 17196 6512 17202
rect 6460 17138 6512 17144
rect 5724 17128 5776 17134
rect 5724 17070 5776 17076
rect 5540 16992 5592 16998
rect 5540 16934 5592 16940
rect 5448 16788 5500 16794
rect 5448 16730 5500 16736
rect 4252 16720 4304 16726
rect 4252 16662 4304 16668
rect 4160 16652 4212 16658
rect 4160 16594 4212 16600
rect 3424 16584 3476 16590
rect 3424 16526 3476 16532
rect 4068 16584 4120 16590
rect 4068 16526 4120 16532
rect 3436 15706 3464 16526
rect 4080 16046 4108 16526
rect 4264 16114 4292 16662
rect 4344 16652 4396 16658
rect 4344 16594 4396 16600
rect 4356 16250 4384 16594
rect 4421 16348 4717 16368
rect 4477 16346 4501 16348
rect 4557 16346 4581 16348
rect 4637 16346 4661 16348
rect 4499 16294 4501 16346
rect 4563 16294 4575 16346
rect 4637 16294 4639 16346
rect 4477 16292 4501 16294
rect 4557 16292 4581 16294
rect 4637 16292 4661 16294
rect 4421 16272 4717 16292
rect 4344 16244 4396 16250
rect 4344 16186 4396 16192
rect 4252 16108 4304 16114
rect 4252 16050 4304 16056
rect 4068 16040 4120 16046
rect 4068 15982 4120 15988
rect 3608 15972 3660 15978
rect 3608 15914 3660 15920
rect 3424 15700 3476 15706
rect 3424 15642 3476 15648
rect 2964 15564 3016 15570
rect 2964 15506 3016 15512
rect 2976 15162 3004 15506
rect 3238 15192 3294 15201
rect 2964 15156 3016 15162
rect 3238 15127 3294 15136
rect 2964 15098 3016 15104
rect 2962 14648 3018 14657
rect 3252 14618 3280 15127
rect 3620 15026 3648 15914
rect 3700 15564 3752 15570
rect 3700 15506 3752 15512
rect 3712 15366 3740 15506
rect 3700 15360 3752 15366
rect 3700 15302 3752 15308
rect 3608 15020 3660 15026
rect 3608 14962 3660 14968
rect 2962 14583 3018 14592
rect 3240 14612 3292 14618
rect 2976 14074 3004 14583
rect 3240 14554 3292 14560
rect 2964 14068 3016 14074
rect 2964 14010 3016 14016
rect 3056 13864 3108 13870
rect 3056 13806 3108 13812
rect 3148 13864 3200 13870
rect 3148 13806 3200 13812
rect 3514 13832 3570 13841
rect 2872 13728 2924 13734
rect 2872 13670 2924 13676
rect 2884 13002 2912 13670
rect 3068 13462 3096 13806
rect 3056 13456 3108 13462
rect 3056 13398 3108 13404
rect 2884 12974 3096 13002
rect 2872 12844 2924 12850
rect 2872 12786 2924 12792
rect 2780 12640 2832 12646
rect 2780 12582 2832 12588
rect 2596 11892 2648 11898
rect 2596 11834 2648 11840
rect 2688 11892 2740 11898
rect 2688 11834 2740 11840
rect 2044 11688 2096 11694
rect 2044 11630 2096 11636
rect 2412 11688 2464 11694
rect 2412 11630 2464 11636
rect 2320 11552 2372 11558
rect 2320 11494 2372 11500
rect 2332 11354 2360 11494
rect 2320 11348 2372 11354
rect 2320 11290 2372 11296
rect 2424 10606 2452 11630
rect 2792 11354 2820 12582
rect 2884 12374 2912 12786
rect 2872 12368 2924 12374
rect 2872 12310 2924 12316
rect 2964 12300 3016 12306
rect 2964 12242 3016 12248
rect 2976 11762 3004 12242
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2976 11218 3004 11698
rect 3068 11354 3096 12974
rect 3160 12442 3188 13806
rect 3514 13767 3570 13776
rect 3528 13530 3556 13767
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 3240 13388 3292 13394
rect 3240 13330 3292 13336
rect 3424 13388 3476 13394
rect 3424 13330 3476 13336
rect 3148 12436 3200 12442
rect 3148 12378 3200 12384
rect 3148 11552 3200 11558
rect 3148 11494 3200 11500
rect 3056 11348 3108 11354
rect 3056 11290 3108 11296
rect 2964 11212 3016 11218
rect 2964 11154 3016 11160
rect 2976 10810 3004 11154
rect 2964 10804 3016 10810
rect 2964 10746 3016 10752
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2964 10532 3016 10538
rect 2964 10474 3016 10480
rect 2688 9988 2740 9994
rect 2688 9930 2740 9936
rect 2700 9518 2728 9930
rect 2976 9654 3004 10474
rect 3160 9994 3188 11494
rect 3148 9988 3200 9994
rect 3148 9930 3200 9936
rect 2964 9648 3016 9654
rect 2964 9590 3016 9596
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 3160 9466 3188 9930
rect 3252 9654 3280 13330
rect 3436 12850 3464 13330
rect 3424 12844 3476 12850
rect 3424 12786 3476 12792
rect 3332 12368 3384 12374
rect 3332 12310 3384 12316
rect 3344 12102 3372 12310
rect 3332 12096 3384 12102
rect 3332 12038 3384 12044
rect 3344 11694 3372 12038
rect 3332 11688 3384 11694
rect 3332 11630 3384 11636
rect 3422 10160 3478 10169
rect 3422 10095 3478 10104
rect 3240 9648 3292 9654
rect 3240 9590 3292 9596
rect 3332 9648 3384 9654
rect 3332 9590 3384 9596
rect 2700 9110 2728 9454
rect 3160 9438 3280 9466
rect 2688 9104 2740 9110
rect 2688 9046 2740 9052
rect 2780 9036 2832 9042
rect 2780 8978 2832 8984
rect 2504 8356 2556 8362
rect 2504 8298 2556 8304
rect 2516 7886 2544 8298
rect 2792 8090 2820 8978
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 2884 8090 2912 8910
rect 3068 8634 3096 8910
rect 3056 8628 3108 8634
rect 3056 8570 3108 8576
rect 3148 8288 3200 8294
rect 3148 8230 3200 8236
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2872 8084 2924 8090
rect 2872 8026 2924 8032
rect 3160 7954 3188 8230
rect 3148 7948 3200 7954
rect 3148 7890 3200 7896
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2516 7546 2544 7822
rect 3056 7812 3108 7818
rect 3056 7754 3108 7760
rect 3068 7546 3096 7754
rect 2504 7540 2556 7546
rect 2504 7482 2556 7488
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 2412 7268 2464 7274
rect 2412 7210 2464 7216
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 2332 5914 2360 6598
rect 2424 6458 2452 7210
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 2872 6860 2924 6866
rect 2872 6802 2924 6808
rect 2884 6662 2912 6802
rect 2872 6656 2924 6662
rect 2872 6598 2924 6604
rect 2412 6452 2464 6458
rect 2412 6394 2464 6400
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 1872 5766 1992 5794
rect 1964 4078 1992 5766
rect 2424 5710 2452 6394
rect 2688 6180 2740 6186
rect 2688 6122 2740 6128
rect 2412 5704 2464 5710
rect 2412 5646 2464 5652
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 1952 4072 2004 4078
rect 1952 4014 2004 4020
rect 1964 3126 1992 4014
rect 2516 4010 2544 4558
rect 2700 4078 2728 6122
rect 2884 6118 2912 6598
rect 2872 6112 2924 6118
rect 2872 6054 2924 6060
rect 2688 4072 2740 4078
rect 2688 4014 2740 4020
rect 2504 4004 2556 4010
rect 2504 3946 2556 3952
rect 2412 3664 2464 3670
rect 2412 3606 2464 3612
rect 1952 3120 2004 3126
rect 1952 3062 2004 3068
rect 1952 2304 2004 2310
rect 1952 2246 2004 2252
rect 1582 2000 1638 2009
rect 1582 1935 1638 1944
rect 1964 800 1992 2246
rect 2424 800 2452 3606
rect 2516 3466 2544 3946
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 2504 3460 2556 3466
rect 2504 3402 2556 3408
rect 2884 3058 2912 3538
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 2884 2854 2912 2994
rect 2872 2848 2924 2854
rect 2872 2790 2924 2796
rect 2884 2689 2912 2790
rect 2870 2680 2926 2689
rect 2870 2615 2926 2624
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 2792 800 2820 2450
rect 202 0 258 800
rect 570 0 626 800
rect 1030 0 1086 800
rect 1490 0 1546 800
rect 1950 0 2006 800
rect 2410 0 2466 800
rect 2778 0 2834 800
rect 2976 241 3004 7142
rect 3056 6928 3108 6934
rect 3056 6870 3108 6876
rect 3068 6322 3096 6870
rect 3056 6316 3108 6322
rect 3056 6258 3108 6264
rect 3056 6112 3108 6118
rect 3056 6054 3108 6060
rect 3068 2553 3096 6054
rect 3160 5574 3188 7890
rect 3252 7410 3280 9438
rect 3344 8362 3372 9590
rect 3332 8356 3384 8362
rect 3332 8298 3384 8304
rect 3332 7948 3384 7954
rect 3332 7890 3384 7896
rect 3344 7546 3372 7890
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 3252 6934 3280 7346
rect 3344 7206 3372 7482
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 3240 6928 3292 6934
rect 3240 6870 3292 6876
rect 3148 5568 3200 5574
rect 3148 5510 3200 5516
rect 3148 4480 3200 4486
rect 3148 4422 3200 4428
rect 3160 3602 3188 4422
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 3252 3505 3280 6870
rect 3436 6866 3464 10095
rect 3514 10024 3570 10033
rect 3514 9959 3570 9968
rect 3528 7449 3556 9959
rect 3608 9920 3660 9926
rect 3608 9862 3660 9868
rect 3620 9518 3648 9862
rect 3712 9654 3740 15302
rect 4080 14770 4108 15982
rect 4356 15434 4384 16186
rect 5552 16114 5580 16934
rect 5736 16658 5764 17070
rect 6276 16992 6328 16998
rect 6276 16934 6328 16940
rect 6288 16794 6316 16934
rect 6276 16788 6328 16794
rect 6276 16730 6328 16736
rect 5908 16720 5960 16726
rect 5908 16662 5960 16668
rect 5724 16652 5776 16658
rect 5724 16594 5776 16600
rect 5540 16108 5592 16114
rect 5540 16050 5592 16056
rect 4988 15904 5040 15910
rect 4988 15846 5040 15852
rect 4896 15632 4948 15638
rect 4896 15574 4948 15580
rect 4344 15428 4396 15434
rect 4344 15370 4396 15376
rect 4160 15360 4212 15366
rect 4160 15302 4212 15308
rect 4172 14958 4200 15302
rect 4421 15260 4717 15280
rect 4477 15258 4501 15260
rect 4557 15258 4581 15260
rect 4637 15258 4661 15260
rect 4499 15206 4501 15258
rect 4563 15206 4575 15258
rect 4637 15206 4639 15258
rect 4477 15204 4501 15206
rect 4557 15204 4581 15206
rect 4637 15204 4661 15206
rect 4421 15184 4717 15204
rect 4908 15094 4936 15574
rect 5000 15552 5028 15846
rect 5080 15564 5132 15570
rect 5000 15524 5080 15552
rect 4896 15088 4948 15094
rect 4896 15030 4948 15036
rect 4160 14952 4212 14958
rect 4160 14894 4212 14900
rect 4436 14952 4488 14958
rect 4436 14894 4488 14900
rect 4080 14742 4200 14770
rect 4172 14414 4200 14742
rect 4448 14414 4476 14894
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 4436 14408 4488 14414
rect 4436 14350 4488 14356
rect 4068 13864 4120 13870
rect 4172 13818 4200 14350
rect 4421 14172 4717 14192
rect 4477 14170 4501 14172
rect 4557 14170 4581 14172
rect 4637 14170 4661 14172
rect 4499 14118 4501 14170
rect 4563 14118 4575 14170
rect 4637 14118 4639 14170
rect 4477 14116 4501 14118
rect 4557 14116 4581 14118
rect 4637 14116 4661 14118
rect 4421 14096 4717 14116
rect 4120 13812 4200 13818
rect 4068 13806 4200 13812
rect 4080 13790 4200 13806
rect 4172 12782 4200 13790
rect 4421 13084 4717 13104
rect 4477 13082 4501 13084
rect 4557 13082 4581 13084
rect 4637 13082 4661 13084
rect 4499 13030 4501 13082
rect 4563 13030 4575 13082
rect 4637 13030 4639 13082
rect 4477 13028 4501 13030
rect 4557 13028 4581 13030
rect 4637 13028 4661 13030
rect 4421 13008 4717 13028
rect 4068 12776 4120 12782
rect 4068 12718 4120 12724
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 3976 12368 4028 12374
rect 3974 12336 3976 12345
rect 4028 12336 4030 12345
rect 3974 12271 4030 12280
rect 3974 11928 4030 11937
rect 3974 11863 4030 11872
rect 3988 11626 4016 11863
rect 3976 11620 4028 11626
rect 3976 11562 4028 11568
rect 3974 11384 4030 11393
rect 3974 11319 4030 11328
rect 3884 11008 3936 11014
rect 3882 10976 3884 10985
rect 3936 10976 3938 10985
rect 3882 10911 3938 10920
rect 3988 10538 4016 11319
rect 3976 10532 4028 10538
rect 3976 10474 4028 10480
rect 3884 10464 3936 10470
rect 3884 10406 3936 10412
rect 3974 10432 4030 10441
rect 3896 10130 3924 10406
rect 3974 10367 4030 10376
rect 3884 10124 3936 10130
rect 3884 10066 3936 10072
rect 3700 9648 3752 9654
rect 3700 9590 3752 9596
rect 3608 9512 3660 9518
rect 3608 9454 3660 9460
rect 3792 9444 3844 9450
rect 3792 9386 3844 9392
rect 3700 9376 3752 9382
rect 3700 9318 3752 9324
rect 3712 9178 3740 9318
rect 3700 9172 3752 9178
rect 3700 9114 3752 9120
rect 3804 8673 3832 9386
rect 3790 8664 3846 8673
rect 3790 8599 3846 8608
rect 3790 8392 3846 8401
rect 3608 8356 3660 8362
rect 3790 8327 3846 8336
rect 3608 8298 3660 8304
rect 3514 7440 3570 7449
rect 3514 7375 3570 7384
rect 3620 6934 3648 8298
rect 3804 7562 3832 8327
rect 3896 8022 3924 10066
rect 3988 9722 4016 10367
rect 3976 9716 4028 9722
rect 3976 9658 4028 9664
rect 4080 9654 4108 12718
rect 4172 12102 4200 12718
rect 4712 12708 4764 12714
rect 4712 12650 4764 12656
rect 4724 12238 4752 12650
rect 4804 12300 4856 12306
rect 4804 12242 4856 12248
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4252 12164 4304 12170
rect 4252 12106 4304 12112
rect 4160 12096 4212 12102
rect 4160 12038 4212 12044
rect 4172 11150 4200 12038
rect 4264 11286 4292 12106
rect 4421 11996 4717 12016
rect 4477 11994 4501 11996
rect 4557 11994 4581 11996
rect 4637 11994 4661 11996
rect 4499 11942 4501 11994
rect 4563 11942 4575 11994
rect 4637 11942 4639 11994
rect 4477 11940 4501 11942
rect 4557 11940 4581 11942
rect 4637 11940 4661 11942
rect 4421 11920 4717 11940
rect 4816 11762 4844 12242
rect 5000 12186 5028 15524
rect 5080 15506 5132 15512
rect 5816 15496 5868 15502
rect 5816 15438 5868 15444
rect 5828 14890 5856 15438
rect 5920 15094 5948 16662
rect 6288 15910 6316 16730
rect 6472 16726 6500 17138
rect 6920 16992 6972 16998
rect 6920 16934 6972 16940
rect 7472 16992 7524 16998
rect 7472 16934 7524 16940
rect 6460 16720 6512 16726
rect 6460 16662 6512 16668
rect 6932 16250 6960 16934
rect 7012 16652 7064 16658
rect 7012 16594 7064 16600
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 7024 15978 7052 16594
rect 7288 16448 7340 16454
rect 7288 16390 7340 16396
rect 7300 16114 7328 16390
rect 7288 16108 7340 16114
rect 7288 16050 7340 16056
rect 7012 15972 7064 15978
rect 7012 15914 7064 15920
rect 6276 15904 6328 15910
rect 6276 15846 6328 15852
rect 6552 15904 6604 15910
rect 6552 15846 6604 15852
rect 7024 15858 7052 15914
rect 7196 15904 7248 15910
rect 5908 15088 5960 15094
rect 5908 15030 5960 15036
rect 5816 14884 5868 14890
rect 5816 14826 5868 14832
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 5264 14476 5316 14482
rect 5264 14418 5316 14424
rect 5276 14074 5304 14418
rect 5644 14074 5672 14758
rect 5828 14618 5856 14826
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 5816 14476 5868 14482
rect 5816 14418 5868 14424
rect 5264 14068 5316 14074
rect 5264 14010 5316 14016
rect 5632 14068 5684 14074
rect 5632 14010 5684 14016
rect 5080 13796 5132 13802
rect 5080 13738 5132 13744
rect 5540 13796 5592 13802
rect 5540 13738 5592 13744
rect 5092 13462 5120 13738
rect 5080 13456 5132 13462
rect 5080 13398 5132 13404
rect 5092 12986 5120 13398
rect 5264 13388 5316 13394
rect 5264 13330 5316 13336
rect 5080 12980 5132 12986
rect 5080 12922 5132 12928
rect 5276 12918 5304 13330
rect 5552 13274 5580 13738
rect 5460 13258 5580 13274
rect 5448 13252 5580 13258
rect 5500 13246 5580 13252
rect 5448 13194 5500 13200
rect 5264 12912 5316 12918
rect 5264 12854 5316 12860
rect 5448 12912 5500 12918
rect 5448 12854 5500 12860
rect 5080 12640 5132 12646
rect 5080 12582 5132 12588
rect 5092 12306 5120 12582
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 5000 12158 5120 12186
rect 4804 11756 4856 11762
rect 4804 11698 4856 11704
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 4252 11280 4304 11286
rect 4252 11222 4304 11228
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 4172 10606 4200 11086
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 4160 10600 4212 10606
rect 4160 10542 4212 10548
rect 4160 10464 4212 10470
rect 4160 10406 4212 10412
rect 4172 10266 4200 10406
rect 4160 10260 4212 10266
rect 4160 10202 4212 10208
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 4172 9926 4200 9998
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 4068 9648 4120 9654
rect 4068 9590 4120 9596
rect 4066 9480 4122 9489
rect 4066 9415 4122 9424
rect 4080 9110 4108 9415
rect 4068 9104 4120 9110
rect 3974 9072 4030 9081
rect 4068 9046 4120 9052
rect 3974 9007 4030 9016
rect 3988 8362 4016 9007
rect 4172 8906 4200 9862
rect 4160 8900 4212 8906
rect 4160 8842 4212 8848
rect 3976 8356 4028 8362
rect 3976 8298 4028 8304
rect 4066 8120 4122 8129
rect 4066 8055 4122 8064
rect 3884 8016 3936 8022
rect 3884 7958 3936 7964
rect 3976 7812 4028 7818
rect 3976 7754 4028 7760
rect 3988 7721 4016 7754
rect 3974 7712 4030 7721
rect 3974 7647 4030 7656
rect 3804 7534 4016 7562
rect 3700 7268 3752 7274
rect 3700 7210 3752 7216
rect 3608 6928 3660 6934
rect 3608 6870 3660 6876
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3608 6656 3660 6662
rect 3608 6598 3660 6604
rect 3620 6254 3648 6598
rect 3608 6248 3660 6254
rect 3514 6216 3570 6225
rect 3608 6190 3660 6196
rect 3514 6151 3570 6160
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3436 5914 3464 6054
rect 3528 5914 3556 6151
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3620 5710 3648 6190
rect 3608 5704 3660 5710
rect 3608 5646 3660 5652
rect 3516 5160 3568 5166
rect 3516 5102 3568 5108
rect 3332 4616 3384 4622
rect 3332 4558 3384 4564
rect 3424 4616 3476 4622
rect 3424 4558 3476 4564
rect 3344 3738 3372 4558
rect 3436 4282 3464 4558
rect 3424 4276 3476 4282
rect 3424 4218 3476 4224
rect 3332 3732 3384 3738
rect 3332 3674 3384 3680
rect 3424 3528 3476 3534
rect 3238 3496 3294 3505
rect 3238 3431 3294 3440
rect 3422 3496 3424 3505
rect 3476 3496 3478 3505
rect 3422 3431 3478 3440
rect 3240 3392 3292 3398
rect 3240 3334 3292 3340
rect 3054 2544 3110 2553
rect 3054 2479 3110 2488
rect 3252 800 3280 3334
rect 3422 2680 3478 2689
rect 3422 2615 3478 2624
rect 3436 2446 3464 2615
rect 3424 2440 3476 2446
rect 3424 2382 3476 2388
rect 2962 232 3018 241
rect 2962 167 3018 176
rect 3238 0 3294 800
rect 3528 649 3556 5102
rect 3608 3528 3660 3534
rect 3608 3470 3660 3476
rect 3620 3194 3648 3470
rect 3608 3188 3660 3194
rect 3608 3130 3660 3136
rect 3712 800 3740 7210
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 3804 6186 3832 6734
rect 3792 6180 3844 6186
rect 3792 6122 3844 6128
rect 3884 6180 3936 6186
rect 3884 6122 3936 6128
rect 3804 5778 3832 6122
rect 3896 5817 3924 6122
rect 3988 6118 4016 7534
rect 4080 7478 4108 8055
rect 4068 7472 4120 7478
rect 4068 7414 4120 7420
rect 4066 6760 4122 6769
rect 4066 6695 4122 6704
rect 4080 6458 4108 6695
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3882 5808 3938 5817
rect 3792 5772 3844 5778
rect 3882 5743 3938 5752
rect 3792 5714 3844 5720
rect 3884 5704 3936 5710
rect 3884 5646 3936 5652
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 3804 1057 3832 5510
rect 3896 5166 3924 5646
rect 3988 5370 4016 6054
rect 3976 5364 4028 5370
rect 3976 5306 4028 5312
rect 4066 5264 4122 5273
rect 4066 5199 4122 5208
rect 3884 5160 3936 5166
rect 3884 5102 3936 5108
rect 3884 5024 3936 5030
rect 3884 4966 3936 4972
rect 3896 1601 3924 4966
rect 4080 4826 4108 5199
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 3976 4752 4028 4758
rect 3976 4694 4028 4700
rect 3988 2514 4016 4694
rect 4068 4548 4120 4554
rect 4068 4490 4120 4496
rect 4080 4457 4108 4490
rect 4066 4448 4122 4457
rect 4066 4383 4122 4392
rect 4172 2961 4200 8842
rect 4264 8838 4292 11018
rect 4356 10606 4384 11494
rect 4421 10908 4717 10928
rect 4477 10906 4501 10908
rect 4557 10906 4581 10908
rect 4637 10906 4661 10908
rect 4499 10854 4501 10906
rect 4563 10854 4575 10906
rect 4637 10854 4639 10906
rect 4477 10852 4501 10854
rect 4557 10852 4581 10854
rect 4637 10852 4661 10854
rect 4421 10832 4717 10852
rect 4344 10600 4396 10606
rect 4344 10542 4396 10548
rect 4356 10062 4384 10542
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4421 9820 4717 9840
rect 4477 9818 4501 9820
rect 4557 9818 4581 9820
rect 4637 9818 4661 9820
rect 4499 9766 4501 9818
rect 4563 9766 4575 9818
rect 4637 9766 4639 9818
rect 4477 9764 4501 9766
rect 4557 9764 4581 9766
rect 4637 9764 4661 9766
rect 4421 9744 4717 9764
rect 4804 9444 4856 9450
rect 4804 9386 4856 9392
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4421 8732 4717 8752
rect 4477 8730 4501 8732
rect 4557 8730 4581 8732
rect 4637 8730 4661 8732
rect 4499 8678 4501 8730
rect 4563 8678 4575 8730
rect 4637 8678 4639 8730
rect 4477 8676 4501 8678
rect 4557 8676 4581 8678
rect 4637 8676 4661 8678
rect 4421 8656 4717 8676
rect 4816 8090 4844 9386
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 4908 9178 4936 9318
rect 5092 9178 5120 12158
rect 5460 11336 5488 12854
rect 5632 12368 5684 12374
rect 5632 12310 5684 12316
rect 5368 11308 5488 11336
rect 5368 10282 5396 11308
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5460 10810 5488 11154
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5460 10674 5488 10746
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5368 10254 5488 10282
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 5368 9382 5396 10066
rect 5460 9738 5488 10254
rect 5644 9994 5672 12310
rect 5828 10810 5856 14418
rect 6000 13728 6052 13734
rect 6000 13670 6052 13676
rect 6012 13530 6040 13670
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 6092 13184 6144 13190
rect 6092 13126 6144 13132
rect 5908 12300 5960 12306
rect 6104 12288 6132 13126
rect 5908 12242 5960 12248
rect 6012 12260 6132 12288
rect 5920 11354 5948 12242
rect 5908 11348 5960 11354
rect 5908 11290 5960 11296
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 5816 10600 5868 10606
rect 5816 10542 5868 10548
rect 5828 10198 5856 10542
rect 5816 10192 5868 10198
rect 5816 10134 5868 10140
rect 5908 10192 5960 10198
rect 5908 10134 5960 10140
rect 5724 10124 5776 10130
rect 5724 10066 5776 10072
rect 5632 9988 5684 9994
rect 5632 9930 5684 9936
rect 5460 9710 5580 9738
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5356 9376 5408 9382
rect 5356 9318 5408 9324
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 4988 8832 5040 8838
rect 4988 8774 5040 8780
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 4804 8084 4856 8090
rect 4804 8026 4856 8032
rect 4421 7644 4717 7664
rect 4477 7642 4501 7644
rect 4557 7642 4581 7644
rect 4637 7642 4661 7644
rect 4499 7590 4501 7642
rect 4563 7590 4575 7642
rect 4637 7590 4639 7642
rect 4477 7588 4501 7590
rect 4557 7588 4581 7590
rect 4637 7588 4661 7590
rect 4421 7568 4717 7588
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 4908 7342 4936 7482
rect 4896 7336 4948 7342
rect 4896 7278 4948 7284
rect 4618 7168 4674 7177
rect 4618 7103 4674 7112
rect 4632 6934 4660 7103
rect 4620 6928 4672 6934
rect 4620 6870 4672 6876
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 4356 6322 4384 6802
rect 4421 6556 4717 6576
rect 4477 6554 4501 6556
rect 4557 6554 4581 6556
rect 4637 6554 4661 6556
rect 4499 6502 4501 6554
rect 4563 6502 4575 6554
rect 4637 6502 4639 6554
rect 4477 6500 4501 6502
rect 4557 6500 4581 6502
rect 4637 6500 4661 6502
rect 4421 6480 4717 6500
rect 4908 6338 4936 7278
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 4724 6310 4936 6338
rect 4724 6254 4752 6310
rect 4712 6248 4764 6254
rect 4712 6190 4764 6196
rect 4894 6216 4950 6225
rect 4894 6151 4950 6160
rect 4252 6112 4304 6118
rect 4252 6054 4304 6060
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 4264 5574 4292 6054
rect 4724 5710 4752 6054
rect 4908 5778 4936 6151
rect 4896 5772 4948 5778
rect 4896 5714 4948 5720
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 4158 2952 4214 2961
rect 4158 2887 4214 2896
rect 3976 2508 4028 2514
rect 3976 2450 4028 2456
rect 3882 1592 3938 1601
rect 3882 1527 3938 1536
rect 3790 1048 3846 1057
rect 3790 983 3846 992
rect 4264 898 4292 5510
rect 4421 5468 4717 5488
rect 4477 5466 4501 5468
rect 4557 5466 4581 5468
rect 4637 5466 4661 5468
rect 4499 5414 4501 5466
rect 4563 5414 4575 5466
rect 4637 5414 4639 5466
rect 4477 5412 4501 5414
rect 4557 5412 4581 5414
rect 4637 5412 4661 5414
rect 4421 5392 4717 5412
rect 4421 4380 4717 4400
rect 4477 4378 4501 4380
rect 4557 4378 4581 4380
rect 4637 4378 4661 4380
rect 4499 4326 4501 4378
rect 4563 4326 4575 4378
rect 4637 4326 4639 4378
rect 4477 4324 4501 4326
rect 4557 4324 4581 4326
rect 4637 4324 4661 4326
rect 4421 4304 4717 4324
rect 4344 3596 4396 3602
rect 4344 3538 4396 3544
rect 4356 2802 4384 3538
rect 4421 3292 4717 3312
rect 4477 3290 4501 3292
rect 4557 3290 4581 3292
rect 4637 3290 4661 3292
rect 4499 3238 4501 3290
rect 4563 3238 4575 3290
rect 4637 3238 4639 3290
rect 4477 3236 4501 3238
rect 4557 3236 4581 3238
rect 4637 3236 4661 3238
rect 4421 3216 4717 3236
rect 4347 2774 4384 2802
rect 4347 2666 4375 2774
rect 4347 2650 4384 2666
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 4421 2204 4717 2224
rect 4477 2202 4501 2204
rect 4557 2202 4581 2204
rect 4637 2202 4661 2204
rect 4499 2150 4501 2202
rect 4563 2150 4575 2202
rect 4637 2150 4639 2202
rect 4477 2148 4501 2150
rect 4557 2148 4581 2150
rect 4637 2148 4661 2150
rect 4421 2128 4717 2148
rect 4816 1034 4844 5646
rect 4908 5030 4936 5714
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4896 4480 4948 4486
rect 4896 4422 4948 4428
rect 4908 4282 4936 4422
rect 4896 4276 4948 4282
rect 4896 4218 4948 4224
rect 4908 3398 4936 4218
rect 4896 3392 4948 3398
rect 4896 3334 4948 3340
rect 4172 870 4292 898
rect 4632 1006 4844 1034
rect 4172 800 4200 870
rect 4632 800 4660 1006
rect 5000 800 5028 8774
rect 5092 8430 5120 8774
rect 5276 8634 5304 8910
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5080 8424 5132 8430
rect 5080 8366 5132 8372
rect 5092 7886 5120 8366
rect 5080 7880 5132 7886
rect 5080 7822 5132 7828
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 5092 5710 5120 7686
rect 5276 7546 5304 8570
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5080 5704 5132 5710
rect 5080 5646 5132 5652
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 5276 4282 5304 4558
rect 5264 4276 5316 4282
rect 5264 4218 5316 4224
rect 5172 4004 5224 4010
rect 5172 3946 5224 3952
rect 5184 3602 5212 3946
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 5080 3392 5132 3398
rect 5080 3334 5132 3340
rect 5092 2990 5120 3334
rect 5184 3194 5212 3538
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5368 3074 5396 9318
rect 5460 8634 5488 9522
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5460 6186 5488 8570
rect 5552 8294 5580 9710
rect 5736 9382 5764 10066
rect 5920 10010 5948 10134
rect 6012 10044 6040 12260
rect 6092 11348 6144 11354
rect 6092 11290 6144 11296
rect 6104 10146 6132 11290
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6196 10266 6224 10406
rect 6184 10260 6236 10266
rect 6184 10202 6236 10208
rect 6288 10169 6316 15846
rect 6564 15638 6592 15846
rect 7024 15830 7144 15858
rect 7196 15846 7248 15852
rect 6552 15632 6604 15638
rect 6552 15574 6604 15580
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6380 12238 6408 12582
rect 6368 12232 6420 12238
rect 6368 12174 6420 12180
rect 6274 10160 6330 10169
rect 6104 10118 6224 10146
rect 6196 10062 6224 10118
rect 6274 10095 6330 10104
rect 6184 10056 6236 10062
rect 6012 10016 6132 10044
rect 5828 9982 5948 10010
rect 5724 9376 5776 9382
rect 5724 9318 5776 9324
rect 5632 9036 5684 9042
rect 5632 8978 5684 8984
rect 5644 8498 5672 8978
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5736 8378 5764 9318
rect 5644 8350 5764 8378
rect 5540 8288 5592 8294
rect 5540 8230 5592 8236
rect 5552 7206 5580 8230
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5552 7002 5580 7142
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 5644 5642 5672 8350
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 5736 7546 5764 7890
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5632 5636 5684 5642
rect 5632 5578 5684 5584
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5552 4146 5580 4218
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 5276 3046 5396 3074
rect 5080 2984 5132 2990
rect 5080 2926 5132 2932
rect 5276 2938 5304 3046
rect 5552 2990 5580 4082
rect 5644 4078 5672 4762
rect 5632 4072 5684 4078
rect 5632 4014 5684 4020
rect 5632 3936 5684 3942
rect 5736 3890 5764 4762
rect 5684 3884 5764 3890
rect 5632 3878 5764 3884
rect 5644 3862 5764 3878
rect 5828 3482 5856 9982
rect 6104 9160 6132 10016
rect 6184 9998 6236 10004
rect 6104 9132 6408 9160
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 6104 8634 6132 8978
rect 6092 8628 6144 8634
rect 6092 8570 6144 8576
rect 6104 7886 6132 8570
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 5920 7274 5948 7822
rect 6104 7410 6132 7822
rect 6092 7404 6144 7410
rect 6092 7346 6144 7352
rect 5908 7268 5960 7274
rect 5908 7210 5960 7216
rect 6092 7200 6144 7206
rect 6092 7142 6144 7148
rect 6104 6866 6132 7142
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 6276 4684 6328 4690
rect 6276 4626 6328 4632
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 5920 3602 5948 4558
rect 5908 3596 5960 3602
rect 5908 3538 5960 3544
rect 5828 3454 5948 3482
rect 5540 2984 5592 2990
rect 5276 2910 5488 2938
rect 5540 2926 5592 2932
rect 5460 800 5488 2910
rect 5920 800 5948 3454
rect 6104 2922 6132 4558
rect 6184 4480 6236 4486
rect 6184 4422 6236 4428
rect 6092 2916 6144 2922
rect 6092 2858 6144 2864
rect 6196 2650 6224 4422
rect 6288 4146 6316 4626
rect 6276 4140 6328 4146
rect 6276 4082 6328 4088
rect 6380 3720 6408 9132
rect 6460 4276 6512 4282
rect 6460 4218 6512 4224
rect 6288 3692 6408 3720
rect 6288 2666 6316 3692
rect 6368 3596 6420 3602
rect 6368 3538 6420 3544
rect 6380 2854 6408 3538
rect 6472 3534 6500 4218
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 6368 2848 6420 2854
rect 6368 2790 6420 2796
rect 6184 2644 6236 2650
rect 6288 2638 6408 2666
rect 6184 2586 6236 2592
rect 6380 800 6408 2638
rect 6564 1170 6592 15574
rect 6920 15360 6972 15366
rect 6920 15302 6972 15308
rect 6932 14482 6960 15302
rect 6920 14476 6972 14482
rect 6920 14418 6972 14424
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6840 12628 6868 13806
rect 6932 13394 6960 14418
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 6920 13388 6972 13394
rect 6920 13330 6972 13336
rect 7024 12986 7052 14010
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 7024 12782 7052 12922
rect 7012 12776 7064 12782
rect 7012 12718 7064 12724
rect 6840 12600 7052 12628
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 6840 11150 6868 12174
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 6918 10160 6974 10169
rect 6918 10095 6920 10104
rect 6972 10095 6974 10104
rect 6920 10066 6972 10072
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6656 8906 6684 9454
rect 6736 9172 6788 9178
rect 6736 9114 6788 9120
rect 6644 8900 6696 8906
rect 6644 8842 6696 8848
rect 6748 5522 6776 9114
rect 6840 8498 6868 9454
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 7024 8401 7052 12600
rect 7010 8392 7066 8401
rect 7010 8327 7066 8336
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6656 5494 6776 5522
rect 6656 4128 6684 5494
rect 6736 5364 6788 5370
rect 6736 5306 6788 5312
rect 6748 4826 6776 5306
rect 6840 5166 6868 6054
rect 7024 5778 7052 7142
rect 7012 5772 7064 5778
rect 6932 5732 7012 5760
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 6932 4706 6960 5732
rect 7012 5714 7064 5720
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 6840 4678 6960 4706
rect 6840 4146 6868 4678
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 6828 4140 6880 4146
rect 6656 4100 6776 4128
rect 6644 4004 6696 4010
rect 6644 3946 6696 3952
rect 6656 3738 6684 3946
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6656 2446 6684 3674
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 6748 2310 6776 4100
rect 6828 4082 6880 4088
rect 6828 2848 6880 2854
rect 6828 2790 6880 2796
rect 6840 2446 6868 2790
rect 6828 2440 6880 2446
rect 6828 2382 6880 2388
rect 6932 2378 6960 4558
rect 7024 3670 7052 4966
rect 7116 4162 7144 15830
rect 7208 15026 7236 15846
rect 7300 15638 7328 16050
rect 7484 15910 7512 16934
rect 7472 15904 7524 15910
rect 7392 15852 7472 15858
rect 7392 15846 7524 15852
rect 7392 15830 7512 15846
rect 7288 15632 7340 15638
rect 7288 15574 7340 15580
rect 7196 15020 7248 15026
rect 7196 14962 7248 14968
rect 7392 12594 7420 15830
rect 7472 15360 7524 15366
rect 7472 15302 7524 15308
rect 7484 15026 7512 15302
rect 7472 15020 7524 15026
rect 7472 14962 7524 14968
rect 7484 14550 7512 14962
rect 7472 14544 7524 14550
rect 7472 14486 7524 14492
rect 7300 12566 7420 12594
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 7208 10266 7236 11154
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7300 9994 7328 12566
rect 7576 11898 7604 17682
rect 8220 17202 8248 17682
rect 8484 17672 8536 17678
rect 8484 17614 8536 17620
rect 8392 17604 8444 17610
rect 8392 17546 8444 17552
rect 8208 17196 8260 17202
rect 8208 17138 8260 17144
rect 7886 16892 8182 16912
rect 7942 16890 7966 16892
rect 8022 16890 8046 16892
rect 8102 16890 8126 16892
rect 7964 16838 7966 16890
rect 8028 16838 8040 16890
rect 8102 16838 8104 16890
rect 7942 16836 7966 16838
rect 8022 16836 8046 16838
rect 8102 16836 8126 16838
rect 7886 16816 8182 16836
rect 7656 15904 7708 15910
rect 7656 15846 7708 15852
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7380 11552 7432 11558
rect 7380 11494 7432 11500
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7392 11354 7420 11494
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7484 10810 7512 11494
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7564 10804 7616 10810
rect 7564 10746 7616 10752
rect 7288 9988 7340 9994
rect 7288 9930 7340 9936
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 7208 8974 7236 9386
rect 7576 9042 7604 10746
rect 7564 9036 7616 9042
rect 7564 8978 7616 8984
rect 7196 8968 7248 8974
rect 7196 8910 7248 8916
rect 7196 8832 7248 8838
rect 7196 8774 7248 8780
rect 7208 7342 7236 8774
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7196 7336 7248 7342
rect 7196 7278 7248 7284
rect 7300 5030 7328 7686
rect 7668 7562 7696 15846
rect 7886 15804 8182 15824
rect 7942 15802 7966 15804
rect 8022 15802 8046 15804
rect 8102 15802 8126 15804
rect 7964 15750 7966 15802
rect 8028 15750 8040 15802
rect 8102 15750 8104 15802
rect 7942 15748 7966 15750
rect 8022 15748 8046 15750
rect 8102 15748 8126 15750
rect 7886 15728 8182 15748
rect 8300 15700 8352 15706
rect 8300 15642 8352 15648
rect 8312 15162 8340 15642
rect 8404 15586 8432 17546
rect 8496 15706 8524 17614
rect 8760 17128 8812 17134
rect 8760 17070 8812 17076
rect 8772 16726 8800 17070
rect 8760 16720 8812 16726
rect 8760 16662 8812 16668
rect 8772 16114 8800 16662
rect 8760 16108 8812 16114
rect 8760 16050 8812 16056
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 8404 15558 8524 15586
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 7886 14716 8182 14736
rect 7942 14714 7966 14716
rect 8022 14714 8046 14716
rect 8102 14714 8126 14716
rect 7964 14662 7966 14714
rect 8028 14662 8040 14714
rect 8102 14662 8104 14714
rect 7942 14660 7966 14662
rect 8022 14660 8046 14662
rect 8102 14660 8126 14662
rect 7886 14640 8182 14660
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 8220 13938 8248 14214
rect 8208 13932 8260 13938
rect 8208 13874 8260 13880
rect 7886 13628 8182 13648
rect 7942 13626 7966 13628
rect 8022 13626 8046 13628
rect 8102 13626 8126 13628
rect 7964 13574 7966 13626
rect 8028 13574 8040 13626
rect 8102 13574 8104 13626
rect 7942 13572 7966 13574
rect 8022 13572 8046 13574
rect 8102 13572 8126 13574
rect 7886 13552 8182 13572
rect 8220 13462 8248 13874
rect 8208 13456 8260 13462
rect 8208 13398 8260 13404
rect 8116 13388 8168 13394
rect 8116 13330 8168 13336
rect 8024 13320 8076 13326
rect 8024 13262 8076 13268
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 7760 10810 7788 12718
rect 8036 12714 8064 13262
rect 8128 12730 8156 13330
rect 8220 12850 8248 13398
rect 8392 13184 8444 13190
rect 8392 13126 8444 13132
rect 8298 12880 8354 12889
rect 8208 12844 8260 12850
rect 8404 12850 8432 13126
rect 8496 12986 8524 15558
rect 8772 14482 8800 16050
rect 8956 15162 8984 19246
rect 10600 19168 10652 19174
rect 10600 19110 10652 19116
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9692 17882 9720 18770
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9312 17672 9364 17678
rect 9312 17614 9364 17620
rect 9680 17672 9732 17678
rect 9680 17614 9732 17620
rect 10324 17672 10376 17678
rect 10324 17614 10376 17620
rect 9324 17066 9352 17614
rect 9312 17060 9364 17066
rect 9312 17002 9364 17008
rect 9324 16794 9352 17002
rect 9692 16794 9720 17614
rect 10232 17060 10284 17066
rect 10232 17002 10284 17008
rect 9312 16788 9364 16794
rect 9312 16730 9364 16736
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 10048 16720 10100 16726
rect 10048 16662 10100 16668
rect 9036 16652 9088 16658
rect 9036 16594 9088 16600
rect 9048 16250 9076 16594
rect 9036 16244 9088 16250
rect 9036 16186 9088 16192
rect 9048 15502 9076 16186
rect 9588 15972 9640 15978
rect 9588 15914 9640 15920
rect 9128 15564 9180 15570
rect 9128 15506 9180 15512
rect 9036 15496 9088 15502
rect 9036 15438 9088 15444
rect 8944 15156 8996 15162
rect 8944 15098 8996 15104
rect 8760 14476 8812 14482
rect 8760 14418 8812 14424
rect 8772 13870 8800 14418
rect 8944 14000 8996 14006
rect 8944 13942 8996 13948
rect 8576 13864 8628 13870
rect 8576 13806 8628 13812
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8484 12980 8536 12986
rect 8484 12922 8536 12928
rect 8298 12815 8354 12824
rect 8392 12844 8444 12850
rect 8208 12786 8260 12792
rect 8024 12708 8076 12714
rect 8128 12702 8248 12730
rect 8024 12650 8076 12656
rect 7886 12540 8182 12560
rect 7942 12538 7966 12540
rect 8022 12538 8046 12540
rect 8102 12538 8126 12540
rect 7964 12486 7966 12538
rect 8028 12486 8040 12538
rect 8102 12486 8104 12538
rect 7942 12484 7966 12486
rect 8022 12484 8046 12486
rect 8102 12484 8126 12486
rect 7886 12464 8182 12484
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 8128 11540 8156 12038
rect 8220 11762 8248 12702
rect 8312 12170 8340 12815
rect 8392 12786 8444 12792
rect 8404 12374 8432 12786
rect 8392 12368 8444 12374
rect 8392 12310 8444 12316
rect 8300 12164 8352 12170
rect 8300 12106 8352 12112
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 8484 11688 8536 11694
rect 8484 11630 8536 11636
rect 8128 11512 8248 11540
rect 7886 11452 8182 11472
rect 7942 11450 7966 11452
rect 8022 11450 8046 11452
rect 8102 11450 8126 11452
rect 7964 11398 7966 11450
rect 8028 11398 8040 11450
rect 8102 11398 8104 11450
rect 7942 11396 7966 11398
rect 8022 11396 8046 11398
rect 8102 11396 8126 11398
rect 7886 11376 8182 11396
rect 8220 11218 8248 11512
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 8220 10674 8248 11154
rect 8496 11082 8524 11630
rect 8484 11076 8536 11082
rect 8484 11018 8536 11024
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 7886 10364 8182 10384
rect 7942 10362 7966 10364
rect 8022 10362 8046 10364
rect 8102 10362 8126 10364
rect 7964 10310 7966 10362
rect 8028 10310 8040 10362
rect 8102 10310 8104 10362
rect 7942 10308 7966 10310
rect 8022 10308 8046 10310
rect 8102 10308 8126 10310
rect 7886 10288 8182 10308
rect 7748 10124 7800 10130
rect 7748 10066 7800 10072
rect 7760 9178 7788 10066
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8220 9382 8248 9998
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 7886 9276 8182 9296
rect 7942 9274 7966 9276
rect 8022 9274 8046 9276
rect 8102 9274 8126 9276
rect 7964 9222 7966 9274
rect 8028 9222 8040 9274
rect 8102 9222 8104 9274
rect 7942 9220 7966 9222
rect 8022 9220 8046 9222
rect 8102 9220 8126 9222
rect 7886 9200 8182 9220
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 8024 8492 8076 8498
rect 8024 8434 8076 8440
rect 8036 8401 8064 8434
rect 8220 8430 8248 9318
rect 8404 9110 8432 9862
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8496 9178 8524 9318
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8392 9104 8444 9110
rect 8392 9046 8444 9052
rect 8208 8424 8260 8430
rect 8022 8392 8078 8401
rect 8208 8366 8260 8372
rect 8022 8327 8078 8336
rect 7886 8188 8182 8208
rect 7942 8186 7966 8188
rect 8022 8186 8046 8188
rect 8102 8186 8126 8188
rect 7964 8134 7966 8186
rect 8028 8134 8040 8186
rect 8102 8134 8104 8186
rect 7942 8132 7966 8134
rect 8022 8132 8046 8134
rect 8102 8132 8126 8134
rect 7886 8112 8182 8132
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 7668 7534 7788 7562
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 7484 5778 7512 6258
rect 7564 5840 7616 5846
rect 7564 5782 7616 5788
rect 7472 5772 7524 5778
rect 7472 5714 7524 5720
rect 7472 5568 7524 5574
rect 7472 5510 7524 5516
rect 7484 5234 7512 5510
rect 7576 5234 7604 5782
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7564 5228 7616 5234
rect 7564 5170 7616 5176
rect 7288 5024 7340 5030
rect 7288 4966 7340 4972
rect 7300 4690 7328 4966
rect 7380 4752 7432 4758
rect 7472 4752 7524 4758
rect 7432 4712 7472 4740
rect 7380 4694 7432 4700
rect 7472 4694 7524 4700
rect 7288 4684 7340 4690
rect 7288 4626 7340 4632
rect 7576 4604 7604 5170
rect 7656 4616 7708 4622
rect 7576 4576 7656 4604
rect 7576 4282 7604 4576
rect 7656 4558 7708 4564
rect 7564 4276 7616 4282
rect 7564 4218 7616 4224
rect 7116 4134 7696 4162
rect 7380 4072 7432 4078
rect 7380 4014 7432 4020
rect 7012 3664 7064 3670
rect 7012 3606 7064 3612
rect 7392 3602 7420 4014
rect 7564 4004 7616 4010
rect 7564 3946 7616 3952
rect 7576 3602 7604 3946
rect 7380 3596 7432 3602
rect 7380 3538 7432 3544
rect 7564 3596 7616 3602
rect 7564 3538 7616 3544
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 7012 2916 7064 2922
rect 7012 2858 7064 2864
rect 6920 2372 6972 2378
rect 6920 2314 6972 2320
rect 6736 2304 6788 2310
rect 6736 2246 6788 2252
rect 7024 2038 7052 2858
rect 7196 2848 7248 2854
rect 7196 2790 7248 2796
rect 7208 2582 7236 2790
rect 7300 2650 7328 3334
rect 7288 2644 7340 2650
rect 7288 2586 7340 2592
rect 7196 2576 7248 2582
rect 7196 2518 7248 2524
rect 7196 2304 7248 2310
rect 7196 2246 7248 2252
rect 7012 2032 7064 2038
rect 7012 1974 7064 1980
rect 6564 1142 6868 1170
rect 6840 800 6868 1142
rect 7208 800 7236 2246
rect 7392 2106 7420 3538
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7484 3058 7512 3470
rect 7576 3058 7604 3538
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 7380 2100 7432 2106
rect 7380 2042 7432 2048
rect 7668 800 7696 4134
rect 7760 2632 7788 7534
rect 7944 7342 7972 7822
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 7886 7100 8182 7120
rect 7942 7098 7966 7100
rect 8022 7098 8046 7100
rect 8102 7098 8126 7100
rect 7964 7046 7966 7098
rect 8028 7046 8040 7098
rect 8102 7046 8104 7098
rect 7942 7044 7966 7046
rect 8022 7044 8046 7046
rect 8102 7044 8126 7046
rect 7886 7024 8182 7044
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8208 6180 8260 6186
rect 8208 6122 8260 6128
rect 7886 6012 8182 6032
rect 7942 6010 7966 6012
rect 8022 6010 8046 6012
rect 8102 6010 8126 6012
rect 7964 5958 7966 6010
rect 8028 5958 8040 6010
rect 8102 5958 8104 6010
rect 7942 5956 7966 5958
rect 8022 5956 8046 5958
rect 8102 5956 8126 5958
rect 7886 5936 8182 5956
rect 8220 5896 8248 6122
rect 8036 5868 8248 5896
rect 8036 5574 8064 5868
rect 8024 5568 8076 5574
rect 8024 5510 8076 5516
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 7886 4924 8182 4944
rect 7942 4922 7966 4924
rect 8022 4922 8046 4924
rect 8102 4922 8126 4924
rect 7964 4870 7966 4922
rect 8028 4870 8040 4922
rect 8102 4870 8104 4922
rect 7942 4868 7966 4870
rect 8022 4868 8046 4870
rect 8102 4868 8126 4870
rect 7886 4848 8182 4868
rect 8220 4826 8248 4966
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8116 4684 8168 4690
rect 8116 4626 8168 4632
rect 8128 4146 8156 4626
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 8220 4078 8248 4558
rect 8392 4480 8444 4486
rect 8496 4468 8524 6598
rect 8444 4440 8524 4468
rect 8392 4422 8444 4428
rect 8404 4078 8432 4422
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 7886 3836 8182 3856
rect 7942 3834 7966 3836
rect 8022 3834 8046 3836
rect 8102 3834 8126 3836
rect 7964 3782 7966 3834
rect 8028 3782 8040 3834
rect 8102 3782 8104 3834
rect 7942 3780 7966 3782
rect 8022 3780 8046 3782
rect 8102 3780 8126 3782
rect 7886 3760 8182 3780
rect 8496 3738 8524 3878
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8392 2916 8444 2922
rect 8392 2858 8444 2864
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 7886 2748 8182 2768
rect 7942 2746 7966 2748
rect 8022 2746 8046 2748
rect 8102 2746 8126 2748
rect 7964 2694 7966 2746
rect 8028 2694 8040 2746
rect 8102 2694 8104 2746
rect 7942 2692 7966 2694
rect 8022 2692 8046 2694
rect 8102 2692 8126 2694
rect 7886 2672 8182 2692
rect 7760 2604 8156 2632
rect 7932 2304 7984 2310
rect 7932 2246 7984 2252
rect 7944 2106 7972 2246
rect 7932 2100 7984 2106
rect 7932 2042 7984 2048
rect 8128 800 8156 2604
rect 8312 2582 8340 2790
rect 8404 2650 8432 2858
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 8300 2576 8352 2582
rect 8300 2518 8352 2524
rect 8404 2310 8432 2586
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 8588 800 8616 13806
rect 8852 12912 8904 12918
rect 8852 12854 8904 12860
rect 8760 12640 8812 12646
rect 8760 12582 8812 12588
rect 8772 10198 8800 12582
rect 8864 12442 8892 12854
rect 8956 12782 8984 13942
rect 9140 13870 9168 15506
rect 9600 15026 9628 15914
rect 10060 15706 10088 16662
rect 10244 16590 10272 17002
rect 10336 16998 10364 17614
rect 10324 16992 10376 16998
rect 10324 16934 10376 16940
rect 10336 16726 10364 16934
rect 10324 16720 10376 16726
rect 10324 16662 10376 16668
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 10232 16584 10284 16590
rect 10232 16526 10284 16532
rect 10152 15978 10180 16526
rect 10140 15972 10192 15978
rect 10140 15914 10192 15920
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 9588 15020 9640 15026
rect 9588 14962 9640 14968
rect 9600 14618 9628 14962
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 9600 13938 9628 14418
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 9128 13864 9180 13870
rect 9128 13806 9180 13812
rect 9404 13864 9456 13870
rect 9404 13806 9456 13812
rect 8944 12776 8996 12782
rect 8944 12718 8996 12724
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 9232 11558 9260 12038
rect 9416 11778 9444 13806
rect 10048 13456 10100 13462
rect 10048 13398 10100 13404
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 9600 12442 9628 12718
rect 9588 12436 9640 12442
rect 9588 12378 9640 12384
rect 9956 12300 10008 12306
rect 10060 12288 10088 13398
rect 10612 12986 10640 19110
rect 10796 18970 10824 21762
rect 11352 20700 11648 20720
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11430 20646 11432 20698
rect 11494 20646 11506 20698
rect 11568 20646 11570 20698
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11352 20624 11648 20644
rect 18282 20700 18578 20720
rect 18338 20698 18362 20700
rect 18418 20698 18442 20700
rect 18498 20698 18522 20700
rect 18360 20646 18362 20698
rect 18424 20646 18436 20698
rect 18498 20646 18500 20698
rect 18338 20644 18362 20646
rect 18418 20644 18442 20646
rect 18498 20644 18522 20646
rect 18282 20624 18578 20644
rect 14817 20156 15113 20176
rect 14873 20154 14897 20156
rect 14953 20154 14977 20156
rect 15033 20154 15057 20156
rect 14895 20102 14897 20154
rect 14959 20102 14971 20154
rect 15033 20102 15035 20154
rect 14873 20100 14897 20102
rect 14953 20100 14977 20102
rect 15033 20100 15057 20102
rect 14817 20080 15113 20100
rect 11352 19612 11648 19632
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11430 19558 11432 19610
rect 11494 19558 11506 19610
rect 11568 19558 11570 19610
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11352 19536 11648 19556
rect 18282 19612 18578 19632
rect 18338 19610 18362 19612
rect 18418 19610 18442 19612
rect 18498 19610 18522 19612
rect 18360 19558 18362 19610
rect 18424 19558 18436 19610
rect 18498 19558 18500 19610
rect 18338 19556 18362 19558
rect 18418 19556 18442 19558
rect 18498 19556 18522 19558
rect 18282 19536 18578 19556
rect 14817 19068 15113 19088
rect 14873 19066 14897 19068
rect 14953 19066 14977 19068
rect 15033 19066 15057 19068
rect 14895 19014 14897 19066
rect 14959 19014 14971 19066
rect 15033 19014 15035 19066
rect 14873 19012 14897 19014
rect 14953 19012 14977 19014
rect 15033 19012 15057 19014
rect 14817 18992 15113 19012
rect 10784 18964 10836 18970
rect 10784 18906 10836 18912
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 11072 18290 11100 18770
rect 11352 18524 11648 18544
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11430 18470 11432 18522
rect 11494 18470 11506 18522
rect 11568 18470 11570 18522
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11352 18448 11648 18468
rect 18282 18524 18578 18544
rect 18338 18522 18362 18524
rect 18418 18522 18442 18524
rect 18498 18522 18522 18524
rect 18360 18470 18362 18522
rect 18424 18470 18436 18522
rect 18498 18470 18500 18522
rect 18338 18468 18362 18470
rect 18418 18468 18442 18470
rect 18498 18468 18522 18470
rect 18282 18448 18578 18468
rect 11060 18284 11112 18290
rect 11060 18226 11112 18232
rect 11428 18216 11480 18222
rect 11428 18158 11480 18164
rect 11440 17882 11468 18158
rect 14817 17980 15113 18000
rect 14873 17978 14897 17980
rect 14953 17978 14977 17980
rect 15033 17978 15057 17980
rect 14895 17926 14897 17978
rect 14959 17926 14971 17978
rect 15033 17926 15035 17978
rect 14873 17924 14897 17926
rect 14953 17924 14977 17926
rect 15033 17924 15057 17926
rect 14817 17904 15113 17924
rect 11428 17876 11480 17882
rect 11428 17818 11480 17824
rect 12440 17740 12492 17746
rect 12440 17682 12492 17688
rect 11888 17672 11940 17678
rect 11888 17614 11940 17620
rect 11352 17436 11648 17456
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11430 17382 11432 17434
rect 11494 17382 11506 17434
rect 11568 17382 11570 17434
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11352 17360 11648 17380
rect 10692 16584 10744 16590
rect 10692 16526 10744 16532
rect 10704 13462 10732 16526
rect 11352 16348 11648 16368
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11430 16294 11432 16346
rect 11494 16294 11506 16346
rect 11568 16294 11570 16346
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11352 16272 11648 16292
rect 11900 16250 11928 17614
rect 12452 17202 12480 17682
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 13740 16794 13768 17614
rect 18282 17436 18578 17456
rect 18338 17434 18362 17436
rect 18418 17434 18442 17436
rect 18498 17434 18522 17436
rect 18360 17382 18362 17434
rect 18424 17382 18436 17434
rect 18498 17382 18500 17434
rect 18338 17380 18362 17382
rect 18418 17380 18442 17382
rect 18498 17380 18522 17382
rect 18282 17360 18578 17380
rect 19246 17232 19302 17241
rect 19246 17167 19302 17176
rect 14817 16892 15113 16912
rect 14873 16890 14897 16892
rect 14953 16890 14977 16892
rect 15033 16890 15057 16892
rect 14895 16838 14897 16890
rect 14959 16838 14971 16890
rect 15033 16838 15035 16890
rect 14873 16836 14897 16838
rect 14953 16836 14977 16838
rect 15033 16836 15057 16838
rect 14817 16816 15113 16836
rect 19260 16794 19288 17167
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 19248 16788 19300 16794
rect 19248 16730 19300 16736
rect 11980 16720 12032 16726
rect 11980 16662 12032 16668
rect 11888 16244 11940 16250
rect 11888 16186 11940 16192
rect 11992 16114 12020 16662
rect 12348 16652 12400 16658
rect 12348 16594 12400 16600
rect 11980 16108 12032 16114
rect 11980 16050 12032 16056
rect 11980 15972 12032 15978
rect 11980 15914 12032 15920
rect 11152 15428 11204 15434
rect 11152 15370 11204 15376
rect 10876 14476 10928 14482
rect 10876 14418 10928 14424
rect 10888 14074 10916 14418
rect 10876 14068 10928 14074
rect 10876 14010 10928 14016
rect 10876 13796 10928 13802
rect 10876 13738 10928 13744
rect 10888 13530 10916 13738
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10692 13456 10744 13462
rect 10692 13398 10744 13404
rect 10600 12980 10652 12986
rect 10600 12922 10652 12928
rect 10888 12918 10916 13466
rect 11060 13388 11112 13394
rect 11060 13330 11112 13336
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 10876 12912 10928 12918
rect 10876 12854 10928 12860
rect 10876 12776 10928 12782
rect 10876 12718 10928 12724
rect 10008 12260 10180 12288
rect 9956 12242 10008 12248
rect 9416 11750 9628 11778
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 9128 10804 9180 10810
rect 9128 10746 9180 10752
rect 8944 10464 8996 10470
rect 8944 10406 8996 10412
rect 8956 10266 8984 10406
rect 8944 10260 8996 10266
rect 8944 10202 8996 10208
rect 8760 10192 8812 10198
rect 8760 10134 8812 10140
rect 8772 9178 8800 10134
rect 8760 9172 8812 9178
rect 8760 9114 8812 9120
rect 8944 8832 8996 8838
rect 8944 8774 8996 8780
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8864 7002 8892 7890
rect 8852 6996 8904 7002
rect 8852 6938 8904 6944
rect 8956 6225 8984 8774
rect 9036 7880 9088 7886
rect 9036 7822 9088 7828
rect 9048 7546 9076 7822
rect 9036 7540 9088 7546
rect 9036 7482 9088 7488
rect 9140 7426 9168 10746
rect 9232 10062 9260 11494
rect 9416 11082 9444 11630
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 9324 10266 9352 10406
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9232 9450 9260 9998
rect 9220 9444 9272 9450
rect 9220 9386 9272 9392
rect 9048 7398 9168 7426
rect 9218 7440 9274 7449
rect 8942 6216 8998 6225
rect 8942 6151 8998 6160
rect 8668 5772 8720 5778
rect 8668 5714 8720 5720
rect 8680 5234 8708 5714
rect 8668 5228 8720 5234
rect 8668 5170 8720 5176
rect 9048 800 9076 7398
rect 9218 7375 9274 7384
rect 9232 5574 9260 7375
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 9324 6662 9352 7278
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9324 6254 9352 6598
rect 9312 6248 9364 6254
rect 9312 6190 9364 6196
rect 9220 5568 9272 5574
rect 9220 5510 9272 5516
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 9324 4010 9352 4558
rect 9312 4004 9364 4010
rect 9312 3946 9364 3952
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 9140 2650 9168 3878
rect 9220 3596 9272 3602
rect 9220 3538 9272 3544
rect 9128 2644 9180 2650
rect 9128 2586 9180 2592
rect 9232 2446 9260 3538
rect 9220 2440 9272 2446
rect 9220 2382 9272 2388
rect 9416 800 9444 11018
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 9508 9382 9536 10610
rect 9600 10130 9628 11750
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9876 11286 9904 11698
rect 10048 11620 10100 11626
rect 10048 11562 10100 11568
rect 10060 11286 10088 11562
rect 10152 11354 10180 12260
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 9864 11280 9916 11286
rect 9864 11222 9916 11228
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9692 11064 9720 11154
rect 9692 11036 9904 11064
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9496 9376 9548 9382
rect 9496 9318 9548 9324
rect 9508 8974 9536 9318
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 9600 8838 9628 10066
rect 9692 9178 9720 10406
rect 9876 9518 9904 11036
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 9864 9512 9916 9518
rect 9864 9454 9916 9460
rect 10336 9450 10364 9998
rect 10508 9512 10560 9518
rect 10508 9454 10560 9460
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 10324 9444 10376 9450
rect 10324 9386 10376 9392
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 10060 8498 10088 8978
rect 10336 8974 10364 9386
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 10520 7954 10548 9454
rect 10600 8900 10652 8906
rect 10600 8842 10652 8848
rect 10612 8430 10640 8842
rect 10796 8838 10824 9454
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10508 7948 10560 7954
rect 10508 7890 10560 7896
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9968 6390 9996 7142
rect 10508 6656 10560 6662
rect 10508 6598 10560 6604
rect 9956 6384 10008 6390
rect 9956 6326 10008 6332
rect 9968 5930 9996 6326
rect 10520 6254 10548 6598
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 9876 5902 9996 5930
rect 9876 5166 9904 5902
rect 9956 5840 10008 5846
rect 9956 5782 10008 5788
rect 9968 5234 9996 5782
rect 10520 5778 10548 6190
rect 10508 5772 10560 5778
rect 10508 5714 10560 5720
rect 9956 5228 10008 5234
rect 9956 5170 10008 5176
rect 9864 5160 9916 5166
rect 9864 5102 9916 5108
rect 10138 5128 10194 5137
rect 10138 5063 10194 5072
rect 9772 5024 9824 5030
rect 9772 4966 9824 4972
rect 9784 4554 9812 4966
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 9772 4548 9824 4554
rect 9772 4490 9824 4496
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9692 3602 9720 4422
rect 9772 4004 9824 4010
rect 9772 3946 9824 3952
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 9508 3194 9536 3538
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 9692 2582 9720 3334
rect 9784 2650 9812 3946
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 9876 2990 9904 3878
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 9968 2836 9996 4762
rect 10152 4690 10180 5063
rect 10140 4684 10192 4690
rect 10140 4626 10192 4632
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10140 4548 10192 4554
rect 10140 4490 10192 4496
rect 10152 3738 10180 4490
rect 10416 4140 10468 4146
rect 10416 4082 10468 4088
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 10048 3596 10100 3602
rect 10048 3538 10100 3544
rect 10060 3398 10088 3538
rect 10048 3392 10100 3398
rect 10048 3334 10100 3340
rect 9876 2808 9996 2836
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 9680 2576 9732 2582
rect 9680 2518 9732 2524
rect 9876 800 9904 2808
rect 10244 2378 10272 3878
rect 10428 3466 10456 4082
rect 10520 4010 10548 4558
rect 10612 4078 10640 8366
rect 10796 7274 10824 8774
rect 10784 7268 10836 7274
rect 10784 7210 10836 7216
rect 10692 7200 10744 7206
rect 10692 7142 10744 7148
rect 10704 5846 10732 7142
rect 10692 5840 10744 5846
rect 10692 5782 10744 5788
rect 10796 5692 10824 7210
rect 10704 5664 10824 5692
rect 10600 4072 10652 4078
rect 10600 4014 10652 4020
rect 10508 4004 10560 4010
rect 10508 3946 10560 3952
rect 10416 3460 10468 3466
rect 10416 3402 10468 3408
rect 10704 3398 10732 5664
rect 10888 4826 10916 12718
rect 10980 12646 11008 13126
rect 11072 12850 11100 13330
rect 11060 12844 11112 12850
rect 11060 12786 11112 12792
rect 10968 12640 11020 12646
rect 10968 12582 11020 12588
rect 11072 12442 11100 12786
rect 11060 12436 11112 12442
rect 11060 12378 11112 12384
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 11072 11694 11100 12242
rect 11060 11688 11112 11694
rect 11060 11630 11112 11636
rect 11072 11354 11100 11630
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 11164 11234 11192 15370
rect 11352 15260 11648 15280
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11430 15206 11432 15258
rect 11494 15206 11506 15258
rect 11568 15206 11570 15258
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11352 15184 11648 15204
rect 11244 14816 11296 14822
rect 11244 14758 11296 14764
rect 11256 14074 11284 14758
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11352 14172 11648 14192
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11430 14118 11432 14170
rect 11494 14118 11506 14170
rect 11568 14118 11570 14170
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11352 14096 11648 14116
rect 11244 14068 11296 14074
rect 11244 14010 11296 14016
rect 11716 13870 11744 14214
rect 11704 13864 11756 13870
rect 11704 13806 11756 13812
rect 11888 13728 11940 13734
rect 11888 13670 11940 13676
rect 11900 13190 11928 13670
rect 11888 13184 11940 13190
rect 11888 13126 11940 13132
rect 11352 13084 11648 13104
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11430 13030 11432 13082
rect 11494 13030 11506 13082
rect 11568 13030 11570 13082
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11352 13008 11648 13028
rect 11704 12368 11756 12374
rect 11704 12310 11756 12316
rect 11352 11996 11648 12016
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11430 11942 11432 11994
rect 11494 11942 11506 11994
rect 11568 11942 11570 11994
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11352 11920 11648 11940
rect 11716 11694 11744 12310
rect 11704 11688 11756 11694
rect 11704 11630 11756 11636
rect 10980 11206 11192 11234
rect 11244 11212 11296 11218
rect 10876 4820 10928 4826
rect 10876 4762 10928 4768
rect 10980 4706 11008 11206
rect 11244 11154 11296 11160
rect 11060 11008 11112 11014
rect 11060 10950 11112 10956
rect 11072 9518 11100 10950
rect 11256 10606 11284 11154
rect 11352 10908 11648 10928
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11430 10854 11432 10906
rect 11494 10854 11506 10906
rect 11568 10854 11570 10906
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11352 10832 11648 10852
rect 11796 10736 11848 10742
rect 11796 10678 11848 10684
rect 11244 10600 11296 10606
rect 11244 10542 11296 10548
rect 11256 10266 11284 10542
rect 11244 10260 11296 10266
rect 11244 10202 11296 10208
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 11072 9178 11100 9454
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 11060 8900 11112 8906
rect 11060 8842 11112 8848
rect 11072 5658 11100 8842
rect 11256 8634 11284 10066
rect 11352 9820 11648 9840
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11430 9766 11432 9818
rect 11494 9766 11506 9818
rect 11568 9766 11570 9818
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11352 9744 11648 9764
rect 11716 9518 11744 10066
rect 11704 9512 11756 9518
rect 11704 9454 11756 9460
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 11716 8974 11744 9114
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11352 8732 11648 8752
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11430 8678 11432 8730
rect 11494 8678 11506 8730
rect 11568 8678 11570 8730
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11352 8656 11648 8676
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 11716 8242 11744 8910
rect 11808 8430 11836 10678
rect 11900 8430 11928 13126
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11992 8242 12020 15914
rect 12164 12436 12216 12442
rect 12164 12378 12216 12384
rect 12176 8786 12204 12378
rect 12360 10810 12388 16594
rect 18282 16348 18578 16368
rect 18338 16346 18362 16348
rect 18418 16346 18442 16348
rect 18498 16346 18522 16348
rect 18360 16294 18362 16346
rect 18424 16294 18436 16346
rect 18498 16294 18500 16346
rect 18338 16292 18362 16294
rect 18418 16292 18442 16294
rect 18498 16292 18522 16294
rect 18282 16272 18578 16292
rect 12440 15904 12492 15910
rect 12440 15846 12492 15852
rect 12452 12442 12480 15846
rect 14817 15804 15113 15824
rect 14873 15802 14897 15804
rect 14953 15802 14977 15804
rect 15033 15802 15057 15804
rect 14895 15750 14897 15802
rect 14959 15750 14971 15802
rect 15033 15750 15035 15802
rect 14873 15748 14897 15750
rect 14953 15748 14977 15750
rect 15033 15748 15057 15750
rect 14817 15728 15113 15748
rect 18282 15260 18578 15280
rect 18338 15258 18362 15260
rect 18418 15258 18442 15260
rect 18498 15258 18522 15260
rect 18360 15206 18362 15258
rect 18424 15206 18436 15258
rect 18498 15206 18500 15258
rect 18338 15204 18362 15206
rect 18418 15204 18442 15206
rect 18498 15204 18522 15206
rect 18282 15184 18578 15204
rect 14817 14716 15113 14736
rect 14873 14714 14897 14716
rect 14953 14714 14977 14716
rect 15033 14714 15057 14716
rect 14895 14662 14897 14714
rect 14959 14662 14971 14714
rect 15033 14662 15035 14714
rect 14873 14660 14897 14662
rect 14953 14660 14977 14662
rect 15033 14660 15057 14662
rect 14817 14640 15113 14660
rect 18282 14172 18578 14192
rect 18338 14170 18362 14172
rect 18418 14170 18442 14172
rect 18498 14170 18522 14172
rect 18360 14118 18362 14170
rect 18424 14118 18436 14170
rect 18498 14118 18500 14170
rect 18338 14116 18362 14118
rect 18418 14116 18442 14118
rect 18498 14116 18522 14118
rect 18282 14096 18578 14116
rect 14817 13628 15113 13648
rect 14873 13626 14897 13628
rect 14953 13626 14977 13628
rect 15033 13626 15057 13628
rect 14895 13574 14897 13626
rect 14959 13574 14971 13626
rect 15033 13574 15035 13626
rect 14873 13572 14897 13574
rect 14953 13572 14977 13574
rect 15033 13572 15057 13574
rect 14817 13552 15113 13572
rect 18282 13084 18578 13104
rect 18338 13082 18362 13084
rect 18418 13082 18442 13084
rect 18498 13082 18522 13084
rect 18360 13030 18362 13082
rect 18424 13030 18436 13082
rect 18498 13030 18500 13082
rect 18338 13028 18362 13030
rect 18418 13028 18442 13030
rect 18498 13028 18522 13030
rect 18282 13008 18578 13028
rect 14817 12540 15113 12560
rect 14873 12538 14897 12540
rect 14953 12538 14977 12540
rect 15033 12538 15057 12540
rect 14895 12486 14897 12538
rect 14959 12486 14971 12538
rect 15033 12486 15035 12538
rect 14873 12484 14897 12486
rect 14953 12484 14977 12486
rect 15033 12484 15057 12486
rect 14817 12464 15113 12484
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 19708 12436 19760 12442
rect 19708 12378 19760 12384
rect 19720 12306 19748 12378
rect 19708 12300 19760 12306
rect 19708 12242 19760 12248
rect 20536 12096 20588 12102
rect 20536 12038 20588 12044
rect 18282 11996 18578 12016
rect 18338 11994 18362 11996
rect 18418 11994 18442 11996
rect 18498 11994 18522 11996
rect 18360 11942 18362 11994
rect 18424 11942 18436 11994
rect 18498 11942 18500 11994
rect 18338 11940 18362 11942
rect 18418 11940 18442 11942
rect 18498 11940 18522 11942
rect 18282 11920 18578 11940
rect 20076 11552 20128 11558
rect 20076 11494 20128 11500
rect 14817 11452 15113 11472
rect 14873 11450 14897 11452
rect 14953 11450 14977 11452
rect 15033 11450 15057 11452
rect 14895 11398 14897 11450
rect 14959 11398 14971 11450
rect 15033 11398 15035 11450
rect 14873 11396 14897 11398
rect 14953 11396 14977 11398
rect 15033 11396 15057 11398
rect 14817 11376 15113 11396
rect 19524 11076 19576 11082
rect 19524 11018 19576 11024
rect 18282 10908 18578 10928
rect 18338 10906 18362 10908
rect 18418 10906 18442 10908
rect 18498 10906 18522 10908
rect 18360 10854 18362 10906
rect 18424 10854 18436 10906
rect 18498 10854 18500 10906
rect 18338 10852 18362 10854
rect 18418 10852 18442 10854
rect 18498 10852 18522 10854
rect 18282 10832 18578 10852
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 12360 9926 12388 10746
rect 19156 10736 19208 10742
rect 19156 10678 19208 10684
rect 14817 10364 15113 10384
rect 14873 10362 14897 10364
rect 14953 10362 14977 10364
rect 15033 10362 15057 10364
rect 14895 10310 14897 10362
rect 14959 10310 14971 10362
rect 15033 10310 15035 10362
rect 14873 10308 14897 10310
rect 14953 10308 14977 10310
rect 15033 10308 15057 10310
rect 14817 10288 15113 10308
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12360 9654 12388 9862
rect 12348 9648 12400 9654
rect 12348 9590 12400 9596
rect 12360 9178 12388 9590
rect 12544 9586 12572 9862
rect 18282 9820 18578 9840
rect 18338 9818 18362 9820
rect 18418 9818 18442 9820
rect 18498 9818 18522 9820
rect 18360 9766 18362 9818
rect 18424 9766 18436 9818
rect 18498 9766 18500 9818
rect 18338 9764 18362 9766
rect 18418 9764 18442 9766
rect 18498 9764 18522 9766
rect 18282 9744 18578 9764
rect 14188 9716 14240 9722
rect 14188 9658 14240 9664
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 12544 9110 12572 9522
rect 12624 9376 12676 9382
rect 12624 9318 12676 9324
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 12532 9104 12584 9110
rect 12532 9046 12584 9052
rect 12176 8758 12388 8786
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 11624 8214 11744 8242
rect 11808 8214 12020 8242
rect 11624 7886 11652 8214
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11612 7880 11664 7886
rect 11612 7822 11664 7828
rect 11352 7644 11648 7664
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11430 7590 11432 7642
rect 11494 7590 11506 7642
rect 11568 7590 11570 7642
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11352 7568 11648 7588
rect 11612 7404 11664 7410
rect 11716 7392 11744 7890
rect 11664 7364 11744 7392
rect 11612 7346 11664 7352
rect 11624 7274 11652 7346
rect 11612 7268 11664 7274
rect 11612 7210 11664 7216
rect 11244 7200 11296 7206
rect 11244 7142 11296 7148
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11256 6866 11284 7142
rect 11348 6934 11376 7142
rect 11336 6928 11388 6934
rect 11336 6870 11388 6876
rect 11244 6860 11296 6866
rect 11244 6802 11296 6808
rect 11352 6556 11648 6576
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11430 6502 11432 6554
rect 11494 6502 11506 6554
rect 11568 6502 11570 6554
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11352 6480 11648 6500
rect 11808 6338 11836 8214
rect 11888 7948 11940 7954
rect 11888 7890 11940 7896
rect 11900 7750 11928 7890
rect 11888 7744 11940 7750
rect 11888 7686 11940 7692
rect 11900 6798 11928 7686
rect 12176 6866 12204 8570
rect 12256 8424 12308 8430
rect 12256 8366 12308 8372
rect 12164 6860 12216 6866
rect 12164 6802 12216 6808
rect 11888 6792 11940 6798
rect 11888 6734 11940 6740
rect 11716 6310 11836 6338
rect 11072 5630 11284 5658
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 11072 5234 11100 5510
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 11072 4758 11100 5170
rect 10796 4678 11008 4706
rect 11060 4752 11112 4758
rect 11060 4694 11112 4700
rect 10692 3392 10744 3398
rect 10692 3334 10744 3340
rect 10324 3188 10376 3194
rect 10324 3130 10376 3136
rect 10232 2372 10284 2378
rect 10232 2314 10284 2320
rect 10336 800 10364 3130
rect 10704 2922 10732 3334
rect 10692 2916 10744 2922
rect 10692 2858 10744 2864
rect 10416 2848 10468 2854
rect 10416 2790 10468 2796
rect 10428 2650 10456 2790
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 10796 800 10824 4678
rect 10876 4276 10928 4282
rect 10876 4218 10928 4224
rect 10888 3534 10916 4218
rect 11256 3942 11284 5630
rect 11352 5468 11648 5488
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11430 5414 11432 5466
rect 11494 5414 11506 5466
rect 11568 5414 11570 5466
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11352 5392 11648 5412
rect 11352 4380 11648 4400
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11430 4326 11432 4378
rect 11494 4326 11506 4378
rect 11568 4326 11570 4378
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11352 4304 11648 4324
rect 11428 4140 11480 4146
rect 11428 4082 11480 4088
rect 10968 3936 11020 3942
rect 10968 3878 11020 3884
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 10980 3670 11008 3878
rect 11440 3738 11468 4082
rect 11428 3732 11480 3738
rect 11428 3674 11480 3680
rect 10968 3664 11020 3670
rect 11716 3618 11744 6310
rect 11796 6180 11848 6186
rect 11796 6122 11848 6128
rect 11808 5710 11836 6122
rect 12164 5840 12216 5846
rect 12164 5782 12216 5788
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11992 5370 12020 5714
rect 12176 5370 12204 5782
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 12164 5364 12216 5370
rect 12164 5306 12216 5312
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 10968 3606 11020 3612
rect 11256 3590 11744 3618
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10888 3058 10916 3470
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 10876 2848 10928 2854
rect 10876 2790 10928 2796
rect 10888 2310 10916 2790
rect 10876 2304 10928 2310
rect 10876 2246 10928 2252
rect 11256 800 11284 3590
rect 11808 3516 11836 4966
rect 12072 4072 12124 4078
rect 12072 4014 12124 4020
rect 11716 3488 11836 3516
rect 11352 3292 11648 3312
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11430 3238 11432 3290
rect 11494 3238 11506 3290
rect 11568 3238 11570 3290
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11352 3216 11648 3236
rect 11352 2204 11648 2224
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11430 2150 11432 2202
rect 11494 2150 11506 2202
rect 11568 2150 11570 2202
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11352 2128 11648 2148
rect 11716 800 11744 3488
rect 11888 2916 11940 2922
rect 11888 2858 11940 2864
rect 11900 2514 11928 2858
rect 11888 2508 11940 2514
rect 11888 2450 11940 2456
rect 12084 800 12112 4014
rect 12176 2854 12204 5306
rect 12268 3194 12296 8366
rect 12360 6338 12388 8758
rect 12636 8566 12664 9318
rect 12624 8560 12676 8566
rect 12624 8502 12676 8508
rect 12820 8498 12848 9318
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 13360 8356 13412 8362
rect 13360 8298 13412 8304
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12992 7200 13044 7206
rect 12992 7142 13044 7148
rect 12452 7002 12480 7142
rect 12440 6996 12492 7002
rect 12440 6938 12492 6944
rect 12440 6792 12492 6798
rect 12440 6734 12492 6740
rect 12452 6458 12480 6734
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12360 6310 12480 6338
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 12360 4078 12388 6190
rect 12452 5030 12480 6310
rect 12544 5846 12572 6598
rect 12532 5840 12584 5846
rect 12532 5782 12584 5788
rect 12716 5772 12768 5778
rect 12716 5714 12768 5720
rect 12728 5234 12756 5714
rect 12808 5568 12860 5574
rect 12808 5510 12860 5516
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 12452 4214 12480 4422
rect 12440 4208 12492 4214
rect 12440 4150 12492 4156
rect 12348 4072 12400 4078
rect 12348 4014 12400 4020
rect 12622 3496 12678 3505
rect 12622 3431 12678 3440
rect 12256 3188 12308 3194
rect 12256 3130 12308 3136
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 12164 2848 12216 2854
rect 12164 2790 12216 2796
rect 12452 2582 12480 2926
rect 12440 2576 12492 2582
rect 12440 2518 12492 2524
rect 12636 2514 12664 3431
rect 12820 2990 12848 5510
rect 13004 5302 13032 7142
rect 13084 6248 13136 6254
rect 13084 6190 13136 6196
rect 13096 5710 13124 6190
rect 13084 5704 13136 5710
rect 13084 5646 13136 5652
rect 13268 5568 13320 5574
rect 13268 5510 13320 5516
rect 13280 5370 13308 5510
rect 13268 5364 13320 5370
rect 13268 5306 13320 5312
rect 12992 5296 13044 5302
rect 12992 5238 13044 5244
rect 13372 5234 13400 8298
rect 14096 8288 14148 8294
rect 14096 8230 14148 8236
rect 13636 7880 13688 7886
rect 13636 7822 13688 7828
rect 13648 7206 13676 7822
rect 14108 7342 14136 8230
rect 14200 8022 14228 9658
rect 14648 9444 14700 9450
rect 14648 9386 14700 9392
rect 14372 9036 14424 9042
rect 14372 8978 14424 8984
rect 14188 8016 14240 8022
rect 14188 7958 14240 7964
rect 14096 7336 14148 7342
rect 14096 7278 14148 7284
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13648 7002 13676 7142
rect 13636 6996 13688 7002
rect 13636 6938 13688 6944
rect 13820 6792 13872 6798
rect 13820 6734 13872 6740
rect 13832 6458 13860 6734
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 14108 6254 14136 7278
rect 14280 6656 14332 6662
rect 14280 6598 14332 6604
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 14292 5778 14320 6598
rect 14280 5772 14332 5778
rect 14280 5714 14332 5720
rect 14384 5234 14412 8978
rect 14660 8974 14688 9386
rect 14817 9276 15113 9296
rect 14873 9274 14897 9276
rect 14953 9274 14977 9276
rect 15033 9274 15057 9276
rect 14895 9222 14897 9274
rect 14959 9222 14971 9274
rect 15033 9222 15035 9274
rect 14873 9220 14897 9222
rect 14953 9220 14977 9222
rect 15033 9220 15057 9222
rect 14817 9200 15113 9220
rect 15108 9036 15160 9042
rect 15108 8978 15160 8984
rect 14556 8968 14608 8974
rect 14556 8910 14608 8916
rect 14648 8968 14700 8974
rect 14648 8910 14700 8916
rect 14464 8356 14516 8362
rect 14464 8298 14516 8304
rect 14476 7886 14504 8298
rect 14568 8090 14596 8910
rect 14660 8634 14688 8910
rect 14648 8628 14700 8634
rect 14648 8570 14700 8576
rect 15120 8498 15148 8978
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 14817 8188 15113 8208
rect 14873 8186 14897 8188
rect 14953 8186 14977 8188
rect 15033 8186 15057 8188
rect 14895 8134 14897 8186
rect 14959 8134 14971 8186
rect 15033 8134 15035 8186
rect 14873 8132 14897 8134
rect 14953 8132 14977 8134
rect 15033 8132 15057 8134
rect 14817 8112 15113 8132
rect 14556 8084 14608 8090
rect 14556 8026 14608 8032
rect 16500 7954 16528 8774
rect 18282 8732 18578 8752
rect 18338 8730 18362 8732
rect 18418 8730 18442 8732
rect 18498 8730 18522 8732
rect 18360 8678 18362 8730
rect 18424 8678 18436 8730
rect 18498 8678 18500 8730
rect 18338 8676 18362 8678
rect 18418 8676 18442 8678
rect 18498 8676 18522 8678
rect 18282 8656 18578 8676
rect 18604 8356 18656 8362
rect 18604 8298 18656 8304
rect 16488 7948 16540 7954
rect 16488 7890 16540 7896
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 17500 7880 17552 7886
rect 17500 7822 17552 7828
rect 14476 7546 14504 7822
rect 14464 7540 14516 7546
rect 14464 7482 14516 7488
rect 14740 7268 14792 7274
rect 14740 7210 14792 7216
rect 14752 6882 14780 7210
rect 14817 7100 15113 7120
rect 14873 7098 14897 7100
rect 14953 7098 14977 7100
rect 15033 7098 15057 7100
rect 14895 7046 14897 7098
rect 14959 7046 14971 7098
rect 15033 7046 15035 7098
rect 14873 7044 14897 7046
rect 14953 7044 14977 7046
rect 15033 7044 15057 7046
rect 14817 7024 15113 7044
rect 15200 6928 15252 6934
rect 14752 6854 14872 6882
rect 15200 6870 15252 6876
rect 14844 6798 14872 6854
rect 14832 6792 14884 6798
rect 14832 6734 14884 6740
rect 14844 6458 14872 6734
rect 14832 6452 14884 6458
rect 14832 6394 14884 6400
rect 14817 6012 15113 6032
rect 14873 6010 14897 6012
rect 14953 6010 14977 6012
rect 15033 6010 15057 6012
rect 14895 5958 14897 6010
rect 14959 5958 14971 6010
rect 15033 5958 15035 6010
rect 14873 5956 14897 5958
rect 14953 5956 14977 5958
rect 15033 5956 15057 5958
rect 14817 5936 15113 5956
rect 15212 5914 15240 6870
rect 15292 6724 15344 6730
rect 15292 6666 15344 6672
rect 15200 5908 15252 5914
rect 15200 5850 15252 5856
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 14096 5228 14148 5234
rect 14096 5170 14148 5176
rect 14372 5228 14424 5234
rect 14372 5170 14424 5176
rect 13176 5024 13228 5030
rect 13176 4966 13228 4972
rect 13188 3738 13216 4966
rect 13636 4684 13688 4690
rect 13636 4626 13688 4632
rect 13648 3942 13676 4626
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 13832 4078 13860 4422
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 13636 3936 13688 3942
rect 13636 3878 13688 3884
rect 13176 3732 13228 3738
rect 13176 3674 13228 3680
rect 13648 3534 13676 3878
rect 14108 3738 14136 5170
rect 14384 4826 14412 5170
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 14188 4480 14240 4486
rect 14188 4422 14240 4428
rect 14200 4078 14228 4422
rect 14188 4072 14240 4078
rect 14188 4014 14240 4020
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14096 3732 14148 3738
rect 14096 3674 14148 3680
rect 14384 3534 14412 4014
rect 13268 3528 13320 3534
rect 13268 3470 13320 3476
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 14372 3528 14424 3534
rect 14372 3470 14424 3476
rect 13280 2990 13308 3470
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13820 3392 13872 3398
rect 13820 3334 13872 3340
rect 13740 3058 13768 3334
rect 13832 3194 13860 3334
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 12808 2984 12860 2990
rect 12808 2926 12860 2932
rect 13268 2984 13320 2990
rect 13268 2926 13320 2932
rect 12716 2916 12768 2922
rect 12716 2858 12768 2864
rect 13728 2916 13780 2922
rect 13728 2858 13780 2864
rect 12728 2514 12756 2858
rect 13740 2514 13768 2858
rect 13912 2848 13964 2854
rect 13912 2790 13964 2796
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 12716 2508 12768 2514
rect 12716 2450 12768 2456
rect 13728 2508 13780 2514
rect 13728 2450 13780 2456
rect 12532 2304 12584 2310
rect 12532 2246 12584 2252
rect 12992 2304 13044 2310
rect 12992 2246 13044 2252
rect 13452 2304 13504 2310
rect 13452 2246 13504 2252
rect 12544 800 12572 2246
rect 13004 800 13032 2246
rect 13464 800 13492 2246
rect 13924 800 13952 2790
rect 14476 2514 14504 5646
rect 14817 4924 15113 4944
rect 14873 4922 14897 4924
rect 14953 4922 14977 4924
rect 15033 4922 15057 4924
rect 14895 4870 14897 4922
rect 14959 4870 14971 4922
rect 15033 4870 15035 4922
rect 14873 4868 14897 4870
rect 14953 4868 14977 4870
rect 15033 4868 15057 4870
rect 14817 4848 15113 4868
rect 14817 3836 15113 3856
rect 14873 3834 14897 3836
rect 14953 3834 14977 3836
rect 15033 3834 15057 3836
rect 14895 3782 14897 3834
rect 14959 3782 14971 3834
rect 15033 3782 15035 3834
rect 14873 3780 14897 3782
rect 14953 3780 14977 3782
rect 15033 3780 15057 3782
rect 14817 3760 15113 3780
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14752 3058 14780 3470
rect 14740 3052 14792 3058
rect 14740 2994 14792 3000
rect 14817 2748 15113 2768
rect 14873 2746 14897 2748
rect 14953 2746 14977 2748
rect 15033 2746 15057 2748
rect 14895 2694 14897 2746
rect 14959 2694 14971 2746
rect 15033 2694 15035 2746
rect 14873 2692 14897 2694
rect 14953 2692 14977 2694
rect 15033 2692 15057 2694
rect 14817 2672 15113 2692
rect 15304 2514 15332 6666
rect 15384 5092 15436 5098
rect 15384 5034 15436 5040
rect 15396 2514 15424 5034
rect 15488 3602 15516 7822
rect 16028 7336 16080 7342
rect 16028 7278 16080 7284
rect 16040 6254 16068 7278
rect 17408 7268 17460 7274
rect 17408 7210 17460 7216
rect 16488 6792 16540 6798
rect 16488 6734 16540 6740
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 16028 6248 16080 6254
rect 16028 6190 16080 6196
rect 16040 5574 16068 6190
rect 16396 5704 16448 5710
rect 16396 5646 16448 5652
rect 16408 5574 16436 5646
rect 16500 5642 16528 6734
rect 17236 6186 17264 6734
rect 17420 6458 17448 7210
rect 17408 6452 17460 6458
rect 17408 6394 17460 6400
rect 17224 6180 17276 6186
rect 17224 6122 17276 6128
rect 16948 6112 17000 6118
rect 16948 6054 17000 6060
rect 16488 5636 16540 5642
rect 16488 5578 16540 5584
rect 16028 5568 16080 5574
rect 16028 5510 16080 5516
rect 16396 5568 16448 5574
rect 16396 5510 16448 5516
rect 16408 5302 16436 5510
rect 16396 5296 16448 5302
rect 16396 5238 16448 5244
rect 16120 5160 16172 5166
rect 16118 5128 16120 5137
rect 16172 5128 16174 5137
rect 16118 5063 16174 5072
rect 15568 5024 15620 5030
rect 15568 4966 15620 4972
rect 16028 5024 16080 5030
rect 16028 4966 16080 4972
rect 15580 4826 15608 4966
rect 15568 4820 15620 4826
rect 15568 4762 15620 4768
rect 16040 4758 16068 4966
rect 16408 4758 16436 5238
rect 16580 5228 16632 5234
rect 16580 5170 16632 5176
rect 16028 4752 16080 4758
rect 16028 4694 16080 4700
rect 16396 4752 16448 4758
rect 16396 4694 16448 4700
rect 16592 4690 16620 5170
rect 15752 4684 15804 4690
rect 15752 4626 15804 4632
rect 16580 4684 16632 4690
rect 16580 4626 16632 4632
rect 15764 4146 15792 4626
rect 16856 4480 16908 4486
rect 16856 4422 16908 4428
rect 15752 4140 15804 4146
rect 15752 4082 15804 4088
rect 15844 4004 15896 4010
rect 15844 3946 15896 3952
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 15660 3392 15712 3398
rect 15660 3334 15712 3340
rect 14464 2508 14516 2514
rect 14464 2450 14516 2456
rect 15292 2508 15344 2514
rect 15292 2450 15344 2456
rect 15384 2508 15436 2514
rect 15384 2450 15436 2456
rect 14280 2304 14332 2310
rect 14280 2246 14332 2252
rect 14740 2304 14792 2310
rect 14740 2246 14792 2252
rect 15200 2304 15252 2310
rect 15200 2246 15252 2252
rect 14292 800 14320 2246
rect 14752 800 14780 2246
rect 15212 800 15240 2246
rect 15672 800 15700 3334
rect 15856 3058 15884 3946
rect 16868 3602 16896 4422
rect 16856 3596 16908 3602
rect 16856 3538 16908 3544
rect 16488 3392 16540 3398
rect 16488 3334 16540 3340
rect 15844 3052 15896 3058
rect 15844 2994 15896 3000
rect 16396 2916 16448 2922
rect 16396 2858 16448 2864
rect 16408 2514 16436 2858
rect 16396 2508 16448 2514
rect 16396 2450 16448 2456
rect 16120 2304 16172 2310
rect 16120 2246 16172 2252
rect 16132 800 16160 2246
rect 16500 800 16528 3334
rect 16960 2990 16988 6054
rect 17236 5574 17264 6122
rect 17316 5772 17368 5778
rect 17316 5714 17368 5720
rect 17224 5568 17276 5574
rect 17224 5510 17276 5516
rect 17236 5234 17264 5510
rect 17224 5228 17276 5234
rect 17224 5170 17276 5176
rect 17132 4684 17184 4690
rect 17132 4626 17184 4632
rect 17144 4282 17172 4626
rect 17328 4554 17356 5714
rect 17316 4548 17368 4554
rect 17316 4490 17368 4496
rect 17132 4276 17184 4282
rect 17132 4218 17184 4224
rect 17512 3602 17540 7822
rect 18282 7644 18578 7664
rect 18338 7642 18362 7644
rect 18418 7642 18442 7644
rect 18498 7642 18522 7644
rect 18360 7590 18362 7642
rect 18424 7590 18436 7642
rect 18498 7590 18500 7642
rect 18338 7588 18362 7590
rect 18418 7588 18442 7590
rect 18498 7588 18522 7590
rect 18282 7568 18578 7588
rect 17684 6656 17736 6662
rect 17684 6598 17736 6604
rect 17696 6254 17724 6598
rect 18282 6556 18578 6576
rect 18338 6554 18362 6556
rect 18418 6554 18442 6556
rect 18498 6554 18522 6556
rect 18360 6502 18362 6554
rect 18424 6502 18436 6554
rect 18498 6502 18500 6554
rect 18338 6500 18362 6502
rect 18418 6500 18442 6502
rect 18498 6500 18522 6502
rect 18282 6480 18578 6500
rect 17684 6248 17736 6254
rect 17684 6190 17736 6196
rect 18144 6112 18196 6118
rect 18144 6054 18196 6060
rect 18156 5370 18184 6054
rect 18282 5468 18578 5488
rect 18338 5466 18362 5468
rect 18418 5466 18442 5468
rect 18498 5466 18522 5468
rect 18360 5414 18362 5466
rect 18424 5414 18436 5466
rect 18498 5414 18500 5466
rect 18338 5412 18362 5414
rect 18418 5412 18442 5414
rect 18498 5412 18522 5414
rect 18282 5392 18578 5412
rect 18144 5364 18196 5370
rect 18144 5306 18196 5312
rect 17960 4684 18012 4690
rect 17960 4626 18012 4632
rect 17972 4146 18000 4626
rect 18282 4380 18578 4400
rect 18338 4378 18362 4380
rect 18418 4378 18442 4380
rect 18498 4378 18522 4380
rect 18360 4326 18362 4378
rect 18424 4326 18436 4378
rect 18498 4326 18500 4378
rect 18338 4324 18362 4326
rect 18418 4324 18442 4326
rect 18498 4324 18522 4326
rect 18282 4304 18578 4324
rect 17960 4140 18012 4146
rect 17960 4082 18012 4088
rect 17500 3596 17552 3602
rect 17500 3538 17552 3544
rect 18052 3528 18104 3534
rect 18052 3470 18104 3476
rect 18064 2990 18092 3470
rect 18144 3392 18196 3398
rect 18144 3334 18196 3340
rect 16948 2984 17000 2990
rect 16948 2926 17000 2932
rect 18052 2984 18104 2990
rect 18052 2926 18104 2932
rect 17408 2916 17460 2922
rect 17408 2858 17460 2864
rect 16948 2848 17000 2854
rect 16948 2790 17000 2796
rect 16960 2650 16988 2790
rect 16948 2644 17000 2650
rect 16948 2586 17000 2592
rect 17420 2514 17448 2858
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 17408 2508 17460 2514
rect 17408 2450 17460 2456
rect 16948 2304 17000 2310
rect 16948 2246 17000 2252
rect 16960 800 16988 2246
rect 17512 1442 17540 2790
rect 17868 2304 17920 2310
rect 17868 2246 17920 2252
rect 17420 1414 17540 1442
rect 17420 800 17448 1414
rect 17880 800 17908 2246
rect 18156 1714 18184 3334
rect 18282 3292 18578 3312
rect 18338 3290 18362 3292
rect 18418 3290 18442 3292
rect 18498 3290 18522 3292
rect 18360 3238 18362 3290
rect 18424 3238 18436 3290
rect 18498 3238 18500 3290
rect 18338 3236 18362 3238
rect 18418 3236 18442 3238
rect 18498 3236 18522 3238
rect 18282 3216 18578 3236
rect 18616 2990 18644 8298
rect 18604 2984 18656 2990
rect 18604 2926 18656 2932
rect 18696 2848 18748 2854
rect 18696 2790 18748 2796
rect 18282 2204 18578 2224
rect 18338 2202 18362 2204
rect 18418 2202 18442 2204
rect 18498 2202 18522 2204
rect 18360 2150 18362 2202
rect 18424 2150 18436 2202
rect 18498 2150 18500 2202
rect 18338 2148 18362 2150
rect 18418 2148 18442 2150
rect 18498 2148 18522 2150
rect 18282 2128 18578 2148
rect 18156 1686 18368 1714
rect 18340 800 18368 1686
rect 18708 800 18736 2790
rect 19168 800 19196 10678
rect 19536 898 19564 11018
rect 19706 3632 19762 3641
rect 19706 3567 19708 3576
rect 19760 3567 19762 3576
rect 19708 3538 19760 3544
rect 19536 870 19656 898
rect 19628 800 19656 870
rect 20088 800 20116 11494
rect 20548 800 20576 12038
rect 20720 10464 20772 10470
rect 20720 10406 20772 10412
rect 20626 5808 20682 5817
rect 20626 5743 20682 5752
rect 20640 5166 20668 5743
rect 20628 5160 20680 5166
rect 20628 5102 20680 5108
rect 20640 4826 20668 5102
rect 20628 4820 20680 4826
rect 20628 4762 20680 4768
rect 20732 3058 20760 10406
rect 21272 5024 21324 5030
rect 21272 4966 21324 4972
rect 20904 3392 20956 3398
rect 20904 3334 20956 3340
rect 20720 3052 20772 3058
rect 20720 2994 20772 3000
rect 20916 800 20944 3334
rect 21284 2122 21312 4966
rect 21824 3936 21876 3942
rect 21824 3878 21876 3884
rect 21836 3602 21864 3878
rect 21824 3596 21876 3602
rect 21824 3538 21876 3544
rect 21364 2984 21416 2990
rect 21364 2926 21416 2932
rect 21376 2310 21404 2926
rect 21364 2304 21416 2310
rect 21364 2246 21416 2252
rect 21284 2094 21404 2122
rect 21376 800 21404 2094
rect 21836 800 21864 3538
rect 22284 3392 22336 3398
rect 22284 3334 22336 3340
rect 22296 800 22324 3334
rect 22744 2304 22796 2310
rect 22744 2246 22796 2252
rect 22756 800 22784 2246
rect 3514 640 3570 649
rect 3514 575 3570 584
rect 3698 0 3754 800
rect 4158 0 4214 800
rect 4618 0 4674 800
rect 4986 0 5042 800
rect 5446 0 5502 800
rect 5906 0 5962 800
rect 6366 0 6422 800
rect 6826 0 6882 800
rect 7194 0 7250 800
rect 7654 0 7710 800
rect 8114 0 8170 800
rect 8574 0 8630 800
rect 9034 0 9090 800
rect 9402 0 9458 800
rect 9862 0 9918 800
rect 10322 0 10378 800
rect 10782 0 10838 800
rect 11242 0 11298 800
rect 11702 0 11758 800
rect 12070 0 12126 800
rect 12530 0 12586 800
rect 12990 0 13046 800
rect 13450 0 13506 800
rect 13910 0 13966 800
rect 14278 0 14334 800
rect 14738 0 14794 800
rect 15198 0 15254 800
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 16486 0 16542 800
rect 16946 0 17002 800
rect 17406 0 17462 800
rect 17866 0 17922 800
rect 18326 0 18382 800
rect 18694 0 18750 800
rect 19154 0 19210 800
rect 19614 0 19670 800
rect 20074 0 20130 800
rect 20534 0 20590 800
rect 20902 0 20958 800
rect 21362 0 21418 800
rect 21822 0 21878 800
rect 22282 0 22338 800
rect 22742 0 22798 800
<< via2 >>
rect 2870 22616 2926 22672
rect 2778 21256 2834 21312
rect 1950 20712 2006 20768
rect 2042 19780 2098 19816
rect 2042 19760 2044 19780
rect 2044 19760 2096 19780
rect 2096 19760 2098 19780
rect 1950 19388 1952 19408
rect 1952 19388 2004 19408
rect 2004 19388 2006 19408
rect 1950 19352 2006 19388
rect 2778 20304 2834 20360
rect 1950 18808 2006 18864
rect 1858 18400 1914 18456
rect 1950 18028 1952 18048
rect 1952 18028 2004 18048
rect 2004 18028 2006 18048
rect 1950 17992 2006 18028
rect 1950 17448 2006 17504
rect 1950 16496 2006 16552
rect 1674 16088 1730 16144
rect 1858 15544 1914 15600
rect 1490 13232 1546 13288
rect 1950 14220 1952 14240
rect 1952 14220 2004 14240
rect 2004 14220 2006 14240
rect 1950 14184 2006 14220
rect 1490 4820 1546 4856
rect 1490 4800 1492 4820
rect 1492 4800 1544 4820
rect 1544 4800 1546 4820
rect 2778 17040 2834 17096
rect 3698 22208 3754 22264
rect 3146 21664 3202 21720
rect 4421 20698 4477 20700
rect 4501 20698 4557 20700
rect 4581 20698 4637 20700
rect 4661 20698 4717 20700
rect 4421 20646 4447 20698
rect 4447 20646 4477 20698
rect 4501 20646 4511 20698
rect 4511 20646 4557 20698
rect 4581 20646 4627 20698
rect 4627 20646 4637 20698
rect 4661 20646 4691 20698
rect 4691 20646 4717 20698
rect 4421 20644 4477 20646
rect 4501 20644 4557 20646
rect 4581 20644 4637 20646
rect 4661 20644 4717 20646
rect 7886 20154 7942 20156
rect 7966 20154 8022 20156
rect 8046 20154 8102 20156
rect 8126 20154 8182 20156
rect 7886 20102 7912 20154
rect 7912 20102 7942 20154
rect 7966 20102 7976 20154
rect 7976 20102 8022 20154
rect 8046 20102 8092 20154
rect 8092 20102 8102 20154
rect 8126 20102 8156 20154
rect 8156 20102 8182 20154
rect 7886 20100 7942 20102
rect 7966 20100 8022 20102
rect 8046 20100 8102 20102
rect 8126 20100 8182 20102
rect 4421 19610 4477 19612
rect 4501 19610 4557 19612
rect 4581 19610 4637 19612
rect 4661 19610 4717 19612
rect 4421 19558 4447 19610
rect 4447 19558 4477 19610
rect 4501 19558 4511 19610
rect 4511 19558 4557 19610
rect 4581 19558 4627 19610
rect 4627 19558 4637 19610
rect 4661 19558 4691 19610
rect 4691 19558 4717 19610
rect 4421 19556 4477 19558
rect 4501 19556 4557 19558
rect 4581 19556 4637 19558
rect 4661 19556 4717 19558
rect 7886 19066 7942 19068
rect 7966 19066 8022 19068
rect 8046 19066 8102 19068
rect 8126 19066 8182 19068
rect 7886 19014 7912 19066
rect 7912 19014 7942 19066
rect 7966 19014 7976 19066
rect 7976 19014 8022 19066
rect 8046 19014 8092 19066
rect 8092 19014 8102 19066
rect 8126 19014 8156 19066
rect 8156 19014 8182 19066
rect 7886 19012 7942 19014
rect 7966 19012 8022 19014
rect 8046 19012 8102 19014
rect 8126 19012 8182 19014
rect 4421 18522 4477 18524
rect 4501 18522 4557 18524
rect 4581 18522 4637 18524
rect 4661 18522 4717 18524
rect 4421 18470 4447 18522
rect 4447 18470 4477 18522
rect 4501 18470 4511 18522
rect 4511 18470 4557 18522
rect 4581 18470 4627 18522
rect 4627 18470 4637 18522
rect 4661 18470 4691 18522
rect 4691 18470 4717 18522
rect 4421 18468 4477 18470
rect 4501 18468 4557 18470
rect 4581 18468 4637 18470
rect 4661 18468 4717 18470
rect 7886 17978 7942 17980
rect 7966 17978 8022 17980
rect 8046 17978 8102 17980
rect 8126 17978 8182 17980
rect 7886 17926 7912 17978
rect 7912 17926 7942 17978
rect 7966 17926 7976 17978
rect 7976 17926 8022 17978
rect 8046 17926 8092 17978
rect 8092 17926 8102 17978
rect 8126 17926 8156 17978
rect 8156 17926 8182 17978
rect 7886 17924 7942 17926
rect 7966 17924 8022 17926
rect 8046 17924 8102 17926
rect 8126 17924 8182 17926
rect 4421 17434 4477 17436
rect 4501 17434 4557 17436
rect 4581 17434 4637 17436
rect 4661 17434 4717 17436
rect 4421 17382 4447 17434
rect 4447 17382 4477 17434
rect 4501 17382 4511 17434
rect 4511 17382 4557 17434
rect 4581 17382 4627 17434
rect 4627 17382 4637 17434
rect 4661 17382 4691 17434
rect 4691 17382 4717 17434
rect 4421 17380 4477 17382
rect 4501 17380 4557 17382
rect 4581 17380 4637 17382
rect 4661 17380 4717 17382
rect 4421 16346 4477 16348
rect 4501 16346 4557 16348
rect 4581 16346 4637 16348
rect 4661 16346 4717 16348
rect 4421 16294 4447 16346
rect 4447 16294 4477 16346
rect 4501 16294 4511 16346
rect 4511 16294 4557 16346
rect 4581 16294 4627 16346
rect 4627 16294 4637 16346
rect 4661 16294 4691 16346
rect 4691 16294 4717 16346
rect 4421 16292 4477 16294
rect 4501 16292 4557 16294
rect 4581 16292 4637 16294
rect 4661 16292 4717 16294
rect 3238 15136 3294 15192
rect 2962 14592 3018 14648
rect 3514 13776 3570 13832
rect 3422 10104 3478 10160
rect 1582 1944 1638 2000
rect 2870 2624 2926 2680
rect 3514 9968 3570 10024
rect 4421 15258 4477 15260
rect 4501 15258 4557 15260
rect 4581 15258 4637 15260
rect 4661 15258 4717 15260
rect 4421 15206 4447 15258
rect 4447 15206 4477 15258
rect 4501 15206 4511 15258
rect 4511 15206 4557 15258
rect 4581 15206 4627 15258
rect 4627 15206 4637 15258
rect 4661 15206 4691 15258
rect 4691 15206 4717 15258
rect 4421 15204 4477 15206
rect 4501 15204 4557 15206
rect 4581 15204 4637 15206
rect 4661 15204 4717 15206
rect 4421 14170 4477 14172
rect 4501 14170 4557 14172
rect 4581 14170 4637 14172
rect 4661 14170 4717 14172
rect 4421 14118 4447 14170
rect 4447 14118 4477 14170
rect 4501 14118 4511 14170
rect 4511 14118 4557 14170
rect 4581 14118 4627 14170
rect 4627 14118 4637 14170
rect 4661 14118 4691 14170
rect 4691 14118 4717 14170
rect 4421 14116 4477 14118
rect 4501 14116 4557 14118
rect 4581 14116 4637 14118
rect 4661 14116 4717 14118
rect 4421 13082 4477 13084
rect 4501 13082 4557 13084
rect 4581 13082 4637 13084
rect 4661 13082 4717 13084
rect 4421 13030 4447 13082
rect 4447 13030 4477 13082
rect 4501 13030 4511 13082
rect 4511 13030 4557 13082
rect 4581 13030 4627 13082
rect 4627 13030 4637 13082
rect 4661 13030 4691 13082
rect 4691 13030 4717 13082
rect 4421 13028 4477 13030
rect 4501 13028 4557 13030
rect 4581 13028 4637 13030
rect 4661 13028 4717 13030
rect 3974 12316 3976 12336
rect 3976 12316 4028 12336
rect 4028 12316 4030 12336
rect 3974 12280 4030 12316
rect 3974 11872 4030 11928
rect 3974 11328 4030 11384
rect 3882 10956 3884 10976
rect 3884 10956 3936 10976
rect 3936 10956 3938 10976
rect 3882 10920 3938 10956
rect 3974 10376 4030 10432
rect 3790 8608 3846 8664
rect 3790 8336 3846 8392
rect 3514 7384 3570 7440
rect 4421 11994 4477 11996
rect 4501 11994 4557 11996
rect 4581 11994 4637 11996
rect 4661 11994 4717 11996
rect 4421 11942 4447 11994
rect 4447 11942 4477 11994
rect 4501 11942 4511 11994
rect 4511 11942 4557 11994
rect 4581 11942 4627 11994
rect 4627 11942 4637 11994
rect 4661 11942 4691 11994
rect 4691 11942 4717 11994
rect 4421 11940 4477 11942
rect 4501 11940 4557 11942
rect 4581 11940 4637 11942
rect 4661 11940 4717 11942
rect 4066 9424 4122 9480
rect 3974 9016 4030 9072
rect 4066 8064 4122 8120
rect 3974 7656 4030 7712
rect 3514 6160 3570 6216
rect 3238 3440 3294 3496
rect 3422 3476 3424 3496
rect 3424 3476 3476 3496
rect 3476 3476 3478 3496
rect 3422 3440 3478 3476
rect 3054 2488 3110 2544
rect 3422 2624 3478 2680
rect 2962 176 3018 232
rect 4066 6704 4122 6760
rect 3882 5752 3938 5808
rect 4066 5208 4122 5264
rect 4066 4392 4122 4448
rect 4421 10906 4477 10908
rect 4501 10906 4557 10908
rect 4581 10906 4637 10908
rect 4661 10906 4717 10908
rect 4421 10854 4447 10906
rect 4447 10854 4477 10906
rect 4501 10854 4511 10906
rect 4511 10854 4557 10906
rect 4581 10854 4627 10906
rect 4627 10854 4637 10906
rect 4661 10854 4691 10906
rect 4691 10854 4717 10906
rect 4421 10852 4477 10854
rect 4501 10852 4557 10854
rect 4581 10852 4637 10854
rect 4661 10852 4717 10854
rect 4421 9818 4477 9820
rect 4501 9818 4557 9820
rect 4581 9818 4637 9820
rect 4661 9818 4717 9820
rect 4421 9766 4447 9818
rect 4447 9766 4477 9818
rect 4501 9766 4511 9818
rect 4511 9766 4557 9818
rect 4581 9766 4627 9818
rect 4627 9766 4637 9818
rect 4661 9766 4691 9818
rect 4691 9766 4717 9818
rect 4421 9764 4477 9766
rect 4501 9764 4557 9766
rect 4581 9764 4637 9766
rect 4661 9764 4717 9766
rect 4421 8730 4477 8732
rect 4501 8730 4557 8732
rect 4581 8730 4637 8732
rect 4661 8730 4717 8732
rect 4421 8678 4447 8730
rect 4447 8678 4477 8730
rect 4501 8678 4511 8730
rect 4511 8678 4557 8730
rect 4581 8678 4627 8730
rect 4627 8678 4637 8730
rect 4661 8678 4691 8730
rect 4691 8678 4717 8730
rect 4421 8676 4477 8678
rect 4501 8676 4557 8678
rect 4581 8676 4637 8678
rect 4661 8676 4717 8678
rect 4421 7642 4477 7644
rect 4501 7642 4557 7644
rect 4581 7642 4637 7644
rect 4661 7642 4717 7644
rect 4421 7590 4447 7642
rect 4447 7590 4477 7642
rect 4501 7590 4511 7642
rect 4511 7590 4557 7642
rect 4581 7590 4627 7642
rect 4627 7590 4637 7642
rect 4661 7590 4691 7642
rect 4691 7590 4717 7642
rect 4421 7588 4477 7590
rect 4501 7588 4557 7590
rect 4581 7588 4637 7590
rect 4661 7588 4717 7590
rect 4618 7112 4674 7168
rect 4421 6554 4477 6556
rect 4501 6554 4557 6556
rect 4581 6554 4637 6556
rect 4661 6554 4717 6556
rect 4421 6502 4447 6554
rect 4447 6502 4477 6554
rect 4501 6502 4511 6554
rect 4511 6502 4557 6554
rect 4581 6502 4627 6554
rect 4627 6502 4637 6554
rect 4661 6502 4691 6554
rect 4691 6502 4717 6554
rect 4421 6500 4477 6502
rect 4501 6500 4557 6502
rect 4581 6500 4637 6502
rect 4661 6500 4717 6502
rect 4894 6160 4950 6216
rect 4158 2896 4214 2952
rect 3882 1536 3938 1592
rect 3790 992 3846 1048
rect 4421 5466 4477 5468
rect 4501 5466 4557 5468
rect 4581 5466 4637 5468
rect 4661 5466 4717 5468
rect 4421 5414 4447 5466
rect 4447 5414 4477 5466
rect 4501 5414 4511 5466
rect 4511 5414 4557 5466
rect 4581 5414 4627 5466
rect 4627 5414 4637 5466
rect 4661 5414 4691 5466
rect 4691 5414 4717 5466
rect 4421 5412 4477 5414
rect 4501 5412 4557 5414
rect 4581 5412 4637 5414
rect 4661 5412 4717 5414
rect 4421 4378 4477 4380
rect 4501 4378 4557 4380
rect 4581 4378 4637 4380
rect 4661 4378 4717 4380
rect 4421 4326 4447 4378
rect 4447 4326 4477 4378
rect 4501 4326 4511 4378
rect 4511 4326 4557 4378
rect 4581 4326 4627 4378
rect 4627 4326 4637 4378
rect 4661 4326 4691 4378
rect 4691 4326 4717 4378
rect 4421 4324 4477 4326
rect 4501 4324 4557 4326
rect 4581 4324 4637 4326
rect 4661 4324 4717 4326
rect 4421 3290 4477 3292
rect 4501 3290 4557 3292
rect 4581 3290 4637 3292
rect 4661 3290 4717 3292
rect 4421 3238 4447 3290
rect 4447 3238 4477 3290
rect 4501 3238 4511 3290
rect 4511 3238 4557 3290
rect 4581 3238 4627 3290
rect 4627 3238 4637 3290
rect 4661 3238 4691 3290
rect 4691 3238 4717 3290
rect 4421 3236 4477 3238
rect 4501 3236 4557 3238
rect 4581 3236 4637 3238
rect 4661 3236 4717 3238
rect 4421 2202 4477 2204
rect 4501 2202 4557 2204
rect 4581 2202 4637 2204
rect 4661 2202 4717 2204
rect 4421 2150 4447 2202
rect 4447 2150 4477 2202
rect 4501 2150 4511 2202
rect 4511 2150 4557 2202
rect 4581 2150 4627 2202
rect 4627 2150 4637 2202
rect 4661 2150 4691 2202
rect 4691 2150 4717 2202
rect 4421 2148 4477 2150
rect 4501 2148 4557 2150
rect 4581 2148 4637 2150
rect 4661 2148 4717 2150
rect 6274 10104 6330 10160
rect 6918 10124 6974 10160
rect 6918 10104 6920 10124
rect 6920 10104 6972 10124
rect 6972 10104 6974 10124
rect 7010 8336 7066 8392
rect 7886 16890 7942 16892
rect 7966 16890 8022 16892
rect 8046 16890 8102 16892
rect 8126 16890 8182 16892
rect 7886 16838 7912 16890
rect 7912 16838 7942 16890
rect 7966 16838 7976 16890
rect 7976 16838 8022 16890
rect 8046 16838 8092 16890
rect 8092 16838 8102 16890
rect 8126 16838 8156 16890
rect 8156 16838 8182 16890
rect 7886 16836 7942 16838
rect 7966 16836 8022 16838
rect 8046 16836 8102 16838
rect 8126 16836 8182 16838
rect 7886 15802 7942 15804
rect 7966 15802 8022 15804
rect 8046 15802 8102 15804
rect 8126 15802 8182 15804
rect 7886 15750 7912 15802
rect 7912 15750 7942 15802
rect 7966 15750 7976 15802
rect 7976 15750 8022 15802
rect 8046 15750 8092 15802
rect 8092 15750 8102 15802
rect 8126 15750 8156 15802
rect 8156 15750 8182 15802
rect 7886 15748 7942 15750
rect 7966 15748 8022 15750
rect 8046 15748 8102 15750
rect 8126 15748 8182 15750
rect 7886 14714 7942 14716
rect 7966 14714 8022 14716
rect 8046 14714 8102 14716
rect 8126 14714 8182 14716
rect 7886 14662 7912 14714
rect 7912 14662 7942 14714
rect 7966 14662 7976 14714
rect 7976 14662 8022 14714
rect 8046 14662 8092 14714
rect 8092 14662 8102 14714
rect 8126 14662 8156 14714
rect 8156 14662 8182 14714
rect 7886 14660 7942 14662
rect 7966 14660 8022 14662
rect 8046 14660 8102 14662
rect 8126 14660 8182 14662
rect 7886 13626 7942 13628
rect 7966 13626 8022 13628
rect 8046 13626 8102 13628
rect 8126 13626 8182 13628
rect 7886 13574 7912 13626
rect 7912 13574 7942 13626
rect 7966 13574 7976 13626
rect 7976 13574 8022 13626
rect 8046 13574 8092 13626
rect 8092 13574 8102 13626
rect 8126 13574 8156 13626
rect 8156 13574 8182 13626
rect 7886 13572 7942 13574
rect 7966 13572 8022 13574
rect 8046 13572 8102 13574
rect 8126 13572 8182 13574
rect 8298 12824 8354 12880
rect 7886 12538 7942 12540
rect 7966 12538 8022 12540
rect 8046 12538 8102 12540
rect 8126 12538 8182 12540
rect 7886 12486 7912 12538
rect 7912 12486 7942 12538
rect 7966 12486 7976 12538
rect 7976 12486 8022 12538
rect 8046 12486 8092 12538
rect 8092 12486 8102 12538
rect 8126 12486 8156 12538
rect 8156 12486 8182 12538
rect 7886 12484 7942 12486
rect 7966 12484 8022 12486
rect 8046 12484 8102 12486
rect 8126 12484 8182 12486
rect 7886 11450 7942 11452
rect 7966 11450 8022 11452
rect 8046 11450 8102 11452
rect 8126 11450 8182 11452
rect 7886 11398 7912 11450
rect 7912 11398 7942 11450
rect 7966 11398 7976 11450
rect 7976 11398 8022 11450
rect 8046 11398 8092 11450
rect 8092 11398 8102 11450
rect 8126 11398 8156 11450
rect 8156 11398 8182 11450
rect 7886 11396 7942 11398
rect 7966 11396 8022 11398
rect 8046 11396 8102 11398
rect 8126 11396 8182 11398
rect 7886 10362 7942 10364
rect 7966 10362 8022 10364
rect 8046 10362 8102 10364
rect 8126 10362 8182 10364
rect 7886 10310 7912 10362
rect 7912 10310 7942 10362
rect 7966 10310 7976 10362
rect 7976 10310 8022 10362
rect 8046 10310 8092 10362
rect 8092 10310 8102 10362
rect 8126 10310 8156 10362
rect 8156 10310 8182 10362
rect 7886 10308 7942 10310
rect 7966 10308 8022 10310
rect 8046 10308 8102 10310
rect 8126 10308 8182 10310
rect 7886 9274 7942 9276
rect 7966 9274 8022 9276
rect 8046 9274 8102 9276
rect 8126 9274 8182 9276
rect 7886 9222 7912 9274
rect 7912 9222 7942 9274
rect 7966 9222 7976 9274
rect 7976 9222 8022 9274
rect 8046 9222 8092 9274
rect 8092 9222 8102 9274
rect 8126 9222 8156 9274
rect 8156 9222 8182 9274
rect 7886 9220 7942 9222
rect 7966 9220 8022 9222
rect 8046 9220 8102 9222
rect 8126 9220 8182 9222
rect 8022 8336 8078 8392
rect 7886 8186 7942 8188
rect 7966 8186 8022 8188
rect 8046 8186 8102 8188
rect 8126 8186 8182 8188
rect 7886 8134 7912 8186
rect 7912 8134 7942 8186
rect 7966 8134 7976 8186
rect 7976 8134 8022 8186
rect 8046 8134 8092 8186
rect 8092 8134 8102 8186
rect 8126 8134 8156 8186
rect 8156 8134 8182 8186
rect 7886 8132 7942 8134
rect 7966 8132 8022 8134
rect 8046 8132 8102 8134
rect 8126 8132 8182 8134
rect 7886 7098 7942 7100
rect 7966 7098 8022 7100
rect 8046 7098 8102 7100
rect 8126 7098 8182 7100
rect 7886 7046 7912 7098
rect 7912 7046 7942 7098
rect 7966 7046 7976 7098
rect 7976 7046 8022 7098
rect 8046 7046 8092 7098
rect 8092 7046 8102 7098
rect 8126 7046 8156 7098
rect 8156 7046 8182 7098
rect 7886 7044 7942 7046
rect 7966 7044 8022 7046
rect 8046 7044 8102 7046
rect 8126 7044 8182 7046
rect 7886 6010 7942 6012
rect 7966 6010 8022 6012
rect 8046 6010 8102 6012
rect 8126 6010 8182 6012
rect 7886 5958 7912 6010
rect 7912 5958 7942 6010
rect 7966 5958 7976 6010
rect 7976 5958 8022 6010
rect 8046 5958 8092 6010
rect 8092 5958 8102 6010
rect 8126 5958 8156 6010
rect 8156 5958 8182 6010
rect 7886 5956 7942 5958
rect 7966 5956 8022 5958
rect 8046 5956 8102 5958
rect 8126 5956 8182 5958
rect 7886 4922 7942 4924
rect 7966 4922 8022 4924
rect 8046 4922 8102 4924
rect 8126 4922 8182 4924
rect 7886 4870 7912 4922
rect 7912 4870 7942 4922
rect 7966 4870 7976 4922
rect 7976 4870 8022 4922
rect 8046 4870 8092 4922
rect 8092 4870 8102 4922
rect 8126 4870 8156 4922
rect 8156 4870 8182 4922
rect 7886 4868 7942 4870
rect 7966 4868 8022 4870
rect 8046 4868 8102 4870
rect 8126 4868 8182 4870
rect 7886 3834 7942 3836
rect 7966 3834 8022 3836
rect 8046 3834 8102 3836
rect 8126 3834 8182 3836
rect 7886 3782 7912 3834
rect 7912 3782 7942 3834
rect 7966 3782 7976 3834
rect 7976 3782 8022 3834
rect 8046 3782 8092 3834
rect 8092 3782 8102 3834
rect 8126 3782 8156 3834
rect 8156 3782 8182 3834
rect 7886 3780 7942 3782
rect 7966 3780 8022 3782
rect 8046 3780 8102 3782
rect 8126 3780 8182 3782
rect 7886 2746 7942 2748
rect 7966 2746 8022 2748
rect 8046 2746 8102 2748
rect 8126 2746 8182 2748
rect 7886 2694 7912 2746
rect 7912 2694 7942 2746
rect 7966 2694 7976 2746
rect 7976 2694 8022 2746
rect 8046 2694 8092 2746
rect 8092 2694 8102 2746
rect 8126 2694 8156 2746
rect 8156 2694 8182 2746
rect 7886 2692 7942 2694
rect 7966 2692 8022 2694
rect 8046 2692 8102 2694
rect 8126 2692 8182 2694
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11378 20698
rect 11378 20646 11408 20698
rect 11432 20646 11442 20698
rect 11442 20646 11488 20698
rect 11512 20646 11558 20698
rect 11558 20646 11568 20698
rect 11592 20646 11622 20698
rect 11622 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 18282 20698 18338 20700
rect 18362 20698 18418 20700
rect 18442 20698 18498 20700
rect 18522 20698 18578 20700
rect 18282 20646 18308 20698
rect 18308 20646 18338 20698
rect 18362 20646 18372 20698
rect 18372 20646 18418 20698
rect 18442 20646 18488 20698
rect 18488 20646 18498 20698
rect 18522 20646 18552 20698
rect 18552 20646 18578 20698
rect 18282 20644 18338 20646
rect 18362 20644 18418 20646
rect 18442 20644 18498 20646
rect 18522 20644 18578 20646
rect 14817 20154 14873 20156
rect 14897 20154 14953 20156
rect 14977 20154 15033 20156
rect 15057 20154 15113 20156
rect 14817 20102 14843 20154
rect 14843 20102 14873 20154
rect 14897 20102 14907 20154
rect 14907 20102 14953 20154
rect 14977 20102 15023 20154
rect 15023 20102 15033 20154
rect 15057 20102 15087 20154
rect 15087 20102 15113 20154
rect 14817 20100 14873 20102
rect 14897 20100 14953 20102
rect 14977 20100 15033 20102
rect 15057 20100 15113 20102
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11378 19610
rect 11378 19558 11408 19610
rect 11432 19558 11442 19610
rect 11442 19558 11488 19610
rect 11512 19558 11558 19610
rect 11558 19558 11568 19610
rect 11592 19558 11622 19610
rect 11622 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 18282 19610 18338 19612
rect 18362 19610 18418 19612
rect 18442 19610 18498 19612
rect 18522 19610 18578 19612
rect 18282 19558 18308 19610
rect 18308 19558 18338 19610
rect 18362 19558 18372 19610
rect 18372 19558 18418 19610
rect 18442 19558 18488 19610
rect 18488 19558 18498 19610
rect 18522 19558 18552 19610
rect 18552 19558 18578 19610
rect 18282 19556 18338 19558
rect 18362 19556 18418 19558
rect 18442 19556 18498 19558
rect 18522 19556 18578 19558
rect 14817 19066 14873 19068
rect 14897 19066 14953 19068
rect 14977 19066 15033 19068
rect 15057 19066 15113 19068
rect 14817 19014 14843 19066
rect 14843 19014 14873 19066
rect 14897 19014 14907 19066
rect 14907 19014 14953 19066
rect 14977 19014 15023 19066
rect 15023 19014 15033 19066
rect 15057 19014 15087 19066
rect 15087 19014 15113 19066
rect 14817 19012 14873 19014
rect 14897 19012 14953 19014
rect 14977 19012 15033 19014
rect 15057 19012 15113 19014
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11378 18522
rect 11378 18470 11408 18522
rect 11432 18470 11442 18522
rect 11442 18470 11488 18522
rect 11512 18470 11558 18522
rect 11558 18470 11568 18522
rect 11592 18470 11622 18522
rect 11622 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 18282 18522 18338 18524
rect 18362 18522 18418 18524
rect 18442 18522 18498 18524
rect 18522 18522 18578 18524
rect 18282 18470 18308 18522
rect 18308 18470 18338 18522
rect 18362 18470 18372 18522
rect 18372 18470 18418 18522
rect 18442 18470 18488 18522
rect 18488 18470 18498 18522
rect 18522 18470 18552 18522
rect 18552 18470 18578 18522
rect 18282 18468 18338 18470
rect 18362 18468 18418 18470
rect 18442 18468 18498 18470
rect 18522 18468 18578 18470
rect 14817 17978 14873 17980
rect 14897 17978 14953 17980
rect 14977 17978 15033 17980
rect 15057 17978 15113 17980
rect 14817 17926 14843 17978
rect 14843 17926 14873 17978
rect 14897 17926 14907 17978
rect 14907 17926 14953 17978
rect 14977 17926 15023 17978
rect 15023 17926 15033 17978
rect 15057 17926 15087 17978
rect 15087 17926 15113 17978
rect 14817 17924 14873 17926
rect 14897 17924 14953 17926
rect 14977 17924 15033 17926
rect 15057 17924 15113 17926
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11378 17434
rect 11378 17382 11408 17434
rect 11432 17382 11442 17434
rect 11442 17382 11488 17434
rect 11512 17382 11558 17434
rect 11558 17382 11568 17434
rect 11592 17382 11622 17434
rect 11622 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11378 16346
rect 11378 16294 11408 16346
rect 11432 16294 11442 16346
rect 11442 16294 11488 16346
rect 11512 16294 11558 16346
rect 11558 16294 11568 16346
rect 11592 16294 11622 16346
rect 11622 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 18282 17434 18338 17436
rect 18362 17434 18418 17436
rect 18442 17434 18498 17436
rect 18522 17434 18578 17436
rect 18282 17382 18308 17434
rect 18308 17382 18338 17434
rect 18362 17382 18372 17434
rect 18372 17382 18418 17434
rect 18442 17382 18488 17434
rect 18488 17382 18498 17434
rect 18522 17382 18552 17434
rect 18552 17382 18578 17434
rect 18282 17380 18338 17382
rect 18362 17380 18418 17382
rect 18442 17380 18498 17382
rect 18522 17380 18578 17382
rect 19246 17176 19302 17232
rect 14817 16890 14873 16892
rect 14897 16890 14953 16892
rect 14977 16890 15033 16892
rect 15057 16890 15113 16892
rect 14817 16838 14843 16890
rect 14843 16838 14873 16890
rect 14897 16838 14907 16890
rect 14907 16838 14953 16890
rect 14977 16838 15023 16890
rect 15023 16838 15033 16890
rect 15057 16838 15087 16890
rect 15087 16838 15113 16890
rect 14817 16836 14873 16838
rect 14897 16836 14953 16838
rect 14977 16836 15033 16838
rect 15057 16836 15113 16838
rect 8942 6160 8998 6216
rect 9218 7384 9274 7440
rect 10138 5072 10194 5128
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11378 15258
rect 11378 15206 11408 15258
rect 11432 15206 11442 15258
rect 11442 15206 11488 15258
rect 11512 15206 11558 15258
rect 11558 15206 11568 15258
rect 11592 15206 11622 15258
rect 11622 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11378 14170
rect 11378 14118 11408 14170
rect 11432 14118 11442 14170
rect 11442 14118 11488 14170
rect 11512 14118 11558 14170
rect 11558 14118 11568 14170
rect 11592 14118 11622 14170
rect 11622 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11378 13082
rect 11378 13030 11408 13082
rect 11432 13030 11442 13082
rect 11442 13030 11488 13082
rect 11512 13030 11558 13082
rect 11558 13030 11568 13082
rect 11592 13030 11622 13082
rect 11622 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11378 11994
rect 11378 11942 11408 11994
rect 11432 11942 11442 11994
rect 11442 11942 11488 11994
rect 11512 11942 11558 11994
rect 11558 11942 11568 11994
rect 11592 11942 11622 11994
rect 11622 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11378 10906
rect 11378 10854 11408 10906
rect 11432 10854 11442 10906
rect 11442 10854 11488 10906
rect 11512 10854 11558 10906
rect 11558 10854 11568 10906
rect 11592 10854 11622 10906
rect 11622 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11378 9818
rect 11378 9766 11408 9818
rect 11432 9766 11442 9818
rect 11442 9766 11488 9818
rect 11512 9766 11558 9818
rect 11558 9766 11568 9818
rect 11592 9766 11622 9818
rect 11622 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11378 8730
rect 11378 8678 11408 8730
rect 11432 8678 11442 8730
rect 11442 8678 11488 8730
rect 11512 8678 11558 8730
rect 11558 8678 11568 8730
rect 11592 8678 11622 8730
rect 11622 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 18282 16346 18338 16348
rect 18362 16346 18418 16348
rect 18442 16346 18498 16348
rect 18522 16346 18578 16348
rect 18282 16294 18308 16346
rect 18308 16294 18338 16346
rect 18362 16294 18372 16346
rect 18372 16294 18418 16346
rect 18442 16294 18488 16346
rect 18488 16294 18498 16346
rect 18522 16294 18552 16346
rect 18552 16294 18578 16346
rect 18282 16292 18338 16294
rect 18362 16292 18418 16294
rect 18442 16292 18498 16294
rect 18522 16292 18578 16294
rect 14817 15802 14873 15804
rect 14897 15802 14953 15804
rect 14977 15802 15033 15804
rect 15057 15802 15113 15804
rect 14817 15750 14843 15802
rect 14843 15750 14873 15802
rect 14897 15750 14907 15802
rect 14907 15750 14953 15802
rect 14977 15750 15023 15802
rect 15023 15750 15033 15802
rect 15057 15750 15087 15802
rect 15087 15750 15113 15802
rect 14817 15748 14873 15750
rect 14897 15748 14953 15750
rect 14977 15748 15033 15750
rect 15057 15748 15113 15750
rect 18282 15258 18338 15260
rect 18362 15258 18418 15260
rect 18442 15258 18498 15260
rect 18522 15258 18578 15260
rect 18282 15206 18308 15258
rect 18308 15206 18338 15258
rect 18362 15206 18372 15258
rect 18372 15206 18418 15258
rect 18442 15206 18488 15258
rect 18488 15206 18498 15258
rect 18522 15206 18552 15258
rect 18552 15206 18578 15258
rect 18282 15204 18338 15206
rect 18362 15204 18418 15206
rect 18442 15204 18498 15206
rect 18522 15204 18578 15206
rect 14817 14714 14873 14716
rect 14897 14714 14953 14716
rect 14977 14714 15033 14716
rect 15057 14714 15113 14716
rect 14817 14662 14843 14714
rect 14843 14662 14873 14714
rect 14897 14662 14907 14714
rect 14907 14662 14953 14714
rect 14977 14662 15023 14714
rect 15023 14662 15033 14714
rect 15057 14662 15087 14714
rect 15087 14662 15113 14714
rect 14817 14660 14873 14662
rect 14897 14660 14953 14662
rect 14977 14660 15033 14662
rect 15057 14660 15113 14662
rect 18282 14170 18338 14172
rect 18362 14170 18418 14172
rect 18442 14170 18498 14172
rect 18522 14170 18578 14172
rect 18282 14118 18308 14170
rect 18308 14118 18338 14170
rect 18362 14118 18372 14170
rect 18372 14118 18418 14170
rect 18442 14118 18488 14170
rect 18488 14118 18498 14170
rect 18522 14118 18552 14170
rect 18552 14118 18578 14170
rect 18282 14116 18338 14118
rect 18362 14116 18418 14118
rect 18442 14116 18498 14118
rect 18522 14116 18578 14118
rect 14817 13626 14873 13628
rect 14897 13626 14953 13628
rect 14977 13626 15033 13628
rect 15057 13626 15113 13628
rect 14817 13574 14843 13626
rect 14843 13574 14873 13626
rect 14897 13574 14907 13626
rect 14907 13574 14953 13626
rect 14977 13574 15023 13626
rect 15023 13574 15033 13626
rect 15057 13574 15087 13626
rect 15087 13574 15113 13626
rect 14817 13572 14873 13574
rect 14897 13572 14953 13574
rect 14977 13572 15033 13574
rect 15057 13572 15113 13574
rect 18282 13082 18338 13084
rect 18362 13082 18418 13084
rect 18442 13082 18498 13084
rect 18522 13082 18578 13084
rect 18282 13030 18308 13082
rect 18308 13030 18338 13082
rect 18362 13030 18372 13082
rect 18372 13030 18418 13082
rect 18442 13030 18488 13082
rect 18488 13030 18498 13082
rect 18522 13030 18552 13082
rect 18552 13030 18578 13082
rect 18282 13028 18338 13030
rect 18362 13028 18418 13030
rect 18442 13028 18498 13030
rect 18522 13028 18578 13030
rect 14817 12538 14873 12540
rect 14897 12538 14953 12540
rect 14977 12538 15033 12540
rect 15057 12538 15113 12540
rect 14817 12486 14843 12538
rect 14843 12486 14873 12538
rect 14897 12486 14907 12538
rect 14907 12486 14953 12538
rect 14977 12486 15023 12538
rect 15023 12486 15033 12538
rect 15057 12486 15087 12538
rect 15087 12486 15113 12538
rect 14817 12484 14873 12486
rect 14897 12484 14953 12486
rect 14977 12484 15033 12486
rect 15057 12484 15113 12486
rect 18282 11994 18338 11996
rect 18362 11994 18418 11996
rect 18442 11994 18498 11996
rect 18522 11994 18578 11996
rect 18282 11942 18308 11994
rect 18308 11942 18338 11994
rect 18362 11942 18372 11994
rect 18372 11942 18418 11994
rect 18442 11942 18488 11994
rect 18488 11942 18498 11994
rect 18522 11942 18552 11994
rect 18552 11942 18578 11994
rect 18282 11940 18338 11942
rect 18362 11940 18418 11942
rect 18442 11940 18498 11942
rect 18522 11940 18578 11942
rect 14817 11450 14873 11452
rect 14897 11450 14953 11452
rect 14977 11450 15033 11452
rect 15057 11450 15113 11452
rect 14817 11398 14843 11450
rect 14843 11398 14873 11450
rect 14897 11398 14907 11450
rect 14907 11398 14953 11450
rect 14977 11398 15023 11450
rect 15023 11398 15033 11450
rect 15057 11398 15087 11450
rect 15087 11398 15113 11450
rect 14817 11396 14873 11398
rect 14897 11396 14953 11398
rect 14977 11396 15033 11398
rect 15057 11396 15113 11398
rect 18282 10906 18338 10908
rect 18362 10906 18418 10908
rect 18442 10906 18498 10908
rect 18522 10906 18578 10908
rect 18282 10854 18308 10906
rect 18308 10854 18338 10906
rect 18362 10854 18372 10906
rect 18372 10854 18418 10906
rect 18442 10854 18488 10906
rect 18488 10854 18498 10906
rect 18522 10854 18552 10906
rect 18552 10854 18578 10906
rect 18282 10852 18338 10854
rect 18362 10852 18418 10854
rect 18442 10852 18498 10854
rect 18522 10852 18578 10854
rect 14817 10362 14873 10364
rect 14897 10362 14953 10364
rect 14977 10362 15033 10364
rect 15057 10362 15113 10364
rect 14817 10310 14843 10362
rect 14843 10310 14873 10362
rect 14897 10310 14907 10362
rect 14907 10310 14953 10362
rect 14977 10310 15023 10362
rect 15023 10310 15033 10362
rect 15057 10310 15087 10362
rect 15087 10310 15113 10362
rect 14817 10308 14873 10310
rect 14897 10308 14953 10310
rect 14977 10308 15033 10310
rect 15057 10308 15113 10310
rect 18282 9818 18338 9820
rect 18362 9818 18418 9820
rect 18442 9818 18498 9820
rect 18522 9818 18578 9820
rect 18282 9766 18308 9818
rect 18308 9766 18338 9818
rect 18362 9766 18372 9818
rect 18372 9766 18418 9818
rect 18442 9766 18488 9818
rect 18488 9766 18498 9818
rect 18522 9766 18552 9818
rect 18552 9766 18578 9818
rect 18282 9764 18338 9766
rect 18362 9764 18418 9766
rect 18442 9764 18498 9766
rect 18522 9764 18578 9766
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11378 7642
rect 11378 7590 11408 7642
rect 11432 7590 11442 7642
rect 11442 7590 11488 7642
rect 11512 7590 11558 7642
rect 11558 7590 11568 7642
rect 11592 7590 11622 7642
rect 11622 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11378 6554
rect 11378 6502 11408 6554
rect 11432 6502 11442 6554
rect 11442 6502 11488 6554
rect 11512 6502 11558 6554
rect 11558 6502 11568 6554
rect 11592 6502 11622 6554
rect 11622 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11378 5466
rect 11378 5414 11408 5466
rect 11432 5414 11442 5466
rect 11442 5414 11488 5466
rect 11512 5414 11558 5466
rect 11558 5414 11568 5466
rect 11592 5414 11622 5466
rect 11622 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11378 4378
rect 11378 4326 11408 4378
rect 11432 4326 11442 4378
rect 11442 4326 11488 4378
rect 11512 4326 11558 4378
rect 11558 4326 11568 4378
rect 11592 4326 11622 4378
rect 11622 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11378 3290
rect 11378 3238 11408 3290
rect 11432 3238 11442 3290
rect 11442 3238 11488 3290
rect 11512 3238 11558 3290
rect 11558 3238 11568 3290
rect 11592 3238 11622 3290
rect 11622 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11378 2202
rect 11378 2150 11408 2202
rect 11432 2150 11442 2202
rect 11442 2150 11488 2202
rect 11512 2150 11558 2202
rect 11558 2150 11568 2202
rect 11592 2150 11622 2202
rect 11622 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 12622 3440 12678 3496
rect 14817 9274 14873 9276
rect 14897 9274 14953 9276
rect 14977 9274 15033 9276
rect 15057 9274 15113 9276
rect 14817 9222 14843 9274
rect 14843 9222 14873 9274
rect 14897 9222 14907 9274
rect 14907 9222 14953 9274
rect 14977 9222 15023 9274
rect 15023 9222 15033 9274
rect 15057 9222 15087 9274
rect 15087 9222 15113 9274
rect 14817 9220 14873 9222
rect 14897 9220 14953 9222
rect 14977 9220 15033 9222
rect 15057 9220 15113 9222
rect 14817 8186 14873 8188
rect 14897 8186 14953 8188
rect 14977 8186 15033 8188
rect 15057 8186 15113 8188
rect 14817 8134 14843 8186
rect 14843 8134 14873 8186
rect 14897 8134 14907 8186
rect 14907 8134 14953 8186
rect 14977 8134 15023 8186
rect 15023 8134 15033 8186
rect 15057 8134 15087 8186
rect 15087 8134 15113 8186
rect 14817 8132 14873 8134
rect 14897 8132 14953 8134
rect 14977 8132 15033 8134
rect 15057 8132 15113 8134
rect 18282 8730 18338 8732
rect 18362 8730 18418 8732
rect 18442 8730 18498 8732
rect 18522 8730 18578 8732
rect 18282 8678 18308 8730
rect 18308 8678 18338 8730
rect 18362 8678 18372 8730
rect 18372 8678 18418 8730
rect 18442 8678 18488 8730
rect 18488 8678 18498 8730
rect 18522 8678 18552 8730
rect 18552 8678 18578 8730
rect 18282 8676 18338 8678
rect 18362 8676 18418 8678
rect 18442 8676 18498 8678
rect 18522 8676 18578 8678
rect 14817 7098 14873 7100
rect 14897 7098 14953 7100
rect 14977 7098 15033 7100
rect 15057 7098 15113 7100
rect 14817 7046 14843 7098
rect 14843 7046 14873 7098
rect 14897 7046 14907 7098
rect 14907 7046 14953 7098
rect 14977 7046 15023 7098
rect 15023 7046 15033 7098
rect 15057 7046 15087 7098
rect 15087 7046 15113 7098
rect 14817 7044 14873 7046
rect 14897 7044 14953 7046
rect 14977 7044 15033 7046
rect 15057 7044 15113 7046
rect 14817 6010 14873 6012
rect 14897 6010 14953 6012
rect 14977 6010 15033 6012
rect 15057 6010 15113 6012
rect 14817 5958 14843 6010
rect 14843 5958 14873 6010
rect 14897 5958 14907 6010
rect 14907 5958 14953 6010
rect 14977 5958 15023 6010
rect 15023 5958 15033 6010
rect 15057 5958 15087 6010
rect 15087 5958 15113 6010
rect 14817 5956 14873 5958
rect 14897 5956 14953 5958
rect 14977 5956 15033 5958
rect 15057 5956 15113 5958
rect 14817 4922 14873 4924
rect 14897 4922 14953 4924
rect 14977 4922 15033 4924
rect 15057 4922 15113 4924
rect 14817 4870 14843 4922
rect 14843 4870 14873 4922
rect 14897 4870 14907 4922
rect 14907 4870 14953 4922
rect 14977 4870 15023 4922
rect 15023 4870 15033 4922
rect 15057 4870 15087 4922
rect 15087 4870 15113 4922
rect 14817 4868 14873 4870
rect 14897 4868 14953 4870
rect 14977 4868 15033 4870
rect 15057 4868 15113 4870
rect 14817 3834 14873 3836
rect 14897 3834 14953 3836
rect 14977 3834 15033 3836
rect 15057 3834 15113 3836
rect 14817 3782 14843 3834
rect 14843 3782 14873 3834
rect 14897 3782 14907 3834
rect 14907 3782 14953 3834
rect 14977 3782 15023 3834
rect 15023 3782 15033 3834
rect 15057 3782 15087 3834
rect 15087 3782 15113 3834
rect 14817 3780 14873 3782
rect 14897 3780 14953 3782
rect 14977 3780 15033 3782
rect 15057 3780 15113 3782
rect 14817 2746 14873 2748
rect 14897 2746 14953 2748
rect 14977 2746 15033 2748
rect 15057 2746 15113 2748
rect 14817 2694 14843 2746
rect 14843 2694 14873 2746
rect 14897 2694 14907 2746
rect 14907 2694 14953 2746
rect 14977 2694 15023 2746
rect 15023 2694 15033 2746
rect 15057 2694 15087 2746
rect 15087 2694 15113 2746
rect 14817 2692 14873 2694
rect 14897 2692 14953 2694
rect 14977 2692 15033 2694
rect 15057 2692 15113 2694
rect 16118 5108 16120 5128
rect 16120 5108 16172 5128
rect 16172 5108 16174 5128
rect 16118 5072 16174 5108
rect 18282 7642 18338 7644
rect 18362 7642 18418 7644
rect 18442 7642 18498 7644
rect 18522 7642 18578 7644
rect 18282 7590 18308 7642
rect 18308 7590 18338 7642
rect 18362 7590 18372 7642
rect 18372 7590 18418 7642
rect 18442 7590 18488 7642
rect 18488 7590 18498 7642
rect 18522 7590 18552 7642
rect 18552 7590 18578 7642
rect 18282 7588 18338 7590
rect 18362 7588 18418 7590
rect 18442 7588 18498 7590
rect 18522 7588 18578 7590
rect 18282 6554 18338 6556
rect 18362 6554 18418 6556
rect 18442 6554 18498 6556
rect 18522 6554 18578 6556
rect 18282 6502 18308 6554
rect 18308 6502 18338 6554
rect 18362 6502 18372 6554
rect 18372 6502 18418 6554
rect 18442 6502 18488 6554
rect 18488 6502 18498 6554
rect 18522 6502 18552 6554
rect 18552 6502 18578 6554
rect 18282 6500 18338 6502
rect 18362 6500 18418 6502
rect 18442 6500 18498 6502
rect 18522 6500 18578 6502
rect 18282 5466 18338 5468
rect 18362 5466 18418 5468
rect 18442 5466 18498 5468
rect 18522 5466 18578 5468
rect 18282 5414 18308 5466
rect 18308 5414 18338 5466
rect 18362 5414 18372 5466
rect 18372 5414 18418 5466
rect 18442 5414 18488 5466
rect 18488 5414 18498 5466
rect 18522 5414 18552 5466
rect 18552 5414 18578 5466
rect 18282 5412 18338 5414
rect 18362 5412 18418 5414
rect 18442 5412 18498 5414
rect 18522 5412 18578 5414
rect 18282 4378 18338 4380
rect 18362 4378 18418 4380
rect 18442 4378 18498 4380
rect 18522 4378 18578 4380
rect 18282 4326 18308 4378
rect 18308 4326 18338 4378
rect 18362 4326 18372 4378
rect 18372 4326 18418 4378
rect 18442 4326 18488 4378
rect 18488 4326 18498 4378
rect 18522 4326 18552 4378
rect 18552 4326 18578 4378
rect 18282 4324 18338 4326
rect 18362 4324 18418 4326
rect 18442 4324 18498 4326
rect 18522 4324 18578 4326
rect 18282 3290 18338 3292
rect 18362 3290 18418 3292
rect 18442 3290 18498 3292
rect 18522 3290 18578 3292
rect 18282 3238 18308 3290
rect 18308 3238 18338 3290
rect 18362 3238 18372 3290
rect 18372 3238 18418 3290
rect 18442 3238 18488 3290
rect 18488 3238 18498 3290
rect 18522 3238 18552 3290
rect 18552 3238 18578 3290
rect 18282 3236 18338 3238
rect 18362 3236 18418 3238
rect 18442 3236 18498 3238
rect 18522 3236 18578 3238
rect 18282 2202 18338 2204
rect 18362 2202 18418 2204
rect 18442 2202 18498 2204
rect 18522 2202 18578 2204
rect 18282 2150 18308 2202
rect 18308 2150 18338 2202
rect 18362 2150 18372 2202
rect 18372 2150 18418 2202
rect 18442 2150 18488 2202
rect 18488 2150 18498 2202
rect 18522 2150 18552 2202
rect 18552 2150 18578 2202
rect 18282 2148 18338 2150
rect 18362 2148 18418 2150
rect 18442 2148 18498 2150
rect 18522 2148 18578 2150
rect 19706 3596 19762 3632
rect 19706 3576 19708 3596
rect 19708 3576 19760 3596
rect 19760 3576 19762 3596
rect 20626 5752 20682 5808
rect 3514 584 3570 640
<< metal3 >>
rect 0 22674 800 22704
rect 2865 22674 2931 22677
rect 0 22672 2931 22674
rect 0 22616 2870 22672
rect 2926 22616 2931 22672
rect 0 22614 2931 22616
rect 0 22584 800 22614
rect 2865 22611 2931 22614
rect 0 22266 800 22296
rect 3693 22266 3759 22269
rect 0 22264 3759 22266
rect 0 22208 3698 22264
rect 3754 22208 3759 22264
rect 0 22206 3759 22208
rect 0 22176 800 22206
rect 3693 22203 3759 22206
rect 0 21722 800 21752
rect 3141 21722 3207 21725
rect 0 21720 3207 21722
rect 0 21664 3146 21720
rect 3202 21664 3207 21720
rect 0 21662 3207 21664
rect 0 21632 800 21662
rect 3141 21659 3207 21662
rect 0 21314 800 21344
rect 2773 21314 2839 21317
rect 0 21312 2839 21314
rect 0 21256 2778 21312
rect 2834 21256 2839 21312
rect 0 21254 2839 21256
rect 0 21224 800 21254
rect 2773 21251 2839 21254
rect 0 20770 800 20800
rect 1945 20770 2011 20773
rect 0 20768 2011 20770
rect 0 20712 1950 20768
rect 2006 20712 2011 20768
rect 0 20710 2011 20712
rect 0 20680 800 20710
rect 1945 20707 2011 20710
rect 4409 20704 4729 20705
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 20639 4729 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 18270 20704 18590 20705
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 18270 20639 18590 20640
rect 0 20362 800 20392
rect 2773 20362 2839 20365
rect 0 20360 2839 20362
rect 0 20304 2778 20360
rect 2834 20304 2839 20360
rect 0 20302 2839 20304
rect 0 20272 800 20302
rect 2773 20299 2839 20302
rect 7874 20160 8194 20161
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8194 20160
rect 7874 20095 8194 20096
rect 14805 20160 15125 20161
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 20095 15125 20096
rect 0 19818 800 19848
rect 2037 19818 2103 19821
rect 0 19816 2103 19818
rect 0 19760 2042 19816
rect 2098 19760 2103 19816
rect 0 19758 2103 19760
rect 0 19728 800 19758
rect 2037 19755 2103 19758
rect 4409 19616 4729 19617
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 19551 4729 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 18270 19616 18590 19617
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 19551 18590 19552
rect 0 19410 800 19440
rect 1945 19410 2011 19413
rect 0 19408 2011 19410
rect 0 19352 1950 19408
rect 2006 19352 2011 19408
rect 0 19350 2011 19352
rect 0 19320 800 19350
rect 1945 19347 2011 19350
rect 7874 19072 8194 19073
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8194 19072
rect 7874 19007 8194 19008
rect 14805 19072 15125 19073
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 19007 15125 19008
rect 0 18866 800 18896
rect 1945 18866 2011 18869
rect 0 18864 2011 18866
rect 0 18808 1950 18864
rect 2006 18808 2011 18864
rect 0 18806 2011 18808
rect 0 18776 800 18806
rect 1945 18803 2011 18806
rect 4409 18528 4729 18529
rect 0 18458 800 18488
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 18463 4729 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 18270 18528 18590 18529
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 18270 18463 18590 18464
rect 1853 18458 1919 18461
rect 0 18456 1919 18458
rect 0 18400 1858 18456
rect 1914 18400 1919 18456
rect 0 18398 1919 18400
rect 0 18368 800 18398
rect 1853 18395 1919 18398
rect 0 18050 800 18080
rect 1945 18050 2011 18053
rect 0 18048 2011 18050
rect 0 17992 1950 18048
rect 2006 17992 2011 18048
rect 0 17990 2011 17992
rect 0 17960 800 17990
rect 1945 17987 2011 17990
rect 7874 17984 8194 17985
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8194 17984
rect 7874 17919 8194 17920
rect 14805 17984 15125 17985
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 17919 15125 17920
rect 0 17506 800 17536
rect 1945 17506 2011 17509
rect 0 17504 2011 17506
rect 0 17448 1950 17504
rect 2006 17448 2011 17504
rect 0 17446 2011 17448
rect 0 17416 800 17446
rect 1945 17443 2011 17446
rect 4409 17440 4729 17441
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 17375 4729 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 18270 17440 18590 17441
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 18270 17375 18590 17376
rect 19241 17234 19307 17237
rect 22200 17234 23000 17264
rect 19241 17232 23000 17234
rect 19241 17176 19246 17232
rect 19302 17176 23000 17232
rect 19241 17174 23000 17176
rect 19241 17171 19307 17174
rect 22200 17144 23000 17174
rect 0 17098 800 17128
rect 2773 17098 2839 17101
rect 0 17096 2839 17098
rect 0 17040 2778 17096
rect 2834 17040 2839 17096
rect 0 17038 2839 17040
rect 0 17008 800 17038
rect 2773 17035 2839 17038
rect 7874 16896 8194 16897
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8194 16896
rect 7874 16831 8194 16832
rect 14805 16896 15125 16897
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 16831 15125 16832
rect 0 16554 800 16584
rect 1945 16554 2011 16557
rect 0 16552 2011 16554
rect 0 16496 1950 16552
rect 2006 16496 2011 16552
rect 0 16494 2011 16496
rect 0 16464 800 16494
rect 1945 16491 2011 16494
rect 4409 16352 4729 16353
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 16287 4729 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 18270 16352 18590 16353
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 16287 18590 16288
rect 0 16146 800 16176
rect 1669 16146 1735 16149
rect 0 16144 1735 16146
rect 0 16088 1674 16144
rect 1730 16088 1735 16144
rect 0 16086 1735 16088
rect 0 16056 800 16086
rect 1669 16083 1735 16086
rect 7874 15808 8194 15809
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8194 15808
rect 7874 15743 8194 15744
rect 14805 15808 15125 15809
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 15743 15125 15744
rect 0 15602 800 15632
rect 1853 15602 1919 15605
rect 0 15600 1919 15602
rect 0 15544 1858 15600
rect 1914 15544 1919 15600
rect 0 15542 1919 15544
rect 0 15512 800 15542
rect 1853 15539 1919 15542
rect 4409 15264 4729 15265
rect 0 15194 800 15224
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 15199 4729 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 18270 15264 18590 15265
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 18270 15199 18590 15200
rect 3233 15194 3299 15197
rect 0 15192 3299 15194
rect 0 15136 3238 15192
rect 3294 15136 3299 15192
rect 0 15134 3299 15136
rect 0 15104 800 15134
rect 3233 15131 3299 15134
rect 7874 14720 8194 14721
rect 0 14650 800 14680
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8194 14720
rect 7874 14655 8194 14656
rect 14805 14720 15125 14721
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 14655 15125 14656
rect 2957 14650 3023 14653
rect 0 14648 3023 14650
rect 0 14592 2962 14648
rect 3018 14592 3023 14648
rect 0 14590 3023 14592
rect 0 14560 800 14590
rect 2957 14587 3023 14590
rect 0 14242 800 14272
rect 1945 14242 2011 14245
rect 0 14240 2011 14242
rect 0 14184 1950 14240
rect 2006 14184 2011 14240
rect 0 14182 2011 14184
rect 0 14152 800 14182
rect 1945 14179 2011 14182
rect 4409 14176 4729 14177
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 14111 4729 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 18270 14176 18590 14177
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 18270 14111 18590 14112
rect 0 13834 800 13864
rect 3509 13834 3575 13837
rect 0 13832 3575 13834
rect 0 13776 3514 13832
rect 3570 13776 3575 13832
rect 0 13774 3575 13776
rect 0 13744 800 13774
rect 3509 13771 3575 13774
rect 7874 13632 8194 13633
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8194 13632
rect 7874 13567 8194 13568
rect 14805 13632 15125 13633
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 13567 15125 13568
rect 0 13290 800 13320
rect 1485 13290 1551 13293
rect 0 13288 1551 13290
rect 0 13232 1490 13288
rect 1546 13232 1551 13288
rect 0 13230 1551 13232
rect 0 13200 800 13230
rect 1485 13227 1551 13230
rect 4409 13088 4729 13089
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 13023 4729 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 18270 13088 18590 13089
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 13023 18590 13024
rect 0 12882 800 12912
rect 8293 12882 8359 12885
rect 0 12880 8359 12882
rect 0 12824 8298 12880
rect 8354 12824 8359 12880
rect 0 12822 8359 12824
rect 0 12792 800 12822
rect 8293 12819 8359 12822
rect 7874 12544 8194 12545
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8194 12544
rect 7874 12479 8194 12480
rect 14805 12544 15125 12545
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 12479 15125 12480
rect 0 12338 800 12368
rect 3969 12338 4035 12341
rect 0 12336 4035 12338
rect 0 12280 3974 12336
rect 4030 12280 4035 12336
rect 0 12278 4035 12280
rect 0 12248 800 12278
rect 3969 12275 4035 12278
rect 4409 12000 4729 12001
rect 0 11930 800 11960
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 11935 4729 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 18270 12000 18590 12001
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 18270 11935 18590 11936
rect 3969 11930 4035 11933
rect 0 11928 4035 11930
rect 0 11872 3974 11928
rect 4030 11872 4035 11928
rect 0 11870 4035 11872
rect 0 11840 800 11870
rect 3969 11867 4035 11870
rect 7874 11456 8194 11457
rect 0 11386 800 11416
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8194 11456
rect 7874 11391 8194 11392
rect 14805 11456 15125 11457
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 11391 15125 11392
rect 3969 11386 4035 11389
rect 0 11384 4035 11386
rect 0 11328 3974 11384
rect 4030 11328 4035 11384
rect 0 11326 4035 11328
rect 0 11296 800 11326
rect 3969 11323 4035 11326
rect 0 10978 800 11008
rect 3877 10978 3943 10981
rect 0 10976 3943 10978
rect 0 10920 3882 10976
rect 3938 10920 3943 10976
rect 0 10918 3943 10920
rect 0 10888 800 10918
rect 3877 10915 3943 10918
rect 4409 10912 4729 10913
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 10847 4729 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 18270 10912 18590 10913
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 18270 10847 18590 10848
rect 0 10434 800 10464
rect 3969 10434 4035 10437
rect 0 10432 4035 10434
rect 0 10376 3974 10432
rect 4030 10376 4035 10432
rect 0 10374 4035 10376
rect 0 10344 800 10374
rect 3969 10371 4035 10374
rect 7874 10368 8194 10369
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8194 10368
rect 7874 10303 8194 10304
rect 14805 10368 15125 10369
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 10303 15125 10304
rect 3417 10162 3483 10165
rect 6269 10162 6335 10165
rect 6913 10162 6979 10165
rect 3417 10160 6979 10162
rect 3417 10104 3422 10160
rect 3478 10104 6274 10160
rect 6330 10104 6918 10160
rect 6974 10104 6979 10160
rect 3417 10102 6979 10104
rect 3417 10099 3483 10102
rect 6269 10099 6335 10102
rect 6913 10099 6979 10102
rect 0 10026 800 10056
rect 3509 10026 3575 10029
rect 0 10024 3575 10026
rect 0 9968 3514 10024
rect 3570 9968 3575 10024
rect 0 9966 3575 9968
rect 0 9936 800 9966
rect 3509 9963 3575 9966
rect 4409 9824 4729 9825
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 9759 4729 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 18270 9824 18590 9825
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 9759 18590 9760
rect 0 9482 800 9512
rect 4061 9482 4127 9485
rect 0 9480 4127 9482
rect 0 9424 4066 9480
rect 4122 9424 4127 9480
rect 0 9422 4127 9424
rect 0 9392 800 9422
rect 4061 9419 4127 9422
rect 7874 9280 8194 9281
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8194 9280
rect 7874 9215 8194 9216
rect 14805 9280 15125 9281
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 9215 15125 9216
rect 0 9074 800 9104
rect 3969 9074 4035 9077
rect 0 9072 4035 9074
rect 0 9016 3974 9072
rect 4030 9016 4035 9072
rect 0 9014 4035 9016
rect 0 8984 800 9014
rect 3969 9011 4035 9014
rect 4409 8736 4729 8737
rect 0 8666 800 8696
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 8671 4729 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 18270 8736 18590 8737
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 8671 18590 8672
rect 3785 8666 3851 8669
rect 0 8664 3851 8666
rect 0 8608 3790 8664
rect 3846 8608 3851 8664
rect 0 8606 3851 8608
rect 0 8576 800 8606
rect 3785 8603 3851 8606
rect 3785 8394 3851 8397
rect 7005 8394 7071 8397
rect 8017 8394 8083 8397
rect 3785 8392 8083 8394
rect 3785 8336 3790 8392
rect 3846 8336 7010 8392
rect 7066 8336 8022 8392
rect 8078 8336 8083 8392
rect 3785 8334 8083 8336
rect 3785 8331 3851 8334
rect 7005 8331 7071 8334
rect 8017 8331 8083 8334
rect 7874 8192 8194 8193
rect 0 8122 800 8152
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8194 8192
rect 7874 8127 8194 8128
rect 14805 8192 15125 8193
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 8127 15125 8128
rect 4061 8122 4127 8125
rect 0 8120 4127 8122
rect 0 8064 4066 8120
rect 4122 8064 4127 8120
rect 0 8062 4127 8064
rect 0 8032 800 8062
rect 4061 8059 4127 8062
rect 0 7714 800 7744
rect 3969 7714 4035 7717
rect 0 7712 4035 7714
rect 0 7656 3974 7712
rect 4030 7656 4035 7712
rect 0 7654 4035 7656
rect 0 7624 800 7654
rect 3969 7651 4035 7654
rect 4409 7648 4729 7649
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 7583 4729 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 18270 7648 18590 7649
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 18270 7583 18590 7584
rect 3509 7442 3575 7445
rect 9213 7442 9279 7445
rect 3509 7440 9279 7442
rect 3509 7384 3514 7440
rect 3570 7384 9218 7440
rect 9274 7384 9279 7440
rect 3509 7382 9279 7384
rect 3509 7379 3575 7382
rect 9213 7379 9279 7382
rect 0 7170 800 7200
rect 4613 7170 4679 7173
rect 0 7168 4679 7170
rect 0 7112 4618 7168
rect 4674 7112 4679 7168
rect 0 7110 4679 7112
rect 0 7080 800 7110
rect 4613 7107 4679 7110
rect 7874 7104 8194 7105
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8194 7104
rect 7874 7039 8194 7040
rect 14805 7104 15125 7105
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 7039 15125 7040
rect 0 6762 800 6792
rect 4061 6762 4127 6765
rect 0 6760 4127 6762
rect 0 6704 4066 6760
rect 4122 6704 4127 6760
rect 0 6702 4127 6704
rect 0 6672 800 6702
rect 4061 6699 4127 6702
rect 4409 6560 4729 6561
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 6495 4729 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 18270 6560 18590 6561
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 18270 6495 18590 6496
rect 0 6218 800 6248
rect 3509 6218 3575 6221
rect 0 6216 3575 6218
rect 0 6160 3514 6216
rect 3570 6160 3575 6216
rect 0 6158 3575 6160
rect 0 6128 800 6158
rect 3509 6155 3575 6158
rect 4889 6218 4955 6221
rect 8937 6218 9003 6221
rect 4889 6216 9003 6218
rect 4889 6160 4894 6216
rect 4950 6160 8942 6216
rect 8998 6160 9003 6216
rect 4889 6158 9003 6160
rect 4889 6155 4955 6158
rect 8937 6155 9003 6158
rect 7874 6016 8194 6017
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8194 6016
rect 7874 5951 8194 5952
rect 14805 6016 15125 6017
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 5951 15125 5952
rect 0 5810 800 5840
rect 3877 5810 3943 5813
rect 0 5808 3943 5810
rect 0 5752 3882 5808
rect 3938 5752 3943 5808
rect 0 5750 3943 5752
rect 0 5720 800 5750
rect 3877 5747 3943 5750
rect 20621 5810 20687 5813
rect 22200 5810 23000 5840
rect 20621 5808 23000 5810
rect 20621 5752 20626 5808
rect 20682 5752 23000 5808
rect 20621 5750 23000 5752
rect 20621 5747 20687 5750
rect 22200 5720 23000 5750
rect 4409 5472 4729 5473
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 5407 4729 5408
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 18270 5472 18590 5473
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 5407 18590 5408
rect 0 5266 800 5296
rect 4061 5266 4127 5269
rect 0 5264 4127 5266
rect 0 5208 4066 5264
rect 4122 5208 4127 5264
rect 0 5206 4127 5208
rect 0 5176 800 5206
rect 4061 5203 4127 5206
rect 10133 5130 10199 5133
rect 16113 5130 16179 5133
rect 10133 5128 16179 5130
rect 10133 5072 10138 5128
rect 10194 5072 16118 5128
rect 16174 5072 16179 5128
rect 10133 5070 16179 5072
rect 10133 5067 10199 5070
rect 16113 5067 16179 5070
rect 7874 4928 8194 4929
rect 0 4858 800 4888
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8194 4928
rect 7874 4863 8194 4864
rect 14805 4928 15125 4929
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 4863 15125 4864
rect 1485 4858 1551 4861
rect 0 4856 1551 4858
rect 0 4800 1490 4856
rect 1546 4800 1551 4856
rect 0 4798 1551 4800
rect 0 4768 800 4798
rect 1485 4795 1551 4798
rect 0 4450 800 4480
rect 4061 4450 4127 4453
rect 0 4448 4127 4450
rect 0 4392 4066 4448
rect 4122 4392 4127 4448
rect 0 4390 4127 4392
rect 0 4360 800 4390
rect 4061 4387 4127 4390
rect 4409 4384 4729 4385
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 4319 4729 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 18270 4384 18590 4385
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 18270 4319 18590 4320
rect 0 3906 800 3936
rect 0 3846 4906 3906
rect 0 3816 800 3846
rect 4846 3634 4906 3846
rect 7874 3840 8194 3841
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8194 3840
rect 7874 3775 8194 3776
rect 14805 3840 15125 3841
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 3775 15125 3776
rect 19701 3634 19767 3637
rect 4846 3632 19767 3634
rect 4846 3576 19706 3632
rect 19762 3576 19767 3632
rect 4846 3574 19767 3576
rect 19701 3571 19767 3574
rect 0 3498 800 3528
rect 3233 3498 3299 3501
rect 0 3496 3299 3498
rect 0 3440 3238 3496
rect 3294 3440 3299 3496
rect 0 3438 3299 3440
rect 0 3408 800 3438
rect 3233 3435 3299 3438
rect 3417 3498 3483 3501
rect 12617 3498 12683 3501
rect 3417 3496 12683 3498
rect 3417 3440 3422 3496
rect 3478 3440 12622 3496
rect 12678 3440 12683 3496
rect 3417 3438 12683 3440
rect 3417 3435 3483 3438
rect 12617 3435 12683 3438
rect 4409 3296 4729 3297
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 3231 4729 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 18270 3296 18590 3297
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 18270 3231 18590 3232
rect 0 2954 800 2984
rect 4153 2954 4219 2957
rect 0 2952 4219 2954
rect 0 2896 4158 2952
rect 4214 2896 4219 2952
rect 0 2894 4219 2896
rect 0 2864 800 2894
rect 4153 2891 4219 2894
rect 7874 2752 8194 2753
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8194 2752
rect 7874 2687 8194 2688
rect 14805 2752 15125 2753
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2687 15125 2688
rect 2865 2682 2931 2685
rect 3417 2682 3483 2685
rect 2865 2680 3483 2682
rect 2865 2624 2870 2680
rect 2926 2624 3422 2680
rect 3478 2624 3483 2680
rect 2865 2622 3483 2624
rect 2865 2619 2931 2622
rect 3417 2619 3483 2622
rect 0 2546 800 2576
rect 3049 2546 3115 2549
rect 0 2544 3115 2546
rect 0 2488 3054 2544
rect 3110 2488 3115 2544
rect 0 2486 3115 2488
rect 0 2456 800 2486
rect 3049 2483 3115 2486
rect 4409 2208 4729 2209
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2143 4729 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 18270 2208 18590 2209
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2143 18590 2144
rect 0 2002 800 2032
rect 1577 2002 1643 2005
rect 0 2000 1643 2002
rect 0 1944 1582 2000
rect 1638 1944 1643 2000
rect 0 1942 1643 1944
rect 0 1912 800 1942
rect 1577 1939 1643 1942
rect 0 1594 800 1624
rect 3877 1594 3943 1597
rect 0 1592 3943 1594
rect 0 1536 3882 1592
rect 3938 1536 3943 1592
rect 0 1534 3943 1536
rect 0 1504 800 1534
rect 3877 1531 3943 1534
rect 0 1050 800 1080
rect 3785 1050 3851 1053
rect 0 1048 3851 1050
rect 0 992 3790 1048
rect 3846 992 3851 1048
rect 0 990 3851 992
rect 0 960 800 990
rect 3785 987 3851 990
rect 0 642 800 672
rect 3509 642 3575 645
rect 0 640 3575 642
rect 0 584 3514 640
rect 3570 584 3575 640
rect 0 582 3575 584
rect 0 552 800 582
rect 3509 579 3575 582
rect 0 234 800 264
rect 2957 234 3023 237
rect 0 232 3023 234
rect 0 176 2962 232
rect 3018 176 3023 232
rect 0 174 3023 176
rect 0 144 800 174
rect 2957 171 3023 174
<< via3 >>
rect 4417 20700 4481 20704
rect 4417 20644 4421 20700
rect 4421 20644 4477 20700
rect 4477 20644 4481 20700
rect 4417 20640 4481 20644
rect 4497 20700 4561 20704
rect 4497 20644 4501 20700
rect 4501 20644 4557 20700
rect 4557 20644 4561 20700
rect 4497 20640 4561 20644
rect 4577 20700 4641 20704
rect 4577 20644 4581 20700
rect 4581 20644 4637 20700
rect 4637 20644 4641 20700
rect 4577 20640 4641 20644
rect 4657 20700 4721 20704
rect 4657 20644 4661 20700
rect 4661 20644 4717 20700
rect 4717 20644 4721 20700
rect 4657 20640 4721 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 18278 20700 18342 20704
rect 18278 20644 18282 20700
rect 18282 20644 18338 20700
rect 18338 20644 18342 20700
rect 18278 20640 18342 20644
rect 18358 20700 18422 20704
rect 18358 20644 18362 20700
rect 18362 20644 18418 20700
rect 18418 20644 18422 20700
rect 18358 20640 18422 20644
rect 18438 20700 18502 20704
rect 18438 20644 18442 20700
rect 18442 20644 18498 20700
rect 18498 20644 18502 20700
rect 18438 20640 18502 20644
rect 18518 20700 18582 20704
rect 18518 20644 18522 20700
rect 18522 20644 18578 20700
rect 18578 20644 18582 20700
rect 18518 20640 18582 20644
rect 7882 20156 7946 20160
rect 7882 20100 7886 20156
rect 7886 20100 7942 20156
rect 7942 20100 7946 20156
rect 7882 20096 7946 20100
rect 7962 20156 8026 20160
rect 7962 20100 7966 20156
rect 7966 20100 8022 20156
rect 8022 20100 8026 20156
rect 7962 20096 8026 20100
rect 8042 20156 8106 20160
rect 8042 20100 8046 20156
rect 8046 20100 8102 20156
rect 8102 20100 8106 20156
rect 8042 20096 8106 20100
rect 8122 20156 8186 20160
rect 8122 20100 8126 20156
rect 8126 20100 8182 20156
rect 8182 20100 8186 20156
rect 8122 20096 8186 20100
rect 14813 20156 14877 20160
rect 14813 20100 14817 20156
rect 14817 20100 14873 20156
rect 14873 20100 14877 20156
rect 14813 20096 14877 20100
rect 14893 20156 14957 20160
rect 14893 20100 14897 20156
rect 14897 20100 14953 20156
rect 14953 20100 14957 20156
rect 14893 20096 14957 20100
rect 14973 20156 15037 20160
rect 14973 20100 14977 20156
rect 14977 20100 15033 20156
rect 15033 20100 15037 20156
rect 14973 20096 15037 20100
rect 15053 20156 15117 20160
rect 15053 20100 15057 20156
rect 15057 20100 15113 20156
rect 15113 20100 15117 20156
rect 15053 20096 15117 20100
rect 4417 19612 4481 19616
rect 4417 19556 4421 19612
rect 4421 19556 4477 19612
rect 4477 19556 4481 19612
rect 4417 19552 4481 19556
rect 4497 19612 4561 19616
rect 4497 19556 4501 19612
rect 4501 19556 4557 19612
rect 4557 19556 4561 19612
rect 4497 19552 4561 19556
rect 4577 19612 4641 19616
rect 4577 19556 4581 19612
rect 4581 19556 4637 19612
rect 4637 19556 4641 19612
rect 4577 19552 4641 19556
rect 4657 19612 4721 19616
rect 4657 19556 4661 19612
rect 4661 19556 4717 19612
rect 4717 19556 4721 19612
rect 4657 19552 4721 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 18278 19612 18342 19616
rect 18278 19556 18282 19612
rect 18282 19556 18338 19612
rect 18338 19556 18342 19612
rect 18278 19552 18342 19556
rect 18358 19612 18422 19616
rect 18358 19556 18362 19612
rect 18362 19556 18418 19612
rect 18418 19556 18422 19612
rect 18358 19552 18422 19556
rect 18438 19612 18502 19616
rect 18438 19556 18442 19612
rect 18442 19556 18498 19612
rect 18498 19556 18502 19612
rect 18438 19552 18502 19556
rect 18518 19612 18582 19616
rect 18518 19556 18522 19612
rect 18522 19556 18578 19612
rect 18578 19556 18582 19612
rect 18518 19552 18582 19556
rect 7882 19068 7946 19072
rect 7882 19012 7886 19068
rect 7886 19012 7942 19068
rect 7942 19012 7946 19068
rect 7882 19008 7946 19012
rect 7962 19068 8026 19072
rect 7962 19012 7966 19068
rect 7966 19012 8022 19068
rect 8022 19012 8026 19068
rect 7962 19008 8026 19012
rect 8042 19068 8106 19072
rect 8042 19012 8046 19068
rect 8046 19012 8102 19068
rect 8102 19012 8106 19068
rect 8042 19008 8106 19012
rect 8122 19068 8186 19072
rect 8122 19012 8126 19068
rect 8126 19012 8182 19068
rect 8182 19012 8186 19068
rect 8122 19008 8186 19012
rect 14813 19068 14877 19072
rect 14813 19012 14817 19068
rect 14817 19012 14873 19068
rect 14873 19012 14877 19068
rect 14813 19008 14877 19012
rect 14893 19068 14957 19072
rect 14893 19012 14897 19068
rect 14897 19012 14953 19068
rect 14953 19012 14957 19068
rect 14893 19008 14957 19012
rect 14973 19068 15037 19072
rect 14973 19012 14977 19068
rect 14977 19012 15033 19068
rect 15033 19012 15037 19068
rect 14973 19008 15037 19012
rect 15053 19068 15117 19072
rect 15053 19012 15057 19068
rect 15057 19012 15113 19068
rect 15113 19012 15117 19068
rect 15053 19008 15117 19012
rect 4417 18524 4481 18528
rect 4417 18468 4421 18524
rect 4421 18468 4477 18524
rect 4477 18468 4481 18524
rect 4417 18464 4481 18468
rect 4497 18524 4561 18528
rect 4497 18468 4501 18524
rect 4501 18468 4557 18524
rect 4557 18468 4561 18524
rect 4497 18464 4561 18468
rect 4577 18524 4641 18528
rect 4577 18468 4581 18524
rect 4581 18468 4637 18524
rect 4637 18468 4641 18524
rect 4577 18464 4641 18468
rect 4657 18524 4721 18528
rect 4657 18468 4661 18524
rect 4661 18468 4717 18524
rect 4717 18468 4721 18524
rect 4657 18464 4721 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 18278 18524 18342 18528
rect 18278 18468 18282 18524
rect 18282 18468 18338 18524
rect 18338 18468 18342 18524
rect 18278 18464 18342 18468
rect 18358 18524 18422 18528
rect 18358 18468 18362 18524
rect 18362 18468 18418 18524
rect 18418 18468 18422 18524
rect 18358 18464 18422 18468
rect 18438 18524 18502 18528
rect 18438 18468 18442 18524
rect 18442 18468 18498 18524
rect 18498 18468 18502 18524
rect 18438 18464 18502 18468
rect 18518 18524 18582 18528
rect 18518 18468 18522 18524
rect 18522 18468 18578 18524
rect 18578 18468 18582 18524
rect 18518 18464 18582 18468
rect 7882 17980 7946 17984
rect 7882 17924 7886 17980
rect 7886 17924 7942 17980
rect 7942 17924 7946 17980
rect 7882 17920 7946 17924
rect 7962 17980 8026 17984
rect 7962 17924 7966 17980
rect 7966 17924 8022 17980
rect 8022 17924 8026 17980
rect 7962 17920 8026 17924
rect 8042 17980 8106 17984
rect 8042 17924 8046 17980
rect 8046 17924 8102 17980
rect 8102 17924 8106 17980
rect 8042 17920 8106 17924
rect 8122 17980 8186 17984
rect 8122 17924 8126 17980
rect 8126 17924 8182 17980
rect 8182 17924 8186 17980
rect 8122 17920 8186 17924
rect 14813 17980 14877 17984
rect 14813 17924 14817 17980
rect 14817 17924 14873 17980
rect 14873 17924 14877 17980
rect 14813 17920 14877 17924
rect 14893 17980 14957 17984
rect 14893 17924 14897 17980
rect 14897 17924 14953 17980
rect 14953 17924 14957 17980
rect 14893 17920 14957 17924
rect 14973 17980 15037 17984
rect 14973 17924 14977 17980
rect 14977 17924 15033 17980
rect 15033 17924 15037 17980
rect 14973 17920 15037 17924
rect 15053 17980 15117 17984
rect 15053 17924 15057 17980
rect 15057 17924 15113 17980
rect 15113 17924 15117 17980
rect 15053 17920 15117 17924
rect 4417 17436 4481 17440
rect 4417 17380 4421 17436
rect 4421 17380 4477 17436
rect 4477 17380 4481 17436
rect 4417 17376 4481 17380
rect 4497 17436 4561 17440
rect 4497 17380 4501 17436
rect 4501 17380 4557 17436
rect 4557 17380 4561 17436
rect 4497 17376 4561 17380
rect 4577 17436 4641 17440
rect 4577 17380 4581 17436
rect 4581 17380 4637 17436
rect 4637 17380 4641 17436
rect 4577 17376 4641 17380
rect 4657 17436 4721 17440
rect 4657 17380 4661 17436
rect 4661 17380 4717 17436
rect 4717 17380 4721 17436
rect 4657 17376 4721 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 18278 17436 18342 17440
rect 18278 17380 18282 17436
rect 18282 17380 18338 17436
rect 18338 17380 18342 17436
rect 18278 17376 18342 17380
rect 18358 17436 18422 17440
rect 18358 17380 18362 17436
rect 18362 17380 18418 17436
rect 18418 17380 18422 17436
rect 18358 17376 18422 17380
rect 18438 17436 18502 17440
rect 18438 17380 18442 17436
rect 18442 17380 18498 17436
rect 18498 17380 18502 17436
rect 18438 17376 18502 17380
rect 18518 17436 18582 17440
rect 18518 17380 18522 17436
rect 18522 17380 18578 17436
rect 18578 17380 18582 17436
rect 18518 17376 18582 17380
rect 7882 16892 7946 16896
rect 7882 16836 7886 16892
rect 7886 16836 7942 16892
rect 7942 16836 7946 16892
rect 7882 16832 7946 16836
rect 7962 16892 8026 16896
rect 7962 16836 7966 16892
rect 7966 16836 8022 16892
rect 8022 16836 8026 16892
rect 7962 16832 8026 16836
rect 8042 16892 8106 16896
rect 8042 16836 8046 16892
rect 8046 16836 8102 16892
rect 8102 16836 8106 16892
rect 8042 16832 8106 16836
rect 8122 16892 8186 16896
rect 8122 16836 8126 16892
rect 8126 16836 8182 16892
rect 8182 16836 8186 16892
rect 8122 16832 8186 16836
rect 14813 16892 14877 16896
rect 14813 16836 14817 16892
rect 14817 16836 14873 16892
rect 14873 16836 14877 16892
rect 14813 16832 14877 16836
rect 14893 16892 14957 16896
rect 14893 16836 14897 16892
rect 14897 16836 14953 16892
rect 14953 16836 14957 16892
rect 14893 16832 14957 16836
rect 14973 16892 15037 16896
rect 14973 16836 14977 16892
rect 14977 16836 15033 16892
rect 15033 16836 15037 16892
rect 14973 16832 15037 16836
rect 15053 16892 15117 16896
rect 15053 16836 15057 16892
rect 15057 16836 15113 16892
rect 15113 16836 15117 16892
rect 15053 16832 15117 16836
rect 4417 16348 4481 16352
rect 4417 16292 4421 16348
rect 4421 16292 4477 16348
rect 4477 16292 4481 16348
rect 4417 16288 4481 16292
rect 4497 16348 4561 16352
rect 4497 16292 4501 16348
rect 4501 16292 4557 16348
rect 4557 16292 4561 16348
rect 4497 16288 4561 16292
rect 4577 16348 4641 16352
rect 4577 16292 4581 16348
rect 4581 16292 4637 16348
rect 4637 16292 4641 16348
rect 4577 16288 4641 16292
rect 4657 16348 4721 16352
rect 4657 16292 4661 16348
rect 4661 16292 4717 16348
rect 4717 16292 4721 16348
rect 4657 16288 4721 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 18278 16348 18342 16352
rect 18278 16292 18282 16348
rect 18282 16292 18338 16348
rect 18338 16292 18342 16348
rect 18278 16288 18342 16292
rect 18358 16348 18422 16352
rect 18358 16292 18362 16348
rect 18362 16292 18418 16348
rect 18418 16292 18422 16348
rect 18358 16288 18422 16292
rect 18438 16348 18502 16352
rect 18438 16292 18442 16348
rect 18442 16292 18498 16348
rect 18498 16292 18502 16348
rect 18438 16288 18502 16292
rect 18518 16348 18582 16352
rect 18518 16292 18522 16348
rect 18522 16292 18578 16348
rect 18578 16292 18582 16348
rect 18518 16288 18582 16292
rect 7882 15804 7946 15808
rect 7882 15748 7886 15804
rect 7886 15748 7942 15804
rect 7942 15748 7946 15804
rect 7882 15744 7946 15748
rect 7962 15804 8026 15808
rect 7962 15748 7966 15804
rect 7966 15748 8022 15804
rect 8022 15748 8026 15804
rect 7962 15744 8026 15748
rect 8042 15804 8106 15808
rect 8042 15748 8046 15804
rect 8046 15748 8102 15804
rect 8102 15748 8106 15804
rect 8042 15744 8106 15748
rect 8122 15804 8186 15808
rect 8122 15748 8126 15804
rect 8126 15748 8182 15804
rect 8182 15748 8186 15804
rect 8122 15744 8186 15748
rect 14813 15804 14877 15808
rect 14813 15748 14817 15804
rect 14817 15748 14873 15804
rect 14873 15748 14877 15804
rect 14813 15744 14877 15748
rect 14893 15804 14957 15808
rect 14893 15748 14897 15804
rect 14897 15748 14953 15804
rect 14953 15748 14957 15804
rect 14893 15744 14957 15748
rect 14973 15804 15037 15808
rect 14973 15748 14977 15804
rect 14977 15748 15033 15804
rect 15033 15748 15037 15804
rect 14973 15744 15037 15748
rect 15053 15804 15117 15808
rect 15053 15748 15057 15804
rect 15057 15748 15113 15804
rect 15113 15748 15117 15804
rect 15053 15744 15117 15748
rect 4417 15260 4481 15264
rect 4417 15204 4421 15260
rect 4421 15204 4477 15260
rect 4477 15204 4481 15260
rect 4417 15200 4481 15204
rect 4497 15260 4561 15264
rect 4497 15204 4501 15260
rect 4501 15204 4557 15260
rect 4557 15204 4561 15260
rect 4497 15200 4561 15204
rect 4577 15260 4641 15264
rect 4577 15204 4581 15260
rect 4581 15204 4637 15260
rect 4637 15204 4641 15260
rect 4577 15200 4641 15204
rect 4657 15260 4721 15264
rect 4657 15204 4661 15260
rect 4661 15204 4717 15260
rect 4717 15204 4721 15260
rect 4657 15200 4721 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 18278 15260 18342 15264
rect 18278 15204 18282 15260
rect 18282 15204 18338 15260
rect 18338 15204 18342 15260
rect 18278 15200 18342 15204
rect 18358 15260 18422 15264
rect 18358 15204 18362 15260
rect 18362 15204 18418 15260
rect 18418 15204 18422 15260
rect 18358 15200 18422 15204
rect 18438 15260 18502 15264
rect 18438 15204 18442 15260
rect 18442 15204 18498 15260
rect 18498 15204 18502 15260
rect 18438 15200 18502 15204
rect 18518 15260 18582 15264
rect 18518 15204 18522 15260
rect 18522 15204 18578 15260
rect 18578 15204 18582 15260
rect 18518 15200 18582 15204
rect 7882 14716 7946 14720
rect 7882 14660 7886 14716
rect 7886 14660 7942 14716
rect 7942 14660 7946 14716
rect 7882 14656 7946 14660
rect 7962 14716 8026 14720
rect 7962 14660 7966 14716
rect 7966 14660 8022 14716
rect 8022 14660 8026 14716
rect 7962 14656 8026 14660
rect 8042 14716 8106 14720
rect 8042 14660 8046 14716
rect 8046 14660 8102 14716
rect 8102 14660 8106 14716
rect 8042 14656 8106 14660
rect 8122 14716 8186 14720
rect 8122 14660 8126 14716
rect 8126 14660 8182 14716
rect 8182 14660 8186 14716
rect 8122 14656 8186 14660
rect 14813 14716 14877 14720
rect 14813 14660 14817 14716
rect 14817 14660 14873 14716
rect 14873 14660 14877 14716
rect 14813 14656 14877 14660
rect 14893 14716 14957 14720
rect 14893 14660 14897 14716
rect 14897 14660 14953 14716
rect 14953 14660 14957 14716
rect 14893 14656 14957 14660
rect 14973 14716 15037 14720
rect 14973 14660 14977 14716
rect 14977 14660 15033 14716
rect 15033 14660 15037 14716
rect 14973 14656 15037 14660
rect 15053 14716 15117 14720
rect 15053 14660 15057 14716
rect 15057 14660 15113 14716
rect 15113 14660 15117 14716
rect 15053 14656 15117 14660
rect 4417 14172 4481 14176
rect 4417 14116 4421 14172
rect 4421 14116 4477 14172
rect 4477 14116 4481 14172
rect 4417 14112 4481 14116
rect 4497 14172 4561 14176
rect 4497 14116 4501 14172
rect 4501 14116 4557 14172
rect 4557 14116 4561 14172
rect 4497 14112 4561 14116
rect 4577 14172 4641 14176
rect 4577 14116 4581 14172
rect 4581 14116 4637 14172
rect 4637 14116 4641 14172
rect 4577 14112 4641 14116
rect 4657 14172 4721 14176
rect 4657 14116 4661 14172
rect 4661 14116 4717 14172
rect 4717 14116 4721 14172
rect 4657 14112 4721 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 18278 14172 18342 14176
rect 18278 14116 18282 14172
rect 18282 14116 18338 14172
rect 18338 14116 18342 14172
rect 18278 14112 18342 14116
rect 18358 14172 18422 14176
rect 18358 14116 18362 14172
rect 18362 14116 18418 14172
rect 18418 14116 18422 14172
rect 18358 14112 18422 14116
rect 18438 14172 18502 14176
rect 18438 14116 18442 14172
rect 18442 14116 18498 14172
rect 18498 14116 18502 14172
rect 18438 14112 18502 14116
rect 18518 14172 18582 14176
rect 18518 14116 18522 14172
rect 18522 14116 18578 14172
rect 18578 14116 18582 14172
rect 18518 14112 18582 14116
rect 7882 13628 7946 13632
rect 7882 13572 7886 13628
rect 7886 13572 7942 13628
rect 7942 13572 7946 13628
rect 7882 13568 7946 13572
rect 7962 13628 8026 13632
rect 7962 13572 7966 13628
rect 7966 13572 8022 13628
rect 8022 13572 8026 13628
rect 7962 13568 8026 13572
rect 8042 13628 8106 13632
rect 8042 13572 8046 13628
rect 8046 13572 8102 13628
rect 8102 13572 8106 13628
rect 8042 13568 8106 13572
rect 8122 13628 8186 13632
rect 8122 13572 8126 13628
rect 8126 13572 8182 13628
rect 8182 13572 8186 13628
rect 8122 13568 8186 13572
rect 14813 13628 14877 13632
rect 14813 13572 14817 13628
rect 14817 13572 14873 13628
rect 14873 13572 14877 13628
rect 14813 13568 14877 13572
rect 14893 13628 14957 13632
rect 14893 13572 14897 13628
rect 14897 13572 14953 13628
rect 14953 13572 14957 13628
rect 14893 13568 14957 13572
rect 14973 13628 15037 13632
rect 14973 13572 14977 13628
rect 14977 13572 15033 13628
rect 15033 13572 15037 13628
rect 14973 13568 15037 13572
rect 15053 13628 15117 13632
rect 15053 13572 15057 13628
rect 15057 13572 15113 13628
rect 15113 13572 15117 13628
rect 15053 13568 15117 13572
rect 4417 13084 4481 13088
rect 4417 13028 4421 13084
rect 4421 13028 4477 13084
rect 4477 13028 4481 13084
rect 4417 13024 4481 13028
rect 4497 13084 4561 13088
rect 4497 13028 4501 13084
rect 4501 13028 4557 13084
rect 4557 13028 4561 13084
rect 4497 13024 4561 13028
rect 4577 13084 4641 13088
rect 4577 13028 4581 13084
rect 4581 13028 4637 13084
rect 4637 13028 4641 13084
rect 4577 13024 4641 13028
rect 4657 13084 4721 13088
rect 4657 13028 4661 13084
rect 4661 13028 4717 13084
rect 4717 13028 4721 13084
rect 4657 13024 4721 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 18278 13084 18342 13088
rect 18278 13028 18282 13084
rect 18282 13028 18338 13084
rect 18338 13028 18342 13084
rect 18278 13024 18342 13028
rect 18358 13084 18422 13088
rect 18358 13028 18362 13084
rect 18362 13028 18418 13084
rect 18418 13028 18422 13084
rect 18358 13024 18422 13028
rect 18438 13084 18502 13088
rect 18438 13028 18442 13084
rect 18442 13028 18498 13084
rect 18498 13028 18502 13084
rect 18438 13024 18502 13028
rect 18518 13084 18582 13088
rect 18518 13028 18522 13084
rect 18522 13028 18578 13084
rect 18578 13028 18582 13084
rect 18518 13024 18582 13028
rect 7882 12540 7946 12544
rect 7882 12484 7886 12540
rect 7886 12484 7942 12540
rect 7942 12484 7946 12540
rect 7882 12480 7946 12484
rect 7962 12540 8026 12544
rect 7962 12484 7966 12540
rect 7966 12484 8022 12540
rect 8022 12484 8026 12540
rect 7962 12480 8026 12484
rect 8042 12540 8106 12544
rect 8042 12484 8046 12540
rect 8046 12484 8102 12540
rect 8102 12484 8106 12540
rect 8042 12480 8106 12484
rect 8122 12540 8186 12544
rect 8122 12484 8126 12540
rect 8126 12484 8182 12540
rect 8182 12484 8186 12540
rect 8122 12480 8186 12484
rect 14813 12540 14877 12544
rect 14813 12484 14817 12540
rect 14817 12484 14873 12540
rect 14873 12484 14877 12540
rect 14813 12480 14877 12484
rect 14893 12540 14957 12544
rect 14893 12484 14897 12540
rect 14897 12484 14953 12540
rect 14953 12484 14957 12540
rect 14893 12480 14957 12484
rect 14973 12540 15037 12544
rect 14973 12484 14977 12540
rect 14977 12484 15033 12540
rect 15033 12484 15037 12540
rect 14973 12480 15037 12484
rect 15053 12540 15117 12544
rect 15053 12484 15057 12540
rect 15057 12484 15113 12540
rect 15113 12484 15117 12540
rect 15053 12480 15117 12484
rect 4417 11996 4481 12000
rect 4417 11940 4421 11996
rect 4421 11940 4477 11996
rect 4477 11940 4481 11996
rect 4417 11936 4481 11940
rect 4497 11996 4561 12000
rect 4497 11940 4501 11996
rect 4501 11940 4557 11996
rect 4557 11940 4561 11996
rect 4497 11936 4561 11940
rect 4577 11996 4641 12000
rect 4577 11940 4581 11996
rect 4581 11940 4637 11996
rect 4637 11940 4641 11996
rect 4577 11936 4641 11940
rect 4657 11996 4721 12000
rect 4657 11940 4661 11996
rect 4661 11940 4717 11996
rect 4717 11940 4721 11996
rect 4657 11936 4721 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 18278 11996 18342 12000
rect 18278 11940 18282 11996
rect 18282 11940 18338 11996
rect 18338 11940 18342 11996
rect 18278 11936 18342 11940
rect 18358 11996 18422 12000
rect 18358 11940 18362 11996
rect 18362 11940 18418 11996
rect 18418 11940 18422 11996
rect 18358 11936 18422 11940
rect 18438 11996 18502 12000
rect 18438 11940 18442 11996
rect 18442 11940 18498 11996
rect 18498 11940 18502 11996
rect 18438 11936 18502 11940
rect 18518 11996 18582 12000
rect 18518 11940 18522 11996
rect 18522 11940 18578 11996
rect 18578 11940 18582 11996
rect 18518 11936 18582 11940
rect 7882 11452 7946 11456
rect 7882 11396 7886 11452
rect 7886 11396 7942 11452
rect 7942 11396 7946 11452
rect 7882 11392 7946 11396
rect 7962 11452 8026 11456
rect 7962 11396 7966 11452
rect 7966 11396 8022 11452
rect 8022 11396 8026 11452
rect 7962 11392 8026 11396
rect 8042 11452 8106 11456
rect 8042 11396 8046 11452
rect 8046 11396 8102 11452
rect 8102 11396 8106 11452
rect 8042 11392 8106 11396
rect 8122 11452 8186 11456
rect 8122 11396 8126 11452
rect 8126 11396 8182 11452
rect 8182 11396 8186 11452
rect 8122 11392 8186 11396
rect 14813 11452 14877 11456
rect 14813 11396 14817 11452
rect 14817 11396 14873 11452
rect 14873 11396 14877 11452
rect 14813 11392 14877 11396
rect 14893 11452 14957 11456
rect 14893 11396 14897 11452
rect 14897 11396 14953 11452
rect 14953 11396 14957 11452
rect 14893 11392 14957 11396
rect 14973 11452 15037 11456
rect 14973 11396 14977 11452
rect 14977 11396 15033 11452
rect 15033 11396 15037 11452
rect 14973 11392 15037 11396
rect 15053 11452 15117 11456
rect 15053 11396 15057 11452
rect 15057 11396 15113 11452
rect 15113 11396 15117 11452
rect 15053 11392 15117 11396
rect 4417 10908 4481 10912
rect 4417 10852 4421 10908
rect 4421 10852 4477 10908
rect 4477 10852 4481 10908
rect 4417 10848 4481 10852
rect 4497 10908 4561 10912
rect 4497 10852 4501 10908
rect 4501 10852 4557 10908
rect 4557 10852 4561 10908
rect 4497 10848 4561 10852
rect 4577 10908 4641 10912
rect 4577 10852 4581 10908
rect 4581 10852 4637 10908
rect 4637 10852 4641 10908
rect 4577 10848 4641 10852
rect 4657 10908 4721 10912
rect 4657 10852 4661 10908
rect 4661 10852 4717 10908
rect 4717 10852 4721 10908
rect 4657 10848 4721 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 18278 10908 18342 10912
rect 18278 10852 18282 10908
rect 18282 10852 18338 10908
rect 18338 10852 18342 10908
rect 18278 10848 18342 10852
rect 18358 10908 18422 10912
rect 18358 10852 18362 10908
rect 18362 10852 18418 10908
rect 18418 10852 18422 10908
rect 18358 10848 18422 10852
rect 18438 10908 18502 10912
rect 18438 10852 18442 10908
rect 18442 10852 18498 10908
rect 18498 10852 18502 10908
rect 18438 10848 18502 10852
rect 18518 10908 18582 10912
rect 18518 10852 18522 10908
rect 18522 10852 18578 10908
rect 18578 10852 18582 10908
rect 18518 10848 18582 10852
rect 7882 10364 7946 10368
rect 7882 10308 7886 10364
rect 7886 10308 7942 10364
rect 7942 10308 7946 10364
rect 7882 10304 7946 10308
rect 7962 10364 8026 10368
rect 7962 10308 7966 10364
rect 7966 10308 8022 10364
rect 8022 10308 8026 10364
rect 7962 10304 8026 10308
rect 8042 10364 8106 10368
rect 8042 10308 8046 10364
rect 8046 10308 8102 10364
rect 8102 10308 8106 10364
rect 8042 10304 8106 10308
rect 8122 10364 8186 10368
rect 8122 10308 8126 10364
rect 8126 10308 8182 10364
rect 8182 10308 8186 10364
rect 8122 10304 8186 10308
rect 14813 10364 14877 10368
rect 14813 10308 14817 10364
rect 14817 10308 14873 10364
rect 14873 10308 14877 10364
rect 14813 10304 14877 10308
rect 14893 10364 14957 10368
rect 14893 10308 14897 10364
rect 14897 10308 14953 10364
rect 14953 10308 14957 10364
rect 14893 10304 14957 10308
rect 14973 10364 15037 10368
rect 14973 10308 14977 10364
rect 14977 10308 15033 10364
rect 15033 10308 15037 10364
rect 14973 10304 15037 10308
rect 15053 10364 15117 10368
rect 15053 10308 15057 10364
rect 15057 10308 15113 10364
rect 15113 10308 15117 10364
rect 15053 10304 15117 10308
rect 4417 9820 4481 9824
rect 4417 9764 4421 9820
rect 4421 9764 4477 9820
rect 4477 9764 4481 9820
rect 4417 9760 4481 9764
rect 4497 9820 4561 9824
rect 4497 9764 4501 9820
rect 4501 9764 4557 9820
rect 4557 9764 4561 9820
rect 4497 9760 4561 9764
rect 4577 9820 4641 9824
rect 4577 9764 4581 9820
rect 4581 9764 4637 9820
rect 4637 9764 4641 9820
rect 4577 9760 4641 9764
rect 4657 9820 4721 9824
rect 4657 9764 4661 9820
rect 4661 9764 4717 9820
rect 4717 9764 4721 9820
rect 4657 9760 4721 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 18278 9820 18342 9824
rect 18278 9764 18282 9820
rect 18282 9764 18338 9820
rect 18338 9764 18342 9820
rect 18278 9760 18342 9764
rect 18358 9820 18422 9824
rect 18358 9764 18362 9820
rect 18362 9764 18418 9820
rect 18418 9764 18422 9820
rect 18358 9760 18422 9764
rect 18438 9820 18502 9824
rect 18438 9764 18442 9820
rect 18442 9764 18498 9820
rect 18498 9764 18502 9820
rect 18438 9760 18502 9764
rect 18518 9820 18582 9824
rect 18518 9764 18522 9820
rect 18522 9764 18578 9820
rect 18578 9764 18582 9820
rect 18518 9760 18582 9764
rect 7882 9276 7946 9280
rect 7882 9220 7886 9276
rect 7886 9220 7942 9276
rect 7942 9220 7946 9276
rect 7882 9216 7946 9220
rect 7962 9276 8026 9280
rect 7962 9220 7966 9276
rect 7966 9220 8022 9276
rect 8022 9220 8026 9276
rect 7962 9216 8026 9220
rect 8042 9276 8106 9280
rect 8042 9220 8046 9276
rect 8046 9220 8102 9276
rect 8102 9220 8106 9276
rect 8042 9216 8106 9220
rect 8122 9276 8186 9280
rect 8122 9220 8126 9276
rect 8126 9220 8182 9276
rect 8182 9220 8186 9276
rect 8122 9216 8186 9220
rect 14813 9276 14877 9280
rect 14813 9220 14817 9276
rect 14817 9220 14873 9276
rect 14873 9220 14877 9276
rect 14813 9216 14877 9220
rect 14893 9276 14957 9280
rect 14893 9220 14897 9276
rect 14897 9220 14953 9276
rect 14953 9220 14957 9276
rect 14893 9216 14957 9220
rect 14973 9276 15037 9280
rect 14973 9220 14977 9276
rect 14977 9220 15033 9276
rect 15033 9220 15037 9276
rect 14973 9216 15037 9220
rect 15053 9276 15117 9280
rect 15053 9220 15057 9276
rect 15057 9220 15113 9276
rect 15113 9220 15117 9276
rect 15053 9216 15117 9220
rect 4417 8732 4481 8736
rect 4417 8676 4421 8732
rect 4421 8676 4477 8732
rect 4477 8676 4481 8732
rect 4417 8672 4481 8676
rect 4497 8732 4561 8736
rect 4497 8676 4501 8732
rect 4501 8676 4557 8732
rect 4557 8676 4561 8732
rect 4497 8672 4561 8676
rect 4577 8732 4641 8736
rect 4577 8676 4581 8732
rect 4581 8676 4637 8732
rect 4637 8676 4641 8732
rect 4577 8672 4641 8676
rect 4657 8732 4721 8736
rect 4657 8676 4661 8732
rect 4661 8676 4717 8732
rect 4717 8676 4721 8732
rect 4657 8672 4721 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 18278 8732 18342 8736
rect 18278 8676 18282 8732
rect 18282 8676 18338 8732
rect 18338 8676 18342 8732
rect 18278 8672 18342 8676
rect 18358 8732 18422 8736
rect 18358 8676 18362 8732
rect 18362 8676 18418 8732
rect 18418 8676 18422 8732
rect 18358 8672 18422 8676
rect 18438 8732 18502 8736
rect 18438 8676 18442 8732
rect 18442 8676 18498 8732
rect 18498 8676 18502 8732
rect 18438 8672 18502 8676
rect 18518 8732 18582 8736
rect 18518 8676 18522 8732
rect 18522 8676 18578 8732
rect 18578 8676 18582 8732
rect 18518 8672 18582 8676
rect 7882 8188 7946 8192
rect 7882 8132 7886 8188
rect 7886 8132 7942 8188
rect 7942 8132 7946 8188
rect 7882 8128 7946 8132
rect 7962 8188 8026 8192
rect 7962 8132 7966 8188
rect 7966 8132 8022 8188
rect 8022 8132 8026 8188
rect 7962 8128 8026 8132
rect 8042 8188 8106 8192
rect 8042 8132 8046 8188
rect 8046 8132 8102 8188
rect 8102 8132 8106 8188
rect 8042 8128 8106 8132
rect 8122 8188 8186 8192
rect 8122 8132 8126 8188
rect 8126 8132 8182 8188
rect 8182 8132 8186 8188
rect 8122 8128 8186 8132
rect 14813 8188 14877 8192
rect 14813 8132 14817 8188
rect 14817 8132 14873 8188
rect 14873 8132 14877 8188
rect 14813 8128 14877 8132
rect 14893 8188 14957 8192
rect 14893 8132 14897 8188
rect 14897 8132 14953 8188
rect 14953 8132 14957 8188
rect 14893 8128 14957 8132
rect 14973 8188 15037 8192
rect 14973 8132 14977 8188
rect 14977 8132 15033 8188
rect 15033 8132 15037 8188
rect 14973 8128 15037 8132
rect 15053 8188 15117 8192
rect 15053 8132 15057 8188
rect 15057 8132 15113 8188
rect 15113 8132 15117 8188
rect 15053 8128 15117 8132
rect 4417 7644 4481 7648
rect 4417 7588 4421 7644
rect 4421 7588 4477 7644
rect 4477 7588 4481 7644
rect 4417 7584 4481 7588
rect 4497 7644 4561 7648
rect 4497 7588 4501 7644
rect 4501 7588 4557 7644
rect 4557 7588 4561 7644
rect 4497 7584 4561 7588
rect 4577 7644 4641 7648
rect 4577 7588 4581 7644
rect 4581 7588 4637 7644
rect 4637 7588 4641 7644
rect 4577 7584 4641 7588
rect 4657 7644 4721 7648
rect 4657 7588 4661 7644
rect 4661 7588 4717 7644
rect 4717 7588 4721 7644
rect 4657 7584 4721 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 18278 7644 18342 7648
rect 18278 7588 18282 7644
rect 18282 7588 18338 7644
rect 18338 7588 18342 7644
rect 18278 7584 18342 7588
rect 18358 7644 18422 7648
rect 18358 7588 18362 7644
rect 18362 7588 18418 7644
rect 18418 7588 18422 7644
rect 18358 7584 18422 7588
rect 18438 7644 18502 7648
rect 18438 7588 18442 7644
rect 18442 7588 18498 7644
rect 18498 7588 18502 7644
rect 18438 7584 18502 7588
rect 18518 7644 18582 7648
rect 18518 7588 18522 7644
rect 18522 7588 18578 7644
rect 18578 7588 18582 7644
rect 18518 7584 18582 7588
rect 7882 7100 7946 7104
rect 7882 7044 7886 7100
rect 7886 7044 7942 7100
rect 7942 7044 7946 7100
rect 7882 7040 7946 7044
rect 7962 7100 8026 7104
rect 7962 7044 7966 7100
rect 7966 7044 8022 7100
rect 8022 7044 8026 7100
rect 7962 7040 8026 7044
rect 8042 7100 8106 7104
rect 8042 7044 8046 7100
rect 8046 7044 8102 7100
rect 8102 7044 8106 7100
rect 8042 7040 8106 7044
rect 8122 7100 8186 7104
rect 8122 7044 8126 7100
rect 8126 7044 8182 7100
rect 8182 7044 8186 7100
rect 8122 7040 8186 7044
rect 14813 7100 14877 7104
rect 14813 7044 14817 7100
rect 14817 7044 14873 7100
rect 14873 7044 14877 7100
rect 14813 7040 14877 7044
rect 14893 7100 14957 7104
rect 14893 7044 14897 7100
rect 14897 7044 14953 7100
rect 14953 7044 14957 7100
rect 14893 7040 14957 7044
rect 14973 7100 15037 7104
rect 14973 7044 14977 7100
rect 14977 7044 15033 7100
rect 15033 7044 15037 7100
rect 14973 7040 15037 7044
rect 15053 7100 15117 7104
rect 15053 7044 15057 7100
rect 15057 7044 15113 7100
rect 15113 7044 15117 7100
rect 15053 7040 15117 7044
rect 4417 6556 4481 6560
rect 4417 6500 4421 6556
rect 4421 6500 4477 6556
rect 4477 6500 4481 6556
rect 4417 6496 4481 6500
rect 4497 6556 4561 6560
rect 4497 6500 4501 6556
rect 4501 6500 4557 6556
rect 4557 6500 4561 6556
rect 4497 6496 4561 6500
rect 4577 6556 4641 6560
rect 4577 6500 4581 6556
rect 4581 6500 4637 6556
rect 4637 6500 4641 6556
rect 4577 6496 4641 6500
rect 4657 6556 4721 6560
rect 4657 6500 4661 6556
rect 4661 6500 4717 6556
rect 4717 6500 4721 6556
rect 4657 6496 4721 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 18278 6556 18342 6560
rect 18278 6500 18282 6556
rect 18282 6500 18338 6556
rect 18338 6500 18342 6556
rect 18278 6496 18342 6500
rect 18358 6556 18422 6560
rect 18358 6500 18362 6556
rect 18362 6500 18418 6556
rect 18418 6500 18422 6556
rect 18358 6496 18422 6500
rect 18438 6556 18502 6560
rect 18438 6500 18442 6556
rect 18442 6500 18498 6556
rect 18498 6500 18502 6556
rect 18438 6496 18502 6500
rect 18518 6556 18582 6560
rect 18518 6500 18522 6556
rect 18522 6500 18578 6556
rect 18578 6500 18582 6556
rect 18518 6496 18582 6500
rect 7882 6012 7946 6016
rect 7882 5956 7886 6012
rect 7886 5956 7942 6012
rect 7942 5956 7946 6012
rect 7882 5952 7946 5956
rect 7962 6012 8026 6016
rect 7962 5956 7966 6012
rect 7966 5956 8022 6012
rect 8022 5956 8026 6012
rect 7962 5952 8026 5956
rect 8042 6012 8106 6016
rect 8042 5956 8046 6012
rect 8046 5956 8102 6012
rect 8102 5956 8106 6012
rect 8042 5952 8106 5956
rect 8122 6012 8186 6016
rect 8122 5956 8126 6012
rect 8126 5956 8182 6012
rect 8182 5956 8186 6012
rect 8122 5952 8186 5956
rect 14813 6012 14877 6016
rect 14813 5956 14817 6012
rect 14817 5956 14873 6012
rect 14873 5956 14877 6012
rect 14813 5952 14877 5956
rect 14893 6012 14957 6016
rect 14893 5956 14897 6012
rect 14897 5956 14953 6012
rect 14953 5956 14957 6012
rect 14893 5952 14957 5956
rect 14973 6012 15037 6016
rect 14973 5956 14977 6012
rect 14977 5956 15033 6012
rect 15033 5956 15037 6012
rect 14973 5952 15037 5956
rect 15053 6012 15117 6016
rect 15053 5956 15057 6012
rect 15057 5956 15113 6012
rect 15113 5956 15117 6012
rect 15053 5952 15117 5956
rect 4417 5468 4481 5472
rect 4417 5412 4421 5468
rect 4421 5412 4477 5468
rect 4477 5412 4481 5468
rect 4417 5408 4481 5412
rect 4497 5468 4561 5472
rect 4497 5412 4501 5468
rect 4501 5412 4557 5468
rect 4557 5412 4561 5468
rect 4497 5408 4561 5412
rect 4577 5468 4641 5472
rect 4577 5412 4581 5468
rect 4581 5412 4637 5468
rect 4637 5412 4641 5468
rect 4577 5408 4641 5412
rect 4657 5468 4721 5472
rect 4657 5412 4661 5468
rect 4661 5412 4717 5468
rect 4717 5412 4721 5468
rect 4657 5408 4721 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 18278 5468 18342 5472
rect 18278 5412 18282 5468
rect 18282 5412 18338 5468
rect 18338 5412 18342 5468
rect 18278 5408 18342 5412
rect 18358 5468 18422 5472
rect 18358 5412 18362 5468
rect 18362 5412 18418 5468
rect 18418 5412 18422 5468
rect 18358 5408 18422 5412
rect 18438 5468 18502 5472
rect 18438 5412 18442 5468
rect 18442 5412 18498 5468
rect 18498 5412 18502 5468
rect 18438 5408 18502 5412
rect 18518 5468 18582 5472
rect 18518 5412 18522 5468
rect 18522 5412 18578 5468
rect 18578 5412 18582 5468
rect 18518 5408 18582 5412
rect 7882 4924 7946 4928
rect 7882 4868 7886 4924
rect 7886 4868 7942 4924
rect 7942 4868 7946 4924
rect 7882 4864 7946 4868
rect 7962 4924 8026 4928
rect 7962 4868 7966 4924
rect 7966 4868 8022 4924
rect 8022 4868 8026 4924
rect 7962 4864 8026 4868
rect 8042 4924 8106 4928
rect 8042 4868 8046 4924
rect 8046 4868 8102 4924
rect 8102 4868 8106 4924
rect 8042 4864 8106 4868
rect 8122 4924 8186 4928
rect 8122 4868 8126 4924
rect 8126 4868 8182 4924
rect 8182 4868 8186 4924
rect 8122 4864 8186 4868
rect 14813 4924 14877 4928
rect 14813 4868 14817 4924
rect 14817 4868 14873 4924
rect 14873 4868 14877 4924
rect 14813 4864 14877 4868
rect 14893 4924 14957 4928
rect 14893 4868 14897 4924
rect 14897 4868 14953 4924
rect 14953 4868 14957 4924
rect 14893 4864 14957 4868
rect 14973 4924 15037 4928
rect 14973 4868 14977 4924
rect 14977 4868 15033 4924
rect 15033 4868 15037 4924
rect 14973 4864 15037 4868
rect 15053 4924 15117 4928
rect 15053 4868 15057 4924
rect 15057 4868 15113 4924
rect 15113 4868 15117 4924
rect 15053 4864 15117 4868
rect 4417 4380 4481 4384
rect 4417 4324 4421 4380
rect 4421 4324 4477 4380
rect 4477 4324 4481 4380
rect 4417 4320 4481 4324
rect 4497 4380 4561 4384
rect 4497 4324 4501 4380
rect 4501 4324 4557 4380
rect 4557 4324 4561 4380
rect 4497 4320 4561 4324
rect 4577 4380 4641 4384
rect 4577 4324 4581 4380
rect 4581 4324 4637 4380
rect 4637 4324 4641 4380
rect 4577 4320 4641 4324
rect 4657 4380 4721 4384
rect 4657 4324 4661 4380
rect 4661 4324 4717 4380
rect 4717 4324 4721 4380
rect 4657 4320 4721 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 18278 4380 18342 4384
rect 18278 4324 18282 4380
rect 18282 4324 18338 4380
rect 18338 4324 18342 4380
rect 18278 4320 18342 4324
rect 18358 4380 18422 4384
rect 18358 4324 18362 4380
rect 18362 4324 18418 4380
rect 18418 4324 18422 4380
rect 18358 4320 18422 4324
rect 18438 4380 18502 4384
rect 18438 4324 18442 4380
rect 18442 4324 18498 4380
rect 18498 4324 18502 4380
rect 18438 4320 18502 4324
rect 18518 4380 18582 4384
rect 18518 4324 18522 4380
rect 18522 4324 18578 4380
rect 18578 4324 18582 4380
rect 18518 4320 18582 4324
rect 7882 3836 7946 3840
rect 7882 3780 7886 3836
rect 7886 3780 7942 3836
rect 7942 3780 7946 3836
rect 7882 3776 7946 3780
rect 7962 3836 8026 3840
rect 7962 3780 7966 3836
rect 7966 3780 8022 3836
rect 8022 3780 8026 3836
rect 7962 3776 8026 3780
rect 8042 3836 8106 3840
rect 8042 3780 8046 3836
rect 8046 3780 8102 3836
rect 8102 3780 8106 3836
rect 8042 3776 8106 3780
rect 8122 3836 8186 3840
rect 8122 3780 8126 3836
rect 8126 3780 8182 3836
rect 8182 3780 8186 3836
rect 8122 3776 8186 3780
rect 14813 3836 14877 3840
rect 14813 3780 14817 3836
rect 14817 3780 14873 3836
rect 14873 3780 14877 3836
rect 14813 3776 14877 3780
rect 14893 3836 14957 3840
rect 14893 3780 14897 3836
rect 14897 3780 14953 3836
rect 14953 3780 14957 3836
rect 14893 3776 14957 3780
rect 14973 3836 15037 3840
rect 14973 3780 14977 3836
rect 14977 3780 15033 3836
rect 15033 3780 15037 3836
rect 14973 3776 15037 3780
rect 15053 3836 15117 3840
rect 15053 3780 15057 3836
rect 15057 3780 15113 3836
rect 15113 3780 15117 3836
rect 15053 3776 15117 3780
rect 4417 3292 4481 3296
rect 4417 3236 4421 3292
rect 4421 3236 4477 3292
rect 4477 3236 4481 3292
rect 4417 3232 4481 3236
rect 4497 3292 4561 3296
rect 4497 3236 4501 3292
rect 4501 3236 4557 3292
rect 4557 3236 4561 3292
rect 4497 3232 4561 3236
rect 4577 3292 4641 3296
rect 4577 3236 4581 3292
rect 4581 3236 4637 3292
rect 4637 3236 4641 3292
rect 4577 3232 4641 3236
rect 4657 3292 4721 3296
rect 4657 3236 4661 3292
rect 4661 3236 4717 3292
rect 4717 3236 4721 3292
rect 4657 3232 4721 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 18278 3292 18342 3296
rect 18278 3236 18282 3292
rect 18282 3236 18338 3292
rect 18338 3236 18342 3292
rect 18278 3232 18342 3236
rect 18358 3292 18422 3296
rect 18358 3236 18362 3292
rect 18362 3236 18418 3292
rect 18418 3236 18422 3292
rect 18358 3232 18422 3236
rect 18438 3292 18502 3296
rect 18438 3236 18442 3292
rect 18442 3236 18498 3292
rect 18498 3236 18502 3292
rect 18438 3232 18502 3236
rect 18518 3292 18582 3296
rect 18518 3236 18522 3292
rect 18522 3236 18578 3292
rect 18578 3236 18582 3292
rect 18518 3232 18582 3236
rect 7882 2748 7946 2752
rect 7882 2692 7886 2748
rect 7886 2692 7942 2748
rect 7942 2692 7946 2748
rect 7882 2688 7946 2692
rect 7962 2748 8026 2752
rect 7962 2692 7966 2748
rect 7966 2692 8022 2748
rect 8022 2692 8026 2748
rect 7962 2688 8026 2692
rect 8042 2748 8106 2752
rect 8042 2692 8046 2748
rect 8046 2692 8102 2748
rect 8102 2692 8106 2748
rect 8042 2688 8106 2692
rect 8122 2748 8186 2752
rect 8122 2692 8126 2748
rect 8126 2692 8182 2748
rect 8182 2692 8186 2748
rect 8122 2688 8186 2692
rect 14813 2748 14877 2752
rect 14813 2692 14817 2748
rect 14817 2692 14873 2748
rect 14873 2692 14877 2748
rect 14813 2688 14877 2692
rect 14893 2748 14957 2752
rect 14893 2692 14897 2748
rect 14897 2692 14953 2748
rect 14953 2692 14957 2748
rect 14893 2688 14957 2692
rect 14973 2748 15037 2752
rect 14973 2692 14977 2748
rect 14977 2692 15033 2748
rect 15033 2692 15037 2748
rect 14973 2688 15037 2692
rect 15053 2748 15117 2752
rect 15053 2692 15057 2748
rect 15057 2692 15113 2748
rect 15113 2692 15117 2748
rect 15053 2688 15117 2692
rect 4417 2204 4481 2208
rect 4417 2148 4421 2204
rect 4421 2148 4477 2204
rect 4477 2148 4481 2204
rect 4417 2144 4481 2148
rect 4497 2204 4561 2208
rect 4497 2148 4501 2204
rect 4501 2148 4557 2204
rect 4557 2148 4561 2204
rect 4497 2144 4561 2148
rect 4577 2204 4641 2208
rect 4577 2148 4581 2204
rect 4581 2148 4637 2204
rect 4637 2148 4641 2204
rect 4577 2144 4641 2148
rect 4657 2204 4721 2208
rect 4657 2148 4661 2204
rect 4661 2148 4717 2204
rect 4717 2148 4721 2204
rect 4657 2144 4721 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 18278 2204 18342 2208
rect 18278 2148 18282 2204
rect 18282 2148 18338 2204
rect 18338 2148 18342 2204
rect 18278 2144 18342 2148
rect 18358 2204 18422 2208
rect 18358 2148 18362 2204
rect 18362 2148 18418 2204
rect 18418 2148 18422 2204
rect 18358 2144 18422 2148
rect 18438 2204 18502 2208
rect 18438 2148 18442 2204
rect 18442 2148 18498 2204
rect 18498 2148 18502 2204
rect 18438 2144 18502 2148
rect 18518 2204 18582 2208
rect 18518 2148 18522 2204
rect 18522 2148 18578 2204
rect 18578 2148 18582 2204
rect 18518 2144 18582 2148
<< metal4 >>
rect 4409 20704 4729 20720
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 19616 4729 20640
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 18528 4729 19552
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 17440 4729 18464
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 16352 4729 17376
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 15264 4729 16288
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 14176 4729 15200
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 13088 4729 14112
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 12000 4729 13024
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 10912 4729 11936
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 9824 4729 10848
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 8736 4729 9760
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 7648 4729 8672
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 6560 4729 7584
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 5472 4729 6496
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 4384 4729 5408
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 3296 4729 4320
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 2208 4729 3232
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2128 4729 2144
rect 7874 20160 8195 20720
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8195 20160
rect 7874 19072 8195 20096
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8195 19072
rect 7874 17984 8195 19008
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8195 17984
rect 7874 16896 8195 17920
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8195 16896
rect 7874 15808 8195 16832
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8195 15808
rect 7874 14720 8195 15744
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8195 14720
rect 7874 13632 8195 14656
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8195 13632
rect 7874 12544 8195 13568
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8195 12544
rect 7874 11456 8195 12480
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8195 11456
rect 7874 10368 8195 11392
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8195 10368
rect 7874 9280 8195 10304
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8195 9280
rect 7874 8192 8195 9216
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8195 8192
rect 7874 7104 8195 8128
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8195 7104
rect 7874 6016 8195 7040
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8195 6016
rect 7874 4928 8195 5952
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8195 4928
rect 7874 3840 8195 4864
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8195 3840
rect 7874 2752 8195 3776
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8195 2752
rect 7874 2128 8195 2688
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 14805 20160 15125 20720
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 19072 15125 20096
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 17984 15125 19008
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 16896 15125 17920
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 15808 15125 16832
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 14720 15125 15744
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 13632 15125 14656
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 12544 15125 13568
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 11456 15125 12480
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 10368 15125 11392
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 9280 15125 10304
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 8192 15125 9216
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 7104 15125 8128
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 6016 15125 7040
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 4928 15125 5952
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 3840 15125 4864
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 2752 15125 3776
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2128 15125 2688
rect 18270 20704 18591 20720
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18591 20704
rect 18270 19616 18591 20640
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18591 19616
rect 18270 18528 18591 19552
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18591 18528
rect 18270 17440 18591 18464
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18591 17440
rect 18270 16352 18591 17376
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18591 16352
rect 18270 15264 18591 16288
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18591 15264
rect 18270 14176 18591 15200
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18591 14176
rect 18270 13088 18591 14112
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18591 13088
rect 18270 12000 18591 13024
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18591 12000
rect 18270 10912 18591 11936
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18591 10912
rect 18270 9824 18591 10848
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18591 9824
rect 18270 8736 18591 9760
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18591 8736
rect 18270 7648 18591 8672
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18591 7648
rect 18270 6560 18591 7584
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18591 6560
rect 18270 5472 18591 6496
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18591 5472
rect 18270 4384 18591 5408
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18591 4384
rect 18270 3296 18591 4320
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18591 3296
rect 18270 2208 18591 3232
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18591 2208
rect 18270 2128 18591 2144
use sky130_fd_sc_hd__fill_2  FILLER_1_7 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1748 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1608910539
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1380 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1564 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608910539
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_11
timestamp 1608910539
transform 1 0 2116 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16
timestamp 1608910539
transform 1 0 2576 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11
timestamp 1608910539
transform 1 0 2116 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 2392 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 2760 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1608910539
transform 1 0 2300 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_40
timestamp 1608910539
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_22
timestamp 1608910539
transform 1 0 3128 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_34 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 4232 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3312 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_1_62 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 6808 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_58
timestamp 1608910539
transform 1 0 6440 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60
timestamp 1608910539
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50
timestamp 1608910539
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46
timestamp 1608910539
transform 1 0 5336 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608910539
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608910539
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1608910539
transform 1 0 5796 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 4968 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_1_72
timestamp 1608910539
transform 1 0 7728 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72
timestamp 1608910539
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1608910539
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1608910539
transform 1 0 6900 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_81
timestamp 1608910539
transform 1 0 8556 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_76
timestamp 1608910539
transform 1 0 8096 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_80
timestamp 1608910539
transform 1 0 8464 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76
timestamp 1608910539
transform 1 0 8096 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8280 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 7912 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1608910539
transform 1 0 8648 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _058_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 8280 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 8740 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_1_99
timestamp 1608910539
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_103 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 10580 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1608910539
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608910539
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1608910539
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10396 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1608910539
transform 1 0 11224 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_109
timestamp 1608910539
transform 1 0 11132 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 11224 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116
timestamp 1608910539
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_112
timestamp 1608910539
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 11408 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _091_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 11868 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_118
timestamp 1608910539
transform 1 0 11960 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_121
timestamp 1608910539
transform 1 0 12236 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608910539
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608910539
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 12420 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1608910539
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_129
timestamp 1608910539
transform 1 0 12972 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_129
timestamp 1608910539
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 13156 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1608910539
transform 1 0 13156 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_137
timestamp 1608910539
transform 1 0 13708 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_135
timestamp 1608910539
transform 1 0 13524 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1608910539
transform 1 0 13708 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_143
timestamp 1608910539
transform 1 0 14260 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1608910539
transform 1 0 14076 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 14444 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1608910539
transform 1 0 14260 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1608910539
transform 1 0 13892 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_151
timestamp 1608910539
transform 1 0 14996 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1608910539
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1608910539
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608910539
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l2_in_0_
timestamp 1608910539
transform 1 0 15180 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1608910539
transform 1 0 14812 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_162
timestamp 1608910539
transform 1 0 16008 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_160
timestamp 1608910539
transform 1 0 15824 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 16192 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1608910539
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1608910539
transform 1 0 16376 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_170
timestamp 1608910539
transform 1 0 16744 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_175
timestamp 1608910539
transform 1 0 17204 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_170
timestamp 1608910539
transform 1 0 16744 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 16928 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1608910539
transform 1 0 17388 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1608910539
transform 1 0 16928 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_182
timestamp 1608910539
transform 1 0 17848 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_178
timestamp 1608910539
transform 1 0 17480 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_185
timestamp 1608910539
transform 1 0 18124 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181
timestamp 1608910539
transform 1 0 17756 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608910539
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608910539
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1608910539
transform 1 0 18032 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1608910539
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_206
timestamp 1608910539
transform 1 0 20056 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_194
timestamp 1608910539
transform 1 0 18952 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_188
timestamp 1608910539
transform 1 0 18400 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1608910539
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1608910539
transform 1 0 18584 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_221
timestamp 1608910539
transform 1 0 21436 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_221
timestamp 1608910539
transform 1 0 21436 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_218
timestamp 1608910539
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1608910539
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1608910539
transform 1 0 21252 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608910539
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608910539
transform -1 0 21896 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608910539
transform -1 0 21896 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 20332 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_20
timestamp 1608910539
transform 1 0 2944 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3
timestamp 1608910539
transform 1 0 1380 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608910539
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 1472 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_2_41
timestamp 1608910539
transform 1 0 4876 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_28
timestamp 1608910539
transform 1 0 3680 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608910539
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 3128 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1608910539
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_60
timestamp 1608910539
transform 1 0 6624 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1608910539
transform 1 0 6808 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 5152 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_2_71
timestamp 1608910539
transform 1 0 7636 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 7912 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_102
timestamp 1608910539
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1608910539
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608910539
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1608910539
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_2_124
timestamp 1608910539
transform 1 0 12512 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_114
timestamp 1608910539
transform 1 0 11592 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_110
timestamp 1608910539
transform 1 0 11224 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_106
timestamp 1608910539
transform 1 0 10856 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 11408 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 11040 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 11960 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_136
timestamp 1608910539
transform 1 0 13616 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_0_
timestamp 1608910539
transform 1 0 13800 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l2_in_0_
timestamp 1608910539
transform 1 0 12788 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_2_164
timestamp 1608910539
transform 1 0 16192 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_158
timestamp 1608910539
transform 1 0 15640 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1608910539
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_147
timestamp 1608910539
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608910539
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1608910539
transform 1 0 15824 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1608910539
transform 1 0 15272 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_182
timestamp 1608910539
transform 1 0 17848 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_176
timestamp 1608910539
transform 1 0 17296 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 16744 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1608910539
transform 1 0 17480 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_204
timestamp 1608910539
transform 1 0 19872 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_194
timestamp 1608910539
transform 1 0 18952 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1608910539
transform 1 0 19688 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1608910539
transform 1 0 20056 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_219
timestamp 1608910539
transform 1 0 21252 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_210
timestamp 1608910539
transform 1 0 20424 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608910539
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608910539
transform -1 0 21896 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1608910539
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_7
timestamp 1608910539
transform 1 0 1748 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1608910539
transform 1 0 1380 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608910539
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 1932 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _069_
timestamp 1608910539
transform 1 0 1472 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_25
timestamp 1608910539
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 3588 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1608910539
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1608910539
transform 1 0 6072 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_43
timestamp 1608910539
transform 1 0 5060 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608910539
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1608910539
transform 1 0 5244 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 6808 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1608910539
transform 1 0 6256 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_82
timestamp 1608910539
transform 1 0 8648 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_78
timestamp 1608910539
transform 1 0 8280 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 8464 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_104
timestamp 1608910539
transform 1 0 10672 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_93
timestamp 1608910539
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1608910539
transform 1 0 9844 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1608910539
transform 1 0 8832 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1608910539
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_116
timestamp 1608910539
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608910539
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10948 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 12420 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_139
timestamp 1608910539
transform 1 0 13892 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 14076 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_157
timestamp 1608910539
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15732 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1608910539
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_180
timestamp 1608910539
transform 1 0 17664 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_175
timestamp 1608910539
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608910539
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1608910539
transform 1 0 17388 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_208
timestamp 1608910539
transform 1 0 20240 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1608910539
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_221
timestamp 1608910539
transform 1 0 21436 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_216
timestamp 1608910539
transform 1 0 20976 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1608910539
transform 1 0 21252 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608910539
transform -1 0 21896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_17
timestamp 1608910539
transform 1 0 2668 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_6
timestamp 1608910539
transform 1 0 1656 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 1608910539
transform 1 0 1380 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 1472 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608910539
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1608910539
transform 1 0 2852 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1608910539
transform 1 0 1840 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_39
timestamp 1608910539
transform 1 0 4692 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_36
timestamp 1608910539
transform 1 0 4416 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_32
timestamp 1608910539
transform 1 0 4048 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_28
timestamp 1608910539
transform 1 0 3680 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 4508 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 4876 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608910539
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_59
timestamp 1608910539
transform 1 0 6532 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_54
timestamp 1608910539
transform 1 0 6072 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_43
timestamp 1608910539
transform 1 0 5060 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6348 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 6716 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1608910539
transform 1 0 5244 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_82
timestamp 1608910539
transform 1 0 8648 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_78
timestamp 1608910539
transform 1 0 8280 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_74
timestamp 1608910539
transform 1 0 7912 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_63
timestamp 1608910539
transform 1 0 6900 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 8464 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 8096 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_1_
timestamp 1608910539
transform 1 0 7084 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_4_99
timestamp 1608910539
transform 1 0 10212 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_95
timestamp 1608910539
transform 1 0 9844 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_89
timestamp 1608910539
transform 1 0 9292 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_86
timestamp 1608910539
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 10028 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9108 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608910539
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 10488 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_4_118
timestamp 1608910539
transform 1 0 11960 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_143
timestamp 1608910539
transform 1 0 14260 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_126
timestamp 1608910539
transform 1 0 12696 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 12788 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_157
timestamp 1608910539
transform 1 0 15548 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_154
timestamp 1608910539
transform 1 0 15272 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_151
timestamp 1608910539
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 15364 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608910539
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 15916 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_4_177
timestamp 1608910539
transform 1 0 17388 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l2_in_0_
timestamp 1608910539
transform 1 0 17572 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_4_200
timestamp 1608910539
transform 1 0 19504 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_188
timestamp 1608910539
transform 1 0 18400 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_221
timestamp 1608910539
transform 1 0 21436 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1608910539
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_212
timestamp 1608910539
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608910539
transform 1 0 21252 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608910539
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608910539
transform -1 0 21896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_15
timestamp 1608910539
transform 1 0 2484 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1608910539
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608910539
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_36
timestamp 1608910539
transform 1 0 4416 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_32
timestamp 1608910539
transform 1 0 4048 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_27
timestamp 1608910539
transform 1 0 3588 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_23
timestamp 1608910539
transform 1 0 3220 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 3404 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 3864 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_62
timestamp 1608910539
transform 1 0 6808 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1608910539
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_48
timestamp 1608910539
transform 1 0 5520 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608910539
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l3_in_0_
timestamp 1608910539
transform 1 0 5704 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_73
timestamp 1608910539
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8004 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_0_
timestamp 1608910539
transform 1 0 6992 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_98
timestamp 1608910539
transform 1 0 10120 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_88
timestamp 1608910539
transform 1 0 9200 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_84
timestamp 1608910539
transform 1 0 8832 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1608910539
transform 1 0 10304 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1608910539
transform 1 0 9292 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_118
timestamp 1608910539
transform 1 0 11960 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_114
timestamp 1608910539
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_109
timestamp 1608910539
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608910539
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1608910539
transform 1 0 11316 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1608910539
transform 1 0 12420 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_138
timestamp 1608910539
transform 1 0 13800 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_134
timestamp 1608910539
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_130
timestamp 1608910539
transform 1 0 13064 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_126
timestamp 1608910539
transform 1 0 12696 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1608910539
transform 1 0 13156 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1608910539
transform 1 0 16376 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_156
timestamp 1608910539
transform 1 0 15456 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_152
timestamp 1608910539
transform 1 0 15088 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_0_
timestamp 1608910539
transform 1 0 15548 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 14536 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_186
timestamp 1608910539
transform 1 0 18216 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_181
timestamp 1608910539
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_177
timestamp 1608910539
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 18032 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608910539
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1608910539
transform 1 0 16560 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_204
timestamp 1608910539
transform 1 0 19872 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_198
timestamp 1608910539
transform 1 0 19320 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 19964 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_221
timestamp 1608910539
transform 1 0 21436 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608910539
transform -1 0 21896 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_19
timestamp 1608910539
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_18
timestamp 1608910539
transform 1 0 2760 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3
timestamp 1608910539
transform 1 0 1380 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608910539
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608910539
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1608910539
transform 1 0 1932 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1608910539
transform 1 0 2944 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 1380 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_36
timestamp 1608910539
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_24
timestamp 1608910539
transform 1 0 3312 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_41
timestamp 1608910539
transform 1 0 4876 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1608910539
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608910539
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1608910539
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1608910539
transform 1 0 3588 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4600 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1608910539
transform 1 0 3036 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1608910539
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_54
timestamp 1608910539
transform 1 0 6072 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_45
timestamp 1608910539
transform 1 0 5244 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 5060 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608910539
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_1_
timestamp 1608910539
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 5980 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_76
timestamp 1608910539
transform 1 0 8096 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_71
timestamp 1608910539
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_69
timestamp 1608910539
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 8280 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 7636 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1608910539
transform 1 0 7820 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_98
timestamp 1608910539
transform 1 0 10120 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_94
timestamp 1608910539
transform 1 0 9752 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1608910539
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_87
timestamp 1608910539
transform 1 0 9108 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608910539
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 10488 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9660 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_7_118
timestamp 1608910539
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_120
timestamp 1608910539
transform 1 0 12144 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_109
timestamp 1608910539
transform 1 0 11132 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608910539
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1608910539
transform 1 0 12328 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1608910539
transform 1 0 11316 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 12420 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_139
timestamp 1608910539
transform 1 0 13892 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_135
timestamp 1608910539
transform 1 0 13524 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_131
timestamp 1608910539
transform 1 0 13156 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 13340 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 14260 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 14076 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_7_161
timestamp 1608910539
transform 1 0 15916 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_157
timestamp 1608910539
transform 1 0 15548 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_162
timestamp 1608910539
transform 1 0 16008 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_157
timestamp 1608910539
transform 1 0 15548 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_149
timestamp 1608910539
transform 1 0 14812 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 15732 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608910539
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 16008 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1608910539
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_182
timestamp 1608910539
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_178
timestamp 1608910539
transform 1 0 17480 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_184
timestamp 1608910539
transform 1 0 18032 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608910539
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1608910539
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 16560 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1608910539
transform 1 0 19964 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1608910539
transform 1 0 18860 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_208
timestamp 1608910539
transform 1 0 20240 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_196
timestamp 1608910539
transform 1 0 19136 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1608910539
transform 1 0 21068 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_215
timestamp 1608910539
transform 1 0 20884 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608910539
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608910539
transform -1 0 21896 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608910539
transform -1 0 21896 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_18
timestamp 1608910539
transform 1 0 2760 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_7
timestamp 1608910539
transform 1 0 1748 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1608910539
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 1564 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608910539
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1608910539
transform 1 0 1932 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1608910539
transform 1 0 2944 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1608910539
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608910539
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 4048 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1608910539
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_52
timestamp 1608910539
transform 1 0 5888 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_48
timestamp 1608910539
transform 1 0 5520 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 6072 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 5704 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1608910539
transform 1 0 8648 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1608910539
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 8464 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_102
timestamp 1608910539
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_99
timestamp 1608910539
transform 1 0 10212 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_93
timestamp 1608910539
transform 1 0 9660 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1608910539
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_87
timestamp 1608910539
transform 1 0 9108 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 10304 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 10672 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608910539
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1608910539
transform 1 0 8832 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_122
timestamp 1608910539
transform 1 0 12328 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_118
timestamp 1608910539
transform 1 0 11960 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_107
timestamp 1608910539
transform 1 0 10948 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 12144 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 12512 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l2_in_0_
timestamp 1608910539
transform 1 0 11132 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_140
timestamp 1608910539
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_127
timestamp 1608910539
transform 1 0 12788 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_0_
timestamp 1608910539
transform 1 0 14168 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l1_in_0_
timestamp 1608910539
transform 1 0 13156 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_164
timestamp 1608910539
transform 1 0 16192 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_160
timestamp 1608910539
transform 1 0 15824 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1608910539
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608910539
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1608910539
transform 1 0 16284 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 15272 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_183
timestamp 1608910539
transform 1 0 17940 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_179
timestamp 1608910539
transform 1 0 17572 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_174
timestamp 1608910539
transform 1 0 17112 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 17756 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _066_
timestamp 1608910539
transform 1 0 17296 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_207
timestamp 1608910539
transform 1 0 20148 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_195
timestamp 1608910539
transform 1 0 19044 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_215
timestamp 1608910539
transform 1 0 20884 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1608910539
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608910539
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608910539
transform -1 0 21896 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1608910539
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608910539
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 1748 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_39
timestamp 1608910539
transform 1 0 4692 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_31
timestamp 1608910539
transform 1 0 3956 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_27
timestamp 1608910539
transform 1 0 3588 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_23
timestamp 1608910539
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 3772 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 4876 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_62
timestamp 1608910539
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1608910539
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_48
timestamp 1608910539
transform 1 0 5520 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_43
timestamp 1608910539
transform 1 0 5060 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 5244 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608910539
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1608910539
transform 1 0 5704 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_67
timestamp 1608910539
transform 1 0 7268 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 6992 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 7636 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_87
timestamp 1608910539
transform 1 0 9108 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 9292 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1608910539
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_116
timestamp 1608910539
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_105
timestamp 1608910539
transform 1 0 10764 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608910539
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10948 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1608910539
transform 1 0 12420 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_138
timestamp 1608910539
transform 1 0 13800 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_135
timestamp 1608910539
transform 1 0 13524 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_131
timestamp 1608910539
transform 1 0 13156 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_126
timestamp 1608910539
transform 1 0 12696 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 12972 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 14076 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_9_157
timestamp 1608910539
transform 1 0 15548 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 16100 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1608910539
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_179
timestamp 1608910539
transform 1 0 17572 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608910539
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1608910539
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1608910539
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_220
timestamp 1608910539
transform 1 0 21344 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608910539
transform -1 0 21896 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_18
timestamp 1608910539
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_7
timestamp 1608910539
transform 1 0 1748 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1608910539
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608910539
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1608910539
transform 1 0 1932 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1608910539
transform 1 0 2944 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_34
timestamp 1608910539
transform 1 0 4232 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1608910539
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608910539
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1608910539
transform 1 0 4416 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_62
timestamp 1608910539
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_56
timestamp 1608910539
transform 1 0 6256 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_45
timestamp 1608910539
transform 1 0 5244 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6624 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1608910539
transform 1 0 5428 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_10_77
timestamp 1608910539
transform 1 0 8188 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_66
timestamp 1608910539
transform 1 0 7176 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 6992 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8464 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_0_
timestamp 1608910539
transform 1 0 7360 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_101
timestamp 1608910539
transform 1 0 10396 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_93
timestamp 1608910539
transform 1 0 9660 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_89
timestamp 1608910539
transform 1 0 9292 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608910539
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 10488 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_118
timestamp 1608910539
transform 1 0 11960 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 12144 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_136
timestamp 1608910539
transform 1 0 13616 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l1_in_0_
timestamp 1608910539
transform 1 0 13800 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_160
timestamp 1608910539
transform 1 0 15824 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1608910539
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_147
timestamp 1608910539
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608910539
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 15272 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_186
timestamp 1608910539
transform 1 0 18216 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_174
timestamp 1608910539
transform 1 0 17112 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 16560 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_198
timestamp 1608910539
transform 1 0 19320 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_215
timestamp 1608910539
transform 1 0 20884 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_210
timestamp 1608910539
transform 1 0 20424 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608910539
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608910539
transform -1 0 21896 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_7
timestamp 1608910539
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1608910539
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 1564 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608910539
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 1932 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_11_33
timestamp 1608910539
transform 1 0 4140 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_25
timestamp 1608910539
transform 1 0 3404 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 4232 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_62
timestamp 1608910539
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_55
timestamp 1608910539
transform 1 0 6164 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_50
timestamp 1608910539
transform 1 0 5704 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608910539
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1608910539
transform 1 0 5888 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_80
timestamp 1608910539
transform 1 0 8464 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 6992 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_11_104
timestamp 1608910539
transform 1 0 10672 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_101
timestamp 1608910539
transform 1 0 10396 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_93
timestamp 1608910539
transform 1 0 9660 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_88
timestamp 1608910539
transform 1 0 9200 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 10488 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1608910539
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_117
timestamp 1608910539
transform 1 0 11868 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_112
timestamp 1608910539
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 11592 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608910539
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _068_
timestamp 1608910539
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_126
timestamp 1608910539
transform 1 0 12696 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 13432 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_11_155
timestamp 1608910539
transform 1 0 15364 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_150
timestamp 1608910539
transform 1 0 14904 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _067_
timestamp 1608910539
transform 1 0 15088 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1608910539
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_177
timestamp 1608910539
transform 1 0 17388 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_167
timestamp 1608910539
transform 1 0 16468 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608910539
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 16836 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1608910539
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1608910539
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_220
timestamp 1608910539
transform 1 0 21344 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608910539
transform -1 0 21896 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_11
timestamp 1608910539
transform 1 0 2116 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3
timestamp 1608910539
transform 1 0 1380 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608910539
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1608910539
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_35
timestamp 1608910539
transform 1 0 4324 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_32
timestamp 1608910539
transform 1 0 4048 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_23
timestamp 1608910539
transform 1 0 3220 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 4140 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608910539
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1608910539
transform 1 0 4508 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_46
timestamp 1608910539
transform 1 0 5336 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 5520 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_81
timestamp 1608910539
transform 1 0 8556 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_69
timestamp 1608910539
transform 1 0 7452 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_64
timestamp 1608910539
transform 1 0 6992 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 8740 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 7176 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1608910539
transform 1 0 7728 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_12_102
timestamp 1608910539
transform 1 0 10488 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1608910539
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_85
timestamp 1608910539
transform 1 0 8924 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608910539
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1608910539
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_111
timestamp 1608910539
transform 1 0 11316 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_107
timestamp 1608910539
transform 1 0 10948 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 11132 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 10764 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 11684 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_139
timestamp 1608910539
transform 1 0 13892 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_131
timestamp 1608910539
transform 1 0 13156 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l2_in_0_
timestamp 1608910539
transform 1 0 14076 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1608910539
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1608910539
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_150
timestamp 1608910539
transform 1 0 14904 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608910539
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1608910539
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1608910539
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_190
timestamp 1608910539
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_215
timestamp 1608910539
transform 1 0 20884 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608910539
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608910539
transform -1 0 21896 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_11
timestamp 1608910539
transform 1 0 2116 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3
timestamp 1608910539
transform 1 0 1380 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1608910539
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 1932 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608910539
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608910539
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1608910539
transform 1 0 2300 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 1564 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1608910539
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_22
timestamp 1608910539
transform 1 0 3128 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_21
timestamp 1608910539
transform 1 0 3036 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1608910539
transform 1 0 3220 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1608910539
transform 1 0 3312 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_36
timestamp 1608910539
transform 1 0 4416 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_32
timestamp 1608910539
transform 1 0 4048 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_36
timestamp 1608910539
transform 1 0 4416 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_32
timestamp 1608910539
transform 1 0 4048 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608910539
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1608910539
transform 1 0 4508 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1608910539
transform 1 0 4600 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1608910539
transform 1 0 4140 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_47
timestamp 1608910539
transform 1 0 5428 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_50
timestamp 1608910539
transform 1 0 5704 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_46
timestamp 1608910539
transform 1 0 5336 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 5888 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1608910539
transform 1 0 5612 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_62
timestamp 1608910539
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_58
timestamp 1608910539
transform 1 0 6440 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_60
timestamp 1608910539
transform 1 0 6624 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_54
timestamp 1608910539
transform 1 0 6072 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 6624 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608910539
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 6808 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_14_77
timestamp 1608910539
transform 1 0 8188 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_66
timestamp 1608910539
transform 1 0 7176 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_83
timestamp 1608910539
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_78
timestamp 1608910539
transform 1 0 8280 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1608910539
transform 1 0 7360 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1608910539
transform 1 0 8372 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1608910539
transform 1 0 8464 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_102
timestamp 1608910539
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_88
timestamp 1608910539
transform 1 0 9200 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_87
timestamp 1608910539
transform 1 0 9108 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 10672 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1608910539
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1608910539
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9292 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_14_125
timestamp 1608910539
transform 1 0 12604 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_107
timestamp 1608910539
transform 1 0 10948 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_116
timestamp 1608910539
transform 1 0 11776 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_105
timestamp 1608910539
transform 1 0 10764 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608910539
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_29.mux_l2_in_0_
timestamp 1608910539
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_29.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10948 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 11132 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_14_137
timestamp 1608910539
transform 1 0 13708 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_132
timestamp 1608910539
transform 1 0 13248 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 13800 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_14_166
timestamp 1608910539
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_154
timestamp 1608910539
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_149
timestamp 1608910539
transform 1 0 14812 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_166
timestamp 1608910539
transform 1 0 16376 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_154
timestamp 1608910539
transform 1 0 15272 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1608910539
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_178
timestamp 1608910539
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1608910539
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_182
timestamp 1608910539
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_178
timestamp 1608910539
transform 1 0 17480 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608910539
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_202
timestamp 1608910539
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_190
timestamp 1608910539
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1608910539
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1608910539
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_215
timestamp 1608910539
transform 1 0 20884 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_220
timestamp 1608910539
transform 1 0 21344 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1608910539
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608910539
transform -1 0 21896 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608910539
transform -1 0 21896 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1608910539
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608910539
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 1656 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_30
timestamp 1608910539
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_22
timestamp 1608910539
transform 1 0 3128 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 3680 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 4048 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_62
timestamp 1608910539
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1608910539
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_48
timestamp 1608910539
transform 1 0 5520 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1608910539
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1608910539
transform 1 0 5704 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_15_82
timestamp 1608910539
transform 1 0 8648 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_77
timestamp 1608910539
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_66
timestamp 1608910539
transform 1 0 7176 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6992 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 8372 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l1_in_0_
timestamp 1608910539
transform 1 0 7360 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_98
timestamp 1608910539
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_94
timestamp 1608910539
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 10304 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8924 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_15_125
timestamp 1608910539
transform 1 0 12604 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1608910539
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_mem_bottom_track_1.prog_clk_A
timestamp 1608910539
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1608910539
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_143
timestamp 1608910539
transform 1 0 14260 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_131
timestamp 1608910539
transform 1 0 13156 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 12880 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_155
timestamp 1608910539
transform 1 0 15364 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_184
timestamp 1608910539
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_179
timestamp 1608910539
transform 1 0 17572 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_167
timestamp 1608910539
transform 1 0 16468 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1608910539
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1608910539
transform 1 0 18308 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_207
timestamp 1608910539
transform 1 0 20148 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_195
timestamp 1608910539
transform 1 0 19044 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_191
timestamp 1608910539
transform 1 0 18676 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1608910539
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_219
timestamp 1608910539
transform 1 0 21252 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608910539
transform -1 0 21896 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_16
timestamp 1608910539
transform 1 0 2576 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_11
timestamp 1608910539
transform 1 0 2116 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3
timestamp 1608910539
transform 1 0 1380 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 1932 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608910539
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1608910539
transform 1 0 2760 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1608910539
transform 1 0 2300 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_34
timestamp 1608910539
transform 1 0 4232 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1608910539
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1608910539
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4600 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_16_54
timestamp 1608910539
transform 1 0 6072 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 6348 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_81
timestamp 1608910539
transform 1 0 8556 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_63
timestamp 1608910539
transform 1 0 6900 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 7084 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1608910539
transform 1 0 8740 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1608910539
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_86
timestamp 1608910539
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1608910539
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9660 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_16_114
timestamp 1608910539
transform 1 0 11592 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_109
timestamp 1608910539
transform 1 0 11132 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 11316 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_138
timestamp 1608910539
transform 1 0 13800 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_126
timestamp 1608910539
transform 1 0 12696 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_166
timestamp 1608910539
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_154
timestamp 1608910539
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_150
timestamp 1608910539
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1608910539
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_178
timestamp 1608910539
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_200
timestamp 1608910539
transform 1 0 19504 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_196
timestamp 1608910539
transform 1 0 19136 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_190
timestamp 1608910539
transform 1 0 18584 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1608910539
transform 1 0 19320 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1608910539
transform 1 0 18768 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_215
timestamp 1608910539
transform 1 0 20884 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_212
timestamp 1608910539
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1608910539
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608910539
transform -1 0 21896 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_19
timestamp 1608910539
transform 1 0 2852 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_8
timestamp 1608910539
transform 1 0 1840 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_3
timestamp 1608910539
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 1656 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608910539
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1608910539
transform 1 0 2024 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_37
timestamp 1608910539
transform 1 0 4508 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 3036 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1608910539
transform 1 0 4692 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_62
timestamp 1608910539
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_60
timestamp 1608910539
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_54
timestamp 1608910539
transform 1 0 6072 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_42
timestamp 1608910539
transform 1 0 4968 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1608910539
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_73
timestamp 1608910539
transform 1 0 7820 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l2_in_0_
timestamp 1608910539
transform 1 0 6992 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 8188 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_17_93
timestamp 1608910539
transform 1 0 9660 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1608910539
transform 1 0 9936 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_17_116
timestamp 1608910539
transform 1 0 11776 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_105
timestamp 1608910539
transform 1 0 10764 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1608910539
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1608910539
transform 1 0 10948 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1608910539
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_138
timestamp 1608910539
transform 1 0 13800 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_126
timestamp 1608910539
transform 1 0 12696 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_162
timestamp 1608910539
transform 1 0 16008 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_150
timestamp 1608910539
transform 1 0 14904 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1608910539
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_182
timestamp 1608910539
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_174
timestamp 1608910539
transform 1 0 17112 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1608910539
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_205
timestamp 1608910539
transform 1 0 19964 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_201
timestamp 1608910539
transform 1 0 19596 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_196
timestamp 1608910539
transform 1 0 19136 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1608910539
transform 1 0 19780 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1608910539
transform 1 0 19228 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1608910539
transform 1 0 21068 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608910539
transform -1 0 21896 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_7
timestamp 1608910539
transform 1 0 1748 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608910539
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 1932 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1608910539
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_41
timestamp 1608910539
transform 1 0 4876 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_25
timestamp 1608910539
transform 1 0 3404 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1608910539
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1608910539
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_18_59
timestamp 1608910539
transform 1 0 6532 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 6808 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 5060 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_18_78
timestamp 1608910539
transform 1 0 8280 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_93
timestamp 1608910539
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1608910539
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_86
timestamp 1608910539
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1608910539
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 9844 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_18_123
timestamp 1608910539
transform 1 0 12420 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_111
timestamp 1608910539
transform 1 0 11316 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_135
timestamp 1608910539
transform 1 0 13524 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_166
timestamp 1608910539
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_154
timestamp 1608910539
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_147
timestamp 1608910539
transform 1 0 14628 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1608910539
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_178
timestamp 1608910539
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_206
timestamp 1608910539
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_190
timestamp 1608910539
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1608910539
transform 1 0 20240 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1608910539
transform 1 0 19688 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_215
timestamp 1608910539
transform 1 0 20884 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_210
timestamp 1608910539
transform 1 0 20424 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1608910539
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608910539
transform -1 0 21896 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_7
timestamp 1608910539
transform 1 0 1748 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1608910539
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1608910539
transform 1 0 1380 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608910539
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608910539
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1840 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_14
timestamp 1608910539
transform 1 0 2392 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_11
timestamp 1608910539
transform 1 0 2116 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1608910539
transform 1 0 2208 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2576 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_20_28
timestamp 1608910539
transform 1 0 3680 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_22
timestamp 1608910539
transform 1 0 3128 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_29
timestamp 1608910539
transform 1 0 3772 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_21
timestamp 1608910539
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1608910539
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 3220 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1608910539
transform 1 0 3312 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_40
timestamp 1608910539
transform 1 0 4784 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_35
timestamp 1608910539
transform 1 0 4324 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_32
timestamp 1608910539
transform 1 0 4048 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 4140 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1608910539
transform 1 0 4508 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4140 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_19_49
timestamp 1608910539
transform 1 0 5612 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 5796 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1608910539
transform 1 0 5060 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_20_56
timestamp 1608910539
transform 1 0 6256 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_52
timestamp 1608910539
transform 1 0 5888 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1608910539
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_54
timestamp 1608910539
transform 1 0 6072 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 6072 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1608910539
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_62
timestamp 1608910539
transform 1 0 6808 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_80
timestamp 1608910539
transform 1 0 8464 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_78
timestamp 1608910539
transform 1 0 8280 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_67
timestamp 1608910539
transform 1 0 7268 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 6992 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8464 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1608910539
transform 1 0 7452 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 6992 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1608910539
transform 1 0 8648 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_93
timestamp 1608910539
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_90
timestamp 1608910539
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1608910539
transform 1 0 8924 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_89
timestamp 1608910539
transform 1 0 9292 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1608910539
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1608910539
transform 1 0 9568 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1608910539
transform 1 0 9108 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_101
timestamp 1608910539
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1608910539
transform 1 0 10580 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9936 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_20_116
timestamp 1608910539
transform 1 0 11776 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_112
timestamp 1608910539
transform 1 0 11408 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1608910539
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_116
timestamp 1608910539
transform 1 0 11776 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_112
timestamp 1608910539
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 11592 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1608910539
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_140
timestamp 1608910539
transform 1 0 13984 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_128
timestamp 1608910539
transform 1 0 12880 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1608910539
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_166
timestamp 1608910539
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1608910539
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1608910539
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_159
timestamp 1608910539
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_147
timestamp 1608910539
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1608910539
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1608910539
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1608910539
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_171
timestamp 1608910539
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1608910539
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_202
timestamp 1608910539
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_190
timestamp 1608910539
transform 1 0 18584 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1608910539
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1608910539
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_215
timestamp 1608910539
transform 1 0 20884 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_220
timestamp 1608910539
transform 1 0 21344 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1608910539
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608910539
transform -1 0 21896 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608910539
transform -1 0 21896 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_19
timestamp 1608910539
transform 1 0 2852 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_11
timestamp 1608910539
transform 1 0 2116 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1608910539
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608910539
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1564 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2300 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_25
timestamp 1608910539
transform 1 0 3404 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 3956 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1608910539
transform 1 0 3036 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_62
timestamp 1608910539
transform 1 0 6808 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_21_58
timestamp 1608910539
transform 1 0 6440 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_47
timestamp 1608910539
transform 1 0 5428 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1608910539
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1608910539
transform 1 0 5612 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_81
timestamp 1608910539
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_70
timestamp 1608910539
transform 1 0 7544 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 7360 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 8740 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1608910539
transform 1 0 7728 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_90
timestamp 1608910539
transform 1 0 9384 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_86
timestamp 1608910539
transform 1 0 9016 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9200 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 9568 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1608910539
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_119
timestamp 1608910539
transform 1 0 12052 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_108
timestamp 1608910539
transform 1 0 11040 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1608910539
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1608910539
transform 1 0 11224 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1608910539
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_159
timestamp 1608910539
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_147
timestamp 1608910539
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1608910539
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_171
timestamp 1608910539
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1608910539
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1608910539
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1608910539
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_220
timestamp 1608910539
transform 1 0 21344 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608910539
transform -1 0 21896 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_19
timestamp 1608910539
transform 1 0 2852 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_11
timestamp 1608910539
transform 1 0 2116 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1608910539
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608910539
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2300 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1608910539
transform 1 0 1748 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_32
timestamp 1608910539
transform 1 0 4048 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_25
timestamp 1608910539
transform 1 0 3404 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1608910539
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4416 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1608910539
transform 1 0 3036 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_60
timestamp 1608910539
transform 1 0 6624 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_52
timestamp 1608910539
transform 1 0 5888 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_79
timestamp 1608910539
transform 1 0 8372 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 6900 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_93
timestamp 1608910539
transform 1 0 9660 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1608910539
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1608910539
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 10028 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_22_117
timestamp 1608910539
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_113
timestamp 1608910539
transform 1 0 11500 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 11684 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1608910539
transform 1 0 14076 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_129
timestamp 1608910539
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1608910539
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1608910539
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1608910539
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1608910539
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_202
timestamp 1608910539
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1608910539
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_215
timestamp 1608910539
transform 1 0 20884 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1608910539
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608910539
transform -1 0 21896 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_18
timestamp 1608910539
transform 1 0 2760 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_10
timestamp 1608910539
transform 1 0 2024 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_3
timestamp 1608910539
transform 1 0 1380 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1608910539
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1608910539
transform 1 0 2944 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2208 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1608910539
transform 1 0 1656 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_39
timestamp 1608910539
transform 1 0 4692 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_34
timestamp 1608910539
transform 1 0 4232 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_29
timestamp 1608910539
transform 1 0 3772 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 4508 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 4876 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1608910539
transform 1 0 3956 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1608910539
transform 1 0 6348 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1608910539
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1608910539
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_23_80
timestamp 1608910539
transform 1 0 8464 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_76
timestamp 1608910539
transform 1 0 8096 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_71
timestamp 1608910539
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8280 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1608910539
transform 1 0 7820 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_100
timestamp 1608910539
transform 1 0 10304 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_95
timestamp 1608910539
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1608910539
transform 1 0 9016 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1608910539
transform 1 0 10028 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1608910539
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1608910539
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_112
timestamp 1608910539
transform 1 0 11408 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1608910539
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1608910539
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_159
timestamp 1608910539
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1608910539
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1608910539
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_171
timestamp 1608910539
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1608910539
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1608910539
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1608910539
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_220
timestamp 1608910539
transform 1 0 21344 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1608910539
transform -1 0 21896 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_16
timestamp 1608910539
transform 1 0 2576 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_8
timestamp 1608910539
transform 1 0 1840 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 1608910539
transform 1 0 1380 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1608910539
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2024 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1608910539
transform 1 0 1472 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_41
timestamp 1608910539
transform 1 0 4876 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1608910539
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_24
timestamp 1608910539
transform 1 0 3312 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1608910539
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1608910539
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_24_58
timestamp 1608910539
transform 1 0 6440 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_54
timestamp 1608910539
transform 1 0 6072 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1608910539
transform 1 0 5244 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 6532 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_24_79
timestamp 1608910539
transform 1 0 8372 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_75
timestamp 1608910539
transform 1 0 8004 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8464 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_24_99
timestamp 1608910539
transform 1 0 10212 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_95
timestamp 1608910539
transform 1 0 9844 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_89
timestamp 1608910539
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 10028 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1608910539
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_123
timestamp 1608910539
transform 1 0 12420 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_111
timestamp 1608910539
transform 1 0 11316 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_135
timestamp 1608910539
transform 1 0 13524 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1608910539
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1608910539
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_147
timestamp 1608910539
transform 1 0 14628 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1608910539
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1608910539
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_202
timestamp 1608910539
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1608910539
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_215
timestamp 1608910539
transform 1 0 20884 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1608910539
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1608910539
transform -1 0 21896 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_17
timestamp 1608910539
transform 1 0 2668 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_11
timestamp 1608910539
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1608910539
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1608910539
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 2944 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1608910539
transform 1 0 2300 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1608910539
transform 1 0 1748 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_41
timestamp 1608910539
transform 1 0 4876 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_36
timestamp 1608910539
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1608910539
transform 1 0 4600 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1608910539
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_49
timestamp 1608910539
transform 1 0 5612 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_45
timestamp 1608910539
transform 1 0 5244 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 5060 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 6808 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1608910539
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1608910539
transform 1 0 5704 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_79
timestamp 1608910539
transform 1 0 8372 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_75
timestamp 1608910539
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_64
timestamp 1608910539
transform 1 0 6992 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1608910539
transform 1 0 7176 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 8740 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_25_104
timestamp 1608910539
transform 1 0 10672 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_99
timestamp 1608910539
transform 1 0 10212 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 10488 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1608910539
transform 1 0 12604 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_120
timestamp 1608910539
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_109
timestamp 1608910539
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 10948 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 12420 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1608910539
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1608910539
transform 1 0 11316 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1608910539
transform 1 0 13708 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_161
timestamp 1608910539
transform 1 0 15916 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1608910539
transform 1 0 14812 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1608910539
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_181
timestamp 1608910539
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_173
timestamp 1608910539
transform 1 0 17020 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1608910539
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1608910539
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1608910539
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_220
timestamp 1608910539
transform 1 0 21344 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1608910539
transform -1 0 21896 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1608910539
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_9
timestamp 1608910539
transform 1 0 1932 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_3
timestamp 1608910539
transform 1 0 1380 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1608910539
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1608910539
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1608910539
transform 1 0 1748 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_11
timestamp 1608910539
transform 1 0 2116 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_16
timestamp 1608910539
transform 1 0 2576 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2024 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2392 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_20
timestamp 1608910539
transform 1 0 2944 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1608910539
transform 1 0 2944 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_27_32
timestamp 1608910539
transform 1 0 4048 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_28
timestamp 1608910539
transform 1 0 3680 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1608910539
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1608910539
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 3128 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4140 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 4048 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_27_58
timestamp 1608910539
transform 1 0 6440 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1608910539
transform 1 0 6072 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_49
timestamp 1608910539
transform 1 0 5612 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_48
timestamp 1608910539
transform 1 0 5520 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6256 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1608910539
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1608910539
transform 1 0 6808 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 5888 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1608910539
transform 1 0 5796 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_71
timestamp 1608910539
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_72
timestamp 1608910539
transform 1 0 7728 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_68
timestamp 1608910539
transform 1 0 7360 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 7544 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_80
timestamp 1608910539
transform 1 0 8464 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_75
timestamp 1608910539
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1608910539
transform 1 0 8188 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 8648 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 7912 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_27_98
timestamp 1608910539
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_102
timestamp 1608910539
transform 1 0 10488 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_90
timestamp 1608910539
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1608910539
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1608910539
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 10672 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 10304 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_27_116
timestamp 1608910539
transform 1 0 11776 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_120
timestamp 1608910539
transform 1 0 12144 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1608910539
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 12328 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1608910539
transform 1 0 12420 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_138
timestamp 1608910539
transform 1 0 13800 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_126
timestamp 1608910539
transform 1 0 12696 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_138
timestamp 1608910539
transform 1 0 13800 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_162
timestamp 1608910539
transform 1 0 16008 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_150
timestamp 1608910539
transform 1 0 14904 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1608910539
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1608910539
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_150
timestamp 1608910539
transform 1 0 14904 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1608910539
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1608910539
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_182
timestamp 1608910539
transform 1 0 17848 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_174
timestamp 1608910539
transform 1 0 17112 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1608910539
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1608910539
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1608910539
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1608910539
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_202
timestamp 1608910539
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_190
timestamp 1608910539
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_220
timestamp 1608910539
transform 1 0 21344 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_215
timestamp 1608910539
transform 1 0 20884 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1608910539
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1608910539
transform -1 0 21896 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1608910539
transform -1 0 21896 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_18
timestamp 1608910539
transform 1 0 2760 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_10
timestamp 1608910539
transform 1 0 2024 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_3
timestamp 1608910539
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1608910539
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2944 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2208 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1608910539
transform 1 0 1656 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_40
timestamp 1608910539
transform 1 0 4784 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_32
timestamp 1608910539
transform 1 0 4048 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_30
timestamp 1608910539
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_26
timestamp 1608910539
transform 1 0 3496 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1608910539
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_59
timestamp 1608910539
transform 1 0 6532 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 5060 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_28_71
timestamp 1608910539
transform 1 0 7636 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8004 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_102
timestamp 1608910539
transform 1 0 10488 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_84
timestamp 1608910539
transform 1 0 8832 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1608910539
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1608910539
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1608910539
transform 1 0 10672 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1608910539
transform 1 0 12236 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_111
timestamp 1608910539
transform 1 0 11316 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_107
timestamp 1608910539
transform 1 0 10948 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1608910539
transform 1 0 11408 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_28_145
timestamp 1608910539
transform 1 0 14444 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_133
timestamp 1608910539
transform 1 0 13340 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1608910539
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1608910539
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1608910539
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1608910539
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1608910539
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1608910539
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_215
timestamp 1608910539
transform 1 0 20884 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1608910539
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1608910539
transform -1 0 21896 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_15
timestamp 1608910539
transform 1 0 2484 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_11
timestamp 1608910539
transform 1 0 2116 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1608910539
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1608910539
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2576 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1608910539
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_34
timestamp 1608910539
transform 1 0 4232 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_22
timestamp 1608910539
transform 1 0 3128 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1608910539
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_58
timestamp 1608910539
transform 1 0 6440 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_46
timestamp 1608910539
transform 1 0 5336 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1608910539
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1608910539
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_98
timestamp 1608910539
transform 1 0 10120 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_86
timestamp 1608910539
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1608910539
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1608910539
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_112
timestamp 1608910539
transform 1 0 11408 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1608910539
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 10856 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1608910539
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_159
timestamp 1608910539
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_147
timestamp 1608910539
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1608910539
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1608910539
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1608910539
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1608910539
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1608910539
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_220
timestamp 1608910539
transform 1 0 21344 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1608910539
transform -1 0 21896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_19
timestamp 1608910539
transform 1 0 2852 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_11
timestamp 1608910539
transform 1 0 2116 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1608910539
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1608910539
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2300 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1608910539
transform 1 0 1748 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1608910539
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1608910539
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1608910539
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 3036 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1608910539
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1608910539
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1608910539
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1608910539
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_101
timestamp 1608910539
transform 1 0 10396 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_93
timestamp 1608910539
transform 1 0 9660 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1608910539
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1608910539
transform 1 0 10580 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_119
timestamp 1608910539
transform 1 0 12052 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_107
timestamp 1608910539
transform 1 0 10948 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_143
timestamp 1608910539
transform 1 0 14260 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_131
timestamp 1608910539
transform 1 0 13156 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1608910539
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1608910539
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_151
timestamp 1608910539
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1608910539
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_178
timestamp 1608910539
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_202
timestamp 1608910539
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_190
timestamp 1608910539
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_215
timestamp 1608910539
transform 1 0 20884 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1608910539
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1608910539
transform -1 0 21896 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_19
timestamp 1608910539
transform 1 0 2852 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_11
timestamp 1608910539
transform 1 0 2116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1608910539
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1608910539
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2300 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1608910539
transform 1 0 1748 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1608910539
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1608910539
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 3036 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1608910539
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1608910539
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1608910539
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1608910539
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1608910539
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1608910539
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1608910539
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1608910539
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1608910539
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1608910539
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1608910539
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_159
timestamp 1608910539
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_147
timestamp 1608910539
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1608910539
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_171
timestamp 1608910539
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1608910539
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1608910539
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1608910539
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_220
timestamp 1608910539
transform 1 0 21344 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1608910539
transform -1 0 21896 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_18
timestamp 1608910539
transform 1 0 2760 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_12
timestamp 1608910539
transform 1 0 2208 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_7
timestamp 1608910539
transform 1 0 1748 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1608910539
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1608910539
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1608910539
transform 1 0 2944 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1608910539
transform 1 0 2392 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1608910539
transform 1 0 1840 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1608910539
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_30
timestamp 1608910539
transform 1 0 3864 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_24
timestamp 1608910539
transform 1 0 3312 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1608910539
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1608910539
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1608910539
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_80
timestamp 1608910539
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1608910539
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1608910539
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1608910539
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_117
timestamp 1608910539
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1608910539
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1608910539
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_129
timestamp 1608910539
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_166
timestamp 1608910539
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_154
timestamp 1608910539
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1608910539
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_178
timestamp 1608910539
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_202
timestamp 1608910539
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_190
timestamp 1608910539
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_215
timestamp 1608910539
transform 1 0 20884 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1608910539
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1608910539
transform -1 0 21896 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_17
timestamp 1608910539
transform 1 0 2668 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_11
timestamp 1608910539
transform 1 0 2116 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1608910539
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1608910539
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1608910539
transform 1 0 2300 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1608910539
transform 1 0 1748 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_32
timestamp 1608910539
transform 1 0 4048 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_29
timestamp 1608910539
transform 1 0 3772 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1608910539
transform 1 0 3956 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_56
timestamp 1608910539
transform 1 0 6256 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_44
timestamp 1608910539
transform 1 0 5152 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1608910539
transform 1 0 6808 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_75
timestamp 1608910539
transform 1 0 8004 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_63
timestamp 1608910539
transform 1 0 6900 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_94
timestamp 1608910539
transform 1 0 9752 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_87
timestamp 1608910539
transform 1 0 9108 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1608910539
transform 1 0 9660 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_125
timestamp 1608910539
transform 1 0 12604 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_118
timestamp 1608910539
transform 1 0 11960 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_106
timestamp 1608910539
transform 1 0 10856 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1608910539
transform 1 0 12512 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_137
timestamp 1608910539
transform 1 0 13708 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_156
timestamp 1608910539
transform 1 0 15456 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_149
timestamp 1608910539
transform 1 0 14812 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1608910539
transform 1 0 15364 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_187
timestamp 1608910539
transform 1 0 18308 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_180
timestamp 1608910539
transform 1 0 17664 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_168
timestamp 1608910539
transform 1 0 16560 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1608910539
transform 1 0 18216 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_199
timestamp 1608910539
transform 1 0 19412 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_222
timestamp 1608910539
transform 1 0 21528 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_218
timestamp 1608910539
transform 1 0 21160 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_211
timestamp 1608910539
transform 1 0 20516 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1608910539
transform 1 0 21068 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1608910539
transform -1 0 21896 0 1 20128
box -38 -48 314 592
<< labels >>
rlabel metal2 s 21822 0 21878 800 6 SC_IN_BOT
port 0 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 SC_OUT_BOT
port 1 nsew signal tristate
rlabel metal2 s 202 0 258 800 6 bottom_left_grid_pin_42_
port 2 nsew signal input
rlabel metal2 s 570 0 626 800 6 bottom_left_grid_pin_43_
port 3 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 bottom_left_grid_pin_44_
port 4 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 bottom_left_grid_pin_45_
port 5 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 bottom_left_grid_pin_46_
port 6 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 bottom_left_grid_pin_47_
port 7 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 bottom_left_grid_pin_48_
port 8 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 bottom_left_grid_pin_49_
port 9 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 bottom_right_grid_pin_1_
port 10 nsew signal input
rlabel metal3 s 22200 5720 23000 5840 6 ccff_head
port 11 nsew signal input
rlabel metal3 s 22200 17144 23000 17264 6 ccff_tail
port 12 nsew signal tristate
rlabel metal3 s 0 3816 800 3936 6 chanx_left_in[0]
port 13 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 chanx_left_in[10]
port 14 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 chanx_left_in[11]
port 15 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 chanx_left_in[12]
port 16 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 chanx_left_in[13]
port 17 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 chanx_left_in[14]
port 18 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 chanx_left_in[15]
port 19 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[16]
port 20 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 chanx_left_in[17]
port 21 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[18]
port 22 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 chanx_left_in[19]
port 23 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 chanx_left_in[1]
port 24 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 chanx_left_in[2]
port 25 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 chanx_left_in[3]
port 26 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 chanx_left_in[4]
port 27 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 chanx_left_in[5]
port 28 nsew signal input
rlabel metal3 s 0 6672 800 6792 6 chanx_left_in[6]
port 29 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 chanx_left_in[7]
port 30 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 chanx_left_in[8]
port 31 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 chanx_left_in[9]
port 32 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 chanx_left_out[0]
port 33 nsew signal tristate
rlabel metal3 s 0 17960 800 18080 6 chanx_left_out[10]
port 34 nsew signal tristate
rlabel metal3 s 0 18368 800 18488 6 chanx_left_out[11]
port 35 nsew signal tristate
rlabel metal3 s 0 18776 800 18896 6 chanx_left_out[12]
port 36 nsew signal tristate
rlabel metal3 s 0 19320 800 19440 6 chanx_left_out[13]
port 37 nsew signal tristate
rlabel metal3 s 0 19728 800 19848 6 chanx_left_out[14]
port 38 nsew signal tristate
rlabel metal3 s 0 20272 800 20392 6 chanx_left_out[15]
port 39 nsew signal tristate
rlabel metal3 s 0 20680 800 20800 6 chanx_left_out[16]
port 40 nsew signal tristate
rlabel metal3 s 0 21224 800 21344 6 chanx_left_out[17]
port 41 nsew signal tristate
rlabel metal3 s 0 21632 800 21752 6 chanx_left_out[18]
port 42 nsew signal tristate
rlabel metal3 s 0 22176 800 22296 6 chanx_left_out[19]
port 43 nsew signal tristate
rlabel metal3 s 0 13744 800 13864 6 chanx_left_out[1]
port 44 nsew signal tristate
rlabel metal3 s 0 14152 800 14272 6 chanx_left_out[2]
port 45 nsew signal tristate
rlabel metal3 s 0 14560 800 14680 6 chanx_left_out[3]
port 46 nsew signal tristate
rlabel metal3 s 0 15104 800 15224 6 chanx_left_out[4]
port 47 nsew signal tristate
rlabel metal3 s 0 15512 800 15632 6 chanx_left_out[5]
port 48 nsew signal tristate
rlabel metal3 s 0 16056 800 16176 6 chanx_left_out[6]
port 49 nsew signal tristate
rlabel metal3 s 0 16464 800 16584 6 chanx_left_out[7]
port 50 nsew signal tristate
rlabel metal3 s 0 17008 800 17128 6 chanx_left_out[8]
port 51 nsew signal tristate
rlabel metal3 s 0 17416 800 17536 6 chanx_left_out[9]
port 52 nsew signal tristate
rlabel metal2 s 3698 0 3754 800 6 chany_bottom_in[0]
port 53 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 chany_bottom_in[10]
port 54 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 chany_bottom_in[11]
port 55 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 chany_bottom_in[12]
port 56 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 chany_bottom_in[13]
port 57 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 chany_bottom_in[14]
port 58 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 chany_bottom_in[15]
port 59 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 chany_bottom_in[16]
port 60 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 chany_bottom_in[17]
port 61 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 chany_bottom_in[18]
port 62 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 chany_bottom_in[19]
port 63 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 chany_bottom_in[1]
port 64 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 chany_bottom_in[2]
port 65 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 chany_bottom_in[3]
port 66 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 chany_bottom_in[4]
port 67 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 chany_bottom_in[5]
port 68 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 chany_bottom_in[6]
port 69 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 chany_bottom_in[7]
port 70 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 chany_bottom_in[8]
port 71 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 chany_bottom_in[9]
port 72 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 chany_bottom_out[0]
port 73 nsew signal tristate
rlabel metal2 s 16946 0 17002 800 6 chany_bottom_out[10]
port 74 nsew signal tristate
rlabel metal2 s 17406 0 17462 800 6 chany_bottom_out[11]
port 75 nsew signal tristate
rlabel metal2 s 17866 0 17922 800 6 chany_bottom_out[12]
port 76 nsew signal tristate
rlabel metal2 s 18326 0 18382 800 6 chany_bottom_out[13]
port 77 nsew signal tristate
rlabel metal2 s 18694 0 18750 800 6 chany_bottom_out[14]
port 78 nsew signal tristate
rlabel metal2 s 19154 0 19210 800 6 chany_bottom_out[15]
port 79 nsew signal tristate
rlabel metal2 s 19614 0 19670 800 6 chany_bottom_out[16]
port 80 nsew signal tristate
rlabel metal2 s 20074 0 20130 800 6 chany_bottom_out[17]
port 81 nsew signal tristate
rlabel metal2 s 20534 0 20590 800 6 chany_bottom_out[18]
port 82 nsew signal tristate
rlabel metal2 s 20902 0 20958 800 6 chany_bottom_out[19]
port 83 nsew signal tristate
rlabel metal2 s 12990 0 13046 800 6 chany_bottom_out[1]
port 84 nsew signal tristate
rlabel metal2 s 13450 0 13506 800 6 chany_bottom_out[2]
port 85 nsew signal tristate
rlabel metal2 s 13910 0 13966 800 6 chany_bottom_out[3]
port 86 nsew signal tristate
rlabel metal2 s 14278 0 14334 800 6 chany_bottom_out[4]
port 87 nsew signal tristate
rlabel metal2 s 14738 0 14794 800 6 chany_bottom_out[5]
port 88 nsew signal tristate
rlabel metal2 s 15198 0 15254 800 6 chany_bottom_out[6]
port 89 nsew signal tristate
rlabel metal2 s 15658 0 15714 800 6 chany_bottom_out[7]
port 90 nsew signal tristate
rlabel metal2 s 16118 0 16174 800 6 chany_bottom_out[8]
port 91 nsew signal tristate
rlabel metal2 s 16486 0 16542 800 6 chany_bottom_out[9]
port 92 nsew signal tristate
rlabel metal3 s 0 144 800 264 6 left_bottom_grid_pin_34_
port 93 nsew signal input
rlabel metal3 s 0 552 800 672 6 left_bottom_grid_pin_35_
port 94 nsew signal input
rlabel metal3 s 0 960 800 1080 6 left_bottom_grid_pin_36_
port 95 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 left_bottom_grid_pin_37_
port 96 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 left_bottom_grid_pin_38_
port 97 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 left_bottom_grid_pin_39_
port 98 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 left_bottom_grid_pin_40_
port 99 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 left_bottom_grid_pin_41_
port 100 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 left_top_grid_pin_1_
port 101 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 prog_clk_0_S_in
port 102 nsew signal input
rlabel metal4 s 18271 2128 18591 20720 6 VPWR
port 103 nsew power bidirectional
rlabel metal4 s 11340 2128 11660 20720 6 VPWR
port 104 nsew power bidirectional
rlabel metal4 s 4409 2128 4729 20720 6 VPWR
port 105 nsew power bidirectional
rlabel metal4 s 14805 2128 15125 20720 6 VGND
port 106 nsew ground bidirectional
rlabel metal4 s 7875 2128 8195 20720 6 VGND
port 107 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 23000 22704
<< end >>
