magic
tech EFS8A
magscale 1 2
timestamp 1604348395
<< locali >>
rect 45753 24735 45787 24905
rect 34529 16099 34563 16201
rect 40601 15895 40635 15997
rect 24961 9367 24995 9469
rect 27353 5219 27387 5321
rect 37933 2499 37967 2601
<< viali >>
rect 46949 45509 46983 45543
rect 46765 45373 46799 45407
rect 47317 45373 47351 45407
rect 46949 44489 46983 44523
rect 47409 44489 47443 44523
rect 46765 44285 46799 44319
rect 46949 41769 46983 41803
rect 46765 41633 46799 41667
rect 46765 40885 46799 40919
rect 46949 38505 46983 38539
rect 46765 38369 46799 38403
rect 46765 37621 46799 37655
rect 46949 35241 46983 35275
rect 46765 35105 46799 35139
rect 46765 34697 46799 34731
rect 46949 31977 46983 32011
rect 46765 31841 46799 31875
rect 42165 31637 42199 31671
rect 41981 31229 42015 31263
rect 42073 31229 42107 31263
rect 42340 31161 42374 31195
rect 43453 31093 43487 31127
rect 46765 31093 46799 31127
rect 44741 30889 44775 30923
rect 42073 30821 42107 30855
rect 42257 30821 42291 30855
rect 43628 30753 43662 30787
rect 46101 30753 46135 30787
rect 42349 30685 42383 30719
rect 43361 30685 43395 30719
rect 45845 30685 45879 30719
rect 47225 30617 47259 30651
rect 41797 30549 41831 30583
rect 45753 30549 45787 30583
rect 41797 30345 41831 30379
rect 42073 30345 42107 30379
rect 42625 30345 42659 30379
rect 45201 30277 45235 30311
rect 42717 30209 42751 30243
rect 42984 30141 43018 30175
rect 46121 30141 46155 30175
rect 46377 30141 46411 30175
rect 41429 30005 41463 30039
rect 44097 30005 44131 30039
rect 45477 30005 45511 30039
rect 45845 30005 45879 30039
rect 47501 30005 47535 30039
rect 42257 29801 42291 29835
rect 42809 29801 42843 29835
rect 43545 29801 43579 29835
rect 43913 29801 43947 29835
rect 44557 29801 44591 29835
rect 46581 29801 46615 29835
rect 39396 29733 39430 29767
rect 42073 29733 42107 29767
rect 45468 29733 45502 29767
rect 45201 29665 45235 29699
rect 39129 29597 39163 29631
rect 41613 29597 41647 29631
rect 42349 29597 42383 29631
rect 40509 29461 40543 29495
rect 41797 29461 41831 29495
rect 39589 29257 39623 29291
rect 41797 29257 41831 29291
rect 44005 29257 44039 29291
rect 45477 29257 45511 29291
rect 45845 29257 45879 29291
rect 46949 29257 46983 29291
rect 40601 29189 40635 29223
rect 42257 29189 42291 29223
rect 44557 29189 44591 29223
rect 45017 29121 45051 29155
rect 42533 29053 42567 29087
rect 43177 29053 43211 29087
rect 44373 29053 44407 29087
rect 46765 29053 46799 29087
rect 39957 28985 39991 29019
rect 40877 28985 40911 29019
rect 41061 28985 41095 29019
rect 41153 28985 41187 29019
rect 42717 28985 42751 29019
rect 42809 28985 42843 29019
rect 43637 28985 43671 29019
rect 45017 28985 45051 29019
rect 45109 28985 45143 29019
rect 47317 28985 47351 29019
rect 39129 28917 39163 28951
rect 40233 28917 40267 28951
rect 40325 28713 40359 28747
rect 40969 28713 41003 28747
rect 41245 28713 41279 28747
rect 42441 28713 42475 28747
rect 42809 28713 42843 28747
rect 41981 28645 42015 28679
rect 45109 28645 45143 28679
rect 38945 28577 38979 28611
rect 39212 28577 39246 28611
rect 42073 28577 42107 28611
rect 43361 28577 43395 28611
rect 44925 28577 44959 28611
rect 46121 28577 46155 28611
rect 46388 28577 46422 28611
rect 41889 28509 41923 28543
rect 45201 28509 45235 28543
rect 41521 28373 41555 28407
rect 43545 28373 43579 28407
rect 44649 28373 44683 28407
rect 47501 28373 47535 28407
rect 39313 28169 39347 28203
rect 44005 28169 44039 28203
rect 44465 28169 44499 28203
rect 46213 28169 46247 28203
rect 43085 28101 43119 28135
rect 44741 28101 44775 28135
rect 45845 28101 45879 28135
rect 43545 28033 43579 28067
rect 46581 28033 46615 28067
rect 47501 28033 47535 28067
rect 40233 27965 40267 27999
rect 40509 27965 40543 27999
rect 42901 27965 42935 27999
rect 44557 27965 44591 27999
rect 45109 27965 45143 27999
rect 45569 27965 45603 27999
rect 47133 27965 47167 27999
rect 40754 27897 40788 27931
rect 43545 27897 43579 27931
rect 43637 27897 43671 27931
rect 46673 27897 46707 27931
rect 46765 27897 46799 27931
rect 47869 27897 47903 27931
rect 39037 27829 39071 27863
rect 39957 27829 39991 27863
rect 41889 27829 41923 27863
rect 42441 27829 42475 27863
rect 40509 27625 40543 27659
rect 41521 27625 41555 27659
rect 42717 27625 42751 27659
rect 43085 27625 43119 27659
rect 44741 27625 44775 27659
rect 46949 27625 46983 27659
rect 39396 27557 39430 27591
rect 42165 27557 42199 27591
rect 41981 27489 42015 27523
rect 44097 27489 44131 27523
rect 45569 27489 45603 27523
rect 45836 27489 45870 27523
rect 37749 27421 37783 27455
rect 39129 27421 39163 27455
rect 41153 27421 41187 27455
rect 42257 27421 42291 27455
rect 41705 27353 41739 27387
rect 38301 27285 38335 27319
rect 43913 27285 43947 27319
rect 44281 27285 44315 27319
rect 45109 27285 45143 27319
rect 38117 27081 38151 27115
rect 38393 27081 38427 27115
rect 39681 27081 39715 27115
rect 43269 27081 43303 27115
rect 44833 27081 44867 27115
rect 45569 27081 45603 27115
rect 46305 27081 46339 27115
rect 43913 27013 43947 27047
rect 38761 26945 38795 26979
rect 44281 26945 44315 26979
rect 35817 26877 35851 26911
rect 39313 26877 39347 26911
rect 41153 26877 41187 26911
rect 41337 26877 41371 26911
rect 36084 26809 36118 26843
rect 38945 26809 38979 26843
rect 40877 26809 40911 26843
rect 41582 26809 41616 26843
rect 44465 26809 44499 26843
rect 35725 26741 35759 26775
rect 37197 26741 37231 26775
rect 38853 26741 38887 26775
rect 42717 26741 42751 26775
rect 43729 26741 43763 26775
rect 44373 26741 44407 26775
rect 45293 26741 45327 26775
rect 35909 26537 35943 26571
rect 38393 26537 38427 26571
rect 39865 26537 39899 26571
rect 41245 26537 41279 26571
rect 41889 26469 41923 26503
rect 45109 26469 45143 26503
rect 38752 26401 38786 26435
rect 40509 26401 40543 26435
rect 43361 26401 43395 26435
rect 43913 26401 43947 26435
rect 44925 26401 44959 26435
rect 46121 26401 46155 26435
rect 46388 26401 46422 26435
rect 38485 26333 38519 26367
rect 41889 26333 41923 26367
rect 41981 26333 42015 26367
rect 44465 26333 44499 26367
rect 45201 26333 45235 26367
rect 41429 26265 41463 26299
rect 43545 26265 43579 26299
rect 36737 26197 36771 26231
rect 42441 26197 42475 26231
rect 44649 26197 44683 26231
rect 47501 26197 47535 26231
rect 38025 25993 38059 26027
rect 38669 25993 38703 26027
rect 38945 25993 38979 26027
rect 41613 25993 41647 26027
rect 43729 25993 43763 26027
rect 45017 25993 45051 26027
rect 45845 25993 45879 26027
rect 40601 25925 40635 25959
rect 42165 25925 42199 25959
rect 46213 25925 46247 25959
rect 41153 25857 41187 25891
rect 42349 25857 42383 25891
rect 36645 25789 36679 25823
rect 36912 25789 36946 25823
rect 39957 25789 39991 25823
rect 44833 25789 44867 25823
rect 46489 25789 46523 25823
rect 47133 25789 47167 25823
rect 39221 25721 39255 25755
rect 40325 25721 40359 25755
rect 40877 25721 40911 25755
rect 41061 25721 41095 25755
rect 42616 25721 42650 25755
rect 45569 25721 45603 25755
rect 46765 25721 46799 25755
rect 36001 25653 36035 25687
rect 36461 25653 36495 25687
rect 44649 25653 44683 25687
rect 46673 25653 46707 25687
rect 47501 25653 47535 25687
rect 36461 25449 36495 25483
rect 40693 25449 40727 25483
rect 41429 25449 41463 25483
rect 44557 25449 44591 25483
rect 44925 25449 44959 25483
rect 46949 25449 46983 25483
rect 38301 25381 38335 25415
rect 38393 25381 38427 25415
rect 39580 25381 39614 25415
rect 41797 25381 41831 25415
rect 43361 25381 43395 25415
rect 45753 25381 45787 25415
rect 36277 25313 36311 25347
rect 39313 25313 39347 25347
rect 42165 25313 42199 25347
rect 43545 25313 43579 25347
rect 46765 25313 46799 25347
rect 47317 25313 47351 25347
rect 35817 25245 35851 25279
rect 36553 25245 36587 25279
rect 38209 25245 38243 25279
rect 43729 25245 43763 25279
rect 45753 25245 45787 25279
rect 45845 25245 45879 25279
rect 36001 25177 36035 25211
rect 37841 25177 37875 25211
rect 45293 25177 45327 25211
rect 42349 25109 42383 25143
rect 46305 25109 46339 25143
rect 46673 25109 46707 25143
rect 36921 24905 36955 24939
rect 37841 24905 37875 24939
rect 38209 24905 38243 24939
rect 39313 24905 39347 24939
rect 39681 24905 39715 24939
rect 41705 24905 41739 24939
rect 43729 24905 43763 24939
rect 45753 24905 45787 24939
rect 45845 24905 45879 24939
rect 42809 24769 42843 24803
rect 44925 24769 44959 24803
rect 35541 24701 35575 24735
rect 38577 24701 38611 24735
rect 38669 24701 38703 24735
rect 42073 24701 42107 24735
rect 45753 24701 45787 24735
rect 46121 24701 46155 24735
rect 35808 24633 35842 24667
rect 42533 24633 42567 24667
rect 42717 24633 42751 24667
rect 45293 24633 45327 24667
rect 46388 24633 46422 24667
rect 35449 24565 35483 24599
rect 38853 24565 38887 24599
rect 42239 24565 42273 24599
rect 43453 24565 43487 24599
rect 47501 24565 47535 24599
rect 35081 24361 35115 24395
rect 36001 24361 36035 24395
rect 38025 24361 38059 24395
rect 41797 24361 41831 24395
rect 42257 24361 42291 24395
rect 42625 24361 42659 24395
rect 45293 24361 45327 24395
rect 46857 24361 46891 24395
rect 36645 24293 36679 24327
rect 36737 24293 36771 24327
rect 35633 24225 35667 24259
rect 41613 24225 41647 24259
rect 45744 24225 45778 24259
rect 36645 24157 36679 24191
rect 45477 24157 45511 24191
rect 36185 24089 36219 24123
rect 31217 24021 31251 24055
rect 41061 24021 41095 24055
rect 31309 23817 31343 23851
rect 35265 23817 35299 23851
rect 41061 23817 41095 23851
rect 42073 23817 42107 23851
rect 42349 23817 42383 23851
rect 35633 23749 35667 23783
rect 41613 23681 41647 23715
rect 36093 23613 36127 23647
rect 36360 23613 36394 23647
rect 42533 23613 42567 23647
rect 42789 23613 42823 23647
rect 31125 23545 31159 23579
rect 31585 23545 31619 23579
rect 31861 23545 31895 23579
rect 40877 23545 40911 23579
rect 41337 23545 41371 23579
rect 31769 23477 31803 23511
rect 35909 23477 35943 23511
rect 37473 23477 37507 23511
rect 38669 23477 38703 23511
rect 40325 23477 40359 23511
rect 41521 23477 41555 23511
rect 43913 23477 43947 23511
rect 45477 23477 45511 23511
rect 45937 23477 45971 23511
rect 32137 23273 32171 23307
rect 36553 23273 36587 23307
rect 38485 23273 38519 23307
rect 41613 23273 41647 23307
rect 42625 23273 42659 23307
rect 46029 23273 46063 23307
rect 47317 23273 47351 23307
rect 31309 23205 31343 23239
rect 34069 23205 34103 23239
rect 38669 23137 38703 23171
rect 39405 23137 39439 23171
rect 44916 23137 44950 23171
rect 47133 23137 47167 23171
rect 34069 23069 34103 23103
rect 34161 23069 34195 23103
rect 38992 23069 39026 23103
rect 39129 23069 39163 23103
rect 44649 23069 44683 23103
rect 33609 23001 33643 23035
rect 36185 22933 36219 22967
rect 40509 22933 40543 22967
rect 41153 22933 41187 22967
rect 43637 22933 43671 22967
rect 46673 22933 46707 22967
rect 46949 22933 46983 22967
rect 34253 22729 34287 22763
rect 38025 22729 38059 22763
rect 39865 22729 39899 22763
rect 42349 22729 42383 22763
rect 44925 22729 44959 22763
rect 46305 22729 46339 22763
rect 34621 22661 34655 22695
rect 38577 22661 38611 22695
rect 47317 22661 47351 22695
rect 34897 22593 34931 22627
rect 35541 22593 35575 22627
rect 39129 22593 39163 22627
rect 40233 22593 40267 22627
rect 46857 22593 46891 22627
rect 32321 22525 32355 22559
rect 32577 22525 32611 22559
rect 36001 22525 36035 22559
rect 36268 22525 36302 22559
rect 39497 22525 39531 22559
rect 40969 22525 41003 22559
rect 43361 22525 43395 22559
rect 43545 22525 43579 22559
rect 45477 22525 45511 22559
rect 38393 22457 38427 22491
rect 38853 22457 38887 22491
rect 41236 22457 41270 22491
rect 43812 22457 43846 22491
rect 45937 22457 45971 22491
rect 46581 22457 46615 22491
rect 29561 22389 29595 22423
rect 32229 22389 32263 22423
rect 33701 22389 33735 22423
rect 35909 22389 35943 22423
rect 37381 22389 37415 22423
rect 39037 22389 39071 22423
rect 40785 22389 40819 22423
rect 46765 22389 46799 22423
rect 30297 22185 30331 22219
rect 34989 22185 35023 22219
rect 36645 22185 36679 22219
rect 39773 22185 39807 22219
rect 45109 22185 45143 22219
rect 32413 22117 32447 22151
rect 33854 22117 33888 22151
rect 41521 22117 41555 22151
rect 43913 22117 43947 22151
rect 44741 22117 44775 22151
rect 28825 22049 28859 22083
rect 29173 22049 29207 22083
rect 36461 22049 36495 22083
rect 36737 22049 36771 22083
rect 40417 22049 40451 22083
rect 40877 22049 40911 22083
rect 41337 22049 41371 22083
rect 43729 22049 43763 22083
rect 44005 22049 44039 22083
rect 46377 22049 46411 22083
rect 27905 21981 27939 22015
rect 28917 21981 28951 22015
rect 33609 21981 33643 22015
rect 37933 21981 37967 22015
rect 38256 21981 38290 22015
rect 38393 21981 38427 22015
rect 38669 21981 38703 22015
rect 41613 21981 41647 22015
rect 46121 21981 46155 22015
rect 41061 21913 41095 21947
rect 47501 21913 47535 21947
rect 27721 21845 27755 21879
rect 31217 21845 31251 21879
rect 33425 21845 33459 21879
rect 36185 21845 36219 21879
rect 43453 21845 43487 21879
rect 29009 21641 29043 21675
rect 32505 21641 32539 21675
rect 37289 21641 37323 21675
rect 37565 21641 37599 21675
rect 38669 21641 38703 21675
rect 42625 21641 42659 21675
rect 43453 21641 43487 21675
rect 44833 21641 44867 21675
rect 45569 21641 45603 21675
rect 47501 21641 47535 21675
rect 27721 21573 27755 21607
rect 29377 21573 29411 21607
rect 43821 21573 43855 21607
rect 28273 21505 28307 21539
rect 29929 21505 29963 21539
rect 40325 21505 40359 21539
rect 41245 21505 41279 21539
rect 44373 21505 44407 21539
rect 45109 21505 45143 21539
rect 45937 21505 45971 21539
rect 46121 21505 46155 21539
rect 27537 21437 27571 21471
rect 27997 21437 28031 21471
rect 30297 21437 30331 21471
rect 31125 21437 31159 21471
rect 31381 21437 31415 21471
rect 33977 21437 34011 21471
rect 35173 21437 35207 21471
rect 35265 21437 35299 21471
rect 40785 21437 40819 21471
rect 41521 21437 41555 21471
rect 27169 21369 27203 21403
rect 28181 21369 28215 21403
rect 29653 21369 29687 21403
rect 31033 21369 31067 21403
rect 33701 21369 33735 21403
rect 35532 21369 35566 21403
rect 37749 21369 37783 21403
rect 39957 21369 39991 21403
rect 44097 21369 44131 21403
rect 46388 21369 46422 21403
rect 29837 21301 29871 21335
rect 36645 21301 36679 21335
rect 38209 21301 38243 21335
rect 41247 21301 41281 21335
rect 44281 21301 44315 21335
rect 29285 21097 29319 21131
rect 36185 21097 36219 21131
rect 36553 21097 36587 21131
rect 41245 21097 41279 21131
rect 41613 21097 41647 21131
rect 42349 21097 42383 21131
rect 43177 21097 43211 21131
rect 43453 21097 43487 21131
rect 44005 21097 44039 21131
rect 46121 21097 46155 21131
rect 46949 21097 46983 21131
rect 30941 21029 30975 21063
rect 31033 21029 31067 21063
rect 35357 21029 35391 21063
rect 45017 21029 45051 21063
rect 28181 20961 28215 20995
rect 32736 20961 32770 20995
rect 44833 20961 44867 20995
rect 46765 20961 46799 20995
rect 27445 20893 27479 20927
rect 27768 20893 27802 20927
rect 27905 20893 27939 20927
rect 30849 20893 30883 20927
rect 32413 20893 32447 20927
rect 32873 20893 32907 20927
rect 33149 20893 33183 20927
rect 40325 20893 40359 20927
rect 45109 20893 45143 20927
rect 46489 20893 46523 20927
rect 30481 20825 30515 20859
rect 44557 20825 44591 20859
rect 29929 20757 29963 20791
rect 34253 20757 34287 20791
rect 38025 20757 38059 20791
rect 38301 20757 38335 20791
rect 40785 20757 40819 20791
rect 44281 20757 44315 20791
rect 28181 20553 28215 20587
rect 31769 20553 31803 20587
rect 33241 20553 33275 20587
rect 37749 20553 37783 20587
rect 40325 20553 40359 20587
rect 40601 20553 40635 20587
rect 42073 20553 42107 20587
rect 44097 20553 44131 20587
rect 45017 20553 45051 20587
rect 46765 20553 46799 20587
rect 31033 20485 31067 20519
rect 32413 20485 32447 20519
rect 44649 20485 44683 20519
rect 27905 20417 27939 20451
rect 37933 20417 37967 20451
rect 40969 20417 41003 20451
rect 42717 20417 42751 20451
rect 42993 20417 43027 20451
rect 29561 20349 29595 20383
rect 29653 20349 29687 20383
rect 29920 20349 29954 20383
rect 38189 20349 38223 20383
rect 42257 20349 42291 20383
rect 42580 20349 42614 20383
rect 32137 20281 32171 20315
rect 33517 20281 33551 20315
rect 33793 20281 33827 20315
rect 41153 20281 41187 20315
rect 27169 20213 27203 20247
rect 27445 20213 27479 20247
rect 33057 20213 33091 20247
rect 33701 20213 33735 20247
rect 35173 20213 35207 20247
rect 36921 20213 36955 20247
rect 39313 20213 39347 20247
rect 39865 20213 39899 20247
rect 41061 20213 41095 20247
rect 41521 20213 41555 20247
rect 29745 20009 29779 20043
rect 30481 20009 30515 20043
rect 31217 20009 31251 20043
rect 32321 20009 32355 20043
rect 33241 20009 33275 20043
rect 33609 20009 33643 20043
rect 39129 20009 39163 20043
rect 41613 20009 41647 20043
rect 42625 20009 42659 20043
rect 44557 20009 44591 20043
rect 46121 20009 46155 20043
rect 47409 20009 47443 20043
rect 32781 19941 32815 19975
rect 40478 19941 40512 19975
rect 42349 19941 42383 19975
rect 32137 19873 32171 19907
rect 34980 19873 35014 19907
rect 37749 19873 37783 19907
rect 38016 19873 38050 19907
rect 45008 19873 45042 19907
rect 47225 19873 47259 19907
rect 29837 19805 29871 19839
rect 30757 19805 30791 19839
rect 34713 19805 34747 19839
rect 40233 19805 40267 19839
rect 43729 19805 43763 19839
rect 44741 19805 44775 19839
rect 34621 19669 34655 19703
rect 36093 19669 36127 19703
rect 43637 19669 43671 19703
rect 31125 19465 31159 19499
rect 37749 19465 37783 19499
rect 40601 19465 40635 19499
rect 43453 19465 43487 19499
rect 47317 19465 47351 19499
rect 31677 19397 31711 19431
rect 29653 19329 29687 19363
rect 29745 19329 29779 19363
rect 35541 19329 35575 19363
rect 38669 19329 38703 19363
rect 41153 19329 41187 19363
rect 44005 19329 44039 19363
rect 44189 19329 44223 19363
rect 45109 19329 45143 19363
rect 32137 19261 32171 19295
rect 32229 19261 32263 19295
rect 34345 19261 34379 19295
rect 34713 19261 34747 19295
rect 35081 19261 35115 19295
rect 35817 19261 35851 19295
rect 38099 19261 38133 19295
rect 41521 19261 41555 19295
rect 41889 19261 41923 19295
rect 43619 19261 43653 19295
rect 29101 19193 29135 19227
rect 29990 19193 30024 19227
rect 32474 19193 32508 19227
rect 38393 19193 38427 19227
rect 39037 19193 39071 19227
rect 39957 19193 39991 19227
rect 40877 19193 40911 19227
rect 41061 19193 41095 19227
rect 33609 19125 33643 19159
rect 35543 19125 35577 19159
rect 36921 19125 36955 19159
rect 38577 19125 38611 19159
rect 39405 19125 39439 19159
rect 40325 19125 40359 19159
rect 43085 19125 43119 19159
rect 44097 19125 44131 19159
rect 44833 19125 44867 19159
rect 34621 18921 34655 18955
rect 38761 18921 38795 18955
rect 40233 18921 40267 18955
rect 40787 18921 40821 18955
rect 42165 18921 42199 18955
rect 45017 18921 45051 18955
rect 30113 18853 30147 18887
rect 30205 18853 30239 18887
rect 34897 18853 34931 18887
rect 35449 18853 35483 18887
rect 35633 18853 35667 18887
rect 35725 18853 35759 18887
rect 38301 18853 38335 18887
rect 29929 18785 29963 18819
rect 38117 18785 38151 18819
rect 41061 18785 41095 18819
rect 43904 18785 43938 18819
rect 46377 18785 46411 18819
rect 34069 18717 34103 18751
rect 38393 18717 38427 18751
rect 40325 18717 40359 18751
rect 40785 18717 40819 18751
rect 43637 18717 43671 18751
rect 46121 18717 46155 18751
rect 29653 18649 29687 18683
rect 37565 18649 37599 18683
rect 37841 18649 37875 18683
rect 29469 18581 29503 18615
rect 32321 18581 32355 18615
rect 35173 18581 35207 18615
rect 42901 18581 42935 18615
rect 47501 18581 47535 18615
rect 29101 18377 29135 18411
rect 34713 18377 34747 18411
rect 37749 18377 37783 18411
rect 38117 18377 38151 18411
rect 39957 18377 39991 18411
rect 40785 18377 40819 18411
rect 41981 18377 42015 18411
rect 43913 18377 43947 18411
rect 44373 18377 44407 18411
rect 45569 18377 45603 18411
rect 45937 18377 45971 18411
rect 35173 18309 35207 18343
rect 40233 18309 40267 18343
rect 42993 18309 43027 18343
rect 44649 18309 44683 18343
rect 35541 18241 35575 18275
rect 35725 18241 35759 18275
rect 43545 18241 43579 18275
rect 46121 18241 46155 18275
rect 29561 18173 29595 18207
rect 29653 18173 29687 18207
rect 35981 18173 36015 18207
rect 41797 18173 41831 18207
rect 44465 18173 44499 18207
rect 45017 18173 45051 18207
rect 29920 18105 29954 18139
rect 42441 18105 42475 18139
rect 43269 18105 43303 18139
rect 46388 18105 46422 18139
rect 28733 18037 28767 18071
rect 31033 18037 31067 18071
rect 34345 18037 34379 18071
rect 37105 18037 37139 18071
rect 38577 18037 38611 18071
rect 41061 18037 41095 18071
rect 42809 18037 42843 18071
rect 43453 18037 43487 18071
rect 47501 18037 47535 18071
rect 29285 17833 29319 17867
rect 33609 17833 33643 17867
rect 36001 17833 36035 17867
rect 41153 17833 41187 17867
rect 43913 17833 43947 17867
rect 46213 17833 46247 17867
rect 29745 17765 29779 17799
rect 30573 17765 30607 17799
rect 30757 17765 30791 17799
rect 30849 17765 30883 17799
rect 35449 17765 35483 17799
rect 44005 17765 44039 17799
rect 45753 17765 45787 17799
rect 46765 17765 46799 17799
rect 46949 17765 46983 17799
rect 47409 17765 47443 17799
rect 29101 17697 29135 17731
rect 30113 17697 30147 17731
rect 32229 17697 32263 17731
rect 32485 17697 32519 17731
rect 40969 17697 41003 17731
rect 42073 17697 42107 17731
rect 43729 17697 43763 17731
rect 45569 17697 45603 17731
rect 46581 17697 46615 17731
rect 35357 17629 35391 17663
rect 35541 17629 35575 17663
rect 45845 17629 45879 17663
rect 30297 17561 30331 17595
rect 34989 17561 35023 17595
rect 43453 17561 43487 17595
rect 45109 17561 45143 17595
rect 31953 17493 31987 17527
rect 41613 17493 41647 17527
rect 42257 17493 42291 17527
rect 42993 17493 43027 17527
rect 45293 17493 45327 17527
rect 47133 17493 47167 17527
rect 30021 17289 30055 17323
rect 30297 17289 30331 17323
rect 31769 17289 31803 17323
rect 34713 17289 34747 17323
rect 35173 17289 35207 17323
rect 41245 17289 41279 17323
rect 42165 17289 42199 17323
rect 42625 17289 42659 17323
rect 42993 17289 43027 17323
rect 43269 17289 43303 17323
rect 43729 17289 43763 17323
rect 44097 17289 44131 17323
rect 44833 17289 44867 17323
rect 45937 17289 45971 17323
rect 47501 17289 47535 17323
rect 26525 17221 26559 17255
rect 30665 17221 30699 17255
rect 35541 17221 35575 17255
rect 31861 17153 31895 17187
rect 41613 17153 41647 17187
rect 46121 17153 46155 17187
rect 23765 17085 23799 17119
rect 26801 17085 26835 17119
rect 30113 17085 30147 17119
rect 32117 17085 32151 17119
rect 37197 17085 37231 17119
rect 37453 17085 37487 17119
rect 40325 17085 40359 17119
rect 41797 17085 41831 17119
rect 43085 17085 43119 17119
rect 44189 17085 44223 17119
rect 23489 17017 23523 17051
rect 24010 17017 24044 17051
rect 25973 17017 26007 17051
rect 27077 17017 27111 17051
rect 31401 17017 31435 17051
rect 37105 17017 37139 17051
rect 40969 17017 41003 17051
rect 41705 17017 41739 17051
rect 45201 17017 45235 17051
rect 45569 17017 45603 17051
rect 46388 17017 46422 17051
rect 25145 16949 25179 16983
rect 26341 16949 26375 16983
rect 26985 16949 27019 16983
rect 29561 16949 29595 16983
rect 33241 16949 33275 16983
rect 38577 16949 38611 16983
rect 44373 16949 44407 16983
rect 29459 16745 29493 16779
rect 31861 16745 31895 16779
rect 33241 16745 33275 16779
rect 35173 16745 35207 16779
rect 37289 16745 37323 16779
rect 39681 16745 39715 16779
rect 40601 16745 40635 16779
rect 42165 16745 42199 16779
rect 43435 16745 43469 16779
rect 44833 16745 44867 16779
rect 46581 16745 46615 16779
rect 47133 16745 47167 16779
rect 27160 16677 27194 16711
rect 29929 16677 29963 16711
rect 32505 16677 32539 16711
rect 38568 16677 38602 16711
rect 41030 16677 41064 16711
rect 43913 16677 43947 16711
rect 23857 16609 23891 16643
rect 26801 16609 26835 16643
rect 28825 16609 28859 16643
rect 30021 16609 30055 16643
rect 30849 16609 30883 16643
rect 30941 16609 30975 16643
rect 32137 16609 32171 16643
rect 32321 16609 32355 16643
rect 33793 16609 33827 16643
rect 34060 16609 34094 16643
rect 43177 16609 43211 16643
rect 43729 16609 43763 16643
rect 45201 16609 45235 16643
rect 45468 16609 45502 16643
rect 26893 16541 26927 16575
rect 29285 16541 29319 16575
rect 29837 16541 29871 16575
rect 38301 16541 38335 16575
rect 40785 16541 40819 16575
rect 44005 16541 44039 16575
rect 28273 16405 28307 16439
rect 30481 16405 30515 16439
rect 31125 16405 31159 16439
rect 31493 16405 31527 16439
rect 33701 16405 33735 16439
rect 44465 16405 44499 16439
rect 25329 16201 25363 16235
rect 26893 16201 26927 16235
rect 29009 16201 29043 16235
rect 29377 16201 29411 16235
rect 30389 16201 30423 16235
rect 30941 16201 30975 16235
rect 32505 16201 32539 16235
rect 34253 16201 34287 16235
rect 34529 16201 34563 16235
rect 34713 16201 34747 16235
rect 36921 16201 36955 16235
rect 38669 16201 38703 16235
rect 38945 16201 38979 16235
rect 43821 16201 43855 16235
rect 44557 16201 44591 16235
rect 45569 16201 45603 16235
rect 33333 16133 33367 16167
rect 46213 16133 46247 16167
rect 25513 16065 25547 16099
rect 31309 16065 31343 16099
rect 31493 16065 31527 16099
rect 33701 16065 33735 16099
rect 34529 16065 34563 16099
rect 35357 16065 35391 16099
rect 35541 16065 35575 16099
rect 39405 16065 39439 16099
rect 42809 16065 42843 16099
rect 45017 16065 45051 16099
rect 25780 15997 25814 16031
rect 33149 15997 33183 16031
rect 38025 15997 38059 16031
rect 40601 15997 40635 16031
rect 40693 15997 40727 16031
rect 40960 15997 40994 16031
rect 43269 15997 43303 16031
rect 47133 15997 47167 16031
rect 28641 15929 28675 15963
rect 29653 15929 29687 15963
rect 29929 15929 29963 15963
rect 33793 15929 33827 15963
rect 33885 15929 33919 15963
rect 35786 15929 35820 15963
rect 39405 15929 39439 15963
rect 39497 15929 39531 15963
rect 45017 15929 45051 15963
rect 45109 15929 45143 15963
rect 46489 15929 46523 15963
rect 46765 15929 46799 15963
rect 47593 15929 47627 15963
rect 27445 15861 27479 15895
rect 28365 15861 28399 15895
rect 29837 15861 29871 15895
rect 30665 15861 30699 15895
rect 31401 15861 31435 15895
rect 32229 15861 32263 15895
rect 38301 15861 38335 15895
rect 39865 15861 39899 15895
rect 40233 15861 40267 15895
rect 40601 15861 40635 15895
rect 42073 15861 42107 15895
rect 43177 15861 43211 15895
rect 43453 15861 43487 15895
rect 44281 15861 44315 15895
rect 45937 15861 45971 15895
rect 46673 15861 46707 15895
rect 25605 15657 25639 15691
rect 26893 15657 26927 15691
rect 29561 15657 29595 15691
rect 31309 15657 31343 15691
rect 38853 15657 38887 15691
rect 39313 15657 39347 15691
rect 40601 15657 40635 15691
rect 41245 15657 41279 15691
rect 43913 15657 43947 15691
rect 44557 15657 44591 15691
rect 45293 15657 45327 15691
rect 47501 15657 47535 15691
rect 28448 15589 28482 15623
rect 33517 15589 33551 15623
rect 34603 15589 34637 15623
rect 35081 15589 35115 15623
rect 38025 15589 38059 15623
rect 41061 15589 41095 15623
rect 43729 15589 43763 15623
rect 28181 15521 28215 15555
rect 30665 15521 30699 15555
rect 34897 15521 34931 15555
rect 35541 15521 35575 15555
rect 46121 15521 46155 15555
rect 46388 15521 46422 15555
rect 33517 15453 33551 15487
rect 33609 15453 33643 15487
rect 35173 15453 35207 15487
rect 41337 15453 41371 15487
rect 44005 15453 44039 15487
rect 31769 15385 31803 15419
rect 43453 15385 43487 15419
rect 30389 15317 30423 15351
rect 30849 15317 30883 15351
rect 32321 15317 32355 15351
rect 33057 15317 33091 15351
rect 34437 15317 34471 15351
rect 40785 15317 40819 15351
rect 41797 15317 41831 15351
rect 44833 15317 44867 15351
rect 28181 15113 28215 15147
rect 28641 15113 28675 15147
rect 30389 15113 30423 15147
rect 31309 15113 31343 15147
rect 31953 15113 31987 15147
rect 32965 15113 32999 15147
rect 33241 15113 33275 15147
rect 36553 15113 36587 15147
rect 40785 15113 40819 15147
rect 41153 15113 41187 15147
rect 43085 15113 43119 15147
rect 44189 15113 44223 15147
rect 46305 15113 46339 15147
rect 47317 15113 47351 15147
rect 40325 15045 40359 15079
rect 41705 15045 41739 15079
rect 43269 15045 43303 15079
rect 46949 15045 46983 15079
rect 29101 14977 29135 15011
rect 30941 14977 30975 15011
rect 32505 14977 32539 15011
rect 43637 14977 43671 15011
rect 44557 14977 44591 15011
rect 30665 14909 30699 14943
rect 32229 14909 32263 14943
rect 33425 14909 33459 14943
rect 35173 14909 35207 14943
rect 37933 14909 37967 14943
rect 38200 14909 38234 14943
rect 42257 14909 42291 14943
rect 43821 14909 43855 14943
rect 44925 14909 44959 14943
rect 46765 14909 46799 14943
rect 30205 14841 30239 14875
rect 30849 14841 30883 14875
rect 34345 14841 34379 14875
rect 34713 14841 34747 14875
rect 35440 14841 35474 14875
rect 41981 14841 42015 14875
rect 45937 14841 45971 14875
rect 27629 14773 27663 14807
rect 29745 14773 29779 14807
rect 31677 14773 31711 14807
rect 32413 14773 32447 14807
rect 33609 14773 33643 14807
rect 37749 14773 37783 14807
rect 39313 14773 39347 14807
rect 41521 14773 41555 14807
rect 42165 14773 42199 14807
rect 42625 14773 42659 14807
rect 43729 14773 43763 14807
rect 28825 14569 28859 14603
rect 30297 14569 30331 14603
rect 31125 14569 31159 14603
rect 31953 14569 31987 14603
rect 32413 14569 32447 14603
rect 33609 14569 33643 14603
rect 34621 14569 34655 14603
rect 39129 14569 39163 14603
rect 40141 14569 40175 14603
rect 41705 14569 41739 14603
rect 42257 14569 42291 14603
rect 43177 14569 43211 14603
rect 46949 14569 46983 14603
rect 29837 14501 29871 14535
rect 29929 14501 29963 14535
rect 40739 14501 40773 14535
rect 40877 14501 40911 14535
rect 44373 14501 44407 14535
rect 44465 14501 44499 14535
rect 26617 14433 26651 14467
rect 26884 14433 26918 14467
rect 29193 14433 29227 14467
rect 29653 14433 29687 14467
rect 30113 14433 30147 14467
rect 30665 14433 30699 14467
rect 30941 14433 30975 14467
rect 32229 14433 32263 14467
rect 38016 14433 38050 14467
rect 42073 14433 42107 14467
rect 46765 14433 46799 14467
rect 37749 14365 37783 14399
rect 40693 14365 40727 14399
rect 44281 14365 44315 14399
rect 8401 14297 8435 14331
rect 29377 14297 29411 14331
rect 32965 14297 32999 14331
rect 40325 14297 40359 14331
rect 43913 14297 43947 14331
rect 46213 14297 46247 14331
rect 19809 14229 19843 14263
rect 27997 14229 28031 14263
rect 31585 14229 31619 14263
rect 33333 14229 33367 14263
rect 33977 14229 34011 14263
rect 35265 14229 35299 14263
rect 43637 14229 43671 14263
rect 46581 14229 46615 14263
rect 26617 14025 26651 14059
rect 26985 14025 27019 14059
rect 29745 14025 29779 14059
rect 31033 14025 31067 14059
rect 31769 14025 31803 14059
rect 36277 14025 36311 14059
rect 39865 14025 39899 14059
rect 41889 14025 41923 14059
rect 42533 14025 42567 14059
rect 43085 14025 43119 14059
rect 45477 14025 45511 14059
rect 46213 14025 46247 14059
rect 47225 14025 47259 14059
rect 19809 13957 19843 13991
rect 27629 13957 27663 13991
rect 33333 13957 33367 13991
rect 19625 13889 19659 13923
rect 20269 13889 20303 13923
rect 28089 13889 28123 13923
rect 30297 13889 30331 13923
rect 32321 13889 32355 13923
rect 33885 13889 33919 13923
rect 40325 13889 40359 13923
rect 46673 13889 46707 13923
rect 8217 13821 8251 13855
rect 8309 13821 8343 13855
rect 8565 13821 8599 13855
rect 19257 13821 19291 13855
rect 20361 13821 20395 13855
rect 28181 13821 28215 13855
rect 29101 13821 29135 13855
rect 30021 13821 30055 13855
rect 32045 13821 32079 13855
rect 32689 13821 32723 13855
rect 33609 13821 33643 13855
rect 34253 13821 34287 13855
rect 34897 13821 34931 13855
rect 35164 13821 35198 13855
rect 37933 13821 37967 13855
rect 39589 13821 39623 13855
rect 40509 13821 40543 13855
rect 43545 13821 43579 13855
rect 43801 13821 43835 13855
rect 20269 13753 20303 13787
rect 28089 13753 28123 13787
rect 34621 13753 34655 13787
rect 40754 13753 40788 13787
rect 46765 13753 46799 13787
rect 4169 13685 4203 13719
rect 9689 13685 9723 13719
rect 27445 13685 27479 13719
rect 28641 13685 28675 13719
rect 29561 13685 29595 13719
rect 30205 13685 30239 13719
rect 31585 13685 31619 13719
rect 32229 13685 32263 13719
rect 33149 13685 33183 13719
rect 33793 13685 33827 13719
rect 37381 13685 37415 13719
rect 38301 13685 38335 13719
rect 43361 13685 43395 13719
rect 44925 13685 44959 13719
rect 45937 13685 45971 13719
rect 46673 13685 46707 13719
rect 4629 13481 4663 13515
rect 29377 13481 29411 13515
rect 31033 13481 31067 13515
rect 33517 13481 33551 13515
rect 35817 13481 35851 13515
rect 40693 13481 40727 13515
rect 41245 13481 41279 13515
rect 43177 13481 43211 13515
rect 44741 13481 44775 13515
rect 47501 13481 47535 13515
rect 4721 13413 4755 13447
rect 6285 13413 6319 13447
rect 19809 13413 19843 13447
rect 27436 13413 27470 13447
rect 29920 13413 29954 13447
rect 32689 13413 32723 13447
rect 32781 13413 32815 13447
rect 35357 13413 35391 13447
rect 37565 13413 37599 13447
rect 38301 13413 38335 13447
rect 39558 13413 39592 13447
rect 43606 13413 43640 13447
rect 6736 13345 6770 13379
rect 19625 13345 19659 13379
rect 27169 13345 27203 13379
rect 31953 13345 31987 13379
rect 32505 13345 32539 13379
rect 33793 13345 33827 13379
rect 35633 13345 35667 13379
rect 46029 13345 46063 13379
rect 46388 13345 46422 13379
rect 2053 13277 2087 13311
rect 3893 13277 3927 13311
rect 4629 13277 4663 13311
rect 6469 13277 6503 13311
rect 19901 13277 19935 13311
rect 29653 13277 29687 13311
rect 38209 13277 38243 13311
rect 38393 13277 38427 13311
rect 39313 13277 39347 13311
rect 43361 13277 43395 13311
rect 46121 13277 46155 13311
rect 32229 13209 32263 13243
rect 37841 13209 37875 13243
rect 1593 13141 1627 13175
rect 4169 13141 4203 13175
rect 7849 13141 7883 13175
rect 19349 13141 19383 13175
rect 20269 13141 20303 13175
rect 28549 13141 28583 13175
rect 33149 13141 33183 13175
rect 36185 13141 36219 13175
rect 36921 13141 36955 13175
rect 5641 12937 5675 12971
rect 6469 12937 6503 12971
rect 7941 12937 7975 12971
rect 9873 12937 9907 12971
rect 19349 12937 19383 12971
rect 27169 12937 27203 12971
rect 27537 12937 27571 12971
rect 30021 12937 30055 12971
rect 34345 12937 34379 12971
rect 36277 12937 36311 12971
rect 38761 12937 38795 12971
rect 39681 12937 39715 12971
rect 41429 12937 41463 12971
rect 44097 12937 44131 12971
rect 45109 12937 45143 12971
rect 47501 12937 47535 12971
rect 6929 12869 6963 12903
rect 39405 12869 39439 12903
rect 42901 12869 42935 12903
rect 43821 12869 43855 12903
rect 7389 12801 7423 12835
rect 20361 12801 20395 12835
rect 41521 12801 41555 12835
rect 44557 12801 44591 12835
rect 1501 12733 1535 12767
rect 1768 12733 1802 12767
rect 4169 12733 4203 12767
rect 4261 12733 4295 12767
rect 7481 12733 7515 12767
rect 8493 12733 8527 12767
rect 8760 12733 8794 12767
rect 19901 12733 19935 12767
rect 20637 12733 20671 12767
rect 32965 12733 32999 12767
rect 33232 12733 33266 12767
rect 34897 12733 34931 12767
rect 36829 12733 36863 12767
rect 37085 12733 37119 12767
rect 41788 12733 41822 12767
rect 43545 12733 43579 12767
rect 44649 12733 44683 12767
rect 46121 12733 46155 12767
rect 46388 12733 46422 12767
rect 3801 12665 3835 12699
rect 4506 12665 4540 12699
rect 31125 12665 31159 12699
rect 32873 12665 32907 12699
rect 35142 12665 35176 12699
rect 41061 12665 41095 12699
rect 2881 12597 2915 12631
rect 7389 12597 7423 12631
rect 8401 12597 8435 12631
rect 18889 12597 18923 12631
rect 19809 12597 19843 12631
rect 20363 12597 20397 12631
rect 21741 12597 21775 12631
rect 29653 12597 29687 12631
rect 31033 12597 31067 12631
rect 38209 12597 38243 12631
rect 44557 12597 44591 12631
rect 45569 12597 45603 12631
rect 45845 12597 45879 12631
rect 5457 12393 5491 12427
rect 6377 12393 6411 12427
rect 7665 12393 7699 12427
rect 8585 12393 8619 12427
rect 19349 12393 19383 12427
rect 19533 12393 19567 12427
rect 20085 12393 20119 12427
rect 22293 12393 22327 12427
rect 29745 12393 29779 12427
rect 31585 12393 31619 12427
rect 33517 12393 33551 12427
rect 36001 12393 36035 12427
rect 37565 12393 37599 12427
rect 41337 12393 41371 12427
rect 44097 12393 44131 12427
rect 47685 12393 47719 12427
rect 1768 12325 1802 12359
rect 3893 12325 3927 12359
rect 4344 12325 4378 12359
rect 7113 12325 7147 12359
rect 18521 12325 18555 12359
rect 21180 12325 21214 12359
rect 31953 12325 31987 12359
rect 32404 12325 32438 12359
rect 34866 12325 34900 12359
rect 36921 12325 36955 12359
rect 38577 12325 38611 12359
rect 40141 12325 40175 12359
rect 1501 12257 1535 12291
rect 6929 12257 6963 12291
rect 9956 12257 9990 12291
rect 18337 12257 18371 12291
rect 28365 12257 28399 12291
rect 28632 12257 28666 12291
rect 38393 12257 38427 12291
rect 41153 12257 41187 12291
rect 44465 12257 44499 12291
rect 45284 12257 45318 12291
rect 47501 12257 47535 12291
rect 4077 12189 4111 12223
rect 7205 12189 7239 12223
rect 9689 12189 9723 12223
rect 18613 12189 18647 12223
rect 20913 12189 20947 12223
rect 32137 12189 32171 12223
rect 34437 12189 34471 12223
rect 34621 12189 34655 12223
rect 38669 12189 38703 12223
rect 40049 12189 40083 12223
rect 40233 12189 40267 12223
rect 45017 12189 45051 12223
rect 38117 12121 38151 12155
rect 46397 12121 46431 12155
rect 46949 12121 46983 12155
rect 2881 12053 2915 12087
rect 3525 12053 3559 12087
rect 6653 12053 6687 12087
rect 11069 12053 11103 12087
rect 13645 12053 13679 12087
rect 16037 12053 16071 12087
rect 18061 12053 18095 12087
rect 19073 12053 19107 12087
rect 20453 12053 20487 12087
rect 23673 12053 23707 12087
rect 34069 12053 34103 12087
rect 39681 12053 39715 12087
rect 40877 12053 40911 12087
rect 1593 11849 1627 11883
rect 2881 11849 2915 11883
rect 4353 11849 4387 11883
rect 4813 11849 4847 11883
rect 5549 11849 5583 11883
rect 6285 11849 6319 11883
rect 10057 11849 10091 11883
rect 16129 11849 16163 11883
rect 17877 11849 17911 11883
rect 18245 11849 18279 11883
rect 21373 11849 21407 11883
rect 25053 11849 25087 11883
rect 28365 11849 28399 11883
rect 28733 11849 28767 11883
rect 32137 11849 32171 11883
rect 32597 11849 32631 11883
rect 34253 11849 34287 11883
rect 34621 11849 34655 11883
rect 35173 11849 35207 11883
rect 39037 11849 39071 11883
rect 39681 11849 39715 11883
rect 40049 11849 40083 11883
rect 45385 11849 45419 11883
rect 47501 11849 47535 11883
rect 1869 11781 1903 11815
rect 3433 11781 3467 11815
rect 6653 11781 6687 11815
rect 7573 11781 7607 11815
rect 11437 11781 11471 11815
rect 21005 11781 21039 11815
rect 23397 11781 23431 11815
rect 35633 11781 35667 11815
rect 2329 11713 2363 11747
rect 8033 11713 8067 11747
rect 9781 11713 9815 11747
rect 13369 11713 13403 11747
rect 13553 11713 13587 11747
rect 16681 11713 16715 11747
rect 23673 11713 23707 11747
rect 37565 11713 37599 11747
rect 37657 11713 37691 11747
rect 5641 11645 5675 11679
rect 11253 11645 11287 11679
rect 11805 11645 11839 11679
rect 13809 11645 13843 11679
rect 18981 11645 19015 11679
rect 35449 11645 35483 11679
rect 40785 11645 40819 11679
rect 41521 11645 41555 11679
rect 2329 11577 2363 11611
rect 2421 11577 2455 11611
rect 3709 11577 3743 11611
rect 3985 11577 4019 11611
rect 8125 11577 8159 11611
rect 16405 11577 16439 11611
rect 16589 11577 16623 11611
rect 19248 11577 19282 11611
rect 23918 11577 23952 11611
rect 37197 11577 37231 11611
rect 37902 11577 37936 11611
rect 40969 11577 41003 11611
rect 3249 11509 3283 11543
rect 3893 11509 3927 11543
rect 5825 11509 5859 11543
rect 7389 11509 7423 11543
rect 8033 11509 8067 11543
rect 14933 11509 14967 11543
rect 15485 11509 15519 11543
rect 15853 11509 15887 11543
rect 18797 11509 18831 11543
rect 20361 11509 20395 11543
rect 36001 11509 36035 11543
rect 41153 11509 41187 11543
rect 41797 11509 41831 11543
rect 45017 11509 45051 11543
rect 2421 11305 2455 11339
rect 2697 11305 2731 11339
rect 3341 11305 3375 11339
rect 5447 11305 5481 11339
rect 5917 11305 5951 11339
rect 7573 11305 7607 11339
rect 12725 11305 12759 11339
rect 13369 11305 13403 11339
rect 14197 11305 14231 11339
rect 37473 11305 37507 11339
rect 37933 11305 37967 11339
rect 38393 11305 38427 11339
rect 38669 11305 38703 11339
rect 39037 11305 39071 11339
rect 42073 11305 42107 11339
rect 1685 11237 1719 11271
rect 2053 11237 2087 11271
rect 15936 11237 15970 11271
rect 26884 11237 26918 11271
rect 34130 11237 34164 11271
rect 43913 11237 43947 11271
rect 4261 11169 4295 11203
rect 10241 11169 10275 11203
rect 11345 11169 11379 11203
rect 11612 11169 11646 11203
rect 15669 11169 15703 11203
rect 18061 11169 18095 11203
rect 18420 11169 18454 11203
rect 22457 11169 22491 11203
rect 26617 11169 26651 11203
rect 29101 11169 29135 11203
rect 29368 11169 29402 11203
rect 33885 11169 33919 11203
rect 37749 11169 37783 11203
rect 38853 11169 38887 11203
rect 40693 11169 40727 11203
rect 40960 11169 40994 11203
rect 43729 11169 43763 11203
rect 5825 11101 5859 11135
rect 6009 11101 6043 11135
rect 18153 11101 18187 11135
rect 22201 11101 22235 11135
rect 44005 11101 44039 11135
rect 5273 11033 5307 11067
rect 6469 11033 6503 11067
rect 10425 11033 10459 11067
rect 17049 11033 17083 11067
rect 19533 11033 19567 11067
rect 20453 11033 20487 11067
rect 23581 11033 23615 11067
rect 27997 11033 28031 11067
rect 30481 11033 30515 11067
rect 39865 11033 39899 11067
rect 43177 11033 43211 11067
rect 4445 10965 4479 10999
rect 6929 10965 6963 10999
rect 7849 10965 7883 10999
rect 8493 10965 8527 10999
rect 35265 10965 35299 10999
rect 35817 10965 35851 10999
rect 39497 10965 39531 10999
rect 43453 10965 43487 10999
rect 4353 10761 4387 10795
rect 4997 10761 5031 10795
rect 5273 10761 5307 10795
rect 6193 10761 6227 10795
rect 11069 10761 11103 10795
rect 11897 10761 11931 10795
rect 12541 10761 12575 10795
rect 15669 10761 15703 10795
rect 16037 10761 16071 10795
rect 19073 10761 19107 10795
rect 22753 10761 22787 10795
rect 25881 10761 25915 10795
rect 27261 10761 27295 10795
rect 28365 10761 28399 10795
rect 30665 10761 30699 10795
rect 33885 10761 33919 10795
rect 34253 10761 34287 10795
rect 38393 10761 38427 10795
rect 39865 10761 39899 10795
rect 41061 10761 41095 10795
rect 41521 10761 41555 10795
rect 44741 10761 44775 10795
rect 6929 10693 6963 10727
rect 11437 10693 11471 10727
rect 18153 10693 18187 10727
rect 34621 10693 34655 10727
rect 37933 10693 37967 10727
rect 38669 10693 38703 10727
rect 38945 10693 38979 10727
rect 40785 10693 40819 10727
rect 1593 10625 1627 10659
rect 7481 10625 7515 10659
rect 7849 10625 7883 10659
rect 12173 10625 12207 10659
rect 13093 10625 13127 10659
rect 20821 10625 20855 10659
rect 21097 10625 21131 10659
rect 28641 10625 28675 10659
rect 29009 10625 29043 10659
rect 29285 10625 29319 10659
rect 34989 10625 35023 10659
rect 1860 10557 1894 10591
rect 5549 10557 5583 10591
rect 7205 10557 7239 10591
rect 8309 10557 8343 10591
rect 8401 10557 8435 10591
rect 8657 10557 8691 10591
rect 11253 10557 11287 10591
rect 12817 10557 12851 10591
rect 13461 10557 13495 10591
rect 18705 10557 18739 10591
rect 19901 10557 19935 10591
rect 20361 10557 20395 10591
rect 37657 10557 37691 10591
rect 37749 10557 37783 10591
rect 43361 10557 43395 10591
rect 4721 10489 4755 10523
rect 5825 10489 5859 10523
rect 13001 10489 13035 10523
rect 17509 10489 17543 10523
rect 18429 10489 18463 10523
rect 18613 10489 18647 10523
rect 25973 10489 26007 10523
rect 29552 10489 29586 10523
rect 35256 10489 35290 10523
rect 39221 10489 39255 10523
rect 39405 10489 39439 10523
rect 39497 10489 39531 10523
rect 41797 10489 41831 10523
rect 42073 10489 42107 10523
rect 42533 10489 42567 10523
rect 42901 10489 42935 10523
rect 43628 10489 43662 10523
rect 2973 10421 3007 10455
rect 5733 10421 5767 10455
rect 6653 10421 6687 10455
rect 7389 10421 7423 10455
rect 9781 10421 9815 10455
rect 10425 10421 10459 10455
rect 17785 10421 17819 10455
rect 20269 10421 20303 10455
rect 20823 10421 20857 10455
rect 22201 10421 22235 10455
rect 23673 10421 23707 10455
rect 36369 10421 36403 10455
rect 41981 10421 42015 10455
rect 43269 10421 43303 10455
rect 1593 10217 1627 10251
rect 2513 10217 2547 10251
rect 4353 10217 4387 10251
rect 5273 10217 5307 10251
rect 5549 10217 5583 10251
rect 5917 10217 5951 10251
rect 8585 10217 8619 10251
rect 12725 10217 12759 10251
rect 13185 10217 13219 10251
rect 17877 10217 17911 10251
rect 18429 10217 18463 10251
rect 18705 10217 18739 10251
rect 20361 10217 20395 10251
rect 20995 10217 21029 10251
rect 23029 10217 23063 10251
rect 25421 10217 25455 10251
rect 26709 10217 26743 10251
rect 29009 10217 29043 10251
rect 35449 10217 35483 10251
rect 38945 10217 38979 10251
rect 39497 10217 39531 10251
rect 40601 10217 40635 10251
rect 41797 10217 41831 10251
rect 42349 10217 42383 10251
rect 43085 10217 43119 10251
rect 46949 10217 46983 10251
rect 2605 10149 2639 10183
rect 7021 10149 7055 10183
rect 12541 10149 12575 10183
rect 15853 10149 15887 10183
rect 21281 10149 21315 10183
rect 21465 10149 21499 10183
rect 21557 10149 21591 10183
rect 22201 10149 22235 10183
rect 26065 10149 26099 10183
rect 28825 10149 28859 10183
rect 38301 10149 38335 10183
rect 41061 10149 41095 10183
rect 43729 10149 43763 10183
rect 43913 10149 43947 10183
rect 4169 10081 4203 10115
rect 5365 10081 5399 10115
rect 8401 10081 8435 10115
rect 9956 10081 9990 10115
rect 15669 10081 15703 10115
rect 35541 10081 35575 10115
rect 38117 10081 38151 10115
rect 39313 10081 39347 10115
rect 40417 10081 40451 10115
rect 42165 10081 42199 10115
rect 45836 10081 45870 10115
rect 2513 10013 2547 10047
rect 7021 10013 7055 10047
rect 7113 10013 7147 10047
rect 8677 10013 8711 10047
rect 9045 10013 9079 10047
rect 9689 10013 9723 10047
rect 12817 10013 12851 10047
rect 15945 10013 15979 10047
rect 23029 10013 23063 10047
rect 23121 10013 23155 10047
rect 25329 10013 25363 10047
rect 25513 10013 25547 10047
rect 29101 10013 29135 10047
rect 35357 10013 35391 10047
rect 38393 10013 38427 10047
rect 44005 10013 44039 10047
rect 45569 10013 45603 10047
rect 6561 9945 6595 9979
rect 7573 9945 7607 9979
rect 12265 9945 12299 9979
rect 24777 9945 24811 9979
rect 37841 9945 37875 9979
rect 43453 9945 43487 9979
rect 2053 9877 2087 9911
rect 4721 9877 4755 9911
rect 8125 9877 8159 9911
rect 11069 9877 11103 9911
rect 15393 9877 15427 9911
rect 22569 9877 22603 9911
rect 24961 9877 24995 9911
rect 28549 9877 28583 9911
rect 29561 9877 29595 9911
rect 34989 9877 35023 9911
rect 41521 9877 41555 9911
rect 44557 9877 44591 9911
rect 5365 9673 5399 9707
rect 5641 9673 5675 9707
rect 7021 9673 7055 9707
rect 8953 9673 8987 9707
rect 12633 9673 12667 9707
rect 13001 9673 13035 9707
rect 21005 9673 21039 9707
rect 21741 9673 21775 9707
rect 22569 9673 22603 9707
rect 23213 9673 23247 9707
rect 27629 9673 27663 9707
rect 28733 9673 28767 9707
rect 29929 9673 29963 9707
rect 34621 9673 34655 9707
rect 35357 9673 35391 9707
rect 37749 9673 37783 9707
rect 40785 9673 40819 9707
rect 43729 9673 43763 9707
rect 2789 9605 2823 9639
rect 3985 9605 4019 9639
rect 4905 9605 4939 9639
rect 11437 9605 11471 9639
rect 16865 9605 16899 9639
rect 21281 9605 21315 9639
rect 22937 9605 22971 9639
rect 24777 9605 24811 9639
rect 27169 9605 27203 9639
rect 29009 9605 29043 9639
rect 34345 9605 34379 9639
rect 42349 9605 42383 9639
rect 43361 9605 43395 9639
rect 44557 9605 44591 9639
rect 46949 9605 46983 9639
rect 47409 9605 47443 9639
rect 3709 9537 3743 9571
rect 12265 9537 12299 9571
rect 30113 9537 30147 9571
rect 35541 9537 35575 9571
rect 1409 9469 1443 9503
rect 1676 9469 1710 9503
rect 5457 9469 5491 9503
rect 6009 9469 6043 9503
rect 7573 9469 7607 9503
rect 7829 9469 7863 9503
rect 10425 9469 10459 9503
rect 11253 9469 11287 9503
rect 11805 9469 11839 9503
rect 14473 9469 14507 9503
rect 14565 9469 14599 9503
rect 24961 9469 24995 9503
rect 25237 9469 25271 9503
rect 28089 9469 28123 9503
rect 41429 9469 41463 9503
rect 42901 9469 42935 9503
rect 46305 9469 46339 9503
rect 46765 9469 46799 9503
rect 3433 9401 3467 9435
rect 4261 9401 4295 9435
rect 4445 9401 4479 9435
rect 4537 9401 4571 9435
rect 7389 9401 7423 9435
rect 10057 9401 10091 9435
rect 10241 9401 10275 9435
rect 14810 9401 14844 9435
rect 24041 9401 24075 9435
rect 24409 9401 24443 9435
rect 25504 9401 25538 9435
rect 30380 9401 30414 9435
rect 35808 9401 35842 9435
rect 41797 9401 41831 9435
rect 42625 9401 42659 9435
rect 44833 9401 44867 9435
rect 45109 9401 45143 9435
rect 6561 9333 6595 9367
rect 9689 9333 9723 9367
rect 10701 9333 10735 9367
rect 15945 9333 15979 9367
rect 16497 9333 16531 9367
rect 24961 9333 24995 9367
rect 25053 9333 25087 9367
rect 26617 9333 26651 9367
rect 27905 9333 27939 9367
rect 28273 9333 28307 9367
rect 31493 9333 31527 9367
rect 36921 9333 36955 9367
rect 38117 9333 38151 9367
rect 38577 9333 38611 9367
rect 39313 9333 39347 9367
rect 42165 9333 42199 9367
rect 42809 9333 42843 9367
rect 44373 9333 44407 9367
rect 45017 9333 45051 9367
rect 45569 9333 45603 9367
rect 1593 9129 1627 9163
rect 2053 9129 2087 9163
rect 2421 9129 2455 9163
rect 2789 9129 2823 9163
rect 7849 9129 7883 9163
rect 8493 9129 8527 9163
rect 8861 9129 8895 9163
rect 10425 9129 10459 9163
rect 16681 9129 16715 9163
rect 26065 9129 26099 9163
rect 27077 9129 27111 9163
rect 29653 9129 29687 9163
rect 30205 9129 30239 9163
rect 33517 9129 33551 9163
rect 34989 9129 35023 9163
rect 35633 9129 35667 9163
rect 36461 9129 36495 9163
rect 40049 9129 40083 9163
rect 41981 9129 42015 9163
rect 42441 9129 42475 9163
rect 44557 9129 44591 9163
rect 46489 9129 46523 9163
rect 4629 9061 4663 9095
rect 10149 9061 10183 9095
rect 12256 9061 12290 9095
rect 24593 9061 24627 9095
rect 24930 9061 24964 9095
rect 27169 9061 27203 9095
rect 27905 9061 27939 9095
rect 28089 9061 28123 9095
rect 29469 9061 29503 9095
rect 38945 9061 38979 9095
rect 39129 9061 39163 9095
rect 40215 9061 40249 9095
rect 40693 9061 40727 9095
rect 40785 9061 40819 9095
rect 45376 9061 45410 9095
rect 4721 8993 4755 9027
rect 6285 8993 6319 9027
rect 6725 8993 6759 9027
rect 15557 8993 15591 9027
rect 18052 8993 18086 9027
rect 22293 8993 22327 9027
rect 22560 8993 22594 9027
rect 28549 8993 28583 9027
rect 28917 8993 28951 9027
rect 29745 8993 29779 9027
rect 30481 8993 30515 9027
rect 32393 8993 32427 9027
rect 38485 8993 38519 9027
rect 40509 8993 40543 9027
rect 41797 8993 41831 9027
rect 4629 8925 4663 8959
rect 6469 8925 6503 8959
rect 11989 8925 12023 8959
rect 15301 8925 15335 8959
rect 17785 8925 17819 8959
rect 20913 8925 20947 8959
rect 24685 8925 24719 8959
rect 27077 8925 27111 8959
rect 28181 8925 28215 8959
rect 32137 8925 32171 8959
rect 36461 8925 36495 8959
rect 36553 8925 36587 8959
rect 39221 8925 39255 8959
rect 45109 8925 45143 8959
rect 4169 8857 4203 8891
rect 15025 8857 15059 8891
rect 27629 8857 27663 8891
rect 36001 8857 36035 8891
rect 38669 8857 38703 8891
rect 13369 8789 13403 8823
rect 14657 8789 14691 8823
rect 17601 8789 17635 8823
rect 19165 8789 19199 8823
rect 23673 8789 23707 8823
rect 26617 8789 26651 8823
rect 29193 8789 29227 8823
rect 31861 8789 31895 8823
rect 43085 8789 43119 8823
rect 43637 8789 43671 8823
rect 2053 8585 2087 8619
rect 3893 8585 3927 8619
rect 4537 8585 4571 8619
rect 4813 8585 4847 8619
rect 6101 8585 6135 8619
rect 8217 8585 8251 8619
rect 15025 8585 15059 8619
rect 15301 8585 15335 8619
rect 17417 8585 17451 8619
rect 17785 8585 17819 8619
rect 22477 8585 22511 8619
rect 22937 8585 22971 8619
rect 25053 8585 25087 8619
rect 28549 8585 28583 8619
rect 29561 8585 29595 8619
rect 31585 8585 31619 8619
rect 33149 8585 33183 8619
rect 36001 8585 36035 8619
rect 38945 8585 38979 8619
rect 41889 8585 41923 8619
rect 42441 8585 42475 8619
rect 43085 8585 43119 8619
rect 2329 8517 2363 8551
rect 5181 8517 5215 8551
rect 16405 8517 16439 8551
rect 23397 8517 23431 8551
rect 27537 8517 27571 8551
rect 28181 8517 28215 8551
rect 29101 8517 29135 8551
rect 30297 8517 30331 8551
rect 42809 8517 42843 8551
rect 46949 8517 46983 8551
rect 2513 8449 2547 8483
rect 15853 8449 15887 8483
rect 16865 8449 16899 8483
rect 18061 8449 18095 8483
rect 25697 8449 25731 8483
rect 30113 8449 30147 8483
rect 30849 8449 30883 8483
rect 31769 8449 31803 8483
rect 43637 8449 43671 8483
rect 47409 8449 47443 8483
rect 2780 8381 2814 8415
rect 6837 8381 6871 8415
rect 7093 8381 7127 8415
rect 12449 8381 12483 8415
rect 20361 8381 20395 8415
rect 20545 8381 20579 8415
rect 20812 8381 20846 8415
rect 23673 8381 23707 8415
rect 25973 8381 26007 8415
rect 26157 8381 26191 8415
rect 36277 8381 36311 8415
rect 36461 8381 36495 8415
rect 36717 8381 36751 8415
rect 40509 8381 40543 8415
rect 46765 8381 46799 8415
rect 6561 8313 6595 8347
rect 11529 8313 11563 8347
rect 12694 8313 12728 8347
rect 16221 8313 16255 8347
rect 16957 8313 16991 8347
rect 18328 8313 18362 8347
rect 23940 8313 23974 8347
rect 26424 8313 26458 8347
rect 30573 8313 30607 8347
rect 30757 8313 30791 8347
rect 32036 8313 32070 8347
rect 35633 8313 35667 8347
rect 39589 8313 39623 8347
rect 39957 8313 39991 8347
rect 40776 8313 40810 8347
rect 43361 8313 43395 8347
rect 43545 8313 43579 8347
rect 11805 8245 11839 8279
rect 12173 8245 12207 8279
rect 13829 8245 13863 8279
rect 16865 8245 16899 8279
rect 19441 8245 19475 8279
rect 21925 8245 21959 8279
rect 37841 8245 37875 8279
rect 38577 8245 38611 8279
rect 40325 8245 40359 8279
rect 45109 8245 45143 8279
rect 45569 8245 45603 8279
rect 1685 8041 1719 8075
rect 2605 8041 2639 8075
rect 5457 8041 5491 8075
rect 6561 8041 6595 8075
rect 12081 8041 12115 8075
rect 17601 8041 17635 8075
rect 19073 8041 19107 8075
rect 20637 8041 20671 8075
rect 24685 8041 24719 8075
rect 25421 8041 25455 8075
rect 26249 8041 26283 8075
rect 28457 8041 28491 8075
rect 30297 8041 30331 8075
rect 31769 8041 31803 8075
rect 32321 8041 32355 8075
rect 36461 8041 36495 8075
rect 40141 8041 40175 8075
rect 41613 8041 41647 8075
rect 43545 8041 43579 8075
rect 46213 8041 46247 8075
rect 4344 7973 4378 8007
rect 9956 7973 9990 8007
rect 13001 7973 13035 8007
rect 16313 7973 16347 8007
rect 16497 7973 16531 8007
rect 16957 7973 16991 8007
rect 17960 7973 17994 8007
rect 26792 7973 26826 8007
rect 28917 7973 28951 8007
rect 29377 7973 29411 8007
rect 29561 7973 29595 8007
rect 29653 7973 29687 8007
rect 36001 7973 36035 8007
rect 37994 7973 38028 8007
rect 1501 7905 1535 7939
rect 11713 7905 11747 7939
rect 17693 7905 17727 7939
rect 21189 7905 21223 7939
rect 25513 7905 25547 7939
rect 26525 7905 26559 7939
rect 30573 7905 30607 7939
rect 40489 7905 40523 7939
rect 45100 7905 45134 7939
rect 4077 7837 4111 7871
rect 9689 7837 9723 7871
rect 12909 7837 12943 7871
rect 13093 7837 13127 7871
rect 16589 7837 16623 7871
rect 21512 7837 21546 7871
rect 21649 7837 21683 7871
rect 21925 7837 21959 7871
rect 25421 7837 25455 7871
rect 37749 7837 37783 7871
rect 40233 7837 40267 7871
rect 44833 7837 44867 7871
rect 23765 7769 23799 7803
rect 29101 7769 29135 7803
rect 6929 7701 6963 7735
rect 11069 7701 11103 7735
rect 12541 7701 12575 7735
rect 15025 7701 15059 7735
rect 16037 7701 16071 7735
rect 23029 7701 23063 7735
rect 24961 7701 24995 7735
rect 27905 7701 27939 7735
rect 30757 7701 30791 7735
rect 39129 7701 39163 7735
rect 43085 7701 43119 7735
rect 4537 7497 4571 7531
rect 11253 7497 11287 7531
rect 12173 7497 12207 7531
rect 16405 7497 16439 7531
rect 17785 7497 17819 7531
rect 20269 7497 20303 7531
rect 20637 7497 20671 7531
rect 22477 7497 22511 7531
rect 24593 7497 24627 7531
rect 24869 7497 24903 7531
rect 26985 7497 27019 7531
rect 29653 7497 29687 7531
rect 30573 7497 30607 7531
rect 31033 7497 31067 7531
rect 32505 7497 32539 7531
rect 37013 7497 37047 7531
rect 37381 7497 37415 7531
rect 37933 7497 37967 7531
rect 39957 7497 39991 7531
rect 42441 7497 42475 7531
rect 5273 7429 5307 7463
rect 15025 7429 15059 7463
rect 16037 7429 16071 7463
rect 18153 7429 18187 7463
rect 20821 7429 20855 7463
rect 21741 7429 21775 7463
rect 22109 7429 22143 7463
rect 27721 7429 27755 7463
rect 11897 7361 11931 7395
rect 17417 7361 17451 7395
rect 18613 7361 18647 7395
rect 21281 7361 21315 7395
rect 21373 7361 21407 7395
rect 28181 7361 28215 7395
rect 28641 7361 28675 7395
rect 30205 7361 30239 7395
rect 31125 7361 31159 7395
rect 38393 7361 38427 7395
rect 38485 7361 38519 7395
rect 38945 7361 38979 7395
rect 9321 7293 9355 7327
rect 12449 7293 12483 7327
rect 14841 7293 14875 7327
rect 18705 7293 18739 7327
rect 19073 7293 19107 7327
rect 19901 7293 19935 7327
rect 22845 7293 22879 7327
rect 25329 7293 25363 7327
rect 25881 7293 25915 7327
rect 29929 7293 29963 7327
rect 33609 7293 33643 7327
rect 34161 7293 34195 7327
rect 40325 7293 40359 7327
rect 40969 7293 41003 7327
rect 41061 7293 41095 7327
rect 43545 7293 43579 7327
rect 43801 7293 43835 7327
rect 46765 7293 46799 7327
rect 5549 7225 5583 7259
rect 5825 7225 5859 7259
rect 9588 7225 9622 7259
rect 12716 7225 12750 7259
rect 15301 7225 15335 7259
rect 15485 7225 15519 7259
rect 15577 7225 15611 7259
rect 18613 7225 18647 7259
rect 21281 7225 21315 7259
rect 28273 7225 28307 7259
rect 31370 7225 31404 7259
rect 41306 7225 41340 7259
rect 43453 7225 43487 7259
rect 1685 7157 1719 7191
rect 4169 7157 4203 7191
rect 5089 7157 5123 7191
rect 5733 7157 5767 7191
rect 8769 7157 8803 7191
rect 9137 7157 9171 7191
rect 10701 7157 10735 7191
rect 13829 7157 13863 7191
rect 16681 7157 16715 7191
rect 23673 7157 23707 7191
rect 25513 7157 25547 7191
rect 26617 7157 26651 7191
rect 27537 7157 27571 7191
rect 28181 7157 28215 7191
rect 29101 7157 29135 7191
rect 30113 7157 30147 7191
rect 33793 7157 33827 7191
rect 37657 7157 37691 7191
rect 38393 7157 38427 7191
rect 44925 7157 44959 7191
rect 45569 7157 45603 7191
rect 46949 7157 46983 7191
rect 47409 7157 47443 7191
rect 9413 6953 9447 6987
rect 10241 6953 10275 6987
rect 11805 6953 11839 6987
rect 12541 6953 12575 6987
rect 12909 6953 12943 6987
rect 18521 6953 18555 6987
rect 29745 6953 29779 6987
rect 30665 6953 30699 6987
rect 38393 6953 38427 6987
rect 41153 6953 41187 6987
rect 21649 6885 21683 6919
rect 34161 6885 34195 6919
rect 34345 6885 34379 6919
rect 2881 6817 2915 6851
rect 6184 6817 6218 6851
rect 10057 6817 10091 6851
rect 11897 6817 11931 6851
rect 14933 6817 14967 6851
rect 15301 6817 15335 6851
rect 16405 6817 16439 6851
rect 18153 6817 18187 6851
rect 21465 6817 21499 6851
rect 24961 6817 24995 6851
rect 26525 6817 26559 6851
rect 27977 6817 28011 6851
rect 32689 6817 32723 6851
rect 43617 6817 43651 6851
rect 46101 6817 46135 6851
rect 5917 6749 5951 6783
rect 10333 6749 10367 6783
rect 11805 6749 11839 6783
rect 19809 6749 19843 6783
rect 21741 6749 21775 6783
rect 23949 6749 23983 6783
rect 27721 6749 27755 6783
rect 34437 6749 34471 6783
rect 35357 6749 35391 6783
rect 37841 6749 37875 6783
rect 43361 6749 43395 6783
rect 45845 6749 45879 6783
rect 3065 6681 3099 6715
rect 5181 6681 5215 6715
rect 8217 6681 8251 6715
rect 21189 6681 21223 6715
rect 27537 6681 27571 6715
rect 5549 6613 5583 6647
rect 7297 6613 7331 6647
rect 9781 6613 9815 6647
rect 11345 6613 11379 6647
rect 13277 6613 13311 6647
rect 15485 6613 15519 6647
rect 16589 6613 16623 6647
rect 23765 6613 23799 6647
rect 26249 6613 26283 6647
rect 26709 6613 26743 6647
rect 29101 6613 29135 6647
rect 30389 6613 30423 6647
rect 31217 6613 31251 6647
rect 32505 6613 32539 6647
rect 32873 6613 32907 6647
rect 33333 6613 33367 6647
rect 33701 6613 33735 6647
rect 33885 6613 33919 6647
rect 35265 6613 35299 6647
rect 44741 6613 44775 6647
rect 45385 6613 45419 6647
rect 47225 6613 47259 6647
rect 6285 6409 6319 6443
rect 9505 6409 9539 6443
rect 11069 6409 11103 6443
rect 11621 6409 11655 6443
rect 11989 6409 12023 6443
rect 16405 6409 16439 6443
rect 19533 6409 19567 6443
rect 21741 6409 21775 6443
rect 22477 6409 22511 6443
rect 25053 6409 25087 6443
rect 25973 6409 26007 6443
rect 27721 6409 27755 6443
rect 29101 6409 29135 6443
rect 31677 6409 31711 6443
rect 33977 6409 34011 6443
rect 42625 6409 42659 6443
rect 43821 6409 43855 6443
rect 46305 6409 46339 6443
rect 8217 6341 8251 6375
rect 13093 6341 13127 6375
rect 15485 6341 15519 6375
rect 26249 6341 26283 6375
rect 33057 6341 33091 6375
rect 35265 6341 35299 6375
rect 37749 6341 37783 6375
rect 43453 6341 43487 6375
rect 3157 6273 3191 6307
rect 8677 6273 8711 6307
rect 9689 6273 9723 6307
rect 14565 6273 14599 6307
rect 16037 6273 16071 6307
rect 19717 6273 19751 6307
rect 23489 6273 23523 6307
rect 23673 6273 23707 6307
rect 32413 6273 32447 6307
rect 33609 6273 33643 6307
rect 34713 6273 34747 6307
rect 35817 6273 35851 6307
rect 37565 6273 37599 6307
rect 43085 6273 43119 6307
rect 44281 6273 44315 6307
rect 7665 6205 7699 6239
rect 8769 6205 8803 6239
rect 9956 6205 9990 6239
rect 13369 6205 13403 6239
rect 14933 6205 14967 6239
rect 15761 6205 15795 6239
rect 23929 6205 23963 6239
rect 26801 6205 26835 6239
rect 30297 6205 30331 6239
rect 32873 6205 32907 6239
rect 35541 6205 35575 6239
rect 36185 6205 36219 6239
rect 37197 6205 37231 6239
rect 38025 6205 38059 6239
rect 39313 6205 39347 6239
rect 39865 6205 39899 6239
rect 44373 6205 44407 6239
rect 2605 6137 2639 6171
rect 3402 6137 3436 6171
rect 8033 6137 8067 6171
rect 8677 6137 8711 6171
rect 9229 6137 9263 6171
rect 13645 6137 13679 6171
rect 15301 6137 15335 6171
rect 15945 6137 15979 6171
rect 19257 6137 19291 6171
rect 19984 6137 20018 6171
rect 22017 6137 22051 6171
rect 26525 6137 26559 6171
rect 28089 6137 28123 6171
rect 30113 6137 30147 6171
rect 30564 6137 30598 6171
rect 33333 6137 33367 6171
rect 33517 6137 33551 6171
rect 36829 6137 36863 6171
rect 38209 6137 38243 6171
rect 38301 6137 38335 6171
rect 2973 6069 3007 6103
rect 4537 6069 4571 6103
rect 5917 6069 5951 6103
rect 12909 6069 12943 6103
rect 13553 6069 13587 6103
rect 14105 6069 14139 6103
rect 18061 6069 18095 6103
rect 21097 6069 21131 6103
rect 26709 6069 26743 6103
rect 27169 6069 27203 6103
rect 29653 6069 29687 6103
rect 35725 6069 35759 6103
rect 39497 6069 39531 6103
rect 44281 6069 44315 6103
rect 45937 6069 45971 6103
rect 3249 5865 3283 5899
rect 4629 5865 4663 5899
rect 7297 5865 7331 5899
rect 9965 5865 9999 5899
rect 11989 5865 12023 5899
rect 13921 5865 13955 5899
rect 14473 5865 14507 5899
rect 15485 5865 15519 5899
rect 23031 5865 23065 5899
rect 26249 5865 26283 5899
rect 33793 5865 33827 5899
rect 36277 5865 36311 5899
rect 38211 5865 38245 5899
rect 42073 5865 42107 5899
rect 43821 5865 43855 5899
rect 44189 5865 44223 5899
rect 6184 5797 6218 5831
rect 11529 5797 11563 5831
rect 12808 5797 12842 5831
rect 16028 5797 16062 5831
rect 20729 5797 20763 5831
rect 21465 5797 21499 5831
rect 21557 5797 21591 5831
rect 26792 5797 26826 5831
rect 29438 5797 29472 5831
rect 8401 5729 8435 5763
rect 10241 5729 10275 5763
rect 11345 5729 11379 5763
rect 12541 5729 12575 5763
rect 15761 5729 15795 5763
rect 18501 5729 18535 5763
rect 21281 5729 21315 5763
rect 22477 5729 22511 5763
rect 23305 5729 23339 5763
rect 26525 5729 26559 5763
rect 29193 5729 29227 5763
rect 32669 5729 32703 5763
rect 35164 5729 35198 5763
rect 37565 5729 37599 5763
rect 40693 5729 40727 5763
rect 40960 5729 40994 5763
rect 4629 5661 4663 5695
rect 4721 5661 4755 5695
rect 5917 5661 5951 5695
rect 11621 5661 11655 5695
rect 18245 5661 18279 5695
rect 22569 5661 22603 5695
rect 23029 5661 23063 5695
rect 32413 5661 32447 5695
rect 34897 5661 34931 5695
rect 37749 5661 37783 5695
rect 38209 5661 38243 5695
rect 38485 5661 38519 5695
rect 11069 5593 11103 5627
rect 21005 5593 21039 5627
rect 22109 5593 22143 5627
rect 4169 5525 4203 5559
rect 8309 5525 8343 5559
rect 8585 5525 8619 5559
rect 8953 5525 8987 5559
rect 9505 5525 9539 5559
rect 17141 5525 17175 5559
rect 18061 5525 18095 5559
rect 19625 5525 19659 5559
rect 24409 5525 24443 5559
rect 27905 5525 27939 5559
rect 30573 5525 30607 5559
rect 34345 5525 34379 5559
rect 39589 5525 39623 5559
rect 40601 5525 40635 5559
rect 3065 5321 3099 5355
rect 4537 5321 4571 5355
rect 6561 5321 6595 5355
rect 7021 5321 7055 5355
rect 9229 5321 9263 5355
rect 11069 5321 11103 5355
rect 11437 5321 11471 5355
rect 11805 5321 11839 5355
rect 13001 5321 13035 5355
rect 13553 5321 13587 5355
rect 15761 5321 15795 5355
rect 17417 5321 17451 5355
rect 17877 5321 17911 5355
rect 19073 5321 19107 5355
rect 20545 5321 20579 5355
rect 23121 5321 23155 5355
rect 23489 5321 23523 5355
rect 23765 5321 23799 5355
rect 26249 5321 26283 5355
rect 27169 5321 27203 5355
rect 27353 5321 27387 5355
rect 27629 5321 27663 5355
rect 28733 5321 28767 5355
rect 33241 5321 33275 5355
rect 35081 5321 35115 5355
rect 35449 5321 35483 5355
rect 36001 5321 36035 5355
rect 38669 5321 38703 5355
rect 8309 5253 8343 5287
rect 12633 5253 12667 5287
rect 18153 5253 18187 5287
rect 20913 5253 20947 5287
rect 29377 5253 29411 5287
rect 3157 5185 3191 5219
rect 8677 5185 8711 5219
rect 13737 5185 13771 5219
rect 18521 5185 18555 5219
rect 24133 5185 24167 5219
rect 24317 5185 24351 5219
rect 25329 5185 25363 5219
rect 26709 5185 26743 5219
rect 26801 5185 26835 5219
rect 27353 5185 27387 5219
rect 29009 5185 29043 5219
rect 29929 5185 29963 5219
rect 36093 5185 36127 5219
rect 5641 5117 5675 5151
rect 6837 5117 6871 5151
rect 7389 5117 7423 5151
rect 10701 5117 10735 5151
rect 11253 5117 11287 5151
rect 12449 5117 12483 5151
rect 14004 5117 14038 5151
rect 19809 5117 19843 5151
rect 21097 5117 21131 5151
rect 25697 5117 25731 5151
rect 31125 5117 31159 5151
rect 31309 5117 31343 5151
rect 40325 5117 40359 5151
rect 40509 5117 40543 5151
rect 3402 5049 3436 5083
rect 8861 5049 8895 5083
rect 18705 5049 18739 5083
rect 21364 5049 21398 5083
rect 26709 5049 26743 5083
rect 29653 5049 29687 5083
rect 30757 5049 30791 5083
rect 31554 5049 31588 5083
rect 33609 5049 33643 5083
rect 36338 5049 36372 5083
rect 38393 5049 38427 5083
rect 38945 5049 38979 5083
rect 39221 5049 39255 5083
rect 40754 5049 40788 5083
rect 5089 4981 5123 5015
rect 5549 4981 5583 5015
rect 5825 4981 5859 5015
rect 6285 4981 6319 5015
rect 8125 4981 8159 5015
rect 8769 4981 8803 5015
rect 10333 4981 10367 5015
rect 12173 4981 12207 5015
rect 15117 4981 15151 5015
rect 16129 4981 16163 5015
rect 18613 4981 18647 5015
rect 19625 4981 19659 5015
rect 19993 4981 20027 5015
rect 22477 4981 22511 5015
rect 24225 4981 24259 5015
rect 24685 4981 24719 5015
rect 25973 4981 26007 5015
rect 29837 4981 29871 5015
rect 30297 4981 30331 5015
rect 32689 4981 32723 5015
rect 37473 4981 37507 5015
rect 38117 4981 38151 5015
rect 39129 4981 39163 5015
rect 39681 4981 39715 5015
rect 41889 4981 41923 5015
rect 3249 4777 3283 4811
rect 4353 4777 4387 4811
rect 6101 4777 6135 4811
rect 7849 4777 7883 4811
rect 11713 4777 11747 4811
rect 12449 4777 12483 4811
rect 14197 4777 14231 4811
rect 15853 4777 15887 4811
rect 18337 4777 18371 4811
rect 20729 4777 20763 4811
rect 21925 4777 21959 4811
rect 22569 4777 22603 4811
rect 23581 4777 23615 4811
rect 24133 4777 24167 4811
rect 24961 4777 24995 4811
rect 30573 4777 30607 4811
rect 31401 4777 31435 4811
rect 32505 4777 32539 4811
rect 33609 4777 33643 4811
rect 36185 4777 36219 4811
rect 37105 4777 37139 4811
rect 38761 4777 38795 4811
rect 40601 4777 40635 4811
rect 40969 4777 41003 4811
rect 5917 4709 5951 4743
rect 8585 4709 8619 4743
rect 17141 4709 17175 4743
rect 21465 4709 21499 4743
rect 23397 4709 23431 4743
rect 23673 4709 23707 4743
rect 26341 4709 26375 4743
rect 26893 4709 26927 4743
rect 27077 4709 27111 4743
rect 27169 4709 27203 4743
rect 29009 4709 29043 4743
rect 38117 4709 38151 4743
rect 38301 4709 38335 4743
rect 6193 4641 6227 4675
rect 8677 4641 8711 4675
rect 10057 4641 10091 4675
rect 11529 4641 11563 4675
rect 15301 4641 15335 4675
rect 17233 4641 17267 4675
rect 18613 4641 18647 4675
rect 19717 4641 19751 4675
rect 24777 4641 24811 4675
rect 29460 4641 29494 4675
rect 32137 4641 32171 4675
rect 32321 4641 32355 4675
rect 33425 4641 33459 4675
rect 38393 4641 38427 4675
rect 8585 4573 8619 4607
rect 11805 4573 11839 4607
rect 14105 4573 14139 4607
rect 14289 4573 14323 4607
rect 17141 4573 17175 4607
rect 19625 4573 19659 4607
rect 21373 4573 21407 4607
rect 21557 4573 21591 4607
rect 25605 4573 25639 4607
rect 29193 4573 29227 4607
rect 5641 4505 5675 4539
rect 8125 4505 8159 4539
rect 11253 4505 11287 4539
rect 13737 4505 13771 4539
rect 20361 4505 20395 4539
rect 21005 4505 21039 4539
rect 23121 4505 23155 4539
rect 26617 4505 26651 4539
rect 31861 4505 31895 4539
rect 37473 4505 37507 4539
rect 2697 4437 2731 4471
rect 4721 4437 4755 4471
rect 5273 4437 5307 4471
rect 7481 4437 7515 4471
rect 10241 4437 10275 4471
rect 11069 4437 11103 4471
rect 12817 4437 12851 4471
rect 13185 4437 13219 4471
rect 13461 4437 13495 4471
rect 14657 4437 14691 4471
rect 15025 4437 15059 4471
rect 15485 4437 15519 4471
rect 16681 4437 16715 4471
rect 19901 4437 19935 4471
rect 24409 4437 24443 4471
rect 25881 4437 25915 4471
rect 27721 4437 27755 4471
rect 28181 4437 28215 4471
rect 32873 4437 32907 4471
rect 33241 4437 33275 4471
rect 37841 4437 37875 4471
rect 41245 4437 41279 4471
rect 6193 4233 6227 4267
rect 7205 4233 7239 4267
rect 9873 4233 9907 4267
rect 10977 4233 11011 4267
rect 11253 4233 11287 4267
rect 12817 4233 12851 4267
rect 16221 4233 16255 4267
rect 16681 4233 16715 4267
rect 17325 4233 17359 4267
rect 21005 4233 21039 4267
rect 22753 4233 22787 4267
rect 23397 4233 23431 4267
rect 24961 4233 24995 4267
rect 29009 4233 29043 4267
rect 33977 4233 34011 4267
rect 37381 4233 37415 4267
rect 38301 4233 38335 4267
rect 5273 4165 5307 4199
rect 8217 4165 8251 4199
rect 11989 4165 12023 4199
rect 5641 4097 5675 4131
rect 7941 4097 7975 4131
rect 9505 4097 9539 4131
rect 11713 4097 11747 4131
rect 13185 4097 13219 4131
rect 13369 4097 13403 4131
rect 13829 4097 13863 4131
rect 18613 4097 18647 4131
rect 19073 4097 19107 4131
rect 20545 4097 20579 4131
rect 21741 4097 21775 4131
rect 25881 4097 25915 4131
rect 28273 4097 28307 4131
rect 31401 4097 31435 4131
rect 33609 4097 33643 4131
rect 38025 4097 38059 4131
rect 39865 4097 39899 4131
rect 40969 4097 41003 4131
rect 2605 4029 2639 4063
rect 7021 4029 7055 4063
rect 8493 4029 8527 4063
rect 9689 4029 9723 4063
rect 11069 4029 11103 4063
rect 14289 4029 14323 4063
rect 14556 4029 14590 4063
rect 16773 4029 16807 4063
rect 18135 4029 18169 4063
rect 18705 4029 18739 4063
rect 19717 4029 19751 4063
rect 19993 4029 20027 4063
rect 21171 4029 21205 4063
rect 23673 4029 23707 4063
rect 24225 4029 24259 4063
rect 24777 4029 24811 4063
rect 25329 4029 25363 4063
rect 27537 4029 27571 4063
rect 29285 4029 29319 4063
rect 29837 4029 29871 4063
rect 30389 4029 30423 4063
rect 30941 4029 30975 4063
rect 40509 4029 40543 4063
rect 41245 4029 41279 4063
rect 2850 3961 2884 3995
rect 4721 3961 4755 3995
rect 5825 3961 5859 3995
rect 8769 3961 8803 3995
rect 13277 3961 13311 3995
rect 14105 3961 14139 3995
rect 21465 3961 21499 3995
rect 26249 3961 26283 3995
rect 27997 3961 28031 3995
rect 32965 3961 32999 3995
rect 33241 3961 33275 3995
rect 2513 3893 2547 3927
rect 3985 3893 4019 3927
rect 5089 3893 5123 3927
rect 5733 3893 5767 3927
rect 7665 3893 7699 3927
rect 8677 3893 8711 3927
rect 9229 3893 9263 3927
rect 10333 3893 10367 3927
rect 15669 3893 15703 3927
rect 16957 3893 16991 3927
rect 17877 3893 17911 3927
rect 18613 3893 18647 3927
rect 20177 3893 20211 3927
rect 21649 3893 21683 3927
rect 22109 3893 22143 3927
rect 23121 3893 23155 3927
rect 23857 3893 23891 3927
rect 24593 3893 24627 3927
rect 26341 3893 26375 3927
rect 26801 3893 26835 3927
rect 27711 3893 27745 3927
rect 28181 3893 28215 3927
rect 28641 3893 28675 3927
rect 29469 3893 29503 3927
rect 30573 3893 30607 3927
rect 31493 3893 31527 3927
rect 32137 3893 32171 3927
rect 32679 3893 32713 3927
rect 33149 3893 33183 3927
rect 34897 3893 34931 3927
rect 37473 3893 37507 3927
rect 39405 3893 39439 3927
rect 40325 3893 40359 3927
rect 40971 3893 41005 3927
rect 42349 3893 42383 3927
rect 2329 3689 2363 3723
rect 2973 3689 3007 3723
rect 3893 3689 3927 3723
rect 5733 3689 5767 3723
rect 6101 3689 6135 3723
rect 8217 3689 8251 3723
rect 13645 3689 13679 3723
rect 15945 3689 15979 3723
rect 17233 3689 17267 3723
rect 19257 3689 19291 3723
rect 19809 3689 19843 3723
rect 20269 3689 20303 3723
rect 21097 3689 21131 3723
rect 21557 3689 21591 3723
rect 22099 3689 22133 3723
rect 24317 3689 24351 3723
rect 25513 3689 25547 3723
rect 27077 3689 27111 3723
rect 29469 3689 29503 3723
rect 30481 3689 30515 3723
rect 32599 3689 32633 3723
rect 33977 3689 34011 3723
rect 34529 3689 34563 3723
rect 35633 3689 35667 3723
rect 37105 3689 37139 3723
rect 38301 3689 38335 3723
rect 40785 3689 40819 3723
rect 3065 3621 3099 3655
rect 5181 3621 5215 3655
rect 6438 3621 6472 3655
rect 10241 3621 10275 3655
rect 15025 3621 15059 3655
rect 16037 3621 16071 3655
rect 18122 3621 18156 3655
rect 21833 3621 21867 3655
rect 22569 3621 22603 3655
rect 23673 3621 23707 3655
rect 24133 3621 24167 3655
rect 26893 3621 26927 3655
rect 35449 3621 35483 3655
rect 37473 3621 37507 3655
rect 40049 3621 40083 3655
rect 40233 3621 40267 3655
rect 4537 3553 4571 3587
rect 5273 3553 5307 3587
rect 9137 3553 9171 3587
rect 10057 3553 10091 3587
rect 11161 3553 11195 3587
rect 11601 3553 11635 3587
rect 13829 3553 13863 3587
rect 14749 3553 14783 3587
rect 15761 3553 15795 3587
rect 17877 3553 17911 3587
rect 20913 3553 20947 3587
rect 22385 3553 22419 3587
rect 24409 3553 24443 3587
rect 25329 3553 25363 3587
rect 25973 3553 26007 3587
rect 27169 3553 27203 3587
rect 28356 3553 28390 3587
rect 30941 3553 30975 3587
rect 31953 3553 31987 3587
rect 32873 3553 32907 3587
rect 38117 3553 38151 3587
rect 39221 3553 39255 3587
rect 41245 3553 41279 3587
rect 2973 3485 3007 3519
rect 5181 3485 5215 3519
rect 6193 3485 6227 3519
rect 10333 3485 10367 3519
rect 10701 3485 10735 3519
rect 11345 3485 11379 3519
rect 22661 3485 22695 3519
rect 26341 3485 26375 3519
rect 28089 3485 28123 3519
rect 32137 3485 32171 3519
rect 32597 3485 32631 3519
rect 34989 3485 35023 3519
rect 35725 3485 35759 3519
rect 38393 3485 38427 3519
rect 39589 3485 39623 3519
rect 40325 3485 40359 3519
rect 2513 3417 2547 3451
rect 4721 3417 4755 3451
rect 9781 3417 9815 3451
rect 15485 3417 15519 3451
rect 20729 3417 20763 3451
rect 23857 3417 23891 3451
rect 26617 3417 26651 3451
rect 27629 3417 27663 3451
rect 31493 3417 31527 3451
rect 41797 3417 41831 3451
rect 1685 3349 1719 3383
rect 3525 3349 3559 3383
rect 7573 3349 7607 3383
rect 8493 3349 8527 3383
rect 9505 3349 9539 3383
rect 12725 3349 12759 3383
rect 13277 3349 13311 3383
rect 14013 3349 14047 3383
rect 16497 3349 16531 3383
rect 16865 3349 16899 3383
rect 17785 3349 17819 3383
rect 23305 3349 23339 3383
rect 24869 3349 24903 3383
rect 25145 3349 25179 3383
rect 30205 3349 30239 3383
rect 31125 3349 31159 3383
rect 35173 3349 35207 3383
rect 37841 3349 37875 3383
rect 39773 3349 39807 3383
rect 41061 3349 41095 3383
rect 41429 3349 41463 3383
rect 2329 3145 2363 3179
rect 4169 3145 4203 3179
rect 4721 3145 4755 3179
rect 5181 3145 5215 3179
rect 5549 3145 5583 3179
rect 5825 3145 5859 3179
rect 11253 3145 11287 3179
rect 14381 3145 14415 3179
rect 16405 3145 16439 3179
rect 18153 3145 18187 3179
rect 21741 3145 21775 3179
rect 23489 3145 23523 3179
rect 26065 3145 26099 3179
rect 28089 3145 28123 3179
rect 28733 3145 28767 3179
rect 29561 3145 29595 3179
rect 31125 3145 31159 3179
rect 33609 3145 33643 3179
rect 34621 3145 34655 3179
rect 36921 3145 36955 3179
rect 39681 3145 39715 3179
rect 40325 3145 40359 3179
rect 41889 3145 41923 3179
rect 16957 3077 16991 3111
rect 17417 3077 17451 3111
rect 17785 3077 17819 3111
rect 19625 3077 19659 3111
rect 22661 3077 22695 3111
rect 29101 3077 29135 3111
rect 30205 3077 30239 3111
rect 36277 3077 36311 3111
rect 18705 3009 18739 3043
rect 19809 3009 19843 3043
rect 23673 3009 23707 3043
rect 26249 3009 26283 3043
rect 26709 3009 26743 3043
rect 30757 3009 30791 3043
rect 34897 3009 34931 3043
rect 37381 3009 37415 3043
rect 40509 3009 40543 3043
rect 2789 2941 2823 2975
rect 5641 2941 5675 2975
rect 6285 2941 6319 2975
rect 7389 2941 7423 2975
rect 7656 2941 7690 2975
rect 9873 2941 9907 2975
rect 11805 2941 11839 2975
rect 12173 2941 12207 2975
rect 12449 2941 12483 2975
rect 12716 2941 12750 2975
rect 15025 2941 15059 2975
rect 15292 2941 15326 2975
rect 18429 2941 18463 2975
rect 19073 2941 19107 2975
rect 20076 2941 20110 2975
rect 22477 2941 22511 2975
rect 23940 2941 23974 2975
rect 26985 2941 27019 2975
rect 30021 2941 30055 2975
rect 30481 2941 30515 2975
rect 31677 2941 31711 2975
rect 31933 2941 31967 2975
rect 37637 2941 37671 2975
rect 3034 2873 3068 2907
rect 9413 2873 9447 2907
rect 10140 2873 10174 2907
rect 14841 2873 14875 2907
rect 18613 2873 18647 2907
rect 22109 2873 22143 2907
rect 22293 2873 22327 2907
rect 22937 2873 22971 2907
rect 31585 2873 31619 2907
rect 34345 2873 34379 2907
rect 35164 2873 35198 2907
rect 37289 2873 37323 2907
rect 40754 2873 40788 2907
rect 1593 2805 1627 2839
rect 2605 2805 2639 2839
rect 6561 2805 6595 2839
rect 7205 2805 7239 2839
rect 8769 2805 8803 2839
rect 9781 2805 9815 2839
rect 13829 2805 13863 2839
rect 21189 2805 21223 2839
rect 25053 2805 25087 2839
rect 25605 2805 25639 2839
rect 26711 2805 26745 2839
rect 30665 2805 30699 2839
rect 33057 2805 33091 2839
rect 38761 2805 38795 2839
rect 39313 2805 39347 2839
rect 2881 2601 2915 2635
rect 5733 2601 5767 2635
rect 6285 2601 6319 2635
rect 7113 2601 7147 2635
rect 7573 2601 7607 2635
rect 7849 2601 7883 2635
rect 8585 2601 8619 2635
rect 9045 2601 9079 2635
rect 11161 2601 11195 2635
rect 13001 2601 13035 2635
rect 14473 2601 14507 2635
rect 17141 2601 17175 2635
rect 17785 2601 17819 2635
rect 18061 2601 18095 2635
rect 19993 2601 20027 2635
rect 20637 2601 20671 2635
rect 22845 2601 22879 2635
rect 23489 2601 23523 2635
rect 23765 2601 23799 2635
rect 25697 2601 25731 2635
rect 26525 2601 26559 2635
rect 27905 2601 27939 2635
rect 29469 2601 29503 2635
rect 31125 2601 31159 2635
rect 31769 2601 31803 2635
rect 32229 2601 32263 2635
rect 34253 2601 34287 2635
rect 35173 2601 35207 2635
rect 37933 2601 37967 2635
rect 38025 2601 38059 2635
rect 39681 2601 39715 2635
rect 40509 2601 40543 2635
rect 1746 2533 1780 2567
rect 3525 2533 3559 2567
rect 4620 2533 4654 2567
rect 8401 2533 8435 2567
rect 10048 2533 10082 2567
rect 11713 2533 11747 2567
rect 12449 2533 12483 2567
rect 12817 2533 12851 2567
rect 14197 2533 14231 2567
rect 18858 2533 18892 2567
rect 20913 2533 20947 2567
rect 21710 2533 21744 2567
rect 24562 2533 24596 2567
rect 27261 2533 27295 2567
rect 27445 2533 27479 2567
rect 28273 2533 28307 2567
rect 29990 2533 30024 2567
rect 33140 2533 33174 2567
rect 36369 2533 36403 2567
rect 37749 2533 37783 2567
rect 38546 2533 38580 2567
rect 40969 2533 41003 2567
rect 41705 2533 41739 2567
rect 1501 2465 1535 2499
rect 3801 2465 3835 2499
rect 4353 2465 4387 2499
rect 6929 2465 6963 2499
rect 8677 2465 8711 2499
rect 12633 2465 12667 2499
rect 14289 2465 14323 2499
rect 15301 2465 15335 2499
rect 15761 2465 15795 2499
rect 16017 2465 16051 2499
rect 18613 2465 18647 2499
rect 21465 2465 21499 2499
rect 24317 2465 24351 2499
rect 27537 2465 27571 2499
rect 28457 2465 28491 2499
rect 29009 2465 29043 2499
rect 29745 2465 29779 2499
rect 32873 2465 32907 2499
rect 35449 2465 35483 2499
rect 36001 2465 36035 2499
rect 36645 2465 36679 2499
rect 37197 2465 37231 2499
rect 37933 2465 37967 2499
rect 38301 2465 38335 2499
rect 41797 2465 41831 2499
rect 42165 2465 42199 2499
rect 42717 2465 42751 2499
rect 43269 2465 43303 2499
rect 44833 2465 44867 2499
rect 6745 2397 6779 2431
rect 9505 2397 9539 2431
rect 9781 2397 9815 2431
rect 13277 2397 13311 2431
rect 41613 2397 41647 2431
rect 8125 2329 8159 2363
rect 26985 2329 27019 2363
rect 28641 2329 28675 2363
rect 36829 2329 36863 2363
rect 41245 2329 41279 2363
rect 42901 2329 42935 2363
rect 45017 2329 45051 2363
rect 14933 2261 14967 2295
rect 35633 2261 35667 2295
rect 45385 2261 45419 2295
<< metal1 >>
rect 1104 47354 48852 47376
rect 1104 47302 19606 47354
rect 19658 47302 19670 47354
rect 19722 47302 19734 47354
rect 19786 47302 19798 47354
rect 19850 47302 48852 47354
rect 1104 47280 48852 47302
rect 1104 46810 48852 46832
rect 1104 46758 4246 46810
rect 4298 46758 4310 46810
rect 4362 46758 4374 46810
rect 4426 46758 4438 46810
rect 4490 46758 34966 46810
rect 35018 46758 35030 46810
rect 35082 46758 35094 46810
rect 35146 46758 35158 46810
rect 35210 46758 48852 46810
rect 1104 46736 48852 46758
rect 1104 46266 48852 46288
rect 1104 46214 19606 46266
rect 19658 46214 19670 46266
rect 19722 46214 19734 46266
rect 19786 46214 19798 46266
rect 19850 46214 48852 46266
rect 1104 46192 48852 46214
rect 1104 45722 48852 45744
rect 1104 45670 4246 45722
rect 4298 45670 4310 45722
rect 4362 45670 4374 45722
rect 4426 45670 4438 45722
rect 4490 45670 34966 45722
rect 35018 45670 35030 45722
rect 35082 45670 35094 45722
rect 35146 45670 35158 45722
rect 35210 45670 48852 45722
rect 1104 45648 48852 45670
rect 46934 45540 46940 45552
rect 46895 45512 46940 45540
rect 46934 45500 46940 45512
rect 46992 45500 46998 45552
rect 46750 45404 46756 45416
rect 46711 45376 46756 45404
rect 46750 45364 46756 45376
rect 46808 45404 46814 45416
rect 47305 45407 47363 45413
rect 47305 45404 47317 45407
rect 46808 45376 47317 45404
rect 46808 45364 46814 45376
rect 47305 45373 47317 45376
rect 47351 45373 47363 45407
rect 47305 45367 47363 45373
rect 1104 45178 48852 45200
rect 1104 45126 19606 45178
rect 19658 45126 19670 45178
rect 19722 45126 19734 45178
rect 19786 45126 19798 45178
rect 19850 45126 48852 45178
rect 1104 45104 48852 45126
rect 1104 44634 48852 44656
rect 1104 44582 4246 44634
rect 4298 44582 4310 44634
rect 4362 44582 4374 44634
rect 4426 44582 4438 44634
rect 4490 44582 34966 44634
rect 35018 44582 35030 44634
rect 35082 44582 35094 44634
rect 35146 44582 35158 44634
rect 35210 44582 48852 44634
rect 1104 44560 48852 44582
rect 46934 44520 46940 44532
rect 46895 44492 46940 44520
rect 46934 44480 46940 44492
rect 46992 44480 46998 44532
rect 47394 44520 47400 44532
rect 47355 44492 47400 44520
rect 47394 44480 47400 44492
rect 47452 44480 47458 44532
rect 46106 44276 46112 44328
rect 46164 44316 46170 44328
rect 46753 44319 46811 44325
rect 46753 44316 46765 44319
rect 46164 44288 46765 44316
rect 46164 44276 46170 44288
rect 46753 44285 46765 44288
rect 46799 44316 46811 44319
rect 47394 44316 47400 44328
rect 46799 44288 47400 44316
rect 46799 44285 46811 44288
rect 46753 44279 46811 44285
rect 47394 44276 47400 44288
rect 47452 44276 47458 44328
rect 1104 44090 48852 44112
rect 1104 44038 19606 44090
rect 19658 44038 19670 44090
rect 19722 44038 19734 44090
rect 19786 44038 19798 44090
rect 19850 44038 48852 44090
rect 1104 44016 48852 44038
rect 1104 43546 48852 43568
rect 1104 43494 4246 43546
rect 4298 43494 4310 43546
rect 4362 43494 4374 43546
rect 4426 43494 4438 43546
rect 4490 43494 34966 43546
rect 35018 43494 35030 43546
rect 35082 43494 35094 43546
rect 35146 43494 35158 43546
rect 35210 43494 48852 43546
rect 1104 43472 48852 43494
rect 1104 43002 48852 43024
rect 1104 42950 19606 43002
rect 19658 42950 19670 43002
rect 19722 42950 19734 43002
rect 19786 42950 19798 43002
rect 19850 42950 48852 43002
rect 1104 42928 48852 42950
rect 1104 42458 48852 42480
rect 1104 42406 4246 42458
rect 4298 42406 4310 42458
rect 4362 42406 4374 42458
rect 4426 42406 4438 42458
rect 4490 42406 34966 42458
rect 35018 42406 35030 42458
rect 35082 42406 35094 42458
rect 35146 42406 35158 42458
rect 35210 42406 48852 42458
rect 1104 42384 48852 42406
rect 1104 41914 48852 41936
rect 1104 41862 19606 41914
rect 19658 41862 19670 41914
rect 19722 41862 19734 41914
rect 19786 41862 19798 41914
rect 19850 41862 48852 41914
rect 1104 41840 48852 41862
rect 46934 41800 46940 41812
rect 46895 41772 46940 41800
rect 46934 41760 46940 41772
rect 46992 41760 46998 41812
rect 46750 41664 46756 41676
rect 46711 41636 46756 41664
rect 46750 41624 46756 41636
rect 46808 41624 46814 41676
rect 1104 41370 48852 41392
rect 1104 41318 4246 41370
rect 4298 41318 4310 41370
rect 4362 41318 4374 41370
rect 4426 41318 4438 41370
rect 4490 41318 34966 41370
rect 35018 41318 35030 41370
rect 35082 41318 35094 41370
rect 35146 41318 35158 41370
rect 35210 41318 48852 41370
rect 1104 41296 48852 41318
rect 46750 40916 46756 40928
rect 46711 40888 46756 40916
rect 46750 40876 46756 40888
rect 46808 40876 46814 40928
rect 1104 40826 48852 40848
rect 1104 40774 19606 40826
rect 19658 40774 19670 40826
rect 19722 40774 19734 40826
rect 19786 40774 19798 40826
rect 19850 40774 48852 40826
rect 1104 40752 48852 40774
rect 1104 40282 48852 40304
rect 1104 40230 4246 40282
rect 4298 40230 4310 40282
rect 4362 40230 4374 40282
rect 4426 40230 4438 40282
rect 4490 40230 34966 40282
rect 35018 40230 35030 40282
rect 35082 40230 35094 40282
rect 35146 40230 35158 40282
rect 35210 40230 48852 40282
rect 1104 40208 48852 40230
rect 46290 40060 46296 40112
rect 46348 40100 46354 40112
rect 46750 40100 46756 40112
rect 46348 40072 46756 40100
rect 46348 40060 46354 40072
rect 46750 40060 46756 40072
rect 46808 40060 46814 40112
rect 1104 39738 48852 39760
rect 1104 39686 19606 39738
rect 19658 39686 19670 39738
rect 19722 39686 19734 39738
rect 19786 39686 19798 39738
rect 19850 39686 48852 39738
rect 1104 39664 48852 39686
rect 1104 39194 48852 39216
rect 1104 39142 4246 39194
rect 4298 39142 4310 39194
rect 4362 39142 4374 39194
rect 4426 39142 4438 39194
rect 4490 39142 34966 39194
rect 35018 39142 35030 39194
rect 35082 39142 35094 39194
rect 35146 39142 35158 39194
rect 35210 39142 48852 39194
rect 1104 39120 48852 39142
rect 1104 38650 48852 38672
rect 1104 38598 19606 38650
rect 19658 38598 19670 38650
rect 19722 38598 19734 38650
rect 19786 38598 19798 38650
rect 19850 38598 48852 38650
rect 1104 38576 48852 38598
rect 46934 38536 46940 38548
rect 46895 38508 46940 38536
rect 46934 38496 46940 38508
rect 46992 38496 46998 38548
rect 46750 38400 46756 38412
rect 46711 38372 46756 38400
rect 46750 38360 46756 38372
rect 46808 38360 46814 38412
rect 1104 38106 48852 38128
rect 1104 38054 4246 38106
rect 4298 38054 4310 38106
rect 4362 38054 4374 38106
rect 4426 38054 4438 38106
rect 4490 38054 34966 38106
rect 35018 38054 35030 38106
rect 35082 38054 35094 38106
rect 35146 38054 35158 38106
rect 35210 38054 48852 38106
rect 1104 38032 48852 38054
rect 45646 37612 45652 37664
rect 45704 37652 45710 37664
rect 46750 37652 46756 37664
rect 45704 37624 46756 37652
rect 45704 37612 45710 37624
rect 46750 37612 46756 37624
rect 46808 37612 46814 37664
rect 1104 37562 48852 37584
rect 1104 37510 19606 37562
rect 19658 37510 19670 37562
rect 19722 37510 19734 37562
rect 19786 37510 19798 37562
rect 19850 37510 48852 37562
rect 1104 37488 48852 37510
rect 1104 37018 48852 37040
rect 1104 36966 4246 37018
rect 4298 36966 4310 37018
rect 4362 36966 4374 37018
rect 4426 36966 4438 37018
rect 4490 36966 34966 37018
rect 35018 36966 35030 37018
rect 35082 36966 35094 37018
rect 35146 36966 35158 37018
rect 35210 36966 48852 37018
rect 1104 36944 48852 36966
rect 1104 36474 48852 36496
rect 1104 36422 19606 36474
rect 19658 36422 19670 36474
rect 19722 36422 19734 36474
rect 19786 36422 19798 36474
rect 19850 36422 48852 36474
rect 1104 36400 48852 36422
rect 1104 35930 48852 35952
rect 1104 35878 4246 35930
rect 4298 35878 4310 35930
rect 4362 35878 4374 35930
rect 4426 35878 4438 35930
rect 4490 35878 34966 35930
rect 35018 35878 35030 35930
rect 35082 35878 35094 35930
rect 35146 35878 35158 35930
rect 35210 35878 48852 35930
rect 1104 35856 48852 35878
rect 1104 35386 48852 35408
rect 1104 35334 19606 35386
rect 19658 35334 19670 35386
rect 19722 35334 19734 35386
rect 19786 35334 19798 35386
rect 19850 35334 48852 35386
rect 1104 35312 48852 35334
rect 46934 35272 46940 35284
rect 46895 35244 46940 35272
rect 46934 35232 46940 35244
rect 46992 35232 46998 35284
rect 46750 35136 46756 35148
rect 46711 35108 46756 35136
rect 46750 35096 46756 35108
rect 46808 35096 46814 35148
rect 1104 34842 48852 34864
rect 1104 34790 4246 34842
rect 4298 34790 4310 34842
rect 4362 34790 4374 34842
rect 4426 34790 4438 34842
rect 4490 34790 34966 34842
rect 35018 34790 35030 34842
rect 35082 34790 35094 34842
rect 35146 34790 35158 34842
rect 35210 34790 48852 34842
rect 1104 34768 48852 34790
rect 46750 34728 46756 34740
rect 46711 34700 46756 34728
rect 46750 34688 46756 34700
rect 46808 34688 46814 34740
rect 1104 34298 48852 34320
rect 1104 34246 19606 34298
rect 19658 34246 19670 34298
rect 19722 34246 19734 34298
rect 19786 34246 19798 34298
rect 19850 34246 48852 34298
rect 1104 34224 48852 34246
rect 1104 33754 48852 33776
rect 1104 33702 4246 33754
rect 4298 33702 4310 33754
rect 4362 33702 4374 33754
rect 4426 33702 4438 33754
rect 4490 33702 34966 33754
rect 35018 33702 35030 33754
rect 35082 33702 35094 33754
rect 35146 33702 35158 33754
rect 35210 33702 48852 33754
rect 1104 33680 48852 33702
rect 1104 33210 48852 33232
rect 1104 33158 19606 33210
rect 19658 33158 19670 33210
rect 19722 33158 19734 33210
rect 19786 33158 19798 33210
rect 19850 33158 48852 33210
rect 1104 33136 48852 33158
rect 1104 32666 48852 32688
rect 1104 32614 4246 32666
rect 4298 32614 4310 32666
rect 4362 32614 4374 32666
rect 4426 32614 4438 32666
rect 4490 32614 34966 32666
rect 35018 32614 35030 32666
rect 35082 32614 35094 32666
rect 35146 32614 35158 32666
rect 35210 32614 48852 32666
rect 1104 32592 48852 32614
rect 1104 32122 48852 32144
rect 1104 32070 19606 32122
rect 19658 32070 19670 32122
rect 19722 32070 19734 32122
rect 19786 32070 19798 32122
rect 19850 32070 48852 32122
rect 1104 32048 48852 32070
rect 46934 32008 46940 32020
rect 46895 31980 46940 32008
rect 46934 31968 46940 31980
rect 46992 31968 46998 32020
rect 46750 31872 46756 31884
rect 46711 31844 46756 31872
rect 46750 31832 46756 31844
rect 46808 31832 46814 31884
rect 42153 31671 42211 31677
rect 42153 31637 42165 31671
rect 42199 31668 42211 31671
rect 42334 31668 42340 31680
rect 42199 31640 42340 31668
rect 42199 31637 42211 31640
rect 42153 31631 42211 31637
rect 42334 31628 42340 31640
rect 42392 31628 42398 31680
rect 1104 31578 48852 31600
rect 1104 31526 4246 31578
rect 4298 31526 4310 31578
rect 4362 31526 4374 31578
rect 4426 31526 4438 31578
rect 4490 31526 34966 31578
rect 35018 31526 35030 31578
rect 35082 31526 35094 31578
rect 35146 31526 35158 31578
rect 35210 31526 48852 31578
rect 1104 31504 48852 31526
rect 41969 31263 42027 31269
rect 41969 31229 41981 31263
rect 42015 31260 42027 31263
rect 42061 31263 42119 31269
rect 42061 31260 42073 31263
rect 42015 31232 42073 31260
rect 42015 31229 42027 31232
rect 41969 31223 42027 31229
rect 42061 31229 42073 31232
rect 42107 31260 42119 31263
rect 42610 31260 42616 31272
rect 42107 31232 42616 31260
rect 42107 31229 42119 31232
rect 42061 31223 42119 31229
rect 42610 31220 42616 31232
rect 42668 31220 42674 31272
rect 42334 31201 42340 31204
rect 42328 31192 42340 31201
rect 42295 31164 42340 31192
rect 42328 31155 42340 31164
rect 42334 31152 42340 31155
rect 42392 31152 42398 31204
rect 43438 31124 43444 31136
rect 43399 31096 43444 31124
rect 43438 31084 43444 31096
rect 43496 31084 43502 31136
rect 46750 31124 46756 31136
rect 46711 31096 46756 31124
rect 46750 31084 46756 31096
rect 46808 31084 46814 31136
rect 1104 31034 48852 31056
rect 1104 30982 19606 31034
rect 19658 30982 19670 31034
rect 19722 30982 19734 31034
rect 19786 30982 19798 31034
rect 19850 30982 48852 31034
rect 1104 30960 48852 30982
rect 42334 30920 42340 30932
rect 42076 30892 42340 30920
rect 42076 30864 42104 30892
rect 42334 30880 42340 30892
rect 42392 30920 42398 30932
rect 44729 30923 44787 30929
rect 44729 30920 44741 30923
rect 42392 30892 44741 30920
rect 42392 30880 42398 30892
rect 44729 30889 44741 30892
rect 44775 30889 44787 30923
rect 44729 30883 44787 30889
rect 42058 30852 42064 30864
rect 41971 30824 42064 30852
rect 42058 30812 42064 30824
rect 42116 30812 42122 30864
rect 42245 30855 42303 30861
rect 42245 30821 42257 30855
rect 42291 30821 42303 30855
rect 42245 30815 42303 30821
rect 41874 30744 41880 30796
rect 41932 30784 41938 30796
rect 42260 30784 42288 30815
rect 43622 30793 43628 30796
rect 43616 30784 43628 30793
rect 41932 30756 43628 30784
rect 41932 30744 41938 30756
rect 43616 30747 43628 30756
rect 43622 30744 43628 30747
rect 43680 30744 43686 30796
rect 45554 30744 45560 30796
rect 45612 30784 45618 30796
rect 46089 30787 46147 30793
rect 46089 30784 46101 30787
rect 45612 30756 46101 30784
rect 45612 30744 45618 30756
rect 46089 30753 46101 30756
rect 46135 30753 46147 30787
rect 46089 30747 46147 30753
rect 42334 30716 42340 30728
rect 42295 30688 42340 30716
rect 42334 30676 42340 30688
rect 42392 30676 42398 30728
rect 42610 30676 42616 30728
rect 42668 30716 42674 30728
rect 43346 30716 43352 30728
rect 42668 30688 43352 30716
rect 42668 30676 42674 30688
rect 43346 30676 43352 30688
rect 43404 30676 43410 30728
rect 45830 30716 45836 30728
rect 45791 30688 45836 30716
rect 45830 30676 45836 30688
rect 45888 30676 45894 30728
rect 47210 30648 47216 30660
rect 47171 30620 47216 30648
rect 47210 30608 47216 30620
rect 47268 30608 47274 30660
rect 41782 30580 41788 30592
rect 41743 30552 41788 30580
rect 41782 30540 41788 30552
rect 41840 30540 41846 30592
rect 45741 30583 45799 30589
rect 45741 30549 45753 30583
rect 45787 30580 45799 30583
rect 46198 30580 46204 30592
rect 45787 30552 46204 30580
rect 45787 30549 45799 30552
rect 45741 30543 45799 30549
rect 46198 30540 46204 30552
rect 46256 30540 46262 30592
rect 1104 30490 48852 30512
rect 1104 30438 4246 30490
rect 4298 30438 4310 30490
rect 4362 30438 4374 30490
rect 4426 30438 4438 30490
rect 4490 30438 34966 30490
rect 35018 30438 35030 30490
rect 35082 30438 35094 30490
rect 35146 30438 35158 30490
rect 35210 30438 48852 30490
rect 1104 30416 48852 30438
rect 41785 30379 41843 30385
rect 41785 30345 41797 30379
rect 41831 30376 41843 30379
rect 41874 30376 41880 30388
rect 41831 30348 41880 30376
rect 41831 30345 41843 30348
rect 41785 30339 41843 30345
rect 41874 30336 41880 30348
rect 41932 30336 41938 30388
rect 42058 30376 42064 30388
rect 42019 30348 42064 30376
rect 42058 30336 42064 30348
rect 42116 30336 42122 30388
rect 42610 30376 42616 30388
rect 42571 30348 42616 30376
rect 42610 30336 42616 30348
rect 42668 30336 42674 30388
rect 45922 30336 45928 30388
rect 45980 30376 45986 30388
rect 46750 30376 46756 30388
rect 45980 30348 46756 30376
rect 45980 30336 45986 30348
rect 46750 30336 46756 30348
rect 46808 30336 46814 30388
rect 41690 30200 41696 30252
rect 41748 30240 41754 30252
rect 42628 30240 42656 30336
rect 45189 30311 45247 30317
rect 45189 30277 45201 30311
rect 45235 30308 45247 30311
rect 45554 30308 45560 30320
rect 45235 30280 45560 30308
rect 45235 30277 45247 30280
rect 45189 30271 45247 30277
rect 45554 30268 45560 30280
rect 45612 30268 45618 30320
rect 42705 30243 42763 30249
rect 42705 30240 42717 30243
rect 41748 30212 42717 30240
rect 41748 30200 41754 30212
rect 42705 30209 42717 30212
rect 42751 30209 42763 30243
rect 42705 30203 42763 30209
rect 42794 30132 42800 30184
rect 42852 30172 42858 30184
rect 42972 30175 43030 30181
rect 42972 30172 42984 30175
rect 42852 30144 42984 30172
rect 42852 30132 42858 30144
rect 42972 30141 42984 30144
rect 43018 30172 43030 30175
rect 43438 30172 43444 30184
rect 43018 30144 43444 30172
rect 43018 30141 43030 30144
rect 42972 30135 43030 30141
rect 43438 30132 43444 30144
rect 43496 30132 43502 30184
rect 45830 30132 45836 30184
rect 45888 30172 45894 30184
rect 46109 30175 46167 30181
rect 46109 30172 46121 30175
rect 45888 30144 46121 30172
rect 45888 30132 45894 30144
rect 46109 30141 46121 30144
rect 46155 30141 46167 30175
rect 46109 30135 46167 30141
rect 46198 30132 46204 30184
rect 46256 30172 46262 30184
rect 46365 30175 46423 30181
rect 46365 30172 46377 30175
rect 46256 30144 46377 30172
rect 46256 30132 46262 30144
rect 46365 30141 46377 30144
rect 46411 30141 46423 30175
rect 46365 30135 46423 30141
rect 41414 29996 41420 30048
rect 41472 30036 41478 30048
rect 44082 30036 44088 30048
rect 41472 30008 41517 30036
rect 44043 30008 44088 30036
rect 41472 29996 41478 30008
rect 44082 29996 44088 30008
rect 44140 29996 44146 30048
rect 45186 29996 45192 30048
rect 45244 30036 45250 30048
rect 45465 30039 45523 30045
rect 45465 30036 45477 30039
rect 45244 30008 45477 30036
rect 45244 29996 45250 30008
rect 45465 30005 45477 30008
rect 45511 30036 45523 30039
rect 45830 30036 45836 30048
rect 45511 30008 45836 30036
rect 45511 30005 45523 30008
rect 45465 29999 45523 30005
rect 45830 29996 45836 30008
rect 45888 29996 45894 30048
rect 47486 30036 47492 30048
rect 47447 30008 47492 30036
rect 47486 29996 47492 30008
rect 47544 29996 47550 30048
rect 1104 29946 48852 29968
rect 1104 29894 19606 29946
rect 19658 29894 19670 29946
rect 19722 29894 19734 29946
rect 19786 29894 19798 29946
rect 19850 29894 48852 29946
rect 1104 29872 48852 29894
rect 41874 29792 41880 29844
rect 41932 29832 41938 29844
rect 42245 29835 42303 29841
rect 42245 29832 42257 29835
rect 41932 29804 42257 29832
rect 41932 29792 41938 29804
rect 42245 29801 42257 29804
rect 42291 29832 42303 29835
rect 42794 29832 42800 29844
rect 42291 29804 42800 29832
rect 42291 29801 42303 29804
rect 42245 29795 42303 29801
rect 42794 29792 42800 29804
rect 42852 29792 42858 29844
rect 43346 29792 43352 29844
rect 43404 29832 43410 29844
rect 43533 29835 43591 29841
rect 43533 29832 43545 29835
rect 43404 29804 43545 29832
rect 43404 29792 43410 29804
rect 43533 29801 43545 29804
rect 43579 29801 43591 29835
rect 43533 29795 43591 29801
rect 43622 29792 43628 29844
rect 43680 29832 43686 29844
rect 43901 29835 43959 29841
rect 43901 29832 43913 29835
rect 43680 29804 43913 29832
rect 43680 29792 43686 29804
rect 43901 29801 43913 29804
rect 43947 29801 43959 29835
rect 43901 29795 43959 29801
rect 44545 29835 44603 29841
rect 44545 29801 44557 29835
rect 44591 29832 44603 29835
rect 45002 29832 45008 29844
rect 44591 29804 45008 29832
rect 44591 29801 44603 29804
rect 44545 29795 44603 29801
rect 45002 29792 45008 29804
rect 45060 29832 45066 29844
rect 45554 29832 45560 29844
rect 45060 29804 45560 29832
rect 45060 29792 45066 29804
rect 45554 29792 45560 29804
rect 45612 29832 45618 29844
rect 46569 29835 46627 29841
rect 46569 29832 46581 29835
rect 45612 29804 46581 29832
rect 45612 29792 45618 29804
rect 46569 29801 46581 29804
rect 46615 29801 46627 29835
rect 46569 29795 46627 29801
rect 39384 29767 39442 29773
rect 39384 29733 39396 29767
rect 39430 29764 39442 29767
rect 39574 29764 39580 29776
rect 39430 29736 39580 29764
rect 39430 29733 39442 29736
rect 39384 29727 39442 29733
rect 39574 29724 39580 29736
rect 39632 29724 39638 29776
rect 42061 29767 42119 29773
rect 42061 29733 42073 29767
rect 42107 29764 42119 29767
rect 42426 29764 42432 29776
rect 42107 29736 42432 29764
rect 42107 29733 42119 29736
rect 42061 29727 42119 29733
rect 42426 29724 42432 29736
rect 42484 29764 42490 29776
rect 44082 29764 44088 29776
rect 42484 29736 44088 29764
rect 42484 29724 42490 29736
rect 44082 29724 44088 29736
rect 44140 29724 44146 29776
rect 45456 29767 45514 29773
rect 45456 29733 45468 29767
rect 45502 29764 45514 29767
rect 45830 29764 45836 29776
rect 45502 29736 45836 29764
rect 45502 29733 45514 29736
rect 45456 29727 45514 29733
rect 45830 29724 45836 29736
rect 45888 29764 45894 29776
rect 47486 29764 47492 29776
rect 45888 29736 47492 29764
rect 45888 29724 45894 29736
rect 47486 29724 47492 29736
rect 47544 29724 47550 29776
rect 43346 29656 43352 29708
rect 43404 29696 43410 29708
rect 45186 29696 45192 29708
rect 43404 29668 45192 29696
rect 43404 29656 43410 29668
rect 45186 29656 45192 29668
rect 45244 29656 45250 29708
rect 39022 29588 39028 29640
rect 39080 29628 39086 29640
rect 39117 29631 39175 29637
rect 39117 29628 39129 29631
rect 39080 29600 39129 29628
rect 39080 29588 39086 29600
rect 39117 29597 39129 29600
rect 39163 29597 39175 29631
rect 39117 29591 39175 29597
rect 41414 29588 41420 29640
rect 41472 29628 41478 29640
rect 41601 29631 41659 29637
rect 41601 29628 41613 29631
rect 41472 29600 41613 29628
rect 41472 29588 41478 29600
rect 41601 29597 41613 29600
rect 41647 29628 41659 29631
rect 42058 29628 42064 29640
rect 41647 29600 42064 29628
rect 41647 29597 41659 29600
rect 41601 29591 41659 29597
rect 42058 29588 42064 29600
rect 42116 29628 42122 29640
rect 42334 29628 42340 29640
rect 42116 29600 42340 29628
rect 42116 29588 42122 29600
rect 42334 29588 42340 29600
rect 42392 29588 42398 29640
rect 40218 29452 40224 29504
rect 40276 29492 40282 29504
rect 40497 29495 40555 29501
rect 40497 29492 40509 29495
rect 40276 29464 40509 29492
rect 40276 29452 40282 29464
rect 40497 29461 40509 29464
rect 40543 29461 40555 29495
rect 40497 29455 40555 29461
rect 41785 29495 41843 29501
rect 41785 29461 41797 29495
rect 41831 29492 41843 29495
rect 42334 29492 42340 29504
rect 41831 29464 42340 29492
rect 41831 29461 41843 29464
rect 41785 29455 41843 29461
rect 42334 29452 42340 29464
rect 42392 29452 42398 29504
rect 1104 29402 48852 29424
rect 1104 29350 4246 29402
rect 4298 29350 4310 29402
rect 4362 29350 4374 29402
rect 4426 29350 4438 29402
rect 4490 29350 34966 29402
rect 35018 29350 35030 29402
rect 35082 29350 35094 29402
rect 35146 29350 35158 29402
rect 35210 29350 48852 29402
rect 1104 29328 48852 29350
rect 39574 29288 39580 29300
rect 39535 29260 39580 29288
rect 39574 29248 39580 29260
rect 39632 29248 39638 29300
rect 41785 29291 41843 29297
rect 41785 29257 41797 29291
rect 41831 29288 41843 29291
rect 41874 29288 41880 29300
rect 41831 29260 41880 29288
rect 41831 29257 41843 29260
rect 41785 29251 41843 29257
rect 41874 29248 41880 29260
rect 41932 29248 41938 29300
rect 42058 29248 42064 29300
rect 42116 29288 42122 29300
rect 43993 29291 44051 29297
rect 43993 29288 44005 29291
rect 42116 29260 44005 29288
rect 42116 29248 42122 29260
rect 43993 29257 44005 29260
rect 44039 29288 44051 29291
rect 45094 29288 45100 29300
rect 44039 29260 45100 29288
rect 44039 29257 44051 29260
rect 43993 29251 44051 29257
rect 45094 29248 45100 29260
rect 45152 29248 45158 29300
rect 45186 29248 45192 29300
rect 45244 29288 45250 29300
rect 45465 29291 45523 29297
rect 45465 29288 45477 29291
rect 45244 29260 45477 29288
rect 45244 29248 45250 29260
rect 45465 29257 45477 29260
rect 45511 29288 45523 29291
rect 45554 29288 45560 29300
rect 45511 29260 45560 29288
rect 45511 29257 45523 29260
rect 45465 29251 45523 29257
rect 45554 29248 45560 29260
rect 45612 29248 45618 29300
rect 45830 29288 45836 29300
rect 45791 29260 45836 29288
rect 45830 29248 45836 29260
rect 45888 29248 45894 29300
rect 46934 29288 46940 29300
rect 46895 29260 46940 29288
rect 46934 29248 46940 29260
rect 46992 29248 46998 29300
rect 40589 29223 40647 29229
rect 40589 29189 40601 29223
rect 40635 29220 40647 29223
rect 41322 29220 41328 29232
rect 40635 29192 41328 29220
rect 40635 29189 40647 29192
rect 40589 29183 40647 29189
rect 41322 29180 41328 29192
rect 41380 29180 41386 29232
rect 42245 29223 42303 29229
rect 42245 29189 42257 29223
rect 42291 29220 42303 29223
rect 42886 29220 42892 29232
rect 42291 29192 42892 29220
rect 42291 29189 42303 29192
rect 42245 29183 42303 29189
rect 42886 29180 42892 29192
rect 42944 29180 42950 29232
rect 44545 29223 44603 29229
rect 44545 29189 44557 29223
rect 44591 29220 44603 29223
rect 44910 29220 44916 29232
rect 44591 29192 44916 29220
rect 44591 29189 44603 29192
rect 44545 29183 44603 29189
rect 44910 29180 44916 29192
rect 44968 29180 44974 29232
rect 41230 29112 41236 29164
rect 41288 29112 41294 29164
rect 42794 29152 42800 29164
rect 42536 29124 42800 29152
rect 40218 29044 40224 29096
rect 40276 29084 40282 29096
rect 41248 29084 41276 29112
rect 40276 29056 41092 29084
rect 41248 29056 41368 29084
rect 40276 29044 40282 29056
rect 39390 28976 39396 29028
rect 39448 29016 39454 29028
rect 39945 29019 40003 29025
rect 39945 29016 39957 29019
rect 39448 28988 39957 29016
rect 39448 28976 39454 28988
rect 39945 28985 39957 28988
rect 39991 29016 40003 29019
rect 40310 29016 40316 29028
rect 39991 28988 40316 29016
rect 39991 28985 40003 28988
rect 39945 28979 40003 28985
rect 40310 28976 40316 28988
rect 40368 29016 40374 29028
rect 41064 29025 41092 29056
rect 40865 29019 40923 29025
rect 40865 29016 40877 29019
rect 40368 28988 40877 29016
rect 40368 28976 40374 28988
rect 40865 28985 40877 28988
rect 40911 28985 40923 29019
rect 40865 28979 40923 28985
rect 41049 29019 41107 29025
rect 41049 28985 41061 29019
rect 41095 28985 41107 29019
rect 41049 28979 41107 28985
rect 41141 29019 41199 29025
rect 41141 28985 41153 29019
rect 41187 29016 41199 29019
rect 41230 29016 41236 29028
rect 41187 28988 41236 29016
rect 41187 28985 41199 28988
rect 41141 28979 41199 28985
rect 41230 28976 41236 28988
rect 41288 28976 41294 29028
rect 41340 29016 41368 29056
rect 42334 29044 42340 29096
rect 42392 29084 42398 29096
rect 42536 29093 42564 29124
rect 42794 29112 42800 29124
rect 42852 29112 42858 29164
rect 45002 29152 45008 29164
rect 44963 29124 45008 29152
rect 45002 29112 45008 29124
rect 45060 29112 45066 29164
rect 42521 29087 42579 29093
rect 42521 29084 42533 29087
rect 42392 29056 42533 29084
rect 42392 29044 42398 29056
rect 42521 29053 42533 29056
rect 42567 29053 42579 29087
rect 43165 29087 43223 29093
rect 43165 29084 43177 29087
rect 42521 29047 42579 29053
rect 42720 29056 43177 29084
rect 41690 29016 41696 29028
rect 41340 28988 41696 29016
rect 41690 28976 41696 28988
rect 41748 28976 41754 29028
rect 41782 28976 41788 29028
rect 41840 29016 41846 29028
rect 42720 29025 42748 29056
rect 43165 29053 43177 29056
rect 43211 29053 43223 29087
rect 43165 29047 43223 29053
rect 44361 29087 44419 29093
rect 44361 29053 44373 29087
rect 44407 29084 44419 29087
rect 45830 29084 45836 29096
rect 44407 29056 45836 29084
rect 44407 29053 44419 29056
rect 44361 29047 44419 29053
rect 45020 29025 45048 29056
rect 45830 29044 45836 29056
rect 45888 29044 45894 29096
rect 46753 29087 46811 29093
rect 46753 29053 46765 29087
rect 46799 29053 46811 29087
rect 46753 29047 46811 29053
rect 42705 29019 42763 29025
rect 42705 29016 42717 29019
rect 41840 28988 42717 29016
rect 41840 28976 41846 28988
rect 42705 28985 42717 28988
rect 42751 28985 42763 29019
rect 42705 28979 42763 28985
rect 42797 29019 42855 29025
rect 42797 28985 42809 29019
rect 42843 29016 42855 29019
rect 43625 29019 43683 29025
rect 43625 29016 43637 29019
rect 42843 28988 43637 29016
rect 42843 28985 42855 28988
rect 42797 28979 42855 28985
rect 43625 28985 43637 28988
rect 43671 29016 43683 29019
rect 45005 29019 45063 29025
rect 43671 28988 44220 29016
rect 43671 28985 43683 28988
rect 43625 28979 43683 28985
rect 39022 28908 39028 28960
rect 39080 28948 39086 28960
rect 39117 28951 39175 28957
rect 39117 28948 39129 28951
rect 39080 28920 39129 28948
rect 39080 28908 39086 28920
rect 39117 28917 39129 28920
rect 39163 28917 39175 28951
rect 39117 28911 39175 28917
rect 39206 28908 39212 28960
rect 39264 28948 39270 28960
rect 40218 28948 40224 28960
rect 39264 28920 40224 28948
rect 39264 28908 39270 28920
rect 40218 28908 40224 28920
rect 40276 28908 40282 28960
rect 44192 28948 44220 28988
rect 45005 28985 45017 29019
rect 45051 28985 45063 29019
rect 45005 28979 45063 28985
rect 45094 28976 45100 29028
rect 45152 29016 45158 29028
rect 45462 29016 45468 29028
rect 45152 28988 45468 29016
rect 45152 28976 45158 28988
rect 45462 28976 45468 28988
rect 45520 28976 45526 29028
rect 45738 28976 45744 29028
rect 45796 29016 45802 29028
rect 46768 29016 46796 29047
rect 47302 29016 47308 29028
rect 45796 28988 47308 29016
rect 45796 28976 45802 28988
rect 47302 28976 47308 28988
rect 47360 28976 47366 29028
rect 45186 28948 45192 28960
rect 44192 28920 45192 28948
rect 45186 28908 45192 28920
rect 45244 28908 45250 28960
rect 1104 28858 48852 28880
rect 1104 28806 19606 28858
rect 19658 28806 19670 28858
rect 19722 28806 19734 28858
rect 19786 28806 19798 28858
rect 19850 28806 48852 28858
rect 1104 28784 48852 28806
rect 40310 28744 40316 28756
rect 40271 28716 40316 28744
rect 40310 28704 40316 28716
rect 40368 28704 40374 28756
rect 40957 28747 41015 28753
rect 40957 28713 40969 28747
rect 41003 28744 41015 28747
rect 41230 28744 41236 28756
rect 41003 28716 41236 28744
rect 41003 28713 41015 28716
rect 40957 28707 41015 28713
rect 41230 28704 41236 28716
rect 41288 28704 41294 28756
rect 42426 28744 42432 28756
rect 42387 28716 42432 28744
rect 42426 28704 42432 28716
rect 42484 28704 42490 28756
rect 42794 28744 42800 28756
rect 42755 28716 42800 28744
rect 42794 28704 42800 28716
rect 42852 28704 42858 28756
rect 41966 28676 41972 28688
rect 41927 28648 41972 28676
rect 41966 28636 41972 28648
rect 42024 28636 42030 28688
rect 45094 28676 45100 28688
rect 45055 28648 45100 28676
rect 45094 28636 45100 28648
rect 45152 28636 45158 28688
rect 38933 28611 38991 28617
rect 38933 28577 38945 28611
rect 38979 28608 38991 28611
rect 39022 28608 39028 28620
rect 38979 28580 39028 28608
rect 38979 28577 38991 28580
rect 38933 28571 38991 28577
rect 39022 28568 39028 28580
rect 39080 28568 39086 28620
rect 39206 28617 39212 28620
rect 39200 28608 39212 28617
rect 39167 28580 39212 28608
rect 39200 28571 39212 28580
rect 39206 28568 39212 28571
rect 39264 28568 39270 28620
rect 42058 28608 42064 28620
rect 42019 28580 42064 28608
rect 42058 28568 42064 28580
rect 42116 28568 42122 28620
rect 42886 28568 42892 28620
rect 42944 28608 42950 28620
rect 43349 28611 43407 28617
rect 43349 28608 43361 28611
rect 42944 28580 43361 28608
rect 42944 28568 42950 28580
rect 43349 28577 43361 28580
rect 43395 28608 43407 28611
rect 43990 28608 43996 28620
rect 43395 28580 43996 28608
rect 43395 28577 43407 28580
rect 43349 28571 43407 28577
rect 43990 28568 43996 28580
rect 44048 28568 44054 28620
rect 44910 28608 44916 28620
rect 44871 28580 44916 28608
rect 44910 28568 44916 28580
rect 44968 28568 44974 28620
rect 45554 28568 45560 28620
rect 45612 28608 45618 28620
rect 46382 28617 46388 28620
rect 46109 28611 46167 28617
rect 46109 28608 46121 28611
rect 45612 28580 46121 28608
rect 45612 28568 45618 28580
rect 46109 28577 46121 28580
rect 46155 28577 46167 28611
rect 46376 28608 46388 28617
rect 46343 28580 46388 28608
rect 46109 28571 46167 28577
rect 46376 28571 46388 28580
rect 46382 28568 46388 28571
rect 46440 28568 46446 28620
rect 41874 28540 41880 28552
rect 41835 28512 41880 28540
rect 41874 28500 41880 28512
rect 41932 28500 41938 28552
rect 45186 28540 45192 28552
rect 45147 28512 45192 28540
rect 45186 28500 45192 28512
rect 45244 28500 45250 28552
rect 40310 28432 40316 28484
rect 40368 28472 40374 28484
rect 45738 28472 45744 28484
rect 40368 28444 45744 28472
rect 40368 28432 40374 28444
rect 45738 28432 45744 28444
rect 45796 28432 45802 28484
rect 41506 28404 41512 28416
rect 41467 28376 41512 28404
rect 41506 28364 41512 28376
rect 41564 28364 41570 28416
rect 43530 28404 43536 28416
rect 43491 28376 43536 28404
rect 43530 28364 43536 28376
rect 43588 28364 43594 28416
rect 44634 28404 44640 28416
rect 44595 28376 44640 28404
rect 44634 28364 44640 28376
rect 44692 28364 44698 28416
rect 47486 28404 47492 28416
rect 47447 28376 47492 28404
rect 47486 28364 47492 28376
rect 47544 28364 47550 28416
rect 1104 28314 48852 28336
rect 1104 28262 4246 28314
rect 4298 28262 4310 28314
rect 4362 28262 4374 28314
rect 4426 28262 4438 28314
rect 4490 28262 34966 28314
rect 35018 28262 35030 28314
rect 35082 28262 35094 28314
rect 35146 28262 35158 28314
rect 35210 28262 48852 28314
rect 1104 28240 48852 28262
rect 39206 28160 39212 28212
rect 39264 28200 39270 28212
rect 39301 28203 39359 28209
rect 39301 28200 39313 28203
rect 39264 28172 39313 28200
rect 39264 28160 39270 28172
rect 39301 28169 39313 28172
rect 39347 28169 39359 28203
rect 43990 28200 43996 28212
rect 43951 28172 43996 28200
rect 39301 28163 39359 28169
rect 43990 28160 43996 28172
rect 44048 28160 44054 28212
rect 44453 28203 44511 28209
rect 44453 28169 44465 28203
rect 44499 28200 44511 28203
rect 45094 28200 45100 28212
rect 44499 28172 45100 28200
rect 44499 28169 44511 28172
rect 44453 28163 44511 28169
rect 45094 28160 45100 28172
rect 45152 28200 45158 28212
rect 46201 28203 46259 28209
rect 46201 28200 46213 28203
rect 45152 28172 46213 28200
rect 45152 28160 45158 28172
rect 46201 28169 46213 28172
rect 46247 28169 46259 28203
rect 46201 28163 46259 28169
rect 42886 28092 42892 28144
rect 42944 28132 42950 28144
rect 43073 28135 43131 28141
rect 43073 28132 43085 28135
rect 42944 28104 43085 28132
rect 42944 28092 42950 28104
rect 43073 28101 43085 28104
rect 43119 28101 43131 28135
rect 44729 28135 44787 28141
rect 44729 28132 44741 28135
rect 43073 28095 43131 28101
rect 43548 28104 44741 28132
rect 43162 28024 43168 28076
rect 43220 28064 43226 28076
rect 43548 28073 43576 28104
rect 44729 28101 44741 28104
rect 44775 28101 44787 28135
rect 44729 28095 44787 28101
rect 45554 28092 45560 28144
rect 45612 28132 45618 28144
rect 45833 28135 45891 28141
rect 45833 28132 45845 28135
rect 45612 28104 45845 28132
rect 45612 28092 45618 28104
rect 45833 28101 45845 28104
rect 45879 28101 45891 28135
rect 45833 28095 45891 28101
rect 43533 28067 43591 28073
rect 43533 28064 43545 28067
rect 43220 28036 43545 28064
rect 43220 28024 43226 28036
rect 43533 28033 43545 28036
rect 43579 28033 43591 28067
rect 43533 28027 43591 28033
rect 46198 28024 46204 28076
rect 46256 28064 46262 28076
rect 46569 28067 46627 28073
rect 46569 28064 46581 28067
rect 46256 28036 46581 28064
rect 46256 28024 46262 28036
rect 46569 28033 46581 28036
rect 46615 28064 46627 28067
rect 47486 28064 47492 28076
rect 46615 28036 47492 28064
rect 46615 28033 46627 28036
rect 46569 28027 46627 28033
rect 47486 28024 47492 28036
rect 47544 28024 47550 28076
rect 39114 27956 39120 28008
rect 39172 27996 39178 28008
rect 40221 27999 40279 28005
rect 40221 27996 40233 27999
rect 39172 27968 40233 27996
rect 39172 27956 39178 27968
rect 40221 27965 40233 27968
rect 40267 27996 40279 27999
rect 40497 27999 40555 28005
rect 40497 27996 40509 27999
rect 40267 27968 40509 27996
rect 40267 27965 40279 27968
rect 40221 27959 40279 27965
rect 40497 27965 40509 27968
rect 40543 27996 40555 27999
rect 41138 27996 41144 28008
rect 40543 27968 41144 27996
rect 40543 27965 40555 27968
rect 40497 27959 40555 27965
rect 41138 27956 41144 27968
rect 41196 27956 41202 28008
rect 42889 27999 42947 28005
rect 42889 27965 42901 27999
rect 42935 27996 42947 27999
rect 44542 27996 44548 28008
rect 42935 27968 43576 27996
rect 44503 27968 44548 27996
rect 42935 27965 42947 27968
rect 42889 27959 42947 27965
rect 43548 27940 43576 27968
rect 44542 27956 44548 27968
rect 44600 27996 44606 28008
rect 45097 27999 45155 28005
rect 45097 27996 45109 27999
rect 44600 27968 45109 27996
rect 44600 27956 44606 27968
rect 45097 27965 45109 27968
rect 45143 27965 45155 27999
rect 45097 27959 45155 27965
rect 45557 27999 45615 28005
rect 45557 27965 45569 27999
rect 45603 27996 45615 27999
rect 46382 27996 46388 28008
rect 45603 27968 46388 27996
rect 45603 27965 45615 27968
rect 45557 27959 45615 27965
rect 46382 27956 46388 27968
rect 46440 27996 46446 28008
rect 46934 27996 46940 28008
rect 46440 27968 46940 27996
rect 46440 27956 46446 27968
rect 40742 27931 40800 27937
rect 40742 27928 40754 27931
rect 39960 27900 40754 27928
rect 39960 27872 39988 27900
rect 40742 27897 40754 27900
rect 40788 27897 40800 27931
rect 43530 27928 43536 27940
rect 43491 27900 43536 27928
rect 40742 27891 40800 27897
rect 43530 27888 43536 27900
rect 43588 27888 43594 27940
rect 43625 27931 43683 27937
rect 43625 27897 43637 27931
rect 43671 27928 43683 27931
rect 44082 27928 44088 27940
rect 43671 27900 44088 27928
rect 43671 27897 43683 27900
rect 43625 27891 43683 27897
rect 39025 27863 39083 27869
rect 39025 27829 39037 27863
rect 39071 27860 39083 27863
rect 39114 27860 39120 27872
rect 39071 27832 39120 27860
rect 39071 27829 39083 27832
rect 39025 27823 39083 27829
rect 39114 27820 39120 27832
rect 39172 27820 39178 27872
rect 39942 27860 39948 27872
rect 39903 27832 39948 27860
rect 39942 27820 39948 27832
rect 40000 27820 40006 27872
rect 41874 27860 41880 27872
rect 41835 27832 41880 27860
rect 41874 27820 41880 27832
rect 41932 27860 41938 27872
rect 42429 27863 42487 27869
rect 42429 27860 42441 27863
rect 41932 27832 42441 27860
rect 41932 27820 41938 27832
rect 42429 27829 42441 27832
rect 42475 27829 42487 27863
rect 42429 27823 42487 27829
rect 42794 27820 42800 27872
rect 42852 27860 42858 27872
rect 43640 27860 43668 27891
rect 44082 27888 44088 27900
rect 44140 27888 44146 27940
rect 46676 27937 46704 27968
rect 46934 27956 46940 27968
rect 46992 27996 46998 28008
rect 47121 27999 47179 28005
rect 47121 27996 47133 27999
rect 46992 27968 47133 27996
rect 46992 27956 46998 27968
rect 47121 27965 47133 27968
rect 47167 27965 47179 27999
rect 47121 27959 47179 27965
rect 46661 27931 46719 27937
rect 46661 27897 46673 27931
rect 46707 27897 46719 27931
rect 46661 27891 46719 27897
rect 46753 27931 46811 27937
rect 46753 27897 46765 27931
rect 46799 27928 46811 27931
rect 47394 27928 47400 27940
rect 46799 27900 47400 27928
rect 46799 27897 46811 27900
rect 46753 27891 46811 27897
rect 42852 27832 43668 27860
rect 42852 27820 42858 27832
rect 45462 27820 45468 27872
rect 45520 27860 45526 27872
rect 46768 27860 46796 27891
rect 47394 27888 47400 27900
rect 47452 27928 47458 27940
rect 47857 27931 47915 27937
rect 47857 27928 47869 27931
rect 47452 27900 47869 27928
rect 47452 27888 47458 27900
rect 47857 27897 47869 27900
rect 47903 27897 47915 27931
rect 47857 27891 47915 27897
rect 45520 27832 46796 27860
rect 45520 27820 45526 27832
rect 1104 27770 48852 27792
rect 1104 27718 19606 27770
rect 19658 27718 19670 27770
rect 19722 27718 19734 27770
rect 19786 27718 19798 27770
rect 19850 27718 48852 27770
rect 1104 27696 48852 27718
rect 39942 27616 39948 27668
rect 40000 27656 40006 27668
rect 40497 27659 40555 27665
rect 40497 27656 40509 27659
rect 40000 27628 40509 27656
rect 40000 27616 40006 27628
rect 40497 27625 40509 27628
rect 40543 27656 40555 27659
rect 41509 27659 41567 27665
rect 41509 27656 41521 27659
rect 40543 27628 41521 27656
rect 40543 27625 40555 27628
rect 40497 27619 40555 27625
rect 41509 27625 41521 27628
rect 41555 27656 41567 27659
rect 41966 27656 41972 27668
rect 41555 27628 41972 27656
rect 41555 27625 41567 27628
rect 41509 27619 41567 27625
rect 41966 27616 41972 27628
rect 42024 27616 42030 27668
rect 42705 27659 42763 27665
rect 42705 27625 42717 27659
rect 42751 27656 42763 27659
rect 42794 27656 42800 27668
rect 42751 27628 42800 27656
rect 42751 27625 42763 27628
rect 42705 27619 42763 27625
rect 42794 27616 42800 27628
rect 42852 27616 42858 27668
rect 43073 27659 43131 27665
rect 43073 27625 43085 27659
rect 43119 27656 43131 27659
rect 43162 27656 43168 27668
rect 43119 27628 43168 27656
rect 43119 27625 43131 27628
rect 43073 27619 43131 27625
rect 43162 27616 43168 27628
rect 43220 27616 43226 27668
rect 44729 27659 44787 27665
rect 44729 27625 44741 27659
rect 44775 27656 44787 27659
rect 44910 27656 44916 27668
rect 44775 27628 44916 27656
rect 44775 27625 44787 27628
rect 44729 27619 44787 27625
rect 44910 27616 44916 27628
rect 44968 27616 44974 27668
rect 46934 27656 46940 27668
rect 46895 27628 46940 27656
rect 46934 27616 46940 27628
rect 46992 27616 46998 27668
rect 39390 27597 39396 27600
rect 39384 27588 39396 27597
rect 39351 27560 39396 27588
rect 39384 27551 39396 27560
rect 39390 27548 39396 27551
rect 39448 27548 39454 27600
rect 41414 27548 41420 27600
rect 41472 27588 41478 27600
rect 42153 27591 42211 27597
rect 42153 27588 42165 27591
rect 41472 27560 42165 27588
rect 41472 27548 41478 27560
rect 42153 27557 42165 27560
rect 42199 27588 42211 27591
rect 43254 27588 43260 27600
rect 42199 27560 43260 27588
rect 42199 27557 42211 27560
rect 42153 27551 42211 27557
rect 43254 27548 43260 27560
rect 43312 27548 43318 27600
rect 41506 27480 41512 27532
rect 41564 27520 41570 27532
rect 41969 27523 42027 27529
rect 41969 27520 41981 27523
rect 41564 27492 41981 27520
rect 41564 27480 41570 27492
rect 41969 27489 41981 27492
rect 42015 27489 42027 27523
rect 41969 27483 42027 27489
rect 44085 27523 44143 27529
rect 44085 27489 44097 27523
rect 44131 27520 44143 27523
rect 44634 27520 44640 27532
rect 44131 27492 44640 27520
rect 44131 27489 44143 27492
rect 44085 27483 44143 27489
rect 44634 27480 44640 27492
rect 44692 27480 44698 27532
rect 45554 27520 45560 27532
rect 45515 27492 45560 27520
rect 45554 27480 45560 27492
rect 45612 27480 45618 27532
rect 45824 27523 45882 27529
rect 45824 27489 45836 27523
rect 45870 27520 45882 27523
rect 46198 27520 46204 27532
rect 45870 27492 46204 27520
rect 45870 27489 45882 27492
rect 45824 27483 45882 27489
rect 46198 27480 46204 27492
rect 46256 27480 46262 27532
rect 37737 27455 37795 27461
rect 37737 27421 37749 27455
rect 37783 27452 37795 27455
rect 38102 27452 38108 27464
rect 37783 27424 38108 27452
rect 37783 27421 37795 27424
rect 37737 27415 37795 27421
rect 38102 27412 38108 27424
rect 38160 27412 38166 27464
rect 39114 27452 39120 27464
rect 39075 27424 39120 27452
rect 39114 27412 39120 27424
rect 39172 27412 39178 27464
rect 41141 27455 41199 27461
rect 41141 27421 41153 27455
rect 41187 27452 41199 27455
rect 42242 27452 42248 27464
rect 41187 27424 42248 27452
rect 41187 27421 41199 27424
rect 41141 27415 41199 27421
rect 42242 27412 42248 27424
rect 42300 27412 42306 27464
rect 41690 27384 41696 27396
rect 41651 27356 41696 27384
rect 41690 27344 41696 27356
rect 41748 27344 41754 27396
rect 38286 27316 38292 27328
rect 38247 27288 38292 27316
rect 38286 27276 38292 27288
rect 38344 27276 38350 27328
rect 43901 27319 43959 27325
rect 43901 27285 43913 27319
rect 43947 27316 43959 27319
rect 44266 27316 44272 27328
rect 43947 27288 44272 27316
rect 43947 27285 43959 27288
rect 43901 27279 43959 27285
rect 44266 27276 44272 27288
rect 44324 27276 44330 27328
rect 45097 27319 45155 27325
rect 45097 27285 45109 27319
rect 45143 27316 45155 27319
rect 45186 27316 45192 27328
rect 45143 27288 45192 27316
rect 45143 27285 45155 27288
rect 45097 27279 45155 27285
rect 45186 27276 45192 27288
rect 45244 27276 45250 27328
rect 1104 27226 48852 27248
rect 1104 27174 4246 27226
rect 4298 27174 4310 27226
rect 4362 27174 4374 27226
rect 4426 27174 4438 27226
rect 4490 27174 34966 27226
rect 35018 27174 35030 27226
rect 35082 27174 35094 27226
rect 35146 27174 35158 27226
rect 35210 27174 48852 27226
rect 1104 27152 48852 27174
rect 38102 27112 38108 27124
rect 38063 27084 38108 27112
rect 38102 27072 38108 27084
rect 38160 27072 38166 27124
rect 38378 27112 38384 27124
rect 38339 27084 38384 27112
rect 38378 27072 38384 27084
rect 38436 27072 38442 27124
rect 39390 27072 39396 27124
rect 39448 27112 39454 27124
rect 39669 27115 39727 27121
rect 39669 27112 39681 27115
rect 39448 27084 39681 27112
rect 39448 27072 39454 27084
rect 39669 27081 39681 27084
rect 39715 27081 39727 27115
rect 43254 27112 43260 27124
rect 43215 27084 43260 27112
rect 39669 27075 39727 27081
rect 43254 27072 43260 27084
rect 43312 27072 43318 27124
rect 44634 27072 44640 27124
rect 44692 27112 44698 27124
rect 44821 27115 44879 27121
rect 44821 27112 44833 27115
rect 44692 27084 44833 27112
rect 44692 27072 44698 27084
rect 44821 27081 44833 27084
rect 44867 27081 44879 27115
rect 45554 27112 45560 27124
rect 45515 27084 45560 27112
rect 44821 27075 44879 27081
rect 45554 27072 45560 27084
rect 45612 27072 45618 27124
rect 46198 27072 46204 27124
rect 46256 27112 46262 27124
rect 46293 27115 46351 27121
rect 46293 27112 46305 27115
rect 46256 27084 46305 27112
rect 46256 27072 46262 27084
rect 46293 27081 46305 27084
rect 46339 27081 46351 27115
rect 46293 27075 46351 27081
rect 38120 26976 38148 27072
rect 43898 27044 43904 27056
rect 43859 27016 43904 27044
rect 43898 27004 43904 27016
rect 43956 27004 43962 27056
rect 38749 26979 38807 26985
rect 38749 26976 38761 26979
rect 38120 26948 38761 26976
rect 38749 26945 38761 26948
rect 38795 26945 38807 26979
rect 44266 26976 44272 26988
rect 44227 26948 44272 26976
rect 38749 26939 38807 26945
rect 44266 26936 44272 26948
rect 44324 26936 44330 26988
rect 35805 26911 35863 26917
rect 35805 26877 35817 26911
rect 35851 26877 35863 26911
rect 35805 26871 35863 26877
rect 35713 26775 35771 26781
rect 35713 26741 35725 26775
rect 35759 26772 35771 26775
rect 35820 26772 35848 26871
rect 38654 26868 38660 26920
rect 38712 26908 38718 26920
rect 39114 26908 39120 26920
rect 38712 26880 39120 26908
rect 38712 26868 38718 26880
rect 39114 26868 39120 26880
rect 39172 26908 39178 26920
rect 39301 26911 39359 26917
rect 39301 26908 39313 26911
rect 39172 26880 39313 26908
rect 39172 26868 39178 26880
rect 39301 26877 39313 26880
rect 39347 26908 39359 26911
rect 41141 26911 41199 26917
rect 41141 26908 41153 26911
rect 39347 26880 41153 26908
rect 39347 26877 39359 26880
rect 39301 26871 39359 26877
rect 41141 26877 41153 26880
rect 41187 26908 41199 26911
rect 41325 26911 41383 26917
rect 41325 26908 41337 26911
rect 41187 26880 41337 26908
rect 41187 26877 41199 26880
rect 41141 26871 41199 26877
rect 41325 26877 41337 26880
rect 41371 26908 41383 26911
rect 41414 26908 41420 26920
rect 41371 26880 41420 26908
rect 41371 26877 41383 26880
rect 41325 26871 41383 26877
rect 41414 26868 41420 26880
rect 41472 26868 41478 26920
rect 35894 26800 35900 26852
rect 35952 26840 35958 26852
rect 36072 26843 36130 26849
rect 36072 26840 36084 26843
rect 35952 26812 36084 26840
rect 35952 26800 35958 26812
rect 36072 26809 36084 26812
rect 36118 26840 36130 26843
rect 38378 26840 38384 26852
rect 36118 26812 38384 26840
rect 36118 26809 36130 26812
rect 36072 26803 36130 26809
rect 38378 26800 38384 26812
rect 38436 26840 38442 26852
rect 38933 26843 38991 26849
rect 38933 26840 38945 26843
rect 38436 26812 38945 26840
rect 38436 26800 38442 26812
rect 38933 26809 38945 26812
rect 38979 26809 38991 26843
rect 38933 26803 38991 26809
rect 40865 26843 40923 26849
rect 40865 26809 40877 26843
rect 40911 26840 40923 26843
rect 41570 26843 41628 26849
rect 41570 26840 41582 26843
rect 40911 26812 41582 26840
rect 40911 26809 40923 26812
rect 40865 26803 40923 26809
rect 41570 26809 41582 26812
rect 41616 26840 41628 26843
rect 41874 26840 41880 26852
rect 41616 26812 41880 26840
rect 41616 26809 41628 26812
rect 41570 26803 41628 26809
rect 41874 26800 41880 26812
rect 41932 26800 41938 26852
rect 44082 26800 44088 26852
rect 44140 26840 44146 26852
rect 44453 26843 44511 26849
rect 44453 26840 44465 26843
rect 44140 26812 44465 26840
rect 44140 26800 44146 26812
rect 44453 26809 44465 26812
rect 44499 26840 44511 26843
rect 44499 26812 45324 26840
rect 44499 26809 44511 26812
rect 44453 26803 44511 26809
rect 45296 26784 45324 26812
rect 35986 26772 35992 26784
rect 35759 26744 35992 26772
rect 35759 26741 35771 26744
rect 35713 26735 35771 26741
rect 35986 26732 35992 26744
rect 36044 26732 36050 26784
rect 37182 26772 37188 26784
rect 37143 26744 37188 26772
rect 37182 26732 37188 26744
rect 37240 26732 37246 26784
rect 38286 26732 38292 26784
rect 38344 26772 38350 26784
rect 38841 26775 38899 26781
rect 38841 26772 38853 26775
rect 38344 26744 38853 26772
rect 38344 26732 38350 26744
rect 38841 26741 38853 26744
rect 38887 26741 38899 26775
rect 38841 26735 38899 26741
rect 42426 26732 42432 26784
rect 42484 26772 42490 26784
rect 42705 26775 42763 26781
rect 42705 26772 42717 26775
rect 42484 26744 42717 26772
rect 42484 26732 42490 26744
rect 42705 26741 42717 26744
rect 42751 26741 42763 26775
rect 42705 26735 42763 26741
rect 43717 26775 43775 26781
rect 43717 26741 43729 26775
rect 43763 26772 43775 26775
rect 44361 26775 44419 26781
rect 44361 26772 44373 26775
rect 43763 26744 44373 26772
rect 43763 26741 43775 26744
rect 43717 26735 43775 26741
rect 44361 26741 44373 26744
rect 44407 26772 44419 26775
rect 45002 26772 45008 26784
rect 44407 26744 45008 26772
rect 44407 26741 44419 26744
rect 44361 26735 44419 26741
rect 45002 26732 45008 26744
rect 45060 26732 45066 26784
rect 45278 26772 45284 26784
rect 45239 26744 45284 26772
rect 45278 26732 45284 26744
rect 45336 26732 45342 26784
rect 1104 26682 48852 26704
rect 1104 26630 19606 26682
rect 19658 26630 19670 26682
rect 19722 26630 19734 26682
rect 19786 26630 19798 26682
rect 19850 26630 48852 26682
rect 1104 26608 48852 26630
rect 35894 26568 35900 26580
rect 35855 26540 35900 26568
rect 35894 26528 35900 26540
rect 35952 26528 35958 26580
rect 38378 26568 38384 26580
rect 38339 26540 38384 26568
rect 38378 26528 38384 26540
rect 38436 26528 38442 26580
rect 38562 26528 38568 26580
rect 38620 26568 38626 26580
rect 39853 26571 39911 26577
rect 39853 26568 39865 26571
rect 38620 26540 39865 26568
rect 38620 26528 38626 26540
rect 39853 26537 39865 26540
rect 39899 26537 39911 26571
rect 39853 26531 39911 26537
rect 41233 26571 41291 26577
rect 41233 26537 41245 26571
rect 41279 26568 41291 26571
rect 41506 26568 41512 26580
rect 41279 26540 41512 26568
rect 41279 26537 41291 26540
rect 41233 26531 41291 26537
rect 41506 26528 41512 26540
rect 41564 26528 41570 26580
rect 41874 26500 41880 26512
rect 41835 26472 41880 26500
rect 41874 26460 41880 26472
rect 41932 26460 41938 26512
rect 44726 26460 44732 26512
rect 44784 26500 44790 26512
rect 45097 26503 45155 26509
rect 45097 26500 45109 26503
rect 44784 26472 45109 26500
rect 44784 26460 44790 26472
rect 45097 26469 45109 26472
rect 45143 26469 45155 26503
rect 45097 26463 45155 26469
rect 38746 26441 38752 26444
rect 38740 26395 38752 26441
rect 38804 26432 38810 26444
rect 40497 26435 40555 26441
rect 40497 26432 40509 26435
rect 38804 26404 40509 26432
rect 38746 26392 38752 26395
rect 38804 26392 38810 26404
rect 40497 26401 40509 26404
rect 40543 26432 40555 26435
rect 40678 26432 40684 26444
rect 40543 26404 40684 26432
rect 40543 26401 40555 26404
rect 40497 26395 40555 26401
rect 40678 26392 40684 26404
rect 40736 26392 40742 26444
rect 43346 26432 43352 26444
rect 43307 26404 43352 26432
rect 43346 26392 43352 26404
rect 43404 26432 43410 26444
rect 43898 26432 43904 26444
rect 43404 26404 43904 26432
rect 43404 26392 43410 26404
rect 43898 26392 43904 26404
rect 43956 26392 43962 26444
rect 44542 26392 44548 26444
rect 44600 26432 44606 26444
rect 44913 26435 44971 26441
rect 44913 26432 44925 26435
rect 44600 26404 44925 26432
rect 44600 26392 44606 26404
rect 44913 26401 44925 26404
rect 44959 26401 44971 26435
rect 44913 26395 44971 26401
rect 45554 26392 45560 26444
rect 45612 26432 45618 26444
rect 46109 26435 46167 26441
rect 46109 26432 46121 26435
rect 45612 26404 46121 26432
rect 45612 26392 45618 26404
rect 46109 26401 46121 26404
rect 46155 26401 46167 26435
rect 46109 26395 46167 26401
rect 46376 26435 46434 26441
rect 46376 26401 46388 26435
rect 46422 26432 46434 26435
rect 46842 26432 46848 26444
rect 46422 26404 46848 26432
rect 46422 26401 46434 26404
rect 46376 26395 46434 26401
rect 46842 26392 46848 26404
rect 46900 26392 46906 26444
rect 38473 26367 38531 26373
rect 38473 26333 38485 26367
rect 38519 26333 38531 26367
rect 38473 26327 38531 26333
rect 41877 26367 41935 26373
rect 41877 26333 41889 26367
rect 41923 26333 41935 26367
rect 41877 26327 41935 26333
rect 38488 26296 38516 26327
rect 37200 26268 38516 26296
rect 36722 26228 36728 26240
rect 36683 26200 36728 26228
rect 36722 26188 36728 26200
rect 36780 26188 36786 26240
rect 37090 26188 37096 26240
rect 37148 26228 37154 26240
rect 37200 26228 37228 26268
rect 37148 26200 37228 26228
rect 38488 26228 38516 26268
rect 41322 26256 41328 26308
rect 41380 26296 41386 26308
rect 41417 26299 41475 26305
rect 41417 26296 41429 26299
rect 41380 26268 41429 26296
rect 41380 26256 41386 26268
rect 41417 26265 41429 26268
rect 41463 26265 41475 26299
rect 41417 26259 41475 26265
rect 41598 26256 41604 26308
rect 41656 26296 41662 26308
rect 41892 26296 41920 26327
rect 41966 26324 41972 26376
rect 42024 26364 42030 26376
rect 44453 26367 44511 26373
rect 42024 26336 42069 26364
rect 42024 26324 42030 26336
rect 44453 26333 44465 26367
rect 44499 26364 44511 26367
rect 45186 26364 45192 26376
rect 44499 26336 45192 26364
rect 44499 26333 44511 26336
rect 44453 26327 44511 26333
rect 45186 26324 45192 26336
rect 45244 26324 45250 26376
rect 43533 26299 43591 26305
rect 43533 26296 43545 26299
rect 41656 26268 43545 26296
rect 41656 26256 41662 26268
rect 43533 26265 43545 26268
rect 43579 26265 43591 26299
rect 43533 26259 43591 26265
rect 38654 26228 38660 26240
rect 38488 26200 38660 26228
rect 37148 26188 37154 26200
rect 38654 26188 38660 26200
rect 38712 26188 38718 26240
rect 42426 26228 42432 26240
rect 42387 26200 42432 26228
rect 42426 26188 42432 26200
rect 42484 26188 42490 26240
rect 44634 26228 44640 26240
rect 44595 26200 44640 26228
rect 44634 26188 44640 26200
rect 44692 26188 44698 26240
rect 47486 26228 47492 26240
rect 47447 26200 47492 26228
rect 47486 26188 47492 26200
rect 47544 26188 47550 26240
rect 1104 26138 48852 26160
rect 1104 26086 4246 26138
rect 4298 26086 4310 26138
rect 4362 26086 4374 26138
rect 4426 26086 4438 26138
rect 4490 26086 34966 26138
rect 35018 26086 35030 26138
rect 35082 26086 35094 26138
rect 35146 26086 35158 26138
rect 35210 26086 48852 26138
rect 1104 26064 48852 26086
rect 38013 26027 38071 26033
rect 38013 25993 38025 26027
rect 38059 26024 38071 26027
rect 38378 26024 38384 26036
rect 38059 25996 38384 26024
rect 38059 25993 38071 25996
rect 38013 25987 38071 25993
rect 38378 25984 38384 25996
rect 38436 25984 38442 26036
rect 38654 26024 38660 26036
rect 38615 25996 38660 26024
rect 38654 25984 38660 25996
rect 38712 25984 38718 26036
rect 38746 25984 38752 26036
rect 38804 26024 38810 26036
rect 38933 26027 38991 26033
rect 38933 26024 38945 26027
rect 38804 25996 38945 26024
rect 38804 25984 38810 25996
rect 38933 25993 38945 25996
rect 38979 25993 38991 26027
rect 41598 26024 41604 26036
rect 41559 25996 41604 26024
rect 38933 25987 38991 25993
rect 41598 25984 41604 25996
rect 41656 25984 41662 26036
rect 41966 25984 41972 26036
rect 42024 26024 42030 26036
rect 43717 26027 43775 26033
rect 43717 26024 43729 26027
rect 42024 25996 43729 26024
rect 42024 25984 42030 25996
rect 43717 25993 43729 25996
rect 43763 25993 43775 26027
rect 45002 26024 45008 26036
rect 44963 25996 45008 26024
rect 43717 25987 43775 25993
rect 45002 25984 45008 25996
rect 45060 25984 45066 26036
rect 45554 25984 45560 26036
rect 45612 26024 45618 26036
rect 45833 26027 45891 26033
rect 45833 26024 45845 26027
rect 45612 25996 45845 26024
rect 45612 25984 45618 25996
rect 45833 25993 45845 25996
rect 45879 25993 45891 26027
rect 45833 25987 45891 25993
rect 40586 25956 40592 25968
rect 40547 25928 40592 25956
rect 40586 25916 40592 25928
rect 40644 25916 40650 25968
rect 41414 25916 41420 25968
rect 41472 25956 41478 25968
rect 42153 25959 42211 25965
rect 42153 25956 42165 25959
rect 41472 25928 42165 25956
rect 41472 25916 41478 25928
rect 42153 25925 42165 25928
rect 42199 25956 42211 25959
rect 42242 25956 42248 25968
rect 42199 25928 42248 25956
rect 42199 25925 42211 25928
rect 42153 25919 42211 25925
rect 42242 25916 42248 25928
rect 42300 25956 42306 25968
rect 42300 25928 42380 25956
rect 42300 25916 42306 25928
rect 40678 25848 40684 25900
rect 40736 25888 40742 25900
rect 42352 25897 42380 25928
rect 44542 25916 44548 25968
rect 44600 25956 44606 25968
rect 46201 25959 46259 25965
rect 46201 25956 46213 25959
rect 44600 25928 46213 25956
rect 44600 25916 44606 25928
rect 46201 25925 46213 25928
rect 46247 25925 46259 25959
rect 46201 25919 46259 25925
rect 41141 25891 41199 25897
rect 41141 25888 41153 25891
rect 40736 25860 41153 25888
rect 40736 25848 40742 25860
rect 41141 25857 41153 25860
rect 41187 25857 41199 25891
rect 41141 25851 41199 25857
rect 42337 25891 42395 25897
rect 42337 25857 42349 25891
rect 42383 25857 42395 25891
rect 42337 25851 42395 25857
rect 35986 25780 35992 25832
rect 36044 25820 36050 25832
rect 36633 25823 36691 25829
rect 36633 25820 36645 25823
rect 36044 25792 36645 25820
rect 36044 25780 36050 25792
rect 36464 25752 36492 25792
rect 36633 25789 36645 25792
rect 36679 25789 36691 25823
rect 36633 25783 36691 25789
rect 36722 25780 36728 25832
rect 36780 25820 36786 25832
rect 36900 25823 36958 25829
rect 36900 25820 36912 25823
rect 36780 25792 36912 25820
rect 36780 25780 36786 25792
rect 36900 25789 36912 25792
rect 36946 25820 36958 25823
rect 38562 25820 38568 25832
rect 36946 25792 38568 25820
rect 36946 25789 36958 25792
rect 36900 25783 36958 25789
rect 38562 25780 38568 25792
rect 38620 25780 38626 25832
rect 39945 25823 40003 25829
rect 39945 25789 39957 25823
rect 39991 25820 40003 25823
rect 39991 25792 41092 25820
rect 39991 25789 40003 25792
rect 39945 25783 40003 25789
rect 37090 25752 37096 25764
rect 36464 25724 37096 25752
rect 35986 25684 35992 25696
rect 35947 25656 35992 25684
rect 35986 25644 35992 25656
rect 36044 25644 36050 25696
rect 36354 25644 36360 25696
rect 36412 25684 36418 25696
rect 36464 25693 36492 25724
rect 37090 25712 37096 25724
rect 37148 25712 37154 25764
rect 41064 25761 41092 25792
rect 44634 25780 44640 25832
rect 44692 25820 44698 25832
rect 44821 25823 44879 25829
rect 44821 25820 44833 25823
rect 44692 25792 44833 25820
rect 44692 25780 44698 25792
rect 44821 25789 44833 25792
rect 44867 25789 44879 25823
rect 44821 25783 44879 25789
rect 46198 25780 46204 25832
rect 46256 25820 46262 25832
rect 46477 25823 46535 25829
rect 46477 25820 46489 25823
rect 46256 25792 46489 25820
rect 46256 25780 46262 25792
rect 46477 25789 46489 25792
rect 46523 25820 46535 25823
rect 47121 25823 47179 25829
rect 47121 25820 47133 25823
rect 46523 25792 47133 25820
rect 46523 25789 46535 25792
rect 46477 25783 46535 25789
rect 47121 25789 47133 25792
rect 47167 25820 47179 25823
rect 47486 25820 47492 25832
rect 47167 25792 47492 25820
rect 47167 25789 47179 25792
rect 47121 25783 47179 25789
rect 47486 25780 47492 25792
rect 47544 25780 47550 25832
rect 39209 25755 39267 25761
rect 39209 25721 39221 25755
rect 39255 25752 39267 25755
rect 40313 25755 40371 25761
rect 40313 25752 40325 25755
rect 39255 25724 40325 25752
rect 39255 25721 39267 25724
rect 39209 25715 39267 25721
rect 40313 25721 40325 25724
rect 40359 25752 40371 25755
rect 40865 25755 40923 25761
rect 40865 25752 40877 25755
rect 40359 25724 40877 25752
rect 40359 25721 40371 25724
rect 40313 25715 40371 25721
rect 40865 25721 40877 25724
rect 40911 25721 40923 25755
rect 40865 25715 40923 25721
rect 41049 25755 41107 25761
rect 41049 25721 41061 25755
rect 41095 25752 41107 25755
rect 41322 25752 41328 25764
rect 41095 25724 41328 25752
rect 41095 25721 41107 25724
rect 41049 25715 41107 25721
rect 41322 25712 41328 25724
rect 41380 25712 41386 25764
rect 42426 25712 42432 25764
rect 42484 25752 42490 25764
rect 42604 25755 42662 25761
rect 42604 25752 42616 25755
rect 42484 25724 42616 25752
rect 42484 25712 42490 25724
rect 42604 25721 42616 25724
rect 42650 25752 42662 25755
rect 43530 25752 43536 25764
rect 42650 25724 43536 25752
rect 42650 25721 42662 25724
rect 42604 25715 42662 25721
rect 43530 25712 43536 25724
rect 43588 25712 43594 25764
rect 45557 25755 45615 25761
rect 45557 25721 45569 25755
rect 45603 25752 45615 25755
rect 46753 25755 46811 25761
rect 45603 25724 46704 25752
rect 45603 25721 45615 25724
rect 45557 25715 45615 25721
rect 36449 25687 36507 25693
rect 36449 25684 36461 25687
rect 36412 25656 36461 25684
rect 36412 25644 36418 25656
rect 36449 25653 36461 25656
rect 36495 25653 36507 25687
rect 36449 25647 36507 25653
rect 44637 25687 44695 25693
rect 44637 25653 44649 25687
rect 44683 25684 44695 25687
rect 44726 25684 44732 25696
rect 44683 25656 44732 25684
rect 44683 25653 44695 25656
rect 44637 25647 44695 25653
rect 44726 25644 44732 25656
rect 44784 25644 44790 25696
rect 46676 25693 46704 25724
rect 46753 25721 46765 25755
rect 46799 25752 46811 25755
rect 46799 25724 47440 25752
rect 46799 25721 46811 25724
rect 46753 25715 46811 25721
rect 47412 25696 47440 25724
rect 46661 25687 46719 25693
rect 46661 25653 46673 25687
rect 46707 25684 46719 25687
rect 46842 25684 46848 25696
rect 46707 25656 46848 25684
rect 46707 25653 46719 25656
rect 46661 25647 46719 25653
rect 46842 25644 46848 25656
rect 46900 25644 46906 25696
rect 47394 25644 47400 25696
rect 47452 25684 47458 25696
rect 47489 25687 47547 25693
rect 47489 25684 47501 25687
rect 47452 25656 47501 25684
rect 47452 25644 47458 25656
rect 47489 25653 47501 25656
rect 47535 25653 47547 25687
rect 47489 25647 47547 25653
rect 1104 25594 48852 25616
rect 1104 25542 19606 25594
rect 19658 25542 19670 25594
rect 19722 25542 19734 25594
rect 19786 25542 19798 25594
rect 19850 25542 48852 25594
rect 1104 25520 48852 25542
rect 35986 25440 35992 25492
rect 36044 25480 36050 25492
rect 36170 25480 36176 25492
rect 36044 25452 36176 25480
rect 36044 25440 36050 25452
rect 36170 25440 36176 25452
rect 36228 25480 36234 25492
rect 36449 25483 36507 25489
rect 36449 25480 36461 25483
rect 36228 25452 36461 25480
rect 36228 25440 36234 25452
rect 36449 25449 36461 25452
rect 36495 25449 36507 25483
rect 40678 25480 40684 25492
rect 40639 25452 40684 25480
rect 36449 25443 36507 25449
rect 40678 25440 40684 25452
rect 40736 25440 40742 25492
rect 41417 25483 41475 25489
rect 41417 25449 41429 25483
rect 41463 25480 41475 25483
rect 41874 25480 41880 25492
rect 41463 25452 41880 25480
rect 41463 25449 41475 25452
rect 41417 25443 41475 25449
rect 41874 25440 41880 25452
rect 41932 25440 41938 25492
rect 44542 25480 44548 25492
rect 44503 25452 44548 25480
rect 44542 25440 44548 25452
rect 44600 25440 44606 25492
rect 44634 25440 44640 25492
rect 44692 25480 44698 25492
rect 44913 25483 44971 25489
rect 44913 25480 44925 25483
rect 44692 25452 44925 25480
rect 44692 25440 44698 25452
rect 44913 25449 44925 25452
rect 44959 25449 44971 25483
rect 46934 25480 46940 25492
rect 46895 25452 46940 25480
rect 44913 25443 44971 25449
rect 46934 25440 46940 25452
rect 46992 25440 46998 25492
rect 37826 25372 37832 25424
rect 37884 25412 37890 25424
rect 38289 25415 38347 25421
rect 38289 25412 38301 25415
rect 37884 25384 38301 25412
rect 37884 25372 37890 25384
rect 38289 25381 38301 25384
rect 38335 25381 38347 25415
rect 38289 25375 38347 25381
rect 38381 25415 38439 25421
rect 38381 25381 38393 25415
rect 38427 25412 38439 25415
rect 38562 25412 38568 25424
rect 38427 25384 38568 25412
rect 38427 25381 38439 25384
rect 38381 25375 38439 25381
rect 38562 25372 38568 25384
rect 38620 25372 38626 25424
rect 39574 25421 39580 25424
rect 39568 25412 39580 25421
rect 39535 25384 39580 25412
rect 39568 25375 39580 25384
rect 39574 25372 39580 25375
rect 39632 25372 39638 25424
rect 41785 25415 41843 25421
rect 41785 25381 41797 25415
rect 41831 25412 41843 25415
rect 41966 25412 41972 25424
rect 41831 25384 41972 25412
rect 41831 25381 41843 25384
rect 41785 25375 41843 25381
rect 41966 25372 41972 25384
rect 42024 25372 42030 25424
rect 43349 25415 43407 25421
rect 43349 25381 43361 25415
rect 43395 25412 43407 25415
rect 43438 25412 43444 25424
rect 43395 25384 43444 25412
rect 43395 25381 43407 25384
rect 43349 25375 43407 25381
rect 43438 25372 43444 25384
rect 43496 25372 43502 25424
rect 45741 25415 45799 25421
rect 45741 25381 45753 25415
rect 45787 25412 45799 25415
rect 46014 25412 46020 25424
rect 45787 25384 46020 25412
rect 45787 25381 45799 25384
rect 45741 25375 45799 25381
rect 46014 25372 46020 25384
rect 46072 25372 46078 25424
rect 36262 25344 36268 25356
rect 36223 25316 36268 25344
rect 36262 25304 36268 25316
rect 36320 25304 36326 25356
rect 38654 25304 38660 25356
rect 38712 25344 38718 25356
rect 39301 25347 39359 25353
rect 39301 25344 39313 25347
rect 38712 25316 39313 25344
rect 38712 25304 38718 25316
rect 39301 25313 39313 25316
rect 39347 25313 39359 25347
rect 39301 25307 39359 25313
rect 42153 25347 42211 25353
rect 42153 25313 42165 25347
rect 42199 25313 42211 25347
rect 43530 25344 43536 25356
rect 43491 25316 43536 25344
rect 42153 25307 42211 25313
rect 35805 25279 35863 25285
rect 35805 25245 35817 25279
rect 35851 25276 35863 25279
rect 36541 25279 36599 25285
rect 36541 25276 36553 25279
rect 35851 25248 36553 25276
rect 35851 25245 35863 25248
rect 35805 25239 35863 25245
rect 36541 25245 36553 25248
rect 36587 25276 36599 25279
rect 36906 25276 36912 25288
rect 36587 25248 36912 25276
rect 36587 25245 36599 25248
rect 36541 25239 36599 25245
rect 36906 25236 36912 25248
rect 36964 25236 36970 25288
rect 38194 25276 38200 25288
rect 38155 25248 38200 25276
rect 38194 25236 38200 25248
rect 38252 25236 38258 25288
rect 42168 25276 42196 25307
rect 43530 25304 43536 25316
rect 43588 25304 43594 25356
rect 46750 25344 46756 25356
rect 46711 25316 46756 25344
rect 46750 25304 46756 25316
rect 46808 25344 46814 25356
rect 47302 25344 47308 25356
rect 46808 25316 47308 25344
rect 46808 25304 46814 25316
rect 47302 25304 47308 25316
rect 47360 25304 47366 25356
rect 42610 25276 42616 25288
rect 42168 25248 42616 25276
rect 42610 25236 42616 25248
rect 42668 25276 42674 25288
rect 43717 25279 43775 25285
rect 43717 25276 43729 25279
rect 42668 25248 43729 25276
rect 42668 25236 42674 25248
rect 43717 25245 43729 25248
rect 43763 25245 43775 25279
rect 43717 25239 43775 25245
rect 45741 25279 45799 25285
rect 45741 25245 45753 25279
rect 45787 25245 45799 25279
rect 45741 25239 45799 25245
rect 35986 25208 35992 25220
rect 35947 25180 35992 25208
rect 35986 25168 35992 25180
rect 36044 25168 36050 25220
rect 37829 25211 37887 25217
rect 37829 25177 37841 25211
rect 37875 25208 37887 25211
rect 38286 25208 38292 25220
rect 37875 25180 38292 25208
rect 37875 25177 37887 25180
rect 37829 25171 37887 25177
rect 38286 25168 38292 25180
rect 38344 25168 38350 25220
rect 44726 25168 44732 25220
rect 44784 25208 44790 25220
rect 45281 25211 45339 25217
rect 45281 25208 45293 25211
rect 44784 25180 45293 25208
rect 44784 25168 44790 25180
rect 45281 25177 45293 25180
rect 45327 25177 45339 25211
rect 45756 25208 45784 25239
rect 45830 25236 45836 25288
rect 45888 25276 45894 25288
rect 47394 25276 47400 25288
rect 45888 25248 47400 25276
rect 45888 25236 45894 25248
rect 47394 25236 47400 25248
rect 47452 25236 47458 25288
rect 45756 25180 46336 25208
rect 45281 25171 45339 25177
rect 42334 25140 42340 25152
rect 42295 25112 42340 25140
rect 42334 25100 42340 25112
rect 42392 25100 42398 25152
rect 46308 25149 46336 25180
rect 46293 25143 46351 25149
rect 46293 25109 46305 25143
rect 46339 25140 46351 25143
rect 46382 25140 46388 25152
rect 46339 25112 46388 25140
rect 46339 25109 46351 25112
rect 46293 25103 46351 25109
rect 46382 25100 46388 25112
rect 46440 25100 46446 25152
rect 46661 25143 46719 25149
rect 46661 25109 46673 25143
rect 46707 25140 46719 25143
rect 46842 25140 46848 25152
rect 46707 25112 46848 25140
rect 46707 25109 46719 25112
rect 46661 25103 46719 25109
rect 46842 25100 46848 25112
rect 46900 25100 46906 25152
rect 1104 25050 48852 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 34966 25050
rect 35018 24998 35030 25050
rect 35082 24998 35094 25050
rect 35146 24998 35158 25050
rect 35210 24998 48852 25050
rect 1104 24976 48852 24998
rect 36906 24936 36912 24948
rect 36867 24908 36912 24936
rect 36906 24896 36912 24908
rect 36964 24896 36970 24948
rect 37826 24936 37832 24948
rect 37787 24908 37832 24936
rect 37826 24896 37832 24908
rect 37884 24896 37890 24948
rect 38194 24936 38200 24948
rect 38155 24908 38200 24936
rect 38194 24896 38200 24908
rect 38252 24896 38258 24948
rect 38654 24896 38660 24948
rect 38712 24936 38718 24948
rect 39301 24939 39359 24945
rect 39301 24936 39313 24939
rect 38712 24908 39313 24936
rect 38712 24896 38718 24908
rect 39301 24905 39313 24908
rect 39347 24905 39359 24939
rect 39301 24899 39359 24905
rect 39574 24896 39580 24948
rect 39632 24936 39638 24948
rect 39669 24939 39727 24945
rect 39669 24936 39681 24939
rect 39632 24908 39681 24936
rect 39632 24896 39638 24908
rect 39669 24905 39681 24908
rect 39715 24905 39727 24939
rect 39669 24899 39727 24905
rect 41693 24939 41751 24945
rect 41693 24905 41705 24939
rect 41739 24936 41751 24939
rect 42334 24936 42340 24948
rect 41739 24908 42340 24936
rect 41739 24905 41751 24908
rect 41693 24899 41751 24905
rect 42334 24896 42340 24908
rect 42392 24896 42398 24948
rect 43530 24896 43536 24948
rect 43588 24936 43594 24948
rect 43717 24939 43775 24945
rect 43717 24936 43729 24939
rect 43588 24908 43729 24936
rect 43588 24896 43594 24908
rect 43717 24905 43729 24908
rect 43763 24905 43775 24939
rect 43717 24899 43775 24905
rect 45554 24896 45560 24948
rect 45612 24936 45618 24948
rect 45741 24939 45799 24945
rect 45741 24936 45753 24939
rect 45612 24908 45753 24936
rect 45612 24896 45618 24908
rect 45741 24905 45753 24908
rect 45787 24936 45799 24939
rect 45833 24939 45891 24945
rect 45833 24936 45845 24939
rect 45787 24908 45845 24936
rect 45787 24905 45799 24908
rect 45741 24899 45799 24905
rect 45833 24905 45845 24908
rect 45879 24905 45891 24939
rect 45833 24899 45891 24905
rect 37844 24800 37872 24896
rect 38746 24800 38752 24812
rect 37844 24772 38752 24800
rect 38746 24760 38752 24772
rect 38804 24760 38810 24812
rect 42352 24800 42380 24896
rect 42797 24803 42855 24809
rect 42797 24800 42809 24803
rect 42352 24772 42809 24800
rect 42797 24769 42809 24772
rect 42843 24769 42855 24803
rect 42797 24763 42855 24769
rect 44913 24803 44971 24809
rect 44913 24769 44925 24803
rect 44959 24800 44971 24803
rect 44959 24772 46244 24800
rect 44959 24769 44971 24772
rect 44913 24763 44971 24769
rect 35529 24735 35587 24741
rect 35529 24732 35541 24735
rect 35452 24704 35541 24732
rect 35452 24608 35480 24704
rect 35529 24701 35541 24704
rect 35575 24732 35587 24735
rect 36354 24732 36360 24744
rect 35575 24704 36360 24732
rect 35575 24701 35587 24704
rect 35529 24695 35587 24701
rect 36354 24692 36360 24704
rect 36412 24692 36418 24744
rect 38565 24735 38623 24741
rect 38565 24701 38577 24735
rect 38611 24732 38623 24735
rect 38654 24732 38660 24744
rect 38611 24704 38660 24732
rect 38611 24701 38623 24704
rect 38565 24695 38623 24701
rect 38654 24692 38660 24704
rect 38712 24692 38718 24744
rect 42061 24735 42119 24741
rect 42061 24701 42073 24735
rect 42107 24732 42119 24735
rect 43346 24732 43352 24744
rect 42107 24704 43352 24732
rect 42107 24701 42119 24704
rect 42061 24695 42119 24701
rect 35802 24673 35808 24676
rect 35796 24664 35808 24673
rect 35763 24636 35808 24664
rect 35796 24627 35808 24636
rect 35802 24624 35808 24627
rect 35860 24624 35866 24676
rect 42720 24673 42748 24704
rect 43346 24692 43352 24704
rect 43404 24692 43410 24744
rect 45741 24735 45799 24741
rect 45741 24701 45753 24735
rect 45787 24732 45799 24735
rect 46109 24735 46167 24741
rect 46109 24732 46121 24735
rect 45787 24704 46121 24732
rect 45787 24701 45799 24704
rect 45741 24695 45799 24701
rect 46109 24701 46121 24704
rect 46155 24701 46167 24735
rect 46109 24695 46167 24701
rect 42521 24667 42579 24673
rect 42521 24633 42533 24667
rect 42567 24633 42579 24667
rect 42521 24627 42579 24633
rect 42705 24667 42763 24673
rect 42705 24633 42717 24667
rect 42751 24633 42763 24667
rect 42705 24627 42763 24633
rect 45281 24667 45339 24673
rect 45281 24633 45293 24667
rect 45327 24664 45339 24667
rect 46014 24664 46020 24676
rect 45327 24636 46020 24664
rect 45327 24633 45339 24636
rect 45281 24627 45339 24633
rect 35434 24596 35440 24608
rect 35395 24568 35440 24596
rect 35434 24556 35440 24568
rect 35492 24556 35498 24608
rect 38841 24599 38899 24605
rect 38841 24565 38853 24599
rect 38887 24596 38899 24599
rect 39114 24596 39120 24608
rect 38887 24568 39120 24596
rect 38887 24565 38899 24568
rect 38841 24559 38899 24565
rect 39114 24556 39120 24568
rect 39172 24556 39178 24608
rect 42058 24556 42064 24608
rect 42116 24596 42122 24608
rect 42227 24599 42285 24605
rect 42227 24596 42239 24599
rect 42116 24568 42239 24596
rect 42116 24556 42122 24568
rect 42227 24565 42239 24568
rect 42273 24565 42285 24599
rect 42227 24559 42285 24565
rect 42334 24556 42340 24608
rect 42392 24596 42398 24608
rect 42536 24596 42564 24627
rect 46014 24624 46020 24636
rect 46072 24624 46078 24676
rect 46216 24664 46244 24772
rect 46382 24673 46388 24676
rect 46376 24664 46388 24673
rect 46216 24636 46388 24664
rect 46376 24627 46388 24636
rect 46440 24664 46446 24676
rect 46842 24664 46848 24676
rect 46440 24636 46848 24664
rect 46382 24624 46388 24627
rect 46440 24624 46446 24636
rect 46842 24624 46848 24636
rect 46900 24624 46906 24676
rect 42886 24596 42892 24608
rect 42392 24568 42892 24596
rect 42392 24556 42398 24568
rect 42886 24556 42892 24568
rect 42944 24556 42950 24608
rect 43438 24596 43444 24608
rect 43399 24568 43444 24596
rect 43438 24556 43444 24568
rect 43496 24556 43502 24608
rect 46934 24556 46940 24608
rect 46992 24596 46998 24608
rect 47489 24599 47547 24605
rect 47489 24596 47501 24599
rect 46992 24568 47501 24596
rect 46992 24556 46998 24568
rect 47489 24565 47501 24568
rect 47535 24565 47547 24599
rect 47489 24559 47547 24565
rect 1104 24506 48852 24528
rect 1104 24454 19606 24506
rect 19658 24454 19670 24506
rect 19722 24454 19734 24506
rect 19786 24454 19798 24506
rect 19850 24454 48852 24506
rect 1104 24432 48852 24454
rect 35069 24395 35127 24401
rect 35069 24361 35081 24395
rect 35115 24392 35127 24395
rect 35989 24395 36047 24401
rect 35989 24392 36001 24395
rect 35115 24364 36001 24392
rect 35115 24361 35127 24364
rect 35069 24355 35127 24361
rect 35989 24361 36001 24364
rect 36035 24392 36047 24395
rect 36262 24392 36268 24404
rect 36035 24364 36268 24392
rect 36035 24361 36047 24364
rect 35989 24355 36047 24361
rect 36262 24352 36268 24364
rect 36320 24352 36326 24404
rect 38013 24395 38071 24401
rect 38013 24361 38025 24395
rect 38059 24392 38071 24395
rect 38562 24392 38568 24404
rect 38059 24364 38568 24392
rect 38059 24361 38071 24364
rect 38013 24355 38071 24361
rect 38562 24352 38568 24364
rect 38620 24352 38626 24404
rect 41785 24395 41843 24401
rect 41785 24361 41797 24395
rect 41831 24392 41843 24395
rect 41874 24392 41880 24404
rect 41831 24364 41880 24392
rect 41831 24361 41843 24364
rect 41785 24355 41843 24361
rect 41874 24352 41880 24364
rect 41932 24352 41938 24404
rect 42245 24395 42303 24401
rect 42245 24361 42257 24395
rect 42291 24392 42303 24395
rect 42334 24392 42340 24404
rect 42291 24364 42340 24392
rect 42291 24361 42303 24364
rect 42245 24355 42303 24361
rect 42334 24352 42340 24364
rect 42392 24352 42398 24404
rect 42610 24392 42616 24404
rect 42571 24364 42616 24392
rect 42610 24352 42616 24364
rect 42668 24352 42674 24404
rect 45281 24395 45339 24401
rect 45281 24361 45293 24395
rect 45327 24392 45339 24395
rect 45830 24392 45836 24404
rect 45327 24364 45836 24392
rect 45327 24361 45339 24364
rect 45281 24355 45339 24361
rect 45830 24352 45836 24364
rect 45888 24352 45894 24404
rect 46842 24392 46848 24404
rect 46803 24364 46848 24392
rect 46842 24352 46848 24364
rect 46900 24352 46906 24404
rect 36630 24324 36636 24336
rect 36591 24296 36636 24324
rect 36630 24284 36636 24296
rect 36688 24284 36694 24336
rect 36725 24327 36783 24333
rect 36725 24293 36737 24327
rect 36771 24324 36783 24327
rect 37182 24324 37188 24336
rect 36771 24296 37188 24324
rect 36771 24293 36783 24296
rect 36725 24287 36783 24293
rect 35621 24259 35679 24265
rect 35621 24225 35633 24259
rect 35667 24256 35679 24259
rect 35802 24256 35808 24268
rect 35667 24228 35808 24256
rect 35667 24225 35679 24228
rect 35621 24219 35679 24225
rect 35802 24216 35808 24228
rect 35860 24256 35866 24268
rect 36740 24256 36768 24287
rect 37182 24284 37188 24296
rect 37240 24284 37246 24336
rect 35860 24228 36768 24256
rect 41601 24259 41659 24265
rect 35860 24216 35866 24228
rect 41601 24225 41613 24259
rect 41647 24256 41659 24259
rect 42058 24256 42064 24268
rect 41647 24228 42064 24256
rect 41647 24225 41659 24228
rect 41601 24219 41659 24225
rect 42058 24216 42064 24228
rect 42116 24216 42122 24268
rect 45732 24259 45790 24265
rect 45732 24225 45744 24259
rect 45778 24256 45790 24259
rect 46014 24256 46020 24268
rect 45778 24228 46020 24256
rect 45778 24225 45790 24228
rect 45732 24219 45790 24225
rect 46014 24216 46020 24228
rect 46072 24216 46078 24268
rect 35710 24148 35716 24200
rect 35768 24188 35774 24200
rect 36633 24191 36691 24197
rect 36633 24188 36645 24191
rect 35768 24160 36645 24188
rect 35768 24148 35774 24160
rect 36633 24157 36645 24160
rect 36679 24188 36691 24191
rect 37182 24188 37188 24200
rect 36679 24160 37188 24188
rect 36679 24157 36691 24160
rect 36633 24151 36691 24157
rect 37182 24148 37188 24160
rect 37240 24148 37246 24200
rect 45462 24188 45468 24200
rect 45423 24160 45468 24188
rect 45462 24148 45468 24160
rect 45520 24148 45526 24200
rect 36170 24120 36176 24132
rect 36131 24092 36176 24120
rect 36170 24080 36176 24092
rect 36228 24080 36234 24132
rect 30466 24012 30472 24064
rect 30524 24052 30530 24064
rect 31205 24055 31263 24061
rect 31205 24052 31217 24055
rect 30524 24024 31217 24052
rect 30524 24012 30530 24024
rect 31205 24021 31217 24024
rect 31251 24021 31263 24055
rect 31205 24015 31263 24021
rect 41049 24055 41107 24061
rect 41049 24021 41061 24055
rect 41095 24052 41107 24055
rect 41598 24052 41604 24064
rect 41095 24024 41604 24052
rect 41095 24021 41107 24024
rect 41049 24015 41107 24021
rect 41598 24012 41604 24024
rect 41656 24012 41662 24064
rect 1104 23962 48852 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 34966 23962
rect 35018 23910 35030 23962
rect 35082 23910 35094 23962
rect 35146 23910 35158 23962
rect 35210 23910 48852 23962
rect 1104 23888 48852 23910
rect 31294 23848 31300 23860
rect 31255 23820 31300 23848
rect 31294 23808 31300 23820
rect 31352 23808 31358 23860
rect 35253 23851 35311 23857
rect 35253 23817 35265 23851
rect 35299 23848 35311 23851
rect 35802 23848 35808 23860
rect 35299 23820 35808 23848
rect 35299 23817 35311 23820
rect 35253 23811 35311 23817
rect 35802 23808 35808 23820
rect 35860 23808 35866 23860
rect 41046 23848 41052 23860
rect 41007 23820 41052 23848
rect 41046 23808 41052 23820
rect 41104 23808 41110 23860
rect 42058 23848 42064 23860
rect 42019 23820 42064 23848
rect 42058 23808 42064 23820
rect 42116 23808 42122 23860
rect 42242 23808 42248 23860
rect 42300 23848 42306 23860
rect 42337 23851 42395 23857
rect 42337 23848 42349 23851
rect 42300 23820 42349 23848
rect 42300 23808 42306 23820
rect 42337 23817 42349 23820
rect 42383 23817 42395 23851
rect 42337 23811 42395 23817
rect 35621 23783 35679 23789
rect 35621 23749 35633 23783
rect 35667 23780 35679 23783
rect 35710 23780 35716 23792
rect 35667 23752 35716 23780
rect 35667 23749 35679 23752
rect 35621 23743 35679 23749
rect 35710 23740 35716 23752
rect 35768 23740 35774 23792
rect 41598 23712 41604 23724
rect 41559 23684 41604 23712
rect 41598 23672 41604 23684
rect 41656 23712 41662 23724
rect 41656 23684 42656 23712
rect 41656 23672 41662 23684
rect 42628 23656 42656 23684
rect 35434 23604 35440 23656
rect 35492 23644 35498 23656
rect 36081 23647 36139 23653
rect 36081 23644 36093 23647
rect 35492 23616 36093 23644
rect 35492 23604 35498 23616
rect 31113 23579 31171 23585
rect 31113 23545 31125 23579
rect 31159 23576 31171 23579
rect 31573 23579 31631 23585
rect 31573 23576 31585 23579
rect 31159 23548 31585 23576
rect 31159 23545 31171 23548
rect 31113 23539 31171 23545
rect 31573 23545 31585 23548
rect 31619 23576 31631 23579
rect 31662 23576 31668 23588
rect 31619 23548 31668 23576
rect 31619 23545 31631 23548
rect 31573 23539 31631 23545
rect 31662 23536 31668 23548
rect 31720 23536 31726 23588
rect 31846 23576 31852 23588
rect 31807 23548 31852 23576
rect 31846 23536 31852 23548
rect 31904 23536 31910 23588
rect 30466 23468 30472 23520
rect 30524 23508 30530 23520
rect 31757 23511 31815 23517
rect 31757 23508 31769 23511
rect 30524 23480 31769 23508
rect 30524 23468 30530 23480
rect 31757 23477 31769 23480
rect 31803 23477 31815 23511
rect 31757 23471 31815 23477
rect 35802 23468 35808 23520
rect 35860 23508 35866 23520
rect 35912 23517 35940 23616
rect 36081 23613 36093 23616
rect 36127 23613 36139 23647
rect 36081 23607 36139 23613
rect 36348 23647 36406 23653
rect 36348 23613 36360 23647
rect 36394 23644 36406 23647
rect 36906 23644 36912 23656
rect 36394 23616 36912 23644
rect 36394 23613 36406 23616
rect 36348 23607 36406 23613
rect 36906 23604 36912 23616
rect 36964 23604 36970 23656
rect 42242 23604 42248 23656
rect 42300 23644 42306 23656
rect 42521 23647 42579 23653
rect 42521 23644 42533 23647
rect 42300 23616 42533 23644
rect 42300 23604 42306 23616
rect 42521 23613 42533 23616
rect 42567 23613 42579 23647
rect 42521 23607 42579 23613
rect 42610 23604 42616 23656
rect 42668 23644 42674 23656
rect 42777 23647 42835 23653
rect 42777 23644 42789 23647
rect 42668 23616 42789 23644
rect 42668 23604 42674 23616
rect 42777 23613 42789 23616
rect 42823 23613 42835 23647
rect 42777 23607 42835 23613
rect 40865 23579 40923 23585
rect 40865 23545 40877 23579
rect 40911 23576 40923 23579
rect 41325 23579 41383 23585
rect 41325 23576 41337 23579
rect 40911 23548 41337 23576
rect 40911 23545 40923 23548
rect 40865 23539 40923 23545
rect 41325 23545 41337 23548
rect 41371 23576 41383 23579
rect 41414 23576 41420 23588
rect 41371 23548 41420 23576
rect 41371 23545 41383 23548
rect 41325 23539 41383 23545
rect 41414 23536 41420 23548
rect 41472 23536 41478 23588
rect 35897 23511 35955 23517
rect 35897 23508 35909 23511
rect 35860 23480 35909 23508
rect 35860 23468 35866 23480
rect 35897 23477 35909 23480
rect 35943 23477 35955 23511
rect 35897 23471 35955 23477
rect 37274 23468 37280 23520
rect 37332 23508 37338 23520
rect 37461 23511 37519 23517
rect 37461 23508 37473 23511
rect 37332 23480 37473 23508
rect 37332 23468 37338 23480
rect 37461 23477 37473 23480
rect 37507 23508 37519 23511
rect 38470 23508 38476 23520
rect 37507 23480 38476 23508
rect 37507 23477 37519 23480
rect 37461 23471 37519 23477
rect 38470 23468 38476 23480
rect 38528 23468 38534 23520
rect 38654 23508 38660 23520
rect 38615 23480 38660 23508
rect 38654 23468 38660 23480
rect 38712 23468 38718 23520
rect 40313 23511 40371 23517
rect 40313 23477 40325 23511
rect 40359 23508 40371 23511
rect 41046 23508 41052 23520
rect 40359 23480 41052 23508
rect 40359 23477 40371 23480
rect 40313 23471 40371 23477
rect 41046 23468 41052 23480
rect 41104 23508 41110 23520
rect 41509 23511 41567 23517
rect 41509 23508 41521 23511
rect 41104 23480 41521 23508
rect 41104 23468 41110 23480
rect 41509 23477 41521 23480
rect 41555 23477 41567 23511
rect 41509 23471 41567 23477
rect 43901 23511 43959 23517
rect 43901 23477 43913 23511
rect 43947 23508 43959 23511
rect 44082 23508 44088 23520
rect 43947 23480 44088 23508
rect 43947 23477 43959 23480
rect 43901 23471 43959 23477
rect 44082 23468 44088 23480
rect 44140 23468 44146 23520
rect 44634 23468 44640 23520
rect 44692 23508 44698 23520
rect 45462 23508 45468 23520
rect 44692 23480 45468 23508
rect 44692 23468 44698 23480
rect 45462 23468 45468 23480
rect 45520 23468 45526 23520
rect 45925 23511 45983 23517
rect 45925 23477 45937 23511
rect 45971 23508 45983 23511
rect 46014 23508 46020 23520
rect 45971 23480 46020 23508
rect 45971 23477 45983 23480
rect 45925 23471 45983 23477
rect 46014 23468 46020 23480
rect 46072 23468 46078 23520
rect 1104 23418 48852 23440
rect 1104 23366 19606 23418
rect 19658 23366 19670 23418
rect 19722 23366 19734 23418
rect 19786 23366 19798 23418
rect 19850 23366 48852 23418
rect 1104 23344 48852 23366
rect 31754 23264 31760 23316
rect 31812 23304 31818 23316
rect 32125 23307 32183 23313
rect 32125 23304 32137 23307
rect 31812 23276 32137 23304
rect 31812 23264 31818 23276
rect 32125 23273 32137 23276
rect 32171 23273 32183 23307
rect 32125 23267 32183 23273
rect 36541 23307 36599 23313
rect 36541 23273 36553 23307
rect 36587 23304 36599 23307
rect 36906 23304 36912 23316
rect 36587 23276 36912 23304
rect 36587 23273 36599 23276
rect 36541 23267 36599 23273
rect 36906 23264 36912 23276
rect 36964 23264 36970 23316
rect 38194 23264 38200 23316
rect 38252 23304 38258 23316
rect 38473 23307 38531 23313
rect 38473 23304 38485 23307
rect 38252 23276 38485 23304
rect 38252 23264 38258 23276
rect 38473 23273 38485 23276
rect 38519 23304 38531 23307
rect 38930 23304 38936 23316
rect 38519 23276 38936 23304
rect 38519 23273 38531 23276
rect 38473 23267 38531 23273
rect 38930 23264 38936 23276
rect 38988 23264 38994 23316
rect 41414 23264 41420 23316
rect 41472 23304 41478 23316
rect 41601 23307 41659 23313
rect 41601 23304 41613 23307
rect 41472 23276 41613 23304
rect 41472 23264 41478 23276
rect 41601 23273 41613 23276
rect 41647 23273 41659 23307
rect 42610 23304 42616 23316
rect 42571 23276 42616 23304
rect 41601 23267 41659 23273
rect 42610 23264 42616 23276
rect 42668 23264 42674 23316
rect 46014 23304 46020 23316
rect 45975 23276 46020 23304
rect 46014 23264 46020 23276
rect 46072 23264 46078 23316
rect 47026 23264 47032 23316
rect 47084 23304 47090 23316
rect 47305 23307 47363 23313
rect 47305 23304 47317 23307
rect 47084 23276 47317 23304
rect 47084 23264 47090 23276
rect 47305 23273 47317 23276
rect 47351 23273 47363 23307
rect 47305 23267 47363 23273
rect 31297 23239 31355 23245
rect 31297 23205 31309 23239
rect 31343 23236 31355 23239
rect 31846 23236 31852 23248
rect 31343 23208 31852 23236
rect 31343 23205 31355 23208
rect 31297 23199 31355 23205
rect 31846 23196 31852 23208
rect 31904 23196 31910 23248
rect 33226 23196 33232 23248
rect 33284 23236 33290 23248
rect 34057 23239 34115 23245
rect 34057 23236 34069 23239
rect 33284 23208 34069 23236
rect 33284 23196 33290 23208
rect 34057 23205 34069 23208
rect 34103 23205 34115 23239
rect 34057 23199 34115 23205
rect 38654 23168 38660 23180
rect 38615 23140 38660 23168
rect 38654 23128 38660 23140
rect 38712 23128 38718 23180
rect 38746 23128 38752 23180
rect 38804 23168 38810 23180
rect 39393 23171 39451 23177
rect 39393 23168 39405 23171
rect 38804 23140 39405 23168
rect 38804 23128 38810 23140
rect 39393 23137 39405 23140
rect 39439 23168 39451 23171
rect 39850 23168 39856 23180
rect 39439 23140 39856 23168
rect 39439 23137 39451 23140
rect 39393 23131 39451 23137
rect 39850 23128 39856 23140
rect 39908 23128 39914 23180
rect 44910 23177 44916 23180
rect 44904 23131 44916 23177
rect 44968 23168 44974 23180
rect 47121 23171 47179 23177
rect 44968 23140 45004 23168
rect 44910 23128 44916 23131
rect 44968 23128 44974 23140
rect 47121 23137 47133 23171
rect 47167 23168 47179 23171
rect 47302 23168 47308 23180
rect 47167 23140 47308 23168
rect 47167 23137 47179 23140
rect 47121 23131 47179 23137
rect 47302 23128 47308 23140
rect 47360 23128 47366 23180
rect 34054 23100 34060 23112
rect 34015 23072 34060 23100
rect 34054 23060 34060 23072
rect 34112 23060 34118 23112
rect 34149 23103 34207 23109
rect 34149 23069 34161 23103
rect 34195 23100 34207 23103
rect 34606 23100 34612 23112
rect 34195 23072 34612 23100
rect 34195 23069 34207 23072
rect 34149 23063 34207 23069
rect 34606 23060 34612 23072
rect 34664 23060 34670 23112
rect 39022 23109 39028 23112
rect 38980 23103 39028 23109
rect 38980 23069 38992 23103
rect 39026 23069 39028 23103
rect 38980 23063 39028 23069
rect 39022 23060 39028 23063
rect 39080 23060 39086 23112
rect 39114 23060 39120 23112
rect 39172 23100 39178 23112
rect 44634 23100 44640 23112
rect 39172 23072 39217 23100
rect 44595 23072 44640 23100
rect 39172 23060 39178 23072
rect 44634 23060 44640 23072
rect 44692 23060 44698 23112
rect 33594 23032 33600 23044
rect 33555 23004 33600 23032
rect 33594 22992 33600 23004
rect 33652 22992 33658 23044
rect 36170 22964 36176 22976
rect 36131 22936 36176 22964
rect 36170 22924 36176 22936
rect 36228 22924 36234 22976
rect 40494 22964 40500 22976
rect 40455 22936 40500 22964
rect 40494 22924 40500 22936
rect 40552 22924 40558 22976
rect 41141 22967 41199 22973
rect 41141 22933 41153 22967
rect 41187 22964 41199 22967
rect 41322 22964 41328 22976
rect 41187 22936 41328 22964
rect 41187 22933 41199 22936
rect 41141 22927 41199 22933
rect 41322 22924 41328 22936
rect 41380 22924 41386 22976
rect 43625 22967 43683 22973
rect 43625 22933 43637 22967
rect 43671 22964 43683 22967
rect 44082 22964 44088 22976
rect 43671 22936 44088 22964
rect 43671 22933 43683 22936
rect 43625 22927 43683 22933
rect 44082 22924 44088 22936
rect 44140 22924 44146 22976
rect 46658 22964 46664 22976
rect 46619 22936 46664 22964
rect 46658 22924 46664 22936
rect 46716 22924 46722 22976
rect 46934 22964 46940 22976
rect 46895 22936 46940 22964
rect 46934 22924 46940 22936
rect 46992 22924 46998 22976
rect 1104 22874 48852 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 34966 22874
rect 35018 22822 35030 22874
rect 35082 22822 35094 22874
rect 35146 22822 35158 22874
rect 35210 22822 48852 22874
rect 1104 22800 48852 22822
rect 34054 22720 34060 22772
rect 34112 22760 34118 22772
rect 34241 22763 34299 22769
rect 34241 22760 34253 22763
rect 34112 22732 34253 22760
rect 34112 22720 34118 22732
rect 34241 22729 34253 22732
rect 34287 22760 34299 22763
rect 34287 22732 34928 22760
rect 34287 22729 34299 22732
rect 34241 22723 34299 22729
rect 34606 22692 34612 22704
rect 34567 22664 34612 22692
rect 34606 22652 34612 22664
rect 34664 22652 34670 22704
rect 31846 22584 31852 22636
rect 31904 22624 31910 22636
rect 34900 22633 34928 22732
rect 37366 22720 37372 22772
rect 37424 22760 37430 22772
rect 38013 22763 38071 22769
rect 38013 22760 38025 22763
rect 37424 22732 38025 22760
rect 37424 22720 37430 22732
rect 38013 22729 38025 22732
rect 38059 22760 38071 22763
rect 39114 22760 39120 22772
rect 38059 22732 39120 22760
rect 38059 22729 38071 22732
rect 38013 22723 38071 22729
rect 39114 22720 39120 22732
rect 39172 22720 39178 22772
rect 39850 22760 39856 22772
rect 39811 22732 39856 22760
rect 39850 22720 39856 22732
rect 39908 22720 39914 22772
rect 42337 22763 42395 22769
rect 42337 22729 42349 22763
rect 42383 22760 42395 22763
rect 42610 22760 42616 22772
rect 42383 22732 42616 22760
rect 42383 22729 42395 22732
rect 42337 22723 42395 22729
rect 42610 22720 42616 22732
rect 42668 22720 42674 22772
rect 44910 22760 44916 22772
rect 44871 22732 44916 22760
rect 44910 22720 44916 22732
rect 44968 22720 44974 22772
rect 46290 22760 46296 22772
rect 46251 22732 46296 22760
rect 46290 22720 46296 22732
rect 46348 22720 46354 22772
rect 38562 22692 38568 22704
rect 38523 22664 38568 22692
rect 38562 22652 38568 22664
rect 38620 22652 38626 22704
rect 47302 22692 47308 22704
rect 47263 22664 47308 22692
rect 47302 22652 47308 22664
rect 47360 22652 47366 22704
rect 34885 22627 34943 22633
rect 31904 22596 32444 22624
rect 31904 22584 31910 22596
rect 32416 22568 32444 22596
rect 34885 22593 34897 22627
rect 34931 22593 34943 22627
rect 34885 22587 34943 22593
rect 35529 22627 35587 22633
rect 35529 22593 35541 22627
rect 35575 22624 35587 22627
rect 35575 22596 36124 22624
rect 35575 22593 35587 22596
rect 35529 22587 35587 22593
rect 32309 22559 32367 22565
rect 32309 22556 32321 22559
rect 32232 22528 32321 22556
rect 32232 22432 32260 22528
rect 32309 22525 32321 22528
rect 32355 22525 32367 22559
rect 32309 22519 32367 22525
rect 32398 22516 32404 22568
rect 32456 22556 32462 22568
rect 32565 22559 32623 22565
rect 32565 22556 32577 22559
rect 32456 22528 32577 22556
rect 32456 22516 32462 22528
rect 32565 22525 32577 22528
rect 32611 22525 32623 22559
rect 35989 22559 36047 22565
rect 35989 22556 36001 22559
rect 32565 22519 32623 22525
rect 35912 22528 36001 22556
rect 29546 22420 29552 22432
rect 29507 22392 29552 22420
rect 29546 22380 29552 22392
rect 29604 22380 29610 22432
rect 32214 22420 32220 22432
rect 32175 22392 32220 22420
rect 32214 22380 32220 22392
rect 32272 22380 32278 22432
rect 33594 22380 33600 22432
rect 33652 22420 33658 22432
rect 33689 22423 33747 22429
rect 33689 22420 33701 22423
rect 33652 22392 33701 22420
rect 33652 22380 33658 22392
rect 33689 22389 33701 22392
rect 33735 22389 33747 22423
rect 33689 22383 33747 22389
rect 35802 22380 35808 22432
rect 35860 22420 35866 22432
rect 35912 22429 35940 22528
rect 35989 22525 36001 22528
rect 36035 22525 36047 22559
rect 36096 22556 36124 22596
rect 38470 22584 38476 22636
rect 38528 22624 38534 22636
rect 39117 22627 39175 22633
rect 39117 22624 39129 22627
rect 38528 22596 39129 22624
rect 38528 22584 38534 22596
rect 39117 22593 39129 22596
rect 39163 22624 39175 22627
rect 40221 22627 40279 22633
rect 40221 22624 40233 22627
rect 39163 22596 40233 22624
rect 39163 22593 39175 22596
rect 39117 22587 39175 22593
rect 40221 22593 40233 22596
rect 40267 22593 40279 22627
rect 40221 22587 40279 22593
rect 46658 22584 46664 22636
rect 46716 22624 46722 22636
rect 46842 22624 46848 22636
rect 46716 22596 46848 22624
rect 46716 22584 46722 22596
rect 46842 22584 46848 22596
rect 46900 22584 46906 22636
rect 36256 22559 36314 22565
rect 36256 22556 36268 22559
rect 36096 22528 36268 22556
rect 35989 22519 36047 22525
rect 36256 22525 36268 22528
rect 36302 22556 36314 22559
rect 37182 22556 37188 22568
rect 36302 22528 37188 22556
rect 36302 22525 36314 22528
rect 36256 22519 36314 22525
rect 37182 22516 37188 22528
rect 37240 22516 37246 22568
rect 38194 22516 38200 22568
rect 38252 22556 38258 22568
rect 39022 22556 39028 22568
rect 38252 22528 39028 22556
rect 38252 22516 38258 22528
rect 39022 22516 39028 22528
rect 39080 22556 39086 22568
rect 39485 22559 39543 22565
rect 39485 22556 39497 22559
rect 39080 22528 39497 22556
rect 39080 22516 39086 22528
rect 39485 22525 39497 22528
rect 39531 22525 39543 22559
rect 40957 22559 41015 22565
rect 40957 22556 40969 22559
rect 39485 22519 39543 22525
rect 40788 22528 40969 22556
rect 38381 22491 38439 22497
rect 38381 22457 38393 22491
rect 38427 22488 38439 22491
rect 38654 22488 38660 22500
rect 38427 22460 38660 22488
rect 38427 22457 38439 22460
rect 38381 22451 38439 22457
rect 38654 22448 38660 22460
rect 38712 22488 38718 22500
rect 38841 22491 38899 22497
rect 38841 22488 38853 22491
rect 38712 22460 38853 22488
rect 38712 22448 38718 22460
rect 38841 22457 38853 22460
rect 38887 22457 38899 22491
rect 38841 22451 38899 22457
rect 35897 22423 35955 22429
rect 35897 22420 35909 22423
rect 35860 22392 35909 22420
rect 35860 22380 35866 22392
rect 35897 22389 35909 22392
rect 35943 22389 35955 22423
rect 35897 22383 35955 22389
rect 37274 22380 37280 22432
rect 37332 22420 37338 22432
rect 37369 22423 37427 22429
rect 37369 22420 37381 22423
rect 37332 22392 37381 22420
rect 37332 22380 37338 22392
rect 37369 22389 37381 22392
rect 37415 22389 37427 22423
rect 37369 22383 37427 22389
rect 38930 22380 38936 22432
rect 38988 22420 38994 22432
rect 39025 22423 39083 22429
rect 39025 22420 39037 22423
rect 38988 22392 39037 22420
rect 38988 22380 38994 22392
rect 39025 22389 39037 22392
rect 39071 22389 39083 22423
rect 39025 22383 39083 22389
rect 40402 22380 40408 22432
rect 40460 22420 40466 22432
rect 40788 22429 40816 22528
rect 40957 22525 40969 22528
rect 41003 22556 41015 22559
rect 43349 22559 43407 22565
rect 43349 22556 43361 22559
rect 41003 22528 43361 22556
rect 41003 22525 41015 22528
rect 40957 22519 41015 22525
rect 43349 22525 43361 22528
rect 43395 22556 43407 22559
rect 43533 22559 43591 22565
rect 43533 22556 43545 22559
rect 43395 22528 43545 22556
rect 43395 22525 43407 22528
rect 43349 22519 43407 22525
rect 43533 22525 43545 22528
rect 43579 22556 43591 22559
rect 44634 22556 44640 22568
rect 43579 22528 44640 22556
rect 43579 22525 43591 22528
rect 43533 22519 43591 22525
rect 44634 22516 44640 22528
rect 44692 22556 44698 22568
rect 45465 22559 45523 22565
rect 45465 22556 45477 22559
rect 44692 22528 45477 22556
rect 44692 22516 44698 22528
rect 45465 22525 45477 22528
rect 45511 22556 45523 22559
rect 46106 22556 46112 22568
rect 45511 22528 46112 22556
rect 45511 22525 45523 22528
rect 45465 22519 45523 22525
rect 46106 22516 46112 22528
rect 46164 22516 46170 22568
rect 41224 22491 41282 22497
rect 41224 22457 41236 22491
rect 41270 22488 41282 22491
rect 41322 22488 41328 22500
rect 41270 22460 41328 22488
rect 41270 22457 41282 22460
rect 41224 22451 41282 22457
rect 41322 22448 41328 22460
rect 41380 22488 41386 22500
rect 41598 22488 41604 22500
rect 41380 22460 41604 22488
rect 41380 22448 41386 22460
rect 41598 22448 41604 22460
rect 41656 22448 41662 22500
rect 43800 22491 43858 22497
rect 43800 22457 43812 22491
rect 43846 22488 43858 22491
rect 44082 22488 44088 22500
rect 43846 22460 44088 22488
rect 43846 22457 43858 22460
rect 43800 22451 43858 22457
rect 44082 22448 44088 22460
rect 44140 22448 44146 22500
rect 45094 22448 45100 22500
rect 45152 22488 45158 22500
rect 45925 22491 45983 22497
rect 45925 22488 45937 22491
rect 45152 22460 45937 22488
rect 45152 22448 45158 22460
rect 45925 22457 45937 22460
rect 45971 22488 45983 22491
rect 46569 22491 46627 22497
rect 46569 22488 46581 22491
rect 45971 22460 46581 22488
rect 45971 22457 45983 22460
rect 45925 22451 45983 22457
rect 46569 22457 46581 22460
rect 46615 22457 46627 22491
rect 46569 22451 46627 22457
rect 40773 22423 40831 22429
rect 40773 22420 40785 22423
rect 40460 22392 40785 22420
rect 40460 22380 40466 22392
rect 40773 22389 40785 22392
rect 40819 22389 40831 22423
rect 40773 22383 40831 22389
rect 45554 22380 45560 22432
rect 45612 22420 45618 22432
rect 46753 22423 46811 22429
rect 46753 22420 46765 22423
rect 45612 22392 46765 22420
rect 45612 22380 45618 22392
rect 46753 22389 46765 22392
rect 46799 22420 46811 22423
rect 46934 22420 46940 22432
rect 46799 22392 46940 22420
rect 46799 22389 46811 22392
rect 46753 22383 46811 22389
rect 46934 22380 46940 22392
rect 46992 22380 46998 22432
rect 1104 22330 48852 22352
rect 1104 22278 19606 22330
rect 19658 22278 19670 22330
rect 19722 22278 19734 22330
rect 19786 22278 19798 22330
rect 19850 22278 48852 22330
rect 1104 22256 48852 22278
rect 29546 22176 29552 22228
rect 29604 22216 29610 22228
rect 29914 22216 29920 22228
rect 29604 22188 29920 22216
rect 29604 22176 29610 22188
rect 29914 22176 29920 22188
rect 29972 22216 29978 22228
rect 30285 22219 30343 22225
rect 30285 22216 30297 22219
rect 29972 22188 30297 22216
rect 29972 22176 29978 22188
rect 30285 22185 30297 22188
rect 30331 22185 30343 22219
rect 30285 22179 30343 22185
rect 31754 22176 31760 22228
rect 31812 22216 31818 22228
rect 32214 22216 32220 22228
rect 31812 22188 32220 22216
rect 31812 22176 31818 22188
rect 32214 22176 32220 22188
rect 32272 22216 32278 22228
rect 33042 22216 33048 22228
rect 32272 22188 33048 22216
rect 32272 22176 32278 22188
rect 33042 22176 33048 22188
rect 33100 22176 33106 22228
rect 34606 22176 34612 22228
rect 34664 22216 34670 22228
rect 34977 22219 35035 22225
rect 34977 22216 34989 22219
rect 34664 22188 34989 22216
rect 34664 22176 34670 22188
rect 34977 22185 34989 22188
rect 35023 22185 35035 22219
rect 34977 22179 35035 22185
rect 36633 22219 36691 22225
rect 36633 22185 36645 22219
rect 36679 22216 36691 22219
rect 37366 22216 37372 22228
rect 36679 22188 37372 22216
rect 36679 22185 36691 22188
rect 36633 22179 36691 22185
rect 37366 22176 37372 22188
rect 37424 22216 37430 22228
rect 38562 22216 38568 22228
rect 37424 22188 38568 22216
rect 37424 22176 37430 22188
rect 38562 22176 38568 22188
rect 38620 22176 38626 22228
rect 38746 22176 38752 22228
rect 38804 22216 38810 22228
rect 39761 22219 39819 22225
rect 38804 22188 39712 22216
rect 38804 22176 38810 22188
rect 32398 22148 32404 22160
rect 32359 22120 32404 22148
rect 32398 22108 32404 22120
rect 32456 22108 32462 22160
rect 33594 22108 33600 22160
rect 33652 22148 33658 22160
rect 33842 22151 33900 22157
rect 33842 22148 33854 22151
rect 33652 22120 33854 22148
rect 33652 22108 33658 22120
rect 33842 22117 33854 22120
rect 33888 22117 33900 22151
rect 39684 22148 39712 22188
rect 39761 22185 39773 22219
rect 39807 22216 39819 22219
rect 39850 22216 39856 22228
rect 39807 22188 39856 22216
rect 39807 22185 39819 22188
rect 39761 22179 39819 22185
rect 39850 22176 39856 22188
rect 39908 22176 39914 22228
rect 45094 22216 45100 22228
rect 45055 22188 45100 22216
rect 45094 22176 45100 22188
rect 45152 22176 45158 22228
rect 41506 22148 41512 22160
rect 39684 22120 39988 22148
rect 41467 22120 41512 22148
rect 33842 22111 33900 22117
rect 28813 22083 28871 22089
rect 28813 22049 28825 22083
rect 28859 22080 28871 22083
rect 29161 22083 29219 22089
rect 29161 22080 29173 22083
rect 28859 22052 29173 22080
rect 28859 22049 28871 22052
rect 28813 22043 28871 22049
rect 29161 22049 29173 22052
rect 29207 22080 29219 22083
rect 30282 22080 30288 22092
rect 29207 22052 30288 22080
rect 29207 22049 29219 22052
rect 29161 22043 29219 22049
rect 30282 22040 30288 22052
rect 30340 22040 30346 22092
rect 36446 22080 36452 22092
rect 36407 22052 36452 22080
rect 36446 22040 36452 22052
rect 36504 22040 36510 22092
rect 36538 22040 36544 22092
rect 36596 22080 36602 22092
rect 36725 22083 36783 22089
rect 36725 22080 36737 22083
rect 36596 22052 36737 22080
rect 36596 22040 36602 22052
rect 36725 22049 36737 22052
rect 36771 22080 36783 22083
rect 37182 22080 37188 22092
rect 36771 22052 37188 22080
rect 36771 22049 36783 22052
rect 36725 22043 36783 22049
rect 37182 22040 37188 22052
rect 37240 22040 37246 22092
rect 37550 22040 37556 22092
rect 37608 22080 37614 22092
rect 39960 22080 39988 22120
rect 41506 22108 41512 22120
rect 41564 22108 41570 22160
rect 43898 22148 43904 22160
rect 43859 22120 43904 22148
rect 43898 22108 43904 22120
rect 43956 22108 43962 22160
rect 44729 22151 44787 22157
rect 44729 22148 44741 22151
rect 44639 22120 44741 22148
rect 44729 22117 44741 22120
rect 44775 22148 44787 22151
rect 44910 22148 44916 22160
rect 44775 22120 44916 22148
rect 44775 22117 44787 22120
rect 44729 22111 44787 22117
rect 40405 22083 40463 22089
rect 40405 22080 40417 22083
rect 37608 22052 38424 22080
rect 39960 22052 40417 22080
rect 37608 22040 37614 22052
rect 27893 22015 27951 22021
rect 27893 21981 27905 22015
rect 27939 22012 27951 22015
rect 27982 22012 27988 22024
rect 27939 21984 27988 22012
rect 27939 21981 27951 21984
rect 27893 21975 27951 21981
rect 27982 21972 27988 21984
rect 28040 21972 28046 22024
rect 28902 22012 28908 22024
rect 28863 21984 28908 22012
rect 28902 21972 28908 21984
rect 28960 21972 28966 22024
rect 33042 21972 33048 22024
rect 33100 22012 33106 22024
rect 33502 22012 33508 22024
rect 33100 21984 33508 22012
rect 33100 21972 33106 21984
rect 33502 21972 33508 21984
rect 33560 22012 33566 22024
rect 33597 22015 33655 22021
rect 33597 22012 33609 22015
rect 33560 21984 33609 22012
rect 33560 21972 33566 21984
rect 33597 21981 33609 21984
rect 33643 21981 33655 22015
rect 33597 21975 33655 21981
rect 37921 22015 37979 22021
rect 37921 21981 37933 22015
rect 37967 21981 37979 22015
rect 37921 21975 37979 21981
rect 27709 21879 27767 21885
rect 27709 21845 27721 21879
rect 27755 21876 27767 21879
rect 28258 21876 28264 21888
rect 27755 21848 28264 21876
rect 27755 21845 27767 21848
rect 27709 21839 27767 21845
rect 28258 21836 28264 21848
rect 28316 21836 28322 21888
rect 31202 21876 31208 21888
rect 31163 21848 31208 21876
rect 31202 21836 31208 21848
rect 31260 21836 31266 21888
rect 33226 21836 33232 21888
rect 33284 21876 33290 21888
rect 33413 21879 33471 21885
rect 33413 21876 33425 21879
rect 33284 21848 33425 21876
rect 33284 21836 33290 21848
rect 33413 21845 33425 21848
rect 33459 21845 33471 21879
rect 33413 21839 33471 21845
rect 36173 21879 36231 21885
rect 36173 21845 36185 21879
rect 36219 21876 36231 21879
rect 37550 21876 37556 21888
rect 36219 21848 37556 21876
rect 36219 21845 36231 21848
rect 36173 21839 36231 21845
rect 37550 21836 37556 21848
rect 37608 21836 37614 21888
rect 37936 21876 37964 21975
rect 38194 21972 38200 22024
rect 38252 22021 38258 22024
rect 38396 22021 38424 22052
rect 40405 22049 40417 22052
rect 40451 22080 40463 22083
rect 40770 22080 40776 22092
rect 40451 22052 40776 22080
rect 40451 22049 40463 22052
rect 40405 22043 40463 22049
rect 40770 22040 40776 22052
rect 40828 22040 40834 22092
rect 40865 22083 40923 22089
rect 40865 22049 40877 22083
rect 40911 22080 40923 22083
rect 41322 22080 41328 22092
rect 40911 22052 41328 22080
rect 40911 22049 40923 22052
rect 40865 22043 40923 22049
rect 41322 22040 41328 22052
rect 41380 22040 41386 22092
rect 43438 22040 43444 22092
rect 43496 22080 43502 22092
rect 43717 22083 43775 22089
rect 43717 22080 43729 22083
rect 43496 22052 43729 22080
rect 43496 22040 43502 22052
rect 43717 22049 43729 22052
rect 43763 22049 43775 22083
rect 43717 22043 43775 22049
rect 43993 22083 44051 22089
rect 43993 22049 44005 22083
rect 44039 22080 44051 22083
rect 44744 22080 44772 22111
rect 44910 22108 44916 22120
rect 44968 22108 44974 22160
rect 44039 22052 44772 22080
rect 44039 22049 44051 22052
rect 43993 22043 44051 22049
rect 45554 22040 45560 22092
rect 45612 22080 45618 22092
rect 46365 22083 46423 22089
rect 46365 22080 46377 22083
rect 45612 22052 46377 22080
rect 45612 22040 45618 22052
rect 46365 22049 46377 22052
rect 46411 22080 46423 22083
rect 46842 22080 46848 22092
rect 46411 22052 46848 22080
rect 46411 22049 46423 22052
rect 46365 22043 46423 22049
rect 46842 22040 46848 22052
rect 46900 22040 46906 22092
rect 38252 22015 38302 22021
rect 38252 21981 38256 22015
rect 38290 21981 38302 22015
rect 38252 21975 38302 21981
rect 38381 22015 38439 22021
rect 38381 21981 38393 22015
rect 38427 21981 38439 22015
rect 38654 22012 38660 22024
rect 38615 21984 38660 22012
rect 38381 21975 38439 21981
rect 38252 21972 38258 21975
rect 38654 21972 38660 21984
rect 38712 21972 38718 22024
rect 41598 22012 41604 22024
rect 41559 21984 41604 22012
rect 41598 21972 41604 21984
rect 41656 21972 41662 22024
rect 46106 22012 46112 22024
rect 46067 21984 46112 22012
rect 46106 21972 46112 21984
rect 46164 21972 46170 22024
rect 41046 21944 41052 21956
rect 41007 21916 41052 21944
rect 41046 21904 41052 21916
rect 41104 21904 41110 21956
rect 47486 21944 47492 21956
rect 47447 21916 47492 21944
rect 47486 21904 47492 21916
rect 47544 21904 47550 21956
rect 38286 21876 38292 21888
rect 37936 21848 38292 21876
rect 38286 21836 38292 21848
rect 38344 21876 38350 21888
rect 38746 21876 38752 21888
rect 38344 21848 38752 21876
rect 38344 21836 38350 21848
rect 38746 21836 38752 21848
rect 38804 21836 38810 21888
rect 42334 21836 42340 21888
rect 42392 21876 42398 21888
rect 43441 21879 43499 21885
rect 43441 21876 43453 21879
rect 42392 21848 43453 21876
rect 42392 21836 42398 21848
rect 43441 21845 43453 21848
rect 43487 21845 43499 21879
rect 43441 21839 43499 21845
rect 1104 21786 48852 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 34966 21786
rect 35018 21734 35030 21786
rect 35082 21734 35094 21786
rect 35146 21734 35158 21786
rect 35210 21734 48852 21786
rect 1104 21712 48852 21734
rect 28902 21632 28908 21684
rect 28960 21672 28966 21684
rect 28997 21675 29055 21681
rect 28997 21672 29009 21675
rect 28960 21644 29009 21672
rect 28960 21632 28966 21644
rect 28997 21641 29009 21644
rect 29043 21672 29055 21675
rect 29730 21672 29736 21684
rect 29043 21644 29736 21672
rect 29043 21641 29055 21644
rect 28997 21635 29055 21641
rect 29730 21632 29736 21644
rect 29788 21632 29794 21684
rect 32398 21632 32404 21684
rect 32456 21672 32462 21684
rect 32493 21675 32551 21681
rect 32493 21672 32505 21675
rect 32456 21644 32505 21672
rect 32456 21632 32462 21644
rect 32493 21641 32505 21644
rect 32539 21641 32551 21675
rect 32493 21635 32551 21641
rect 37277 21675 37335 21681
rect 37277 21641 37289 21675
rect 37323 21672 37335 21675
rect 37366 21672 37372 21684
rect 37323 21644 37372 21672
rect 37323 21641 37335 21644
rect 37277 21635 37335 21641
rect 37366 21632 37372 21644
rect 37424 21632 37430 21684
rect 37550 21672 37556 21684
rect 37511 21644 37556 21672
rect 37550 21632 37556 21644
rect 37608 21632 37614 21684
rect 38654 21672 38660 21684
rect 38567 21644 38660 21672
rect 38654 21632 38660 21644
rect 38712 21672 38718 21684
rect 41414 21672 41420 21684
rect 38712 21644 41420 21672
rect 38712 21632 38718 21644
rect 41414 21632 41420 21644
rect 41472 21672 41478 21684
rect 42613 21675 42671 21681
rect 42613 21672 42625 21675
rect 41472 21644 42625 21672
rect 41472 21632 41478 21644
rect 42613 21641 42625 21644
rect 42659 21641 42671 21675
rect 43438 21672 43444 21684
rect 43399 21644 43444 21672
rect 42613 21635 42671 21641
rect 43438 21632 43444 21644
rect 43496 21632 43502 21684
rect 44821 21675 44879 21681
rect 44821 21641 44833 21675
rect 44867 21672 44879 21675
rect 44910 21672 44916 21684
rect 44867 21644 44916 21672
rect 44867 21641 44879 21644
rect 44821 21635 44879 21641
rect 44910 21632 44916 21644
rect 44968 21632 44974 21684
rect 45554 21672 45560 21684
rect 45515 21644 45560 21672
rect 45554 21632 45560 21644
rect 45612 21632 45618 21684
rect 46842 21632 46848 21684
rect 46900 21672 46906 21684
rect 47489 21675 47547 21681
rect 47489 21672 47501 21675
rect 46900 21644 47501 21672
rect 46900 21632 46906 21644
rect 47489 21641 47501 21644
rect 47535 21641 47547 21675
rect 47489 21635 47547 21641
rect 27709 21607 27767 21613
rect 27709 21573 27721 21607
rect 27755 21604 27767 21607
rect 27890 21604 27896 21616
rect 27755 21576 27896 21604
rect 27755 21573 27767 21576
rect 27709 21567 27767 21573
rect 27890 21564 27896 21576
rect 27948 21564 27954 21616
rect 29365 21607 29423 21613
rect 29365 21573 29377 21607
rect 29411 21573 29423 21607
rect 29365 21567 29423 21573
rect 28258 21536 28264 21548
rect 28219 21508 28264 21536
rect 28258 21496 28264 21508
rect 28316 21496 28322 21548
rect 27525 21471 27583 21477
rect 27525 21437 27537 21471
rect 27571 21468 27583 21471
rect 27982 21468 27988 21480
rect 27571 21440 27988 21468
rect 27571 21437 27583 21440
rect 27525 21431 27583 21437
rect 27982 21428 27988 21440
rect 28040 21428 28046 21480
rect 29380 21468 29408 21567
rect 43162 21564 43168 21616
rect 43220 21604 43226 21616
rect 43809 21607 43867 21613
rect 43809 21604 43821 21607
rect 43220 21576 43821 21604
rect 43220 21564 43226 21576
rect 43809 21573 43821 21576
rect 43855 21604 43867 21607
rect 43898 21604 43904 21616
rect 43855 21576 43904 21604
rect 43855 21573 43867 21576
rect 43809 21567 43867 21573
rect 43898 21564 43904 21576
rect 43956 21564 43962 21616
rect 29914 21536 29920 21548
rect 29875 21508 29920 21536
rect 29914 21496 29920 21508
rect 29972 21496 29978 21548
rect 40313 21539 40371 21545
rect 40313 21505 40325 21539
rect 40359 21536 40371 21539
rect 41233 21539 41291 21545
rect 41233 21536 41245 21539
rect 40359 21508 41245 21536
rect 40359 21505 40371 21508
rect 40313 21499 40371 21505
rect 41233 21505 41245 21508
rect 41279 21536 41291 21539
rect 41322 21536 41328 21548
rect 41279 21508 41328 21536
rect 41279 21505 41291 21508
rect 41233 21499 41291 21505
rect 41322 21496 41328 21508
rect 41380 21536 41386 21548
rect 41966 21536 41972 21548
rect 41380 21508 41972 21536
rect 41380 21496 41386 21508
rect 41966 21496 41972 21508
rect 42024 21496 42030 21548
rect 44174 21496 44180 21548
rect 44232 21536 44238 21548
rect 44361 21539 44419 21545
rect 44361 21536 44373 21539
rect 44232 21508 44373 21536
rect 44232 21496 44238 21508
rect 44361 21505 44373 21508
rect 44407 21536 44419 21539
rect 45097 21539 45155 21545
rect 45097 21536 45109 21539
rect 44407 21508 45109 21536
rect 44407 21505 44419 21508
rect 44361 21499 44419 21505
rect 45097 21505 45109 21508
rect 45143 21505 45155 21539
rect 45097 21499 45155 21505
rect 45925 21539 45983 21545
rect 45925 21505 45937 21539
rect 45971 21536 45983 21539
rect 46106 21536 46112 21548
rect 45971 21508 46112 21536
rect 45971 21505 45983 21508
rect 45925 21499 45983 21505
rect 46106 21496 46112 21508
rect 46164 21496 46170 21548
rect 30285 21471 30343 21477
rect 30285 21468 30297 21471
rect 28184 21440 29408 21468
rect 29656 21440 30297 21468
rect 28184 21409 28212 21440
rect 29656 21412 29684 21440
rect 30285 21437 30297 21440
rect 30331 21437 30343 21471
rect 30285 21431 30343 21437
rect 31113 21471 31171 21477
rect 31113 21437 31125 21471
rect 31159 21437 31171 21471
rect 31113 21431 31171 21437
rect 27157 21403 27215 21409
rect 27157 21369 27169 21403
rect 27203 21400 27215 21403
rect 28169 21403 28227 21409
rect 28169 21400 28181 21403
rect 27203 21372 28181 21400
rect 27203 21369 27215 21372
rect 27157 21363 27215 21369
rect 28169 21369 28181 21372
rect 28215 21369 28227 21403
rect 29638 21400 29644 21412
rect 29599 21372 29644 21400
rect 28169 21363 28227 21369
rect 29638 21360 29644 21372
rect 29696 21360 29702 21412
rect 29730 21360 29736 21412
rect 29788 21400 29794 21412
rect 31021 21403 31079 21409
rect 31021 21400 31033 21403
rect 29788 21372 31033 21400
rect 29788 21360 29794 21372
rect 31021 21369 31033 21372
rect 31067 21400 31079 21403
rect 31128 21400 31156 21431
rect 31202 21428 31208 21480
rect 31260 21468 31266 21480
rect 31369 21471 31427 21477
rect 31369 21468 31381 21471
rect 31260 21440 31381 21468
rect 31260 21428 31266 21440
rect 31369 21437 31381 21440
rect 31415 21437 31427 21471
rect 31369 21431 31427 21437
rect 33594 21428 33600 21480
rect 33652 21468 33658 21480
rect 33965 21471 34023 21477
rect 33965 21468 33977 21471
rect 33652 21440 33977 21468
rect 33652 21428 33658 21440
rect 33965 21437 33977 21440
rect 34011 21437 34023 21471
rect 33965 21431 34023 21437
rect 35161 21471 35219 21477
rect 35161 21437 35173 21471
rect 35207 21468 35219 21471
rect 35253 21471 35311 21477
rect 35253 21468 35265 21471
rect 35207 21440 35265 21468
rect 35207 21437 35219 21440
rect 35161 21431 35219 21437
rect 35253 21437 35265 21440
rect 35299 21468 35311 21471
rect 35802 21468 35808 21480
rect 35299 21440 35808 21468
rect 35299 21437 35311 21440
rect 35253 21431 35311 21437
rect 31662 21400 31668 21412
rect 31067 21372 31668 21400
rect 31067 21369 31079 21372
rect 31021 21363 31079 21369
rect 31662 21360 31668 21372
rect 31720 21360 31726 21412
rect 33502 21360 33508 21412
rect 33560 21400 33566 21412
rect 33689 21403 33747 21409
rect 33689 21400 33701 21403
rect 33560 21372 33701 21400
rect 33560 21360 33566 21372
rect 33689 21369 33701 21372
rect 33735 21400 33747 21403
rect 35176 21400 35204 21431
rect 35802 21428 35808 21440
rect 35860 21428 35866 21480
rect 40770 21468 40776 21480
rect 40731 21440 40776 21468
rect 40770 21428 40776 21440
rect 40828 21428 40834 21480
rect 41509 21471 41567 21477
rect 41509 21468 41521 21471
rect 40880 21440 41521 21468
rect 35526 21409 35532 21412
rect 35520 21400 35532 21409
rect 33735 21372 35204 21400
rect 35487 21372 35532 21400
rect 33735 21369 33747 21372
rect 33689 21363 33747 21369
rect 35520 21363 35532 21372
rect 35526 21360 35532 21363
rect 35584 21360 35590 21412
rect 36446 21360 36452 21412
rect 36504 21400 36510 21412
rect 37737 21403 37795 21409
rect 37737 21400 37749 21403
rect 36504 21372 37749 21400
rect 36504 21360 36510 21372
rect 37737 21369 37749 21372
rect 37783 21369 37795 21403
rect 37737 21363 37795 21369
rect 39945 21403 40003 21409
rect 39945 21369 39957 21403
rect 39991 21400 40003 21403
rect 40880 21400 40908 21440
rect 41509 21437 41521 21440
rect 41555 21468 41567 21471
rect 42794 21468 42800 21480
rect 41555 21440 42800 21468
rect 41555 21437 41567 21440
rect 41509 21431 41567 21437
rect 42794 21428 42800 21440
rect 42852 21428 42858 21480
rect 44082 21400 44088 21412
rect 39991 21372 40908 21400
rect 44043 21372 44088 21400
rect 39991 21369 40003 21372
rect 39945 21363 40003 21369
rect 44082 21360 44088 21372
rect 44140 21360 44146 21412
rect 46382 21409 46388 21412
rect 46376 21400 46388 21409
rect 46343 21372 46388 21400
rect 46376 21363 46388 21372
rect 46382 21360 46388 21363
rect 46440 21360 46446 21412
rect 29822 21332 29828 21344
rect 29783 21304 29828 21332
rect 29822 21292 29828 21304
rect 29880 21292 29886 21344
rect 36630 21332 36636 21344
rect 36591 21304 36636 21332
rect 36630 21292 36636 21304
rect 36688 21292 36694 21344
rect 38194 21332 38200 21344
rect 38155 21304 38200 21332
rect 38194 21292 38200 21304
rect 38252 21292 38258 21344
rect 40770 21292 40776 21344
rect 40828 21332 40834 21344
rect 41235 21335 41293 21341
rect 41235 21332 41247 21335
rect 40828 21304 41247 21332
rect 40828 21292 40834 21304
rect 41235 21301 41247 21304
rect 41281 21301 41293 21335
rect 41235 21295 41293 21301
rect 44174 21292 44180 21344
rect 44232 21332 44238 21344
rect 44269 21335 44327 21341
rect 44269 21332 44281 21335
rect 44232 21304 44281 21332
rect 44232 21292 44238 21304
rect 44269 21301 44281 21304
rect 44315 21301 44327 21335
rect 44269 21295 44327 21301
rect 1104 21242 48852 21264
rect 1104 21190 19606 21242
rect 19658 21190 19670 21242
rect 19722 21190 19734 21242
rect 19786 21190 19798 21242
rect 19850 21190 48852 21242
rect 1104 21168 48852 21190
rect 29273 21131 29331 21137
rect 29273 21097 29285 21131
rect 29319 21097 29331 21131
rect 29273 21091 29331 21097
rect 36173 21131 36231 21137
rect 36173 21097 36185 21131
rect 36219 21128 36231 21131
rect 36446 21128 36452 21140
rect 36219 21100 36452 21128
rect 36219 21097 36231 21100
rect 36173 21091 36231 21097
rect 29288 21060 29316 21091
rect 36446 21088 36452 21100
rect 36504 21088 36510 21140
rect 36538 21088 36544 21140
rect 36596 21128 36602 21140
rect 41233 21131 41291 21137
rect 36596 21100 36641 21128
rect 36596 21088 36602 21100
rect 41233 21097 41245 21131
rect 41279 21128 41291 21131
rect 41414 21128 41420 21140
rect 41279 21100 41420 21128
rect 41279 21097 41291 21100
rect 41233 21091 41291 21097
rect 41414 21088 41420 21100
rect 41472 21088 41478 21140
rect 41598 21128 41604 21140
rect 41559 21100 41604 21128
rect 41598 21088 41604 21100
rect 41656 21088 41662 21140
rect 42334 21128 42340 21140
rect 42295 21100 42340 21128
rect 42334 21088 42340 21100
rect 42392 21088 42398 21140
rect 43162 21128 43168 21140
rect 43123 21100 43168 21128
rect 43162 21088 43168 21100
rect 43220 21088 43226 21140
rect 43438 21128 43444 21140
rect 43399 21100 43444 21128
rect 43438 21088 43444 21100
rect 43496 21088 43502 21140
rect 43993 21131 44051 21137
rect 43993 21097 44005 21131
rect 44039 21128 44051 21131
rect 44082 21128 44088 21140
rect 44039 21100 44088 21128
rect 44039 21097 44051 21100
rect 43993 21091 44051 21097
rect 44082 21088 44088 21100
rect 44140 21088 44146 21140
rect 46106 21128 46112 21140
rect 46067 21100 46112 21128
rect 46106 21088 46112 21100
rect 46164 21088 46170 21140
rect 46937 21131 46995 21137
rect 46937 21097 46949 21131
rect 46983 21128 46995 21131
rect 47210 21128 47216 21140
rect 46983 21100 47216 21128
rect 46983 21097 46995 21100
rect 46937 21091 46995 21097
rect 47210 21088 47216 21100
rect 47268 21088 47274 21140
rect 30926 21060 30932 21072
rect 29288 21032 30932 21060
rect 30926 21020 30932 21032
rect 30984 21020 30990 21072
rect 31021 21063 31079 21069
rect 31021 21029 31033 21063
rect 31067 21060 31079 21063
rect 31202 21060 31208 21072
rect 31067 21032 31208 21060
rect 31067 21029 31079 21032
rect 31021 21023 31079 21029
rect 31202 21020 31208 21032
rect 31260 21020 31266 21072
rect 35345 21063 35403 21069
rect 35345 21029 35357 21063
rect 35391 21060 35403 21063
rect 35526 21060 35532 21072
rect 35391 21032 35532 21060
rect 35391 21029 35403 21032
rect 35345 21023 35403 21029
rect 35526 21020 35532 21032
rect 35584 21060 35590 21072
rect 36556 21060 36584 21088
rect 35584 21032 36584 21060
rect 35584 21020 35590 21032
rect 44634 21020 44640 21072
rect 44692 21060 44698 21072
rect 45005 21063 45063 21069
rect 45005 21060 45017 21063
rect 44692 21032 45017 21060
rect 44692 21020 44698 21032
rect 45005 21029 45017 21032
rect 45051 21029 45063 21063
rect 45005 21023 45063 21029
rect 28074 20952 28080 21004
rect 28132 20992 28138 21004
rect 28169 20995 28227 21001
rect 28169 20992 28181 20995
rect 28132 20964 28181 20992
rect 28132 20952 28138 20964
rect 28169 20961 28181 20964
rect 28215 20961 28227 20995
rect 28169 20955 28227 20961
rect 32490 20952 32496 21004
rect 32548 20992 32554 21004
rect 32724 20995 32782 21001
rect 32724 20992 32736 20995
rect 32548 20964 32736 20992
rect 32548 20952 32554 20964
rect 32724 20961 32736 20964
rect 32770 20961 32782 20995
rect 32724 20955 32782 20961
rect 44174 20952 44180 21004
rect 44232 20992 44238 21004
rect 44821 20995 44879 21001
rect 44821 20992 44833 20995
rect 44232 20964 44833 20992
rect 44232 20952 44238 20964
rect 44821 20961 44833 20964
rect 44867 20961 44879 20995
rect 46750 20992 46756 21004
rect 46711 20964 46756 20992
rect 44821 20955 44879 20961
rect 46750 20952 46756 20964
rect 46808 20952 46814 21004
rect 27246 20884 27252 20936
rect 27304 20924 27310 20936
rect 27433 20927 27491 20933
rect 27433 20924 27445 20927
rect 27304 20896 27445 20924
rect 27304 20884 27310 20896
rect 27433 20893 27445 20896
rect 27479 20893 27491 20927
rect 27433 20887 27491 20893
rect 27614 20884 27620 20936
rect 27672 20924 27678 20936
rect 27756 20927 27814 20933
rect 27756 20924 27768 20927
rect 27672 20896 27768 20924
rect 27672 20884 27678 20896
rect 27756 20893 27768 20896
rect 27802 20893 27814 20927
rect 27890 20924 27896 20936
rect 27851 20896 27896 20924
rect 27756 20887 27814 20893
rect 27890 20884 27896 20896
rect 27948 20884 27954 20936
rect 30837 20927 30895 20933
rect 30837 20924 30849 20927
rect 30576 20896 30849 20924
rect 30466 20856 30472 20868
rect 30427 20828 30472 20856
rect 30466 20816 30472 20828
rect 30524 20816 30530 20868
rect 29822 20748 29828 20800
rect 29880 20788 29886 20800
rect 29917 20791 29975 20797
rect 29917 20788 29929 20791
rect 29880 20760 29929 20788
rect 29880 20748 29886 20760
rect 29917 20757 29929 20760
rect 29963 20788 29975 20791
rect 30374 20788 30380 20800
rect 29963 20760 30380 20788
rect 29963 20757 29975 20760
rect 29917 20751 29975 20757
rect 30374 20748 30380 20760
rect 30432 20788 30438 20800
rect 30576 20788 30604 20896
rect 30837 20893 30849 20896
rect 30883 20893 30895 20927
rect 30837 20887 30895 20893
rect 32401 20927 32459 20933
rect 32401 20893 32413 20927
rect 32447 20893 32459 20927
rect 32858 20924 32864 20936
rect 32819 20896 32864 20924
rect 32401 20887 32459 20893
rect 30432 20760 30604 20788
rect 32416 20788 32444 20887
rect 32858 20884 32864 20896
rect 32916 20884 32922 20936
rect 33042 20884 33048 20936
rect 33100 20924 33106 20936
rect 33137 20927 33195 20933
rect 33137 20924 33149 20927
rect 33100 20896 33149 20924
rect 33100 20884 33106 20896
rect 33137 20893 33149 20896
rect 33183 20893 33195 20927
rect 40310 20924 40316 20936
rect 40271 20896 40316 20924
rect 33137 20887 33195 20893
rect 40310 20884 40316 20896
rect 40368 20884 40374 20936
rect 45094 20924 45100 20936
rect 45055 20896 45100 20924
rect 45094 20884 45100 20896
rect 45152 20924 45158 20936
rect 46382 20924 46388 20936
rect 45152 20896 46388 20924
rect 45152 20884 45158 20896
rect 46382 20884 46388 20896
rect 46440 20924 46446 20936
rect 46477 20927 46535 20933
rect 46477 20924 46489 20927
rect 46440 20896 46489 20924
rect 46440 20884 46446 20896
rect 46477 20893 46489 20896
rect 46523 20893 46535 20927
rect 46477 20887 46535 20893
rect 44545 20859 44603 20865
rect 44545 20825 44557 20859
rect 44591 20856 44603 20859
rect 45462 20856 45468 20868
rect 44591 20828 45468 20856
rect 44591 20825 44603 20828
rect 44545 20819 44603 20825
rect 45462 20816 45468 20828
rect 45520 20816 45526 20868
rect 32766 20788 32772 20800
rect 32416 20760 32772 20788
rect 30432 20748 30438 20760
rect 32766 20748 32772 20760
rect 32824 20748 32830 20800
rect 34238 20788 34244 20800
rect 34199 20760 34244 20788
rect 34238 20748 34244 20760
rect 34296 20748 34302 20800
rect 38010 20788 38016 20800
rect 37971 20760 38016 20788
rect 38010 20748 38016 20760
rect 38068 20748 38074 20800
rect 38286 20788 38292 20800
rect 38247 20760 38292 20788
rect 38286 20748 38292 20760
rect 38344 20748 38350 20800
rect 40770 20788 40776 20800
rect 40731 20760 40776 20788
rect 40770 20748 40776 20760
rect 40828 20788 40834 20800
rect 41322 20788 41328 20800
rect 40828 20760 41328 20788
rect 40828 20748 40834 20760
rect 41322 20748 41328 20760
rect 41380 20748 41386 20800
rect 44174 20748 44180 20800
rect 44232 20788 44238 20800
rect 44269 20791 44327 20797
rect 44269 20788 44281 20791
rect 44232 20760 44281 20788
rect 44232 20748 44238 20760
rect 44269 20757 44281 20760
rect 44315 20757 44327 20791
rect 44269 20751 44327 20757
rect 1104 20698 48852 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 34966 20698
rect 35018 20646 35030 20698
rect 35082 20646 35094 20698
rect 35146 20646 35158 20698
rect 35210 20646 48852 20698
rect 1104 20624 48852 20646
rect 27890 20544 27896 20596
rect 27948 20584 27954 20596
rect 28169 20587 28227 20593
rect 28169 20584 28181 20587
rect 27948 20556 28181 20584
rect 27948 20544 27954 20556
rect 28169 20553 28181 20556
rect 28215 20553 28227 20587
rect 28169 20547 28227 20553
rect 30926 20544 30932 20596
rect 30984 20584 30990 20596
rect 31757 20587 31815 20593
rect 31757 20584 31769 20587
rect 30984 20556 31769 20584
rect 30984 20544 30990 20556
rect 31757 20553 31769 20556
rect 31803 20584 31815 20587
rect 33042 20584 33048 20596
rect 31803 20556 33048 20584
rect 31803 20553 31815 20556
rect 31757 20547 31815 20553
rect 33042 20544 33048 20556
rect 33100 20544 33106 20596
rect 33226 20584 33232 20596
rect 33187 20556 33232 20584
rect 33226 20544 33232 20556
rect 33284 20544 33290 20596
rect 34698 20544 34704 20596
rect 34756 20584 34762 20596
rect 35802 20584 35808 20596
rect 34756 20556 35808 20584
rect 34756 20544 34762 20556
rect 35802 20544 35808 20556
rect 35860 20584 35866 20596
rect 37737 20587 37795 20593
rect 37737 20584 37749 20587
rect 35860 20556 37749 20584
rect 35860 20544 35866 20556
rect 37737 20553 37749 20556
rect 37783 20553 37795 20587
rect 40310 20584 40316 20596
rect 40271 20556 40316 20584
rect 37737 20547 37795 20553
rect 31018 20516 31024 20528
rect 30979 20488 31024 20516
rect 31018 20476 31024 20488
rect 31076 20476 31082 20528
rect 32398 20516 32404 20528
rect 32359 20488 32404 20516
rect 32398 20476 32404 20488
rect 32456 20476 32462 20528
rect 37752 20460 37780 20547
rect 40310 20544 40316 20556
rect 40368 20544 40374 20596
rect 40586 20584 40592 20596
rect 40547 20556 40592 20584
rect 40586 20544 40592 20556
rect 40644 20544 40650 20596
rect 41414 20544 41420 20596
rect 41472 20584 41478 20596
rect 42061 20587 42119 20593
rect 42061 20584 42073 20587
rect 41472 20556 42073 20584
rect 41472 20544 41478 20556
rect 42061 20553 42073 20556
rect 42107 20553 42119 20587
rect 42061 20547 42119 20553
rect 27893 20451 27951 20457
rect 27893 20417 27905 20451
rect 27939 20448 27951 20451
rect 28074 20448 28080 20460
rect 27939 20420 28080 20448
rect 27939 20417 27951 20420
rect 27893 20411 27951 20417
rect 28074 20408 28080 20420
rect 28132 20408 28138 20460
rect 37734 20448 37740 20460
rect 37647 20420 37740 20448
rect 37734 20408 37740 20420
rect 37792 20448 37798 20460
rect 37921 20451 37979 20457
rect 37921 20448 37933 20451
rect 37792 20420 37933 20448
rect 37792 20408 37798 20420
rect 37921 20417 37933 20420
rect 37967 20417 37979 20451
rect 40328 20448 40356 20544
rect 40957 20451 41015 20457
rect 40957 20448 40969 20451
rect 40328 20420 40969 20448
rect 37921 20411 37979 20417
rect 40957 20417 40969 20420
rect 41003 20417 41015 20451
rect 42076 20448 42104 20547
rect 42794 20544 42800 20596
rect 42852 20584 42858 20596
rect 44085 20587 44143 20593
rect 44085 20584 44097 20587
rect 42852 20556 44097 20584
rect 42852 20544 42858 20556
rect 44085 20553 44097 20556
rect 44131 20553 44143 20587
rect 44085 20547 44143 20553
rect 44100 20516 44128 20547
rect 44174 20544 44180 20596
rect 44232 20584 44238 20596
rect 45005 20587 45063 20593
rect 45005 20584 45017 20587
rect 44232 20556 45017 20584
rect 44232 20544 44238 20556
rect 45005 20553 45017 20556
rect 45051 20553 45063 20587
rect 46750 20584 46756 20596
rect 46711 20556 46756 20584
rect 45005 20547 45063 20553
rect 46750 20544 46756 20556
rect 46808 20544 46814 20596
rect 44634 20516 44640 20528
rect 44100 20488 44640 20516
rect 44634 20476 44640 20488
rect 44692 20476 44698 20528
rect 42076 20420 42380 20448
rect 40957 20411 41015 20417
rect 29549 20383 29607 20389
rect 29549 20349 29561 20383
rect 29595 20380 29607 20383
rect 29641 20383 29699 20389
rect 29641 20380 29653 20383
rect 29595 20352 29653 20380
rect 29595 20349 29607 20352
rect 29549 20343 29607 20349
rect 29641 20349 29653 20352
rect 29687 20380 29699 20383
rect 29730 20380 29736 20392
rect 29687 20352 29736 20380
rect 29687 20349 29699 20352
rect 29641 20343 29699 20349
rect 29730 20340 29736 20352
rect 29788 20340 29794 20392
rect 29914 20389 29920 20392
rect 29908 20380 29920 20389
rect 29875 20352 29920 20380
rect 29908 20343 29920 20352
rect 29914 20340 29920 20343
rect 29972 20340 29978 20392
rect 38010 20340 38016 20392
rect 38068 20380 38074 20392
rect 38177 20383 38235 20389
rect 38177 20380 38189 20383
rect 38068 20352 38189 20380
rect 38068 20340 38074 20352
rect 38177 20349 38189 20352
rect 38223 20349 38235 20383
rect 38177 20343 38235 20349
rect 40678 20340 40684 20392
rect 40736 20380 40742 20392
rect 42242 20380 42248 20392
rect 40736 20352 42248 20380
rect 40736 20340 40742 20352
rect 42242 20340 42248 20352
rect 42300 20340 42306 20392
rect 42352 20380 42380 20420
rect 42426 20408 42432 20460
rect 42484 20448 42490 20460
rect 42705 20451 42763 20457
rect 42705 20448 42717 20451
rect 42484 20420 42717 20448
rect 42484 20408 42490 20420
rect 42705 20417 42717 20420
rect 42751 20417 42763 20451
rect 42978 20448 42984 20460
rect 42891 20420 42984 20448
rect 42705 20411 42763 20417
rect 42978 20408 42984 20420
rect 43036 20448 43042 20460
rect 43990 20448 43996 20460
rect 43036 20420 43996 20448
rect 43036 20408 43042 20420
rect 43990 20408 43996 20420
rect 44048 20408 44054 20460
rect 42568 20383 42626 20389
rect 42568 20380 42580 20383
rect 42352 20352 42580 20380
rect 42568 20349 42580 20352
rect 42614 20349 42626 20383
rect 42568 20343 42626 20349
rect 32125 20315 32183 20321
rect 32125 20281 32137 20315
rect 32171 20312 32183 20315
rect 32858 20312 32864 20324
rect 32171 20284 32864 20312
rect 32171 20281 32183 20284
rect 32125 20275 32183 20281
rect 32858 20272 32864 20284
rect 32916 20312 32922 20324
rect 33226 20312 33232 20324
rect 32916 20284 33232 20312
rect 32916 20272 32922 20284
rect 33226 20272 33232 20284
rect 33284 20312 33290 20324
rect 33505 20315 33563 20321
rect 33505 20312 33517 20315
rect 33284 20284 33517 20312
rect 33284 20272 33290 20284
rect 33505 20281 33517 20284
rect 33551 20281 33563 20315
rect 33505 20275 33563 20281
rect 33594 20272 33600 20324
rect 33652 20312 33658 20324
rect 33781 20315 33839 20321
rect 33781 20312 33793 20315
rect 33652 20284 33793 20312
rect 33652 20272 33658 20284
rect 33781 20281 33793 20284
rect 33827 20281 33839 20315
rect 41141 20315 41199 20321
rect 41141 20312 41153 20315
rect 33781 20275 33839 20281
rect 39868 20284 41153 20312
rect 39868 20256 39896 20284
rect 41141 20281 41153 20284
rect 41187 20312 41199 20315
rect 41598 20312 41604 20324
rect 41187 20284 41604 20312
rect 41187 20281 41199 20284
rect 41141 20275 41199 20281
rect 41598 20272 41604 20284
rect 41656 20272 41662 20324
rect 27157 20247 27215 20253
rect 27157 20213 27169 20247
rect 27203 20244 27215 20247
rect 27246 20244 27252 20256
rect 27203 20216 27252 20244
rect 27203 20213 27215 20216
rect 27157 20207 27215 20213
rect 27246 20204 27252 20216
rect 27304 20204 27310 20256
rect 27430 20244 27436 20256
rect 27391 20216 27436 20244
rect 27430 20204 27436 20216
rect 27488 20204 27494 20256
rect 33045 20247 33103 20253
rect 33045 20213 33057 20247
rect 33091 20244 33103 20247
rect 33689 20247 33747 20253
rect 33689 20244 33701 20247
rect 33091 20216 33701 20244
rect 33091 20213 33103 20216
rect 33045 20207 33103 20213
rect 33689 20213 33701 20216
rect 33735 20244 33747 20247
rect 34238 20244 34244 20256
rect 33735 20216 34244 20244
rect 33735 20213 33747 20216
rect 33689 20207 33747 20213
rect 34238 20204 34244 20216
rect 34296 20244 34302 20256
rect 34514 20244 34520 20256
rect 34296 20216 34520 20244
rect 34296 20204 34302 20216
rect 34514 20204 34520 20216
rect 34572 20204 34578 20256
rect 35161 20247 35219 20253
rect 35161 20213 35173 20247
rect 35207 20244 35219 20247
rect 35434 20244 35440 20256
rect 35207 20216 35440 20244
rect 35207 20213 35219 20216
rect 35161 20207 35219 20213
rect 35434 20204 35440 20216
rect 35492 20204 35498 20256
rect 36909 20247 36967 20253
rect 36909 20213 36921 20247
rect 36955 20244 36967 20247
rect 37182 20244 37188 20256
rect 36955 20216 37188 20244
rect 36955 20213 36967 20216
rect 36909 20207 36967 20213
rect 37182 20204 37188 20216
rect 37240 20204 37246 20256
rect 39298 20244 39304 20256
rect 39259 20216 39304 20244
rect 39298 20204 39304 20216
rect 39356 20204 39362 20256
rect 39850 20244 39856 20256
rect 39811 20216 39856 20244
rect 39850 20204 39856 20216
rect 39908 20204 39914 20256
rect 40586 20204 40592 20256
rect 40644 20244 40650 20256
rect 41049 20247 41107 20253
rect 41049 20244 41061 20247
rect 40644 20216 41061 20244
rect 40644 20204 40650 20216
rect 41049 20213 41061 20216
rect 41095 20244 41107 20247
rect 41509 20247 41567 20253
rect 41509 20244 41521 20247
rect 41095 20216 41521 20244
rect 41095 20213 41107 20216
rect 41049 20207 41107 20213
rect 41509 20213 41521 20216
rect 41555 20213 41567 20247
rect 41509 20207 41567 20213
rect 1104 20154 48852 20176
rect 1104 20102 19606 20154
rect 19658 20102 19670 20154
rect 19722 20102 19734 20154
rect 19786 20102 19798 20154
rect 19850 20102 48852 20154
rect 1104 20080 48852 20102
rect 29733 20043 29791 20049
rect 29733 20009 29745 20043
rect 29779 20040 29791 20043
rect 29914 20040 29920 20052
rect 29779 20012 29920 20040
rect 29779 20009 29791 20012
rect 29733 20003 29791 20009
rect 29914 20000 29920 20012
rect 29972 20000 29978 20052
rect 30469 20043 30527 20049
rect 30469 20009 30481 20043
rect 30515 20040 30527 20043
rect 30926 20040 30932 20052
rect 30515 20012 30932 20040
rect 30515 20009 30527 20012
rect 30469 20003 30527 20009
rect 30926 20000 30932 20012
rect 30984 20000 30990 20052
rect 31202 20040 31208 20052
rect 31163 20012 31208 20040
rect 31202 20000 31208 20012
rect 31260 20000 31266 20052
rect 32309 20043 32367 20049
rect 32309 20009 32321 20043
rect 32355 20040 32367 20043
rect 33226 20040 33232 20052
rect 32355 20012 33232 20040
rect 32355 20009 32367 20012
rect 32309 20003 32367 20009
rect 33226 20000 33232 20012
rect 33284 20000 33290 20052
rect 33594 20040 33600 20052
rect 33555 20012 33600 20040
rect 33594 20000 33600 20012
rect 33652 20000 33658 20052
rect 38010 20000 38016 20052
rect 38068 20040 38074 20052
rect 38654 20040 38660 20052
rect 38068 20012 38660 20040
rect 38068 20000 38074 20012
rect 38654 20000 38660 20012
rect 38712 20040 38718 20052
rect 39117 20043 39175 20049
rect 39117 20040 39129 20043
rect 38712 20012 39129 20040
rect 38712 20000 38718 20012
rect 39117 20009 39129 20012
rect 39163 20009 39175 20043
rect 41598 20040 41604 20052
rect 41559 20012 41604 20040
rect 39117 20003 39175 20009
rect 41598 20000 41604 20012
rect 41656 20000 41662 20052
rect 42242 20000 42248 20052
rect 42300 20040 42306 20052
rect 42613 20043 42671 20049
rect 42613 20040 42625 20043
rect 42300 20012 42625 20040
rect 42300 20000 42306 20012
rect 42613 20009 42625 20012
rect 42659 20009 42671 20043
rect 42613 20003 42671 20009
rect 44545 20043 44603 20049
rect 44545 20009 44557 20043
rect 44591 20040 44603 20043
rect 45094 20040 45100 20052
rect 44591 20012 45100 20040
rect 44591 20009 44603 20012
rect 44545 20003 44603 20009
rect 45094 20000 45100 20012
rect 45152 20040 45158 20052
rect 46109 20043 46167 20049
rect 46109 20040 46121 20043
rect 45152 20012 46121 20040
rect 45152 20000 45158 20012
rect 46109 20009 46121 20012
rect 46155 20009 46167 20043
rect 47394 20040 47400 20052
rect 47355 20012 47400 20040
rect 46109 20003 46167 20009
rect 47394 20000 47400 20012
rect 47452 20000 47458 20052
rect 32766 19972 32772 19984
rect 32727 19944 32772 19972
rect 32766 19932 32772 19944
rect 32824 19932 32830 19984
rect 39298 19932 39304 19984
rect 39356 19972 39362 19984
rect 40218 19972 40224 19984
rect 39356 19944 40224 19972
rect 39356 19932 39362 19944
rect 40218 19932 40224 19944
rect 40276 19972 40282 19984
rect 40466 19975 40524 19981
rect 40466 19972 40478 19975
rect 40276 19944 40478 19972
rect 40276 19932 40282 19944
rect 40466 19941 40478 19944
rect 40512 19941 40524 19975
rect 40466 19935 40524 19941
rect 42150 19932 42156 19984
rect 42208 19972 42214 19984
rect 42337 19975 42395 19981
rect 42337 19972 42349 19975
rect 42208 19944 42349 19972
rect 42208 19932 42214 19944
rect 42337 19941 42349 19944
rect 42383 19972 42395 19975
rect 42978 19972 42984 19984
rect 42383 19944 42984 19972
rect 42383 19941 42395 19944
rect 42337 19935 42395 19941
rect 42978 19932 42984 19944
rect 43036 19932 43042 19984
rect 32122 19904 32128 19916
rect 32083 19876 32128 19904
rect 32122 19864 32128 19876
rect 32180 19864 32186 19916
rect 34606 19864 34612 19916
rect 34664 19904 34670 19916
rect 34974 19913 34980 19916
rect 34968 19904 34980 19913
rect 34664 19876 34980 19904
rect 34664 19864 34670 19876
rect 34968 19867 34980 19876
rect 34974 19864 34980 19867
rect 35032 19864 35038 19916
rect 37734 19904 37740 19916
rect 37695 19876 37740 19904
rect 37734 19864 37740 19876
rect 37792 19864 37798 19916
rect 38004 19907 38062 19913
rect 38004 19873 38016 19907
rect 38050 19904 38062 19907
rect 38378 19904 38384 19916
rect 38050 19876 38384 19904
rect 38050 19873 38062 19876
rect 38004 19867 38062 19873
rect 38378 19864 38384 19876
rect 38436 19864 38442 19916
rect 45002 19913 45008 19916
rect 44996 19904 45008 19913
rect 44963 19876 45008 19904
rect 44996 19867 45008 19876
rect 45002 19864 45008 19867
rect 45060 19864 45066 19916
rect 47213 19907 47271 19913
rect 47213 19873 47225 19907
rect 47259 19904 47271 19907
rect 47302 19904 47308 19916
rect 47259 19876 47308 19904
rect 47259 19873 47271 19876
rect 47213 19867 47271 19873
rect 47302 19864 47308 19876
rect 47360 19864 47366 19916
rect 29825 19839 29883 19845
rect 29825 19805 29837 19839
rect 29871 19836 29883 19839
rect 29914 19836 29920 19848
rect 29871 19808 29920 19836
rect 29871 19805 29883 19808
rect 29825 19799 29883 19805
rect 29914 19796 29920 19808
rect 29972 19796 29978 19848
rect 30374 19796 30380 19848
rect 30432 19836 30438 19848
rect 30745 19839 30803 19845
rect 30745 19836 30757 19839
rect 30432 19808 30757 19836
rect 30432 19796 30438 19808
rect 30745 19805 30757 19808
rect 30791 19805 30803 19839
rect 30745 19799 30803 19805
rect 34422 19796 34428 19848
rect 34480 19836 34486 19848
rect 34698 19836 34704 19848
rect 34480 19808 34704 19836
rect 34480 19796 34486 19808
rect 34698 19796 34704 19808
rect 34756 19796 34762 19848
rect 40221 19839 40279 19845
rect 40221 19805 40233 19839
rect 40267 19805 40279 19839
rect 43714 19836 43720 19848
rect 43675 19808 43720 19836
rect 40221 19799 40279 19805
rect 34609 19703 34667 19709
rect 34609 19669 34621 19703
rect 34655 19700 34667 19703
rect 34698 19700 34704 19712
rect 34655 19672 34704 19700
rect 34655 19669 34667 19672
rect 34609 19663 34667 19669
rect 34698 19660 34704 19672
rect 34756 19660 34762 19712
rect 36078 19700 36084 19712
rect 36039 19672 36084 19700
rect 36078 19660 36084 19672
rect 36136 19660 36142 19712
rect 40236 19700 40264 19799
rect 43714 19796 43720 19808
rect 43772 19796 43778 19848
rect 44726 19836 44732 19848
rect 44687 19808 44732 19836
rect 44726 19796 44732 19808
rect 44784 19796 44790 19848
rect 40402 19700 40408 19712
rect 40236 19672 40408 19700
rect 40402 19660 40408 19672
rect 40460 19660 40466 19712
rect 43625 19703 43683 19709
rect 43625 19669 43637 19703
rect 43671 19700 43683 19703
rect 44174 19700 44180 19712
rect 43671 19672 44180 19700
rect 43671 19669 43683 19672
rect 43625 19663 43683 19669
rect 44174 19660 44180 19672
rect 44232 19660 44238 19712
rect 1104 19610 48852 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 34966 19610
rect 35018 19558 35030 19610
rect 35082 19558 35094 19610
rect 35146 19558 35158 19610
rect 35210 19558 48852 19610
rect 1104 19536 48852 19558
rect 31113 19499 31171 19505
rect 31113 19465 31125 19499
rect 31159 19496 31171 19499
rect 31202 19496 31208 19508
rect 31159 19468 31208 19496
rect 31159 19465 31171 19468
rect 31113 19459 31171 19465
rect 31202 19456 31208 19468
rect 31260 19456 31266 19508
rect 37734 19496 37740 19508
rect 37695 19468 37740 19496
rect 37734 19456 37740 19468
rect 37792 19456 37798 19508
rect 40586 19496 40592 19508
rect 40547 19468 40592 19496
rect 40586 19456 40592 19468
rect 40644 19456 40650 19508
rect 43441 19499 43499 19505
rect 43441 19465 43453 19499
rect 43487 19496 43499 19499
rect 43714 19496 43720 19508
rect 43487 19468 43720 19496
rect 43487 19465 43499 19468
rect 43441 19459 43499 19465
rect 43714 19456 43720 19468
rect 43772 19456 43778 19508
rect 47302 19496 47308 19508
rect 47263 19468 47308 19496
rect 47302 19456 47308 19468
rect 47360 19456 47366 19508
rect 31018 19388 31024 19440
rect 31076 19428 31082 19440
rect 31665 19431 31723 19437
rect 31665 19428 31677 19431
rect 31076 19400 31677 19428
rect 31076 19388 31082 19400
rect 31665 19397 31677 19400
rect 31711 19397 31723 19431
rect 31665 19391 31723 19397
rect 29641 19363 29699 19369
rect 29641 19329 29653 19363
rect 29687 19360 29699 19363
rect 29730 19360 29736 19372
rect 29687 19332 29736 19360
rect 29687 19329 29699 19332
rect 29641 19323 29699 19329
rect 29730 19320 29736 19332
rect 29788 19320 29794 19372
rect 31680 19292 31708 19391
rect 35434 19320 35440 19372
rect 35492 19360 35498 19372
rect 35529 19363 35587 19369
rect 35529 19360 35541 19363
rect 35492 19332 35541 19360
rect 35492 19320 35498 19332
rect 35529 19329 35541 19332
rect 35575 19329 35587 19363
rect 38654 19360 38660 19372
rect 38615 19332 38660 19360
rect 35529 19323 35587 19329
rect 38654 19320 38660 19332
rect 38712 19320 38718 19372
rect 40218 19320 40224 19372
rect 40276 19360 40282 19372
rect 41141 19363 41199 19369
rect 41141 19360 41153 19363
rect 40276 19332 41153 19360
rect 40276 19320 40282 19332
rect 41141 19329 41153 19332
rect 41187 19360 41199 19363
rect 43732 19360 43760 19456
rect 43993 19363 44051 19369
rect 43993 19360 44005 19363
rect 41187 19332 41644 19360
rect 43732 19332 44005 19360
rect 41187 19329 41199 19332
rect 41141 19323 41199 19329
rect 32125 19295 32183 19301
rect 31680 19264 32076 19292
rect 29089 19227 29147 19233
rect 29089 19193 29101 19227
rect 29135 19224 29147 19227
rect 29978 19227 30036 19233
rect 29978 19224 29990 19227
rect 29135 19196 29990 19224
rect 29135 19193 29147 19196
rect 29089 19187 29147 19193
rect 29978 19193 29990 19196
rect 30024 19224 30036 19227
rect 30190 19224 30196 19236
rect 30024 19196 30196 19224
rect 30024 19193 30036 19196
rect 29978 19187 30036 19193
rect 30190 19184 30196 19196
rect 30248 19184 30254 19236
rect 32048 19224 32076 19264
rect 32125 19261 32137 19295
rect 32171 19292 32183 19295
rect 32214 19292 32220 19304
rect 32171 19264 32220 19292
rect 32171 19261 32183 19264
rect 32125 19255 32183 19261
rect 32214 19252 32220 19264
rect 32272 19292 32278 19304
rect 34333 19295 34391 19301
rect 34333 19292 34345 19295
rect 32272 19264 34345 19292
rect 32272 19252 32278 19264
rect 34333 19261 34345 19264
rect 34379 19292 34391 19295
rect 34422 19292 34428 19304
rect 34379 19264 34428 19292
rect 34379 19261 34391 19264
rect 34333 19255 34391 19261
rect 34422 19252 34428 19264
rect 34480 19252 34486 19304
rect 34698 19292 34704 19304
rect 34659 19264 34704 19292
rect 34698 19252 34704 19264
rect 34756 19252 34762 19304
rect 34790 19252 34796 19304
rect 34848 19292 34854 19304
rect 35069 19295 35127 19301
rect 35069 19292 35081 19295
rect 34848 19264 35081 19292
rect 34848 19252 34854 19264
rect 35069 19261 35081 19264
rect 35115 19261 35127 19295
rect 35069 19255 35127 19261
rect 35342 19252 35348 19304
rect 35400 19292 35406 19304
rect 35805 19295 35863 19301
rect 35805 19292 35817 19295
rect 35400 19264 35817 19292
rect 35400 19252 35406 19264
rect 35805 19261 35817 19264
rect 35851 19261 35863 19295
rect 35805 19255 35863 19261
rect 38087 19295 38145 19301
rect 38087 19261 38099 19295
rect 38133 19292 38145 19295
rect 38562 19292 38568 19304
rect 38133 19264 38568 19292
rect 38133 19261 38145 19264
rect 38087 19255 38145 19261
rect 38562 19252 38568 19264
rect 38620 19252 38626 19304
rect 41509 19295 41567 19301
rect 41509 19292 41521 19295
rect 40972 19264 41521 19292
rect 32462 19227 32520 19233
rect 32462 19224 32474 19227
rect 32048 19196 32474 19224
rect 32462 19193 32474 19196
rect 32508 19193 32520 19227
rect 32462 19187 32520 19193
rect 33594 19156 33600 19168
rect 33555 19128 33600 19156
rect 33594 19116 33600 19128
rect 33652 19116 33658 19168
rect 34716 19156 34744 19252
rect 40972 19236 41000 19264
rect 41509 19261 41521 19264
rect 41555 19261 41567 19295
rect 41616 19292 41644 19332
rect 43993 19329 44005 19332
rect 44039 19329 44051 19363
rect 44174 19360 44180 19372
rect 44135 19332 44180 19360
rect 43993 19323 44051 19329
rect 44174 19320 44180 19332
rect 44232 19360 44238 19372
rect 45002 19360 45008 19372
rect 44232 19332 45008 19360
rect 44232 19320 44238 19332
rect 45002 19320 45008 19332
rect 45060 19360 45066 19372
rect 45097 19363 45155 19369
rect 45097 19360 45109 19363
rect 45060 19332 45109 19360
rect 45060 19320 45066 19332
rect 45097 19329 45109 19332
rect 45143 19329 45155 19363
rect 45097 19323 45155 19329
rect 41877 19295 41935 19301
rect 41877 19292 41889 19295
rect 41616 19264 41889 19292
rect 41509 19255 41567 19261
rect 41877 19261 41889 19264
rect 41923 19261 41935 19295
rect 41877 19255 41935 19261
rect 43607 19295 43665 19301
rect 43607 19261 43619 19295
rect 43653 19292 43665 19295
rect 44082 19292 44088 19304
rect 43653 19264 44088 19292
rect 43653 19261 43665 19264
rect 43607 19255 43665 19261
rect 44082 19252 44088 19264
rect 44140 19252 44146 19304
rect 37182 19184 37188 19236
rect 37240 19224 37246 19236
rect 38381 19227 38439 19233
rect 38381 19224 38393 19227
rect 37240 19196 38393 19224
rect 37240 19184 37246 19196
rect 38381 19193 38393 19196
rect 38427 19224 38439 19227
rect 39025 19227 39083 19233
rect 39025 19224 39037 19227
rect 38427 19196 39037 19224
rect 38427 19193 38439 19196
rect 38381 19187 38439 19193
rect 39025 19193 39037 19196
rect 39071 19193 39083 19227
rect 39025 19187 39083 19193
rect 39945 19227 40003 19233
rect 39945 19193 39957 19227
rect 39991 19224 40003 19227
rect 40865 19227 40923 19233
rect 39991 19196 40816 19224
rect 39991 19193 40003 19196
rect 39945 19187 40003 19193
rect 35531 19159 35589 19165
rect 35531 19156 35543 19159
rect 34716 19128 35543 19156
rect 35531 19125 35543 19128
rect 35577 19156 35589 19159
rect 35618 19156 35624 19168
rect 35577 19128 35624 19156
rect 35577 19125 35589 19128
rect 35531 19119 35589 19125
rect 35618 19116 35624 19128
rect 35676 19116 35682 19168
rect 36906 19156 36912 19168
rect 36867 19128 36912 19156
rect 36906 19116 36912 19128
rect 36964 19116 36970 19168
rect 37826 19116 37832 19168
rect 37884 19156 37890 19168
rect 38565 19159 38623 19165
rect 38565 19156 38577 19159
rect 37884 19128 38577 19156
rect 37884 19116 37890 19128
rect 38565 19125 38577 19128
rect 38611 19125 38623 19159
rect 38565 19119 38623 19125
rect 39114 19116 39120 19168
rect 39172 19156 39178 19168
rect 39393 19159 39451 19165
rect 39393 19156 39405 19159
rect 39172 19128 39405 19156
rect 39172 19116 39178 19128
rect 39393 19125 39405 19128
rect 39439 19125 39451 19159
rect 39393 19119 39451 19125
rect 40313 19159 40371 19165
rect 40313 19125 40325 19159
rect 40359 19156 40371 19159
rect 40402 19156 40408 19168
rect 40359 19128 40408 19156
rect 40359 19125 40371 19128
rect 40313 19119 40371 19125
rect 40402 19116 40408 19128
rect 40460 19116 40466 19168
rect 40788 19156 40816 19196
rect 40865 19193 40877 19227
rect 40911 19224 40923 19227
rect 40954 19224 40960 19236
rect 40911 19196 40960 19224
rect 40911 19193 40923 19196
rect 40865 19187 40923 19193
rect 40954 19184 40960 19196
rect 41012 19184 41018 19236
rect 41049 19227 41107 19233
rect 41049 19193 41061 19227
rect 41095 19224 41107 19227
rect 42150 19224 42156 19236
rect 41095 19196 42156 19224
rect 41095 19193 41107 19196
rect 41049 19187 41107 19193
rect 41064 19156 41092 19187
rect 42150 19184 42156 19196
rect 42208 19184 42214 19236
rect 40788 19128 41092 19156
rect 43073 19159 43131 19165
rect 43073 19125 43085 19159
rect 43119 19156 43131 19159
rect 43438 19156 43444 19168
rect 43119 19128 43444 19156
rect 43119 19125 43131 19128
rect 43073 19119 43131 19125
rect 43438 19116 43444 19128
rect 43496 19156 43502 19168
rect 44085 19159 44143 19165
rect 44085 19156 44097 19159
rect 43496 19128 44097 19156
rect 43496 19116 43502 19128
rect 44085 19125 44097 19128
rect 44131 19125 44143 19159
rect 44085 19119 44143 19125
rect 44726 19116 44732 19168
rect 44784 19156 44790 19168
rect 44821 19159 44879 19165
rect 44821 19156 44833 19159
rect 44784 19128 44833 19156
rect 44784 19116 44790 19128
rect 44821 19125 44833 19128
rect 44867 19156 44879 19159
rect 46106 19156 46112 19168
rect 44867 19128 46112 19156
rect 44867 19125 44879 19128
rect 44821 19119 44879 19125
rect 46106 19116 46112 19128
rect 46164 19116 46170 19168
rect 1104 19066 48852 19088
rect 1104 19014 19606 19066
rect 19658 19014 19670 19066
rect 19722 19014 19734 19066
rect 19786 19014 19798 19066
rect 19850 19014 48852 19066
rect 1104 18992 48852 19014
rect 34606 18952 34612 18964
rect 34567 18924 34612 18952
rect 34606 18912 34612 18924
rect 34664 18912 34670 18964
rect 38654 18912 38660 18964
rect 38712 18952 38718 18964
rect 38749 18955 38807 18961
rect 38749 18952 38761 18955
rect 38712 18924 38761 18952
rect 38712 18912 38718 18924
rect 38749 18921 38761 18924
rect 38795 18921 38807 18955
rect 40218 18952 40224 18964
rect 40179 18924 40224 18952
rect 38749 18915 38807 18921
rect 40218 18912 40224 18924
rect 40276 18912 40282 18964
rect 40770 18912 40776 18964
rect 40828 18952 40834 18964
rect 42150 18952 42156 18964
rect 40828 18924 40873 18952
rect 42111 18924 42156 18952
rect 40828 18912 40834 18924
rect 42150 18912 42156 18924
rect 42208 18912 42214 18964
rect 45002 18952 45008 18964
rect 44963 18924 45008 18952
rect 45002 18912 45008 18924
rect 45060 18912 45066 18964
rect 29362 18844 29368 18896
rect 29420 18884 29426 18896
rect 30101 18887 30159 18893
rect 30101 18884 30113 18887
rect 29420 18856 30113 18884
rect 29420 18844 29426 18856
rect 30101 18853 30113 18856
rect 30147 18853 30159 18887
rect 30101 18847 30159 18853
rect 30190 18844 30196 18896
rect 30248 18884 30254 18896
rect 30248 18856 30293 18884
rect 30248 18844 30254 18856
rect 34514 18844 34520 18896
rect 34572 18884 34578 18896
rect 34885 18887 34943 18893
rect 34885 18884 34897 18887
rect 34572 18856 34897 18884
rect 34572 18844 34578 18856
rect 34885 18853 34897 18856
rect 34931 18884 34943 18887
rect 35342 18884 35348 18896
rect 34931 18856 35348 18884
rect 34931 18853 34943 18856
rect 34885 18847 34943 18853
rect 35342 18844 35348 18856
rect 35400 18884 35406 18896
rect 35437 18887 35495 18893
rect 35437 18884 35449 18887
rect 35400 18856 35449 18884
rect 35400 18844 35406 18856
rect 35437 18853 35449 18856
rect 35483 18853 35495 18887
rect 35618 18884 35624 18896
rect 35579 18856 35624 18884
rect 35437 18847 35495 18853
rect 35618 18844 35624 18856
rect 35676 18844 35682 18896
rect 35713 18887 35771 18893
rect 35713 18853 35725 18887
rect 35759 18884 35771 18887
rect 36078 18884 36084 18896
rect 35759 18856 36084 18884
rect 35759 18853 35771 18856
rect 35713 18847 35771 18853
rect 36078 18844 36084 18856
rect 36136 18844 36142 18896
rect 36906 18844 36912 18896
rect 36964 18884 36970 18896
rect 38289 18887 38347 18893
rect 38289 18884 38301 18887
rect 36964 18856 38301 18884
rect 36964 18844 36970 18856
rect 38289 18853 38301 18856
rect 38335 18853 38347 18887
rect 38289 18847 38347 18853
rect 29914 18816 29920 18828
rect 29875 18788 29920 18816
rect 29914 18776 29920 18788
rect 29972 18776 29978 18828
rect 38102 18816 38108 18828
rect 38063 18788 38108 18816
rect 38102 18776 38108 18788
rect 38160 18776 38166 18828
rect 40218 18776 40224 18828
rect 40276 18816 40282 18828
rect 41049 18819 41107 18825
rect 41049 18816 41061 18819
rect 40276 18788 41061 18816
rect 40276 18776 40282 18788
rect 41049 18785 41061 18788
rect 41095 18785 41107 18819
rect 41049 18779 41107 18785
rect 43892 18819 43950 18825
rect 43892 18785 43904 18819
rect 43938 18816 43950 18819
rect 44358 18816 44364 18828
rect 43938 18788 44364 18816
rect 43938 18785 43950 18788
rect 43892 18779 43950 18785
rect 44358 18776 44364 18788
rect 44416 18776 44422 18828
rect 45554 18776 45560 18828
rect 45612 18816 45618 18828
rect 46365 18819 46423 18825
rect 46365 18816 46377 18819
rect 45612 18788 46377 18816
rect 45612 18776 45618 18788
rect 46365 18785 46377 18788
rect 46411 18816 46423 18819
rect 46934 18816 46940 18828
rect 46411 18788 46940 18816
rect 46411 18785 46423 18788
rect 46365 18779 46423 18785
rect 46934 18776 46940 18788
rect 46992 18776 46998 18828
rect 34057 18751 34115 18757
rect 34057 18717 34069 18751
rect 34103 18748 34115 18751
rect 34514 18748 34520 18760
rect 34103 18720 34520 18748
rect 34103 18717 34115 18720
rect 34057 18711 34115 18717
rect 34514 18708 34520 18720
rect 34572 18708 34578 18760
rect 38378 18748 38384 18760
rect 38339 18720 38384 18748
rect 38378 18708 38384 18720
rect 38436 18708 38442 18760
rect 39942 18708 39948 18760
rect 40000 18748 40006 18760
rect 40313 18751 40371 18757
rect 40313 18748 40325 18751
rect 40000 18720 40325 18748
rect 40000 18708 40006 18720
rect 40313 18717 40325 18720
rect 40359 18748 40371 18751
rect 40678 18748 40684 18760
rect 40359 18720 40684 18748
rect 40359 18717 40371 18720
rect 40313 18711 40371 18717
rect 40678 18708 40684 18720
rect 40736 18708 40742 18760
rect 40773 18751 40831 18757
rect 40773 18717 40785 18751
rect 40819 18748 40831 18751
rect 40954 18748 40960 18760
rect 40819 18720 40960 18748
rect 40819 18717 40831 18720
rect 40773 18711 40831 18717
rect 40954 18708 40960 18720
rect 41012 18708 41018 18760
rect 43622 18748 43628 18760
rect 42996 18720 43628 18748
rect 29641 18683 29699 18689
rect 29641 18649 29653 18683
rect 29687 18680 29699 18683
rect 30282 18680 30288 18692
rect 29687 18652 30288 18680
rect 29687 18649 29699 18652
rect 29641 18643 29699 18649
rect 30282 18640 30288 18652
rect 30340 18640 30346 18692
rect 37553 18683 37611 18689
rect 37553 18649 37565 18683
rect 37599 18680 37611 18683
rect 37826 18680 37832 18692
rect 37599 18652 37832 18680
rect 37599 18649 37611 18652
rect 37553 18643 37611 18649
rect 37826 18640 37832 18652
rect 37884 18640 37890 18692
rect 42996 18680 43024 18720
rect 43622 18708 43628 18720
rect 43680 18708 43686 18760
rect 46106 18748 46112 18760
rect 46067 18720 46112 18748
rect 46106 18708 46112 18720
rect 46164 18708 46170 18760
rect 42720 18652 43024 18680
rect 29457 18615 29515 18621
rect 29457 18581 29469 18615
rect 29503 18612 29515 18615
rect 30098 18612 30104 18624
rect 29503 18584 30104 18612
rect 29503 18581 29515 18584
rect 29457 18575 29515 18581
rect 30098 18572 30104 18584
rect 30156 18572 30162 18624
rect 31754 18572 31760 18624
rect 31812 18612 31818 18624
rect 32122 18612 32128 18624
rect 31812 18584 32128 18612
rect 31812 18572 31818 18584
rect 32122 18572 32128 18584
rect 32180 18612 32186 18624
rect 32309 18615 32367 18621
rect 32309 18612 32321 18615
rect 32180 18584 32321 18612
rect 32180 18572 32186 18584
rect 32309 18581 32321 18584
rect 32355 18581 32367 18615
rect 32309 18575 32367 18581
rect 35161 18615 35219 18621
rect 35161 18581 35173 18615
rect 35207 18612 35219 18615
rect 35250 18612 35256 18624
rect 35207 18584 35256 18612
rect 35207 18581 35219 18584
rect 35161 18575 35219 18581
rect 35250 18572 35256 18584
rect 35308 18572 35314 18624
rect 40494 18572 40500 18624
rect 40552 18612 40558 18624
rect 42720 18612 42748 18652
rect 42886 18612 42892 18624
rect 40552 18584 42748 18612
rect 42847 18584 42892 18612
rect 40552 18572 40558 18584
rect 42886 18572 42892 18584
rect 42944 18572 42950 18624
rect 47486 18612 47492 18624
rect 47447 18584 47492 18612
rect 47486 18572 47492 18584
rect 47544 18572 47550 18624
rect 1104 18522 48852 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 34966 18522
rect 35018 18470 35030 18522
rect 35082 18470 35094 18522
rect 35146 18470 35158 18522
rect 35210 18470 48852 18522
rect 1104 18448 48852 18470
rect 29089 18411 29147 18417
rect 29089 18377 29101 18411
rect 29135 18408 29147 18411
rect 29914 18408 29920 18420
rect 29135 18380 29920 18408
rect 29135 18377 29147 18380
rect 29089 18371 29147 18377
rect 29914 18368 29920 18380
rect 29972 18368 29978 18420
rect 34701 18411 34759 18417
rect 34701 18377 34713 18411
rect 34747 18408 34759 18411
rect 35618 18408 35624 18420
rect 34747 18380 35624 18408
rect 34747 18377 34759 18380
rect 34701 18371 34759 18377
rect 35618 18368 35624 18380
rect 35676 18368 35682 18420
rect 36906 18368 36912 18420
rect 36964 18408 36970 18420
rect 37737 18411 37795 18417
rect 37737 18408 37749 18411
rect 36964 18380 37749 18408
rect 36964 18368 36970 18380
rect 37737 18377 37749 18380
rect 37783 18377 37795 18411
rect 37737 18371 37795 18377
rect 35161 18343 35219 18349
rect 35161 18309 35173 18343
rect 35207 18340 35219 18343
rect 35342 18340 35348 18352
rect 35207 18312 35348 18340
rect 35207 18309 35219 18312
rect 35161 18303 35219 18309
rect 35342 18300 35348 18312
rect 35400 18300 35406 18352
rect 37752 18340 37780 18371
rect 37826 18368 37832 18420
rect 37884 18408 37890 18420
rect 38102 18408 38108 18420
rect 37884 18380 38108 18408
rect 37884 18368 37890 18380
rect 38102 18368 38108 18380
rect 38160 18368 38166 18420
rect 39942 18408 39948 18420
rect 39903 18380 39948 18408
rect 39942 18368 39948 18380
rect 40000 18368 40006 18420
rect 40770 18408 40776 18420
rect 40731 18380 40776 18408
rect 40770 18368 40776 18380
rect 40828 18368 40834 18420
rect 41966 18408 41972 18420
rect 41927 18380 41972 18408
rect 41966 18368 41972 18380
rect 42024 18368 42030 18420
rect 43622 18368 43628 18420
rect 43680 18408 43686 18420
rect 43901 18411 43959 18417
rect 43901 18408 43913 18411
rect 43680 18380 43913 18408
rect 43680 18368 43686 18380
rect 43901 18377 43913 18380
rect 43947 18377 43959 18411
rect 43901 18371 43959 18377
rect 43990 18368 43996 18420
rect 44048 18408 44054 18420
rect 44358 18408 44364 18420
rect 44048 18380 44364 18408
rect 44048 18368 44054 18380
rect 44358 18368 44364 18380
rect 44416 18368 44422 18420
rect 45554 18408 45560 18420
rect 45515 18380 45560 18408
rect 45554 18368 45560 18380
rect 45612 18368 45618 18420
rect 45925 18411 45983 18417
rect 45925 18377 45937 18411
rect 45971 18408 45983 18411
rect 46106 18408 46112 18420
rect 45971 18380 46112 18408
rect 45971 18377 45983 18380
rect 45925 18371 45983 18377
rect 46106 18368 46112 18380
rect 46164 18368 46170 18420
rect 40218 18340 40224 18352
rect 37752 18312 40224 18340
rect 40218 18300 40224 18312
rect 40276 18300 40282 18352
rect 42981 18343 43039 18349
rect 42981 18309 42993 18343
rect 43027 18340 43039 18343
rect 43027 18312 44036 18340
rect 43027 18309 43039 18312
rect 42981 18303 43039 18309
rect 34422 18232 34428 18284
rect 34480 18272 34486 18284
rect 35529 18275 35587 18281
rect 35529 18272 35541 18275
rect 34480 18244 35541 18272
rect 34480 18232 34486 18244
rect 35529 18241 35541 18244
rect 35575 18272 35587 18275
rect 35713 18275 35771 18281
rect 35713 18272 35725 18275
rect 35575 18244 35725 18272
rect 35575 18241 35587 18244
rect 35529 18235 35587 18241
rect 35713 18241 35725 18244
rect 35759 18241 35771 18275
rect 35713 18235 35771 18241
rect 42886 18232 42892 18284
rect 42944 18272 42950 18284
rect 43533 18275 43591 18281
rect 43533 18272 43545 18275
rect 42944 18244 43545 18272
rect 42944 18232 42950 18244
rect 43533 18241 43545 18244
rect 43579 18241 43591 18275
rect 43533 18235 43591 18241
rect 29549 18207 29607 18213
rect 29549 18173 29561 18207
rect 29595 18204 29607 18207
rect 29641 18207 29699 18213
rect 29641 18204 29653 18207
rect 29595 18176 29653 18204
rect 29595 18173 29607 18176
rect 29549 18167 29607 18173
rect 29641 18173 29653 18176
rect 29687 18204 29699 18207
rect 29730 18204 29736 18216
rect 29687 18176 29736 18204
rect 29687 18173 29699 18176
rect 29641 18167 29699 18173
rect 29730 18164 29736 18176
rect 29788 18164 29794 18216
rect 34790 18164 34796 18216
rect 34848 18204 34854 18216
rect 35342 18204 35348 18216
rect 34848 18176 35348 18204
rect 34848 18164 34854 18176
rect 35342 18164 35348 18176
rect 35400 18164 35406 18216
rect 35802 18164 35808 18216
rect 35860 18204 35866 18216
rect 35986 18213 35992 18216
rect 35969 18207 35992 18213
rect 35969 18204 35981 18207
rect 35860 18176 35981 18204
rect 35860 18164 35866 18176
rect 35969 18173 35981 18176
rect 36044 18204 36050 18216
rect 41785 18207 41843 18213
rect 36044 18176 36117 18204
rect 35969 18167 35992 18173
rect 35986 18164 35992 18167
rect 36044 18164 36050 18176
rect 41785 18173 41797 18207
rect 41831 18204 41843 18207
rect 44008 18204 44036 18312
rect 44082 18300 44088 18352
rect 44140 18340 44146 18352
rect 44637 18343 44695 18349
rect 44637 18340 44649 18343
rect 44140 18312 44649 18340
rect 44140 18300 44146 18312
rect 44637 18309 44649 18312
rect 44683 18309 44695 18343
rect 44637 18303 44695 18309
rect 46124 18281 46152 18368
rect 46109 18275 46167 18281
rect 46109 18241 46121 18275
rect 46155 18241 46167 18275
rect 46109 18235 46167 18241
rect 44453 18207 44511 18213
rect 44453 18204 44465 18207
rect 41831 18176 42472 18204
rect 44008 18176 44465 18204
rect 41831 18173 41843 18176
rect 41785 18167 41843 18173
rect 29908 18139 29966 18145
rect 29908 18105 29920 18139
rect 29954 18136 29966 18139
rect 30098 18136 30104 18148
rect 29954 18108 30104 18136
rect 29954 18105 29966 18108
rect 29908 18099 29966 18105
rect 30098 18096 30104 18108
rect 30156 18096 30162 18148
rect 42444 18145 42472 18176
rect 44453 18173 44465 18176
rect 44499 18204 44511 18207
rect 45005 18207 45063 18213
rect 45005 18204 45017 18207
rect 44499 18176 45017 18204
rect 44499 18173 44511 18176
rect 44453 18167 44511 18173
rect 45005 18173 45017 18176
rect 45051 18173 45063 18207
rect 45005 18167 45063 18173
rect 42429 18139 42487 18145
rect 42429 18105 42441 18139
rect 42475 18136 42487 18139
rect 43254 18136 43260 18148
rect 42475 18108 43260 18136
rect 42475 18105 42487 18108
rect 42429 18099 42487 18105
rect 43254 18096 43260 18108
rect 43312 18096 43318 18148
rect 46382 18145 46388 18148
rect 46376 18136 46388 18145
rect 46343 18108 46388 18136
rect 46376 18099 46388 18108
rect 46382 18096 46388 18099
rect 46440 18096 46446 18148
rect 28721 18071 28779 18077
rect 28721 18037 28733 18071
rect 28767 18068 28779 18071
rect 29362 18068 29368 18080
rect 28767 18040 29368 18068
rect 28767 18037 28779 18040
rect 28721 18031 28779 18037
rect 29362 18028 29368 18040
rect 29420 18028 29426 18080
rect 30190 18028 30196 18080
rect 30248 18068 30254 18080
rect 31021 18071 31079 18077
rect 31021 18068 31033 18071
rect 30248 18040 31033 18068
rect 30248 18028 30254 18040
rect 31021 18037 31033 18040
rect 31067 18037 31079 18071
rect 31021 18031 31079 18037
rect 34333 18071 34391 18077
rect 34333 18037 34345 18071
rect 34379 18068 34391 18071
rect 35802 18068 35808 18080
rect 34379 18040 35808 18068
rect 34379 18037 34391 18040
rect 34333 18031 34391 18037
rect 35802 18028 35808 18040
rect 35860 18028 35866 18080
rect 37093 18071 37151 18077
rect 37093 18037 37105 18071
rect 37139 18068 37151 18071
rect 37182 18068 37188 18080
rect 37139 18040 37188 18068
rect 37139 18037 37151 18040
rect 37093 18031 37151 18037
rect 37182 18028 37188 18040
rect 37240 18028 37246 18080
rect 38378 18028 38384 18080
rect 38436 18068 38442 18080
rect 38565 18071 38623 18077
rect 38565 18068 38577 18071
rect 38436 18040 38577 18068
rect 38436 18028 38442 18040
rect 38565 18037 38577 18040
rect 38611 18068 38623 18071
rect 39114 18068 39120 18080
rect 38611 18040 39120 18068
rect 38611 18037 38623 18040
rect 38565 18031 38623 18037
rect 39114 18028 39120 18040
rect 39172 18028 39178 18080
rect 41046 18068 41052 18080
rect 41007 18040 41052 18068
rect 41046 18028 41052 18040
rect 41104 18028 41110 18080
rect 42797 18071 42855 18077
rect 42797 18037 42809 18071
rect 42843 18068 42855 18071
rect 42978 18068 42984 18080
rect 42843 18040 42984 18068
rect 42843 18037 42855 18040
rect 42797 18031 42855 18037
rect 42978 18028 42984 18040
rect 43036 18068 43042 18080
rect 43441 18071 43499 18077
rect 43441 18068 43453 18071
rect 43036 18040 43453 18068
rect 43036 18028 43042 18040
rect 43441 18037 43453 18040
rect 43487 18037 43499 18071
rect 43441 18031 43499 18037
rect 46934 18028 46940 18080
rect 46992 18068 46998 18080
rect 47489 18071 47547 18077
rect 47489 18068 47501 18071
rect 46992 18040 47501 18068
rect 46992 18028 46998 18040
rect 47489 18037 47501 18040
rect 47535 18037 47547 18071
rect 47489 18031 47547 18037
rect 1104 17978 48852 18000
rect 1104 17926 19606 17978
rect 19658 17926 19670 17978
rect 19722 17926 19734 17978
rect 19786 17926 19798 17978
rect 19850 17926 48852 17978
rect 1104 17904 48852 17926
rect 29273 17867 29331 17873
rect 29273 17833 29285 17867
rect 29319 17864 29331 17867
rect 33597 17867 33655 17873
rect 33597 17864 33609 17867
rect 29319 17836 30604 17864
rect 29319 17833 29331 17836
rect 29273 17827 29331 17833
rect 30576 17808 30604 17836
rect 30852 17836 33609 17864
rect 29733 17799 29791 17805
rect 29733 17765 29745 17799
rect 29779 17796 29791 17799
rect 30190 17796 30196 17808
rect 29779 17768 30196 17796
rect 29779 17765 29791 17768
rect 29733 17759 29791 17765
rect 30190 17756 30196 17768
rect 30248 17756 30254 17808
rect 30558 17796 30564 17808
rect 30471 17768 30564 17796
rect 30558 17756 30564 17768
rect 30616 17756 30622 17808
rect 30742 17796 30748 17808
rect 30703 17768 30748 17796
rect 30742 17756 30748 17768
rect 30800 17756 30806 17808
rect 30852 17805 30880 17836
rect 33597 17833 33609 17836
rect 33643 17833 33655 17867
rect 35986 17864 35992 17876
rect 35947 17836 35992 17864
rect 33597 17827 33655 17833
rect 35986 17824 35992 17836
rect 36044 17824 36050 17876
rect 41138 17864 41144 17876
rect 41099 17836 41144 17864
rect 41138 17824 41144 17836
rect 41196 17824 41202 17876
rect 43901 17867 43959 17873
rect 43901 17833 43913 17867
rect 43947 17864 43959 17867
rect 44082 17864 44088 17876
rect 43947 17836 44088 17864
rect 43947 17833 43959 17836
rect 43901 17827 43959 17833
rect 44082 17824 44088 17836
rect 44140 17824 44146 17876
rect 46106 17824 46112 17876
rect 46164 17864 46170 17876
rect 46201 17867 46259 17873
rect 46201 17864 46213 17867
rect 46164 17836 46213 17864
rect 46164 17824 46170 17836
rect 46201 17833 46213 17836
rect 46247 17833 46259 17867
rect 46201 17827 46259 17833
rect 30837 17799 30895 17805
rect 30837 17765 30849 17799
rect 30883 17765 30895 17799
rect 30837 17759 30895 17765
rect 29086 17728 29092 17740
rect 29047 17700 29092 17728
rect 29086 17688 29092 17700
rect 29144 17688 29150 17740
rect 30098 17728 30104 17740
rect 30011 17700 30104 17728
rect 30098 17688 30104 17700
rect 30156 17728 30162 17740
rect 30852 17728 30880 17759
rect 34698 17756 34704 17808
rect 34756 17796 34762 17808
rect 35250 17796 35256 17808
rect 34756 17768 35256 17796
rect 34756 17756 34762 17768
rect 35250 17756 35256 17768
rect 35308 17796 35314 17808
rect 35437 17799 35495 17805
rect 35437 17796 35449 17799
rect 35308 17768 35449 17796
rect 35308 17756 35314 17768
rect 35437 17765 35449 17768
rect 35483 17765 35495 17799
rect 35437 17759 35495 17765
rect 43162 17756 43168 17808
rect 43220 17796 43226 17808
rect 43990 17796 43996 17808
rect 43220 17768 43996 17796
rect 43220 17756 43226 17768
rect 43990 17756 43996 17768
rect 44048 17756 44054 17808
rect 45738 17796 45744 17808
rect 45699 17768 45744 17796
rect 45738 17756 45744 17768
rect 45796 17756 45802 17808
rect 46750 17796 46756 17808
rect 46711 17768 46756 17796
rect 46750 17756 46756 17768
rect 46808 17756 46814 17808
rect 46934 17796 46940 17808
rect 46895 17768 46940 17796
rect 46934 17756 46940 17768
rect 46992 17796 46998 17808
rect 47397 17799 47455 17805
rect 47397 17796 47409 17799
rect 46992 17768 47409 17796
rect 46992 17756 46998 17768
rect 47397 17765 47409 17768
rect 47443 17765 47455 17799
rect 47397 17759 47455 17765
rect 32214 17728 32220 17740
rect 30156 17700 30880 17728
rect 32175 17700 32220 17728
rect 30156 17688 30162 17700
rect 32214 17688 32220 17700
rect 32272 17688 32278 17740
rect 32306 17688 32312 17740
rect 32364 17728 32370 17740
rect 32473 17731 32531 17737
rect 32473 17728 32485 17731
rect 32364 17700 32485 17728
rect 32364 17688 32370 17700
rect 32473 17697 32485 17700
rect 32519 17697 32531 17731
rect 32473 17691 32531 17697
rect 40957 17731 41015 17737
rect 40957 17697 40969 17731
rect 41003 17697 41015 17731
rect 42058 17728 42064 17740
rect 42019 17700 42064 17728
rect 40957 17691 41015 17697
rect 34514 17620 34520 17672
rect 34572 17660 34578 17672
rect 35250 17660 35256 17672
rect 34572 17632 35256 17660
rect 34572 17620 34578 17632
rect 35250 17620 35256 17632
rect 35308 17660 35314 17672
rect 35345 17663 35403 17669
rect 35345 17660 35357 17663
rect 35308 17632 35357 17660
rect 35308 17620 35314 17632
rect 35345 17629 35357 17632
rect 35391 17629 35403 17663
rect 35526 17660 35532 17672
rect 35487 17632 35532 17660
rect 35345 17623 35403 17629
rect 35526 17620 35532 17632
rect 35584 17620 35590 17672
rect 40972 17660 41000 17691
rect 42058 17688 42064 17700
rect 42116 17688 42122 17740
rect 43714 17728 43720 17740
rect 43675 17700 43720 17728
rect 43714 17688 43720 17700
rect 43772 17688 43778 17740
rect 45554 17728 45560 17740
rect 45515 17700 45560 17728
rect 45554 17688 45560 17700
rect 45612 17728 45618 17740
rect 46382 17728 46388 17740
rect 45612 17700 46388 17728
rect 45612 17688 45618 17700
rect 46382 17688 46388 17700
rect 46440 17728 46446 17740
rect 46569 17731 46627 17737
rect 46569 17728 46581 17731
rect 46440 17700 46581 17728
rect 46440 17688 46446 17700
rect 46569 17697 46581 17700
rect 46615 17697 46627 17731
rect 46569 17691 46627 17697
rect 42610 17660 42616 17672
rect 40972 17632 42616 17660
rect 42610 17620 42616 17632
rect 42668 17620 42674 17672
rect 45833 17663 45891 17669
rect 45833 17629 45845 17663
rect 45879 17660 45891 17663
rect 45879 17632 45913 17660
rect 45879 17629 45891 17632
rect 45833 17623 45891 17629
rect 29362 17552 29368 17604
rect 29420 17592 29426 17604
rect 30285 17595 30343 17601
rect 30285 17592 30297 17595
rect 29420 17564 30297 17592
rect 29420 17552 29426 17564
rect 30285 17561 30297 17564
rect 30331 17561 30343 17595
rect 30285 17555 30343 17561
rect 34977 17595 35035 17601
rect 34977 17561 34989 17595
rect 35023 17592 35035 17595
rect 35434 17592 35440 17604
rect 35023 17564 35440 17592
rect 35023 17561 35035 17564
rect 34977 17555 35035 17561
rect 35434 17552 35440 17564
rect 35492 17552 35498 17604
rect 43438 17592 43444 17604
rect 43399 17564 43444 17592
rect 43438 17552 43444 17564
rect 43496 17552 43502 17604
rect 45097 17595 45155 17601
rect 45097 17561 45109 17595
rect 45143 17592 45155 17595
rect 45848 17592 45876 17623
rect 46474 17592 46480 17604
rect 45143 17564 46480 17592
rect 45143 17561 45155 17564
rect 45097 17555 45155 17561
rect 46474 17552 46480 17564
rect 46532 17552 46538 17604
rect 31938 17524 31944 17536
rect 31899 17496 31944 17524
rect 31938 17484 31944 17496
rect 31996 17484 32002 17536
rect 41598 17524 41604 17536
rect 41559 17496 41604 17524
rect 41598 17484 41604 17496
rect 41656 17484 41662 17536
rect 42242 17524 42248 17536
rect 42203 17496 42248 17524
rect 42242 17484 42248 17496
rect 42300 17484 42306 17536
rect 42981 17527 43039 17533
rect 42981 17493 42993 17527
rect 43027 17524 43039 17527
rect 43254 17524 43260 17536
rect 43027 17496 43260 17524
rect 43027 17493 43039 17496
rect 42981 17487 43039 17493
rect 43254 17484 43260 17496
rect 43312 17484 43318 17536
rect 45278 17524 45284 17536
rect 45239 17496 45284 17524
rect 45278 17484 45284 17496
rect 45336 17484 45342 17536
rect 47118 17524 47124 17536
rect 47079 17496 47124 17524
rect 47118 17484 47124 17496
rect 47176 17484 47182 17536
rect 1104 17434 48852 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 34966 17434
rect 35018 17382 35030 17434
rect 35082 17382 35094 17434
rect 35146 17382 35158 17434
rect 35210 17382 48852 17434
rect 1104 17360 48852 17382
rect 30009 17323 30067 17329
rect 30009 17289 30021 17323
rect 30055 17320 30067 17323
rect 30285 17323 30343 17329
rect 30285 17320 30297 17323
rect 30055 17292 30297 17320
rect 30055 17289 30067 17292
rect 30009 17283 30067 17289
rect 30285 17289 30297 17292
rect 30331 17320 30343 17323
rect 30742 17320 30748 17332
rect 30331 17292 30748 17320
rect 30331 17289 30343 17292
rect 30285 17283 30343 17289
rect 30742 17280 30748 17292
rect 30800 17280 30806 17332
rect 31757 17323 31815 17329
rect 31757 17289 31769 17323
rect 31803 17320 31815 17323
rect 32214 17320 32220 17332
rect 31803 17292 32220 17320
rect 31803 17289 31815 17292
rect 31757 17283 31815 17289
rect 26510 17252 26516 17264
rect 26471 17224 26516 17252
rect 26510 17212 26516 17224
rect 26568 17212 26574 17264
rect 30558 17212 30564 17264
rect 30616 17252 30622 17264
rect 30653 17255 30711 17261
rect 30653 17252 30665 17255
rect 30616 17224 30665 17252
rect 30616 17212 30622 17224
rect 30653 17221 30665 17224
rect 30699 17221 30711 17255
rect 30653 17215 30711 17221
rect 31864 17196 31892 17292
rect 32214 17280 32220 17292
rect 32272 17280 32278 17332
rect 34698 17320 34704 17332
rect 34659 17292 34704 17320
rect 34698 17280 34704 17292
rect 34756 17280 34762 17332
rect 35161 17323 35219 17329
rect 35161 17289 35173 17323
rect 35207 17320 35219 17323
rect 35250 17320 35256 17332
rect 35207 17292 35256 17320
rect 35207 17289 35219 17292
rect 35161 17283 35219 17289
rect 35250 17280 35256 17292
rect 35308 17280 35314 17332
rect 41233 17323 41291 17329
rect 41233 17289 41245 17323
rect 41279 17320 41291 17323
rect 42058 17320 42064 17332
rect 41279 17292 42064 17320
rect 41279 17289 41291 17292
rect 41233 17283 41291 17289
rect 42058 17280 42064 17292
rect 42116 17320 42122 17332
rect 42153 17323 42211 17329
rect 42153 17320 42165 17323
rect 42116 17292 42165 17320
rect 42116 17280 42122 17292
rect 42153 17289 42165 17292
rect 42199 17289 42211 17323
rect 42610 17320 42616 17332
rect 42571 17292 42616 17320
rect 42153 17283 42211 17289
rect 42610 17280 42616 17292
rect 42668 17280 42674 17332
rect 42978 17320 42984 17332
rect 42939 17292 42984 17320
rect 42978 17280 42984 17292
rect 43036 17280 43042 17332
rect 43257 17323 43315 17329
rect 43257 17289 43269 17323
rect 43303 17320 43315 17323
rect 43714 17320 43720 17332
rect 43303 17292 43720 17320
rect 43303 17289 43315 17292
rect 43257 17283 43315 17289
rect 43714 17280 43720 17292
rect 43772 17280 43778 17332
rect 44082 17320 44088 17332
rect 44043 17292 44088 17320
rect 44082 17280 44088 17292
rect 44140 17280 44146 17332
rect 44821 17323 44879 17329
rect 44821 17289 44833 17323
rect 44867 17320 44879 17323
rect 45554 17320 45560 17332
rect 44867 17292 45560 17320
rect 44867 17289 44879 17292
rect 44821 17283 44879 17289
rect 45554 17280 45560 17292
rect 45612 17280 45618 17332
rect 45925 17323 45983 17329
rect 45925 17289 45937 17323
rect 45971 17320 45983 17323
rect 46106 17320 46112 17332
rect 45971 17292 46112 17320
rect 45971 17289 45983 17292
rect 45925 17283 45983 17289
rect 46106 17280 46112 17292
rect 46164 17280 46170 17332
rect 46382 17280 46388 17332
rect 46440 17320 46446 17332
rect 47489 17323 47547 17329
rect 47489 17320 47501 17323
rect 46440 17292 47501 17320
rect 46440 17280 46446 17292
rect 47489 17289 47501 17292
rect 47535 17289 47547 17323
rect 47489 17283 47547 17289
rect 35526 17252 35532 17264
rect 35487 17224 35532 17252
rect 35526 17212 35532 17224
rect 35584 17212 35590 17264
rect 31846 17184 31852 17196
rect 31759 17156 31852 17184
rect 31846 17144 31852 17156
rect 31904 17144 31910 17196
rect 41322 17144 41328 17196
rect 41380 17184 41386 17196
rect 41598 17184 41604 17196
rect 41380 17156 41604 17184
rect 41380 17144 41386 17156
rect 41598 17144 41604 17156
rect 41656 17144 41662 17196
rect 46124 17193 46152 17280
rect 46109 17187 46167 17193
rect 46109 17153 46121 17187
rect 46155 17153 46167 17187
rect 46109 17147 46167 17153
rect 23750 17116 23756 17128
rect 23711 17088 23756 17116
rect 23750 17076 23756 17088
rect 23808 17076 23814 17128
rect 26786 17116 26792 17128
rect 26699 17088 26792 17116
rect 26786 17076 26792 17088
rect 26844 17116 26850 17128
rect 27154 17116 27160 17128
rect 26844 17088 27160 17116
rect 26844 17076 26850 17088
rect 27154 17076 27160 17088
rect 27212 17076 27218 17128
rect 30101 17119 30159 17125
rect 30101 17085 30113 17119
rect 30147 17116 30159 17119
rect 30466 17116 30472 17128
rect 30147 17088 30472 17116
rect 30147 17085 30159 17088
rect 30101 17079 30159 17085
rect 30466 17076 30472 17088
rect 30524 17076 30530 17128
rect 31938 17076 31944 17128
rect 31996 17116 32002 17128
rect 32105 17119 32163 17125
rect 32105 17116 32117 17119
rect 31996 17088 32117 17116
rect 31996 17076 32002 17088
rect 32105 17085 32117 17088
rect 32151 17085 32163 17119
rect 32105 17079 32163 17085
rect 37185 17119 37243 17125
rect 37185 17085 37197 17119
rect 37231 17085 37243 17119
rect 37185 17079 37243 17085
rect 23474 17048 23480 17060
rect 23435 17020 23480 17048
rect 23474 17008 23480 17020
rect 23532 17048 23538 17060
rect 23998 17051 24056 17057
rect 23998 17048 24010 17051
rect 23532 17020 24010 17048
rect 23532 17008 23538 17020
rect 23998 17017 24010 17020
rect 24044 17017 24056 17051
rect 23998 17011 24056 17017
rect 25961 17051 26019 17057
rect 25961 17017 25973 17051
rect 26007 17048 26019 17051
rect 26804 17048 26832 17076
rect 26007 17020 26832 17048
rect 26007 17017 26019 17020
rect 25961 17011 26019 17017
rect 26878 17008 26884 17060
rect 26936 17048 26942 17060
rect 27065 17051 27123 17057
rect 27065 17048 27077 17051
rect 26936 17020 27077 17048
rect 26936 17008 26942 17020
rect 27065 17017 27077 17020
rect 27111 17017 27123 17051
rect 27065 17011 27123 17017
rect 31389 17051 31447 17057
rect 31389 17017 31401 17051
rect 31435 17048 31447 17051
rect 37093 17051 37151 17057
rect 31435 17020 32076 17048
rect 31435 17017 31447 17020
rect 31389 17011 31447 17017
rect 25133 16983 25191 16989
rect 25133 16949 25145 16983
rect 25179 16980 25191 16983
rect 25774 16980 25780 16992
rect 25179 16952 25780 16980
rect 25179 16949 25191 16952
rect 25133 16943 25191 16949
rect 25774 16940 25780 16952
rect 25832 16980 25838 16992
rect 26329 16983 26387 16989
rect 26329 16980 26341 16983
rect 25832 16952 26341 16980
rect 25832 16940 25838 16952
rect 26329 16949 26341 16952
rect 26375 16980 26387 16983
rect 26973 16983 27031 16989
rect 26973 16980 26985 16983
rect 26375 16952 26985 16980
rect 26375 16949 26387 16952
rect 26329 16943 26387 16949
rect 26973 16949 26985 16952
rect 27019 16949 27031 16983
rect 26973 16943 27031 16949
rect 29086 16940 29092 16992
rect 29144 16980 29150 16992
rect 29549 16983 29607 16989
rect 29549 16980 29561 16983
rect 29144 16952 29561 16980
rect 29144 16940 29150 16952
rect 29549 16949 29561 16952
rect 29595 16980 29607 16983
rect 30558 16980 30564 16992
rect 29595 16952 30564 16980
rect 29595 16949 29607 16952
rect 29549 16943 29607 16949
rect 30558 16940 30564 16952
rect 30616 16940 30622 16992
rect 32048 16980 32076 17020
rect 37093 17017 37105 17051
rect 37139 17048 37151 17051
rect 37200 17048 37228 17079
rect 37274 17076 37280 17128
rect 37332 17116 37338 17128
rect 37441 17119 37499 17125
rect 37441 17116 37453 17119
rect 37332 17088 37453 17116
rect 37332 17076 37338 17088
rect 37441 17085 37453 17088
rect 37487 17085 37499 17119
rect 37441 17079 37499 17085
rect 40313 17119 40371 17125
rect 40313 17085 40325 17119
rect 40359 17116 40371 17119
rect 41785 17119 41843 17125
rect 41785 17116 41797 17119
rect 40359 17088 41797 17116
rect 40359 17085 40371 17088
rect 40313 17079 40371 17085
rect 41785 17085 41797 17088
rect 41831 17116 41843 17119
rect 42702 17116 42708 17128
rect 41831 17088 42708 17116
rect 41831 17085 41843 17088
rect 41785 17079 41843 17085
rect 42702 17076 42708 17088
rect 42760 17076 42766 17128
rect 42978 17076 42984 17128
rect 43036 17116 43042 17128
rect 43073 17119 43131 17125
rect 43073 17116 43085 17119
rect 43036 17088 43085 17116
rect 43036 17076 43042 17088
rect 43073 17085 43085 17088
rect 43119 17085 43131 17119
rect 43073 17079 43131 17085
rect 44177 17119 44235 17125
rect 44177 17085 44189 17119
rect 44223 17116 44235 17119
rect 44542 17116 44548 17128
rect 44223 17088 44548 17116
rect 44223 17085 44235 17088
rect 44177 17079 44235 17085
rect 44542 17076 44548 17088
rect 44600 17076 44606 17128
rect 37734 17048 37740 17060
rect 37139 17020 37740 17048
rect 37139 17017 37151 17020
rect 37093 17011 37151 17017
rect 37734 17008 37740 17020
rect 37792 17008 37798 17060
rect 40034 17008 40040 17060
rect 40092 17048 40098 17060
rect 40957 17051 41015 17057
rect 40957 17048 40969 17051
rect 40092 17020 40969 17048
rect 40092 17008 40098 17020
rect 40957 17017 40969 17020
rect 41003 17048 41015 17051
rect 41693 17051 41751 17057
rect 41693 17048 41705 17051
rect 41003 17020 41705 17048
rect 41003 17017 41015 17020
rect 40957 17011 41015 17017
rect 41693 17017 41705 17020
rect 41739 17017 41751 17051
rect 41693 17011 41751 17017
rect 45189 17051 45247 17057
rect 45189 17017 45201 17051
rect 45235 17048 45247 17051
rect 45557 17051 45615 17057
rect 45557 17048 45569 17051
rect 45235 17020 45569 17048
rect 45235 17017 45247 17020
rect 45189 17011 45247 17017
rect 45557 17017 45569 17020
rect 45603 17048 45615 17051
rect 45738 17048 45744 17060
rect 45603 17020 45744 17048
rect 45603 17017 45615 17020
rect 45557 17011 45615 17017
rect 45738 17008 45744 17020
rect 45796 17048 45802 17060
rect 46376 17051 46434 17057
rect 46376 17048 46388 17051
rect 45796 17020 46388 17048
rect 45796 17008 45802 17020
rect 46376 17017 46388 17020
rect 46422 17048 46434 17051
rect 46566 17048 46572 17060
rect 46422 17020 46572 17048
rect 46422 17017 46434 17020
rect 46376 17011 46434 17017
rect 46566 17008 46572 17020
rect 46624 17008 46630 17060
rect 32306 16980 32312 16992
rect 32048 16952 32312 16980
rect 32306 16940 32312 16952
rect 32364 16980 32370 16992
rect 33229 16983 33287 16989
rect 33229 16980 33241 16983
rect 32364 16952 33241 16980
rect 32364 16940 32370 16952
rect 33229 16949 33241 16952
rect 33275 16949 33287 16983
rect 33229 16943 33287 16949
rect 38565 16983 38623 16989
rect 38565 16949 38577 16983
rect 38611 16980 38623 16983
rect 38654 16980 38660 16992
rect 38611 16952 38660 16980
rect 38611 16949 38623 16952
rect 38565 16943 38623 16949
rect 38654 16940 38660 16952
rect 38712 16940 38718 16992
rect 44174 16940 44180 16992
rect 44232 16980 44238 16992
rect 44361 16983 44419 16989
rect 44361 16980 44373 16983
rect 44232 16952 44373 16980
rect 44232 16940 44238 16952
rect 44361 16949 44373 16952
rect 44407 16949 44419 16983
rect 44361 16943 44419 16949
rect 1104 16890 48852 16912
rect 1104 16838 19606 16890
rect 19658 16838 19670 16890
rect 19722 16838 19734 16890
rect 19786 16838 19798 16890
rect 19850 16838 48852 16890
rect 1104 16816 48852 16838
rect 29447 16779 29505 16785
rect 29447 16745 29459 16779
rect 29493 16776 29505 16779
rect 31846 16776 31852 16788
rect 29493 16748 30328 16776
rect 31807 16748 31852 16776
rect 29493 16745 29505 16748
rect 29447 16739 29505 16745
rect 26878 16668 26884 16720
rect 26936 16668 26942 16720
rect 27154 16717 27160 16720
rect 27148 16671 27160 16717
rect 27212 16708 27218 16720
rect 29914 16708 29920 16720
rect 27212 16680 27248 16708
rect 29875 16680 29920 16708
rect 27154 16668 27160 16671
rect 27212 16668 27218 16680
rect 29914 16668 29920 16680
rect 29972 16668 29978 16720
rect 23750 16600 23756 16652
rect 23808 16640 23814 16652
rect 23845 16643 23903 16649
rect 23845 16640 23857 16643
rect 23808 16612 23857 16640
rect 23808 16600 23814 16612
rect 23845 16609 23857 16612
rect 23891 16640 23903 16643
rect 26789 16643 26847 16649
rect 23891 16612 24900 16640
rect 23891 16609 23903 16612
rect 23845 16603 23903 16609
rect 24872 16572 24900 16612
rect 26789 16609 26801 16643
rect 26835 16640 26847 16643
rect 26896 16640 26924 16668
rect 28810 16640 28816 16652
rect 26835 16612 28816 16640
rect 26835 16609 26847 16612
rect 26789 16603 26847 16609
rect 28810 16600 28816 16612
rect 28868 16600 28874 16652
rect 30006 16640 30012 16652
rect 29967 16612 30012 16640
rect 30006 16600 30012 16612
rect 30064 16600 30070 16652
rect 25314 16572 25320 16584
rect 24872 16544 25320 16572
rect 25314 16532 25320 16544
rect 25372 16532 25378 16584
rect 26878 16572 26884 16584
rect 26839 16544 26884 16572
rect 26878 16532 26884 16544
rect 26936 16532 26942 16584
rect 29273 16575 29331 16581
rect 29273 16541 29285 16575
rect 29319 16572 29331 16575
rect 29362 16572 29368 16584
rect 29319 16544 29368 16572
rect 29319 16541 29331 16544
rect 29273 16535 29331 16541
rect 29362 16532 29368 16544
rect 29420 16572 29426 16584
rect 29825 16575 29883 16581
rect 29825 16572 29837 16575
rect 29420 16544 29837 16572
rect 29420 16532 29426 16544
rect 29825 16541 29837 16544
rect 29871 16541 29883 16575
rect 30300 16572 30328 16748
rect 31846 16736 31852 16748
rect 31904 16736 31910 16788
rect 31938 16736 31944 16788
rect 31996 16776 32002 16788
rect 33229 16779 33287 16785
rect 33229 16776 33241 16779
rect 31996 16748 33241 16776
rect 31996 16736 32002 16748
rect 33229 16745 33241 16748
rect 33275 16776 33287 16779
rect 33686 16776 33692 16788
rect 33275 16748 33692 16776
rect 33275 16745 33287 16748
rect 33229 16739 33287 16745
rect 33686 16736 33692 16748
rect 33744 16776 33750 16788
rect 35161 16779 35219 16785
rect 35161 16776 35173 16779
rect 33744 16748 35173 16776
rect 33744 16736 33750 16748
rect 35161 16745 35173 16748
rect 35207 16745 35219 16779
rect 37274 16776 37280 16788
rect 37235 16748 37280 16776
rect 35161 16739 35219 16745
rect 37274 16736 37280 16748
rect 37332 16736 37338 16788
rect 39390 16736 39396 16788
rect 39448 16776 39454 16788
rect 39669 16779 39727 16785
rect 39669 16776 39681 16779
rect 39448 16748 39681 16776
rect 39448 16736 39454 16748
rect 39669 16745 39681 16748
rect 39715 16776 39727 16779
rect 40589 16779 40647 16785
rect 40589 16776 40601 16779
rect 39715 16748 40601 16776
rect 39715 16745 39727 16748
rect 39669 16739 39727 16745
rect 40589 16745 40601 16748
rect 40635 16745 40647 16779
rect 40589 16739 40647 16745
rect 32493 16711 32551 16717
rect 32493 16708 32505 16711
rect 30944 16680 32505 16708
rect 30944 16649 30972 16680
rect 32493 16677 32505 16680
rect 32539 16677 32551 16711
rect 34422 16708 34428 16720
rect 32493 16671 32551 16677
rect 33796 16680 34428 16708
rect 33796 16652 33824 16680
rect 34422 16668 34428 16680
rect 34480 16668 34486 16720
rect 38562 16717 38568 16720
rect 38556 16708 38568 16717
rect 38523 16680 38568 16708
rect 38556 16671 38568 16680
rect 38562 16668 38568 16671
rect 38620 16668 38626 16720
rect 40604 16708 40632 16739
rect 41414 16736 41420 16788
rect 41472 16776 41478 16788
rect 42153 16779 42211 16785
rect 42153 16776 42165 16779
rect 41472 16748 42165 16776
rect 41472 16736 41478 16748
rect 42153 16745 42165 16748
rect 42199 16745 42211 16779
rect 42153 16739 42211 16745
rect 42978 16736 42984 16788
rect 43036 16776 43042 16788
rect 43423 16779 43481 16785
rect 43423 16776 43435 16779
rect 43036 16748 43435 16776
rect 43036 16736 43042 16748
rect 43423 16745 43435 16748
rect 43469 16745 43481 16779
rect 43423 16739 43481 16745
rect 44821 16779 44879 16785
rect 44821 16745 44833 16779
rect 44867 16776 44879 16779
rect 45278 16776 45284 16788
rect 44867 16748 45284 16776
rect 44867 16745 44879 16748
rect 44821 16739 44879 16745
rect 45278 16736 45284 16748
rect 45336 16736 45342 16788
rect 46566 16776 46572 16788
rect 46527 16748 46572 16776
rect 46566 16736 46572 16748
rect 46624 16736 46630 16788
rect 46750 16736 46756 16788
rect 46808 16776 46814 16788
rect 47121 16779 47179 16785
rect 47121 16776 47133 16779
rect 46808 16748 47133 16776
rect 46808 16736 46814 16748
rect 47121 16745 47133 16748
rect 47167 16745 47179 16779
rect 47121 16739 47179 16745
rect 41018 16711 41076 16717
rect 41018 16708 41030 16711
rect 40604 16680 41030 16708
rect 41018 16677 41030 16680
rect 41064 16677 41076 16711
rect 41018 16671 41076 16677
rect 42242 16668 42248 16720
rect 42300 16708 42306 16720
rect 43806 16708 43812 16720
rect 42300 16680 43812 16708
rect 42300 16668 42306 16680
rect 43806 16668 43812 16680
rect 43864 16708 43870 16720
rect 43901 16711 43959 16717
rect 43901 16708 43913 16711
rect 43864 16680 43913 16708
rect 43864 16668 43870 16680
rect 43901 16677 43913 16680
rect 43947 16677 43959 16711
rect 45554 16708 45560 16720
rect 43901 16671 43959 16677
rect 45204 16680 45560 16708
rect 30837 16643 30895 16649
rect 30837 16609 30849 16643
rect 30883 16640 30895 16643
rect 30929 16643 30987 16649
rect 30929 16640 30941 16643
rect 30883 16612 30941 16640
rect 30883 16609 30895 16612
rect 30837 16603 30895 16609
rect 30929 16609 30941 16612
rect 30975 16609 30987 16643
rect 32122 16640 32128 16652
rect 32083 16612 32128 16640
rect 30929 16603 30987 16609
rect 32122 16600 32128 16612
rect 32180 16600 32186 16652
rect 32306 16640 32312 16652
rect 32267 16612 32312 16640
rect 32306 16600 32312 16612
rect 32364 16600 32370 16652
rect 33778 16640 33784 16652
rect 33691 16612 33784 16640
rect 33778 16600 33784 16612
rect 33836 16600 33842 16652
rect 34054 16649 34060 16652
rect 34048 16603 34060 16649
rect 34112 16640 34118 16652
rect 43162 16640 43168 16652
rect 34112 16612 34148 16640
rect 43123 16612 43168 16640
rect 34054 16600 34060 16603
rect 34112 16600 34118 16612
rect 43162 16600 43168 16612
rect 43220 16600 43226 16652
rect 43714 16640 43720 16652
rect 43675 16612 43720 16640
rect 43714 16600 43720 16612
rect 43772 16600 43778 16652
rect 45204 16649 45232 16680
rect 45554 16668 45560 16680
rect 45612 16708 45618 16720
rect 46106 16708 46112 16720
rect 45612 16680 46112 16708
rect 45612 16668 45618 16680
rect 46106 16668 46112 16680
rect 46164 16668 46170 16720
rect 45462 16649 45468 16652
rect 45189 16643 45247 16649
rect 45189 16609 45201 16643
rect 45235 16609 45247 16643
rect 45189 16603 45247 16609
rect 45456 16603 45468 16649
rect 45520 16640 45526 16652
rect 45520 16612 45556 16640
rect 45462 16600 45468 16603
rect 45520 16600 45526 16612
rect 30650 16572 30656 16584
rect 30300 16544 30656 16572
rect 29825 16535 29883 16541
rect 30650 16532 30656 16544
rect 30708 16532 30714 16584
rect 38286 16572 38292 16584
rect 38247 16544 38292 16572
rect 38286 16532 38292 16544
rect 38344 16532 38350 16584
rect 40402 16532 40408 16584
rect 40460 16572 40466 16584
rect 40770 16572 40776 16584
rect 40460 16544 40776 16572
rect 40460 16532 40466 16544
rect 40770 16532 40776 16544
rect 40828 16532 40834 16584
rect 43990 16572 43996 16584
rect 43951 16544 43996 16572
rect 43990 16532 43996 16544
rect 44048 16532 44054 16584
rect 28261 16439 28319 16445
rect 28261 16405 28273 16439
rect 28307 16436 28319 16439
rect 28994 16436 29000 16448
rect 28307 16408 29000 16436
rect 28307 16405 28319 16408
rect 28261 16399 28319 16405
rect 28994 16396 29000 16408
rect 29052 16396 29058 16448
rect 30466 16436 30472 16448
rect 30427 16408 30472 16436
rect 30466 16396 30472 16408
rect 30524 16396 30530 16448
rect 31113 16439 31171 16445
rect 31113 16405 31125 16439
rect 31159 16436 31171 16439
rect 31478 16436 31484 16448
rect 31159 16408 31484 16436
rect 31159 16405 31171 16408
rect 31113 16399 31171 16405
rect 31478 16396 31484 16408
rect 31536 16396 31542 16448
rect 33689 16439 33747 16445
rect 33689 16405 33701 16439
rect 33735 16436 33747 16439
rect 33962 16436 33968 16448
rect 33735 16408 33968 16436
rect 33735 16405 33747 16408
rect 33689 16399 33747 16405
rect 33962 16396 33968 16408
rect 34020 16396 34026 16448
rect 44453 16439 44511 16445
rect 44453 16405 44465 16439
rect 44499 16436 44511 16439
rect 44542 16436 44548 16448
rect 44499 16408 44548 16436
rect 44499 16405 44511 16408
rect 44453 16399 44511 16405
rect 44542 16396 44548 16408
rect 44600 16396 44606 16448
rect 1104 16346 48852 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 34966 16346
rect 35018 16294 35030 16346
rect 35082 16294 35094 16346
rect 35146 16294 35158 16346
rect 35210 16294 48852 16346
rect 1104 16272 48852 16294
rect 25314 16232 25320 16244
rect 25275 16204 25320 16232
rect 25314 16192 25320 16204
rect 25372 16192 25378 16244
rect 26786 16192 26792 16244
rect 26844 16232 26850 16244
rect 26881 16235 26939 16241
rect 26881 16232 26893 16235
rect 26844 16204 26893 16232
rect 26844 16192 26850 16204
rect 26881 16201 26893 16204
rect 26927 16201 26939 16235
rect 28994 16232 29000 16244
rect 28955 16204 29000 16232
rect 26881 16195 26939 16201
rect 28994 16192 29000 16204
rect 29052 16192 29058 16244
rect 29362 16232 29368 16244
rect 29323 16204 29368 16232
rect 29362 16192 29368 16204
rect 29420 16192 29426 16244
rect 30374 16232 30380 16244
rect 30335 16204 30380 16232
rect 30374 16192 30380 16204
rect 30432 16192 30438 16244
rect 30466 16192 30472 16244
rect 30524 16232 30530 16244
rect 30929 16235 30987 16241
rect 30929 16232 30941 16235
rect 30524 16204 30941 16232
rect 30524 16192 30530 16204
rect 30929 16201 30941 16204
rect 30975 16201 30987 16235
rect 30929 16195 30987 16201
rect 32306 16192 32312 16244
rect 32364 16232 32370 16244
rect 32493 16235 32551 16241
rect 32493 16232 32505 16235
rect 32364 16204 32505 16232
rect 32364 16192 32370 16204
rect 32493 16201 32505 16204
rect 32539 16201 32551 16235
rect 32493 16195 32551 16201
rect 33778 16192 33784 16244
rect 33836 16232 33842 16244
rect 34241 16235 34299 16241
rect 34241 16232 34253 16235
rect 33836 16204 34253 16232
rect 33836 16192 33842 16204
rect 34241 16201 34253 16204
rect 34287 16232 34299 16235
rect 34517 16235 34575 16241
rect 34517 16232 34529 16235
rect 34287 16204 34529 16232
rect 34287 16201 34299 16204
rect 34241 16195 34299 16201
rect 34517 16201 34529 16204
rect 34563 16201 34575 16235
rect 34517 16195 34575 16201
rect 34701 16235 34759 16241
rect 34701 16201 34713 16235
rect 34747 16232 34759 16235
rect 36909 16235 36967 16241
rect 36909 16232 36921 16235
rect 34747 16204 36921 16232
rect 34747 16201 34759 16204
rect 34701 16195 34759 16201
rect 36909 16201 36921 16204
rect 36955 16201 36967 16235
rect 38654 16232 38660 16244
rect 38615 16204 38660 16232
rect 36909 16195 36967 16201
rect 25332 16096 25360 16192
rect 31754 16164 31760 16176
rect 31312 16136 31760 16164
rect 31312 16108 31340 16136
rect 31754 16124 31760 16136
rect 31812 16124 31818 16176
rect 33321 16167 33379 16173
rect 33321 16133 33333 16167
rect 33367 16164 33379 16167
rect 33502 16164 33508 16176
rect 33367 16136 33508 16164
rect 33367 16133 33379 16136
rect 33321 16127 33379 16133
rect 33502 16124 33508 16136
rect 33560 16124 33566 16176
rect 34054 16164 34060 16176
rect 33888 16136 34060 16164
rect 25501 16099 25559 16105
rect 25501 16096 25513 16099
rect 25332 16068 25513 16096
rect 25501 16065 25513 16068
rect 25547 16065 25559 16099
rect 31294 16096 31300 16108
rect 31207 16068 31300 16096
rect 25501 16059 25559 16065
rect 25516 15892 25544 16059
rect 31294 16056 31300 16068
rect 31352 16056 31358 16108
rect 31478 16096 31484 16108
rect 31439 16068 31484 16096
rect 31478 16056 31484 16068
rect 31536 16056 31542 16108
rect 33686 16096 33692 16108
rect 33647 16068 33692 16096
rect 33686 16056 33692 16068
rect 33744 16056 33750 16108
rect 25774 16037 25780 16040
rect 25768 16028 25780 16037
rect 25735 16000 25780 16028
rect 25768 15991 25780 16000
rect 25774 15988 25780 15991
rect 25832 15988 25838 16040
rect 28810 15988 28816 16040
rect 28868 16028 28874 16040
rect 33137 16031 33195 16037
rect 28868 16000 29960 16028
rect 28868 15988 28874 16000
rect 27614 15920 27620 15972
rect 27672 15960 27678 15972
rect 28629 15963 28687 15969
rect 28629 15960 28641 15963
rect 27672 15932 28641 15960
rect 27672 15920 27678 15932
rect 28629 15929 28641 15932
rect 28675 15960 28687 15963
rect 29546 15960 29552 15972
rect 28675 15932 29552 15960
rect 28675 15929 28687 15932
rect 28629 15923 28687 15929
rect 29546 15920 29552 15932
rect 29604 15960 29610 15972
rect 29932 15969 29960 16000
rect 33137 15997 33149 16031
rect 33183 16028 33195 16031
rect 33888 16028 33916 16136
rect 34054 16124 34060 16136
rect 34112 16164 34118 16176
rect 34716 16164 34744 16195
rect 38654 16192 38660 16204
rect 38712 16192 38718 16244
rect 38933 16235 38991 16241
rect 38933 16201 38945 16235
rect 38979 16232 38991 16235
rect 39942 16232 39948 16244
rect 38979 16204 39948 16232
rect 38979 16201 38991 16204
rect 38933 16195 38991 16201
rect 39942 16192 39948 16204
rect 40000 16192 40006 16244
rect 43806 16232 43812 16244
rect 43767 16204 43812 16232
rect 43806 16192 43812 16204
rect 43864 16192 43870 16244
rect 44542 16232 44548 16244
rect 44503 16204 44548 16232
rect 44542 16192 44548 16204
rect 44600 16192 44606 16244
rect 45554 16232 45560 16244
rect 45515 16204 45560 16232
rect 45554 16192 45560 16204
rect 45612 16192 45618 16244
rect 34112 16136 34744 16164
rect 46201 16167 46259 16173
rect 34112 16124 34118 16136
rect 46201 16133 46213 16167
rect 46247 16133 46259 16167
rect 46201 16127 46259 16133
rect 34517 16099 34575 16105
rect 34517 16065 34529 16099
rect 34563 16096 34575 16099
rect 35345 16099 35403 16105
rect 35345 16096 35357 16099
rect 34563 16068 35357 16096
rect 34563 16065 34575 16068
rect 34517 16059 34575 16065
rect 35345 16065 35357 16068
rect 35391 16096 35403 16099
rect 35529 16099 35587 16105
rect 35529 16096 35541 16099
rect 35391 16068 35541 16096
rect 35391 16065 35403 16068
rect 35345 16059 35403 16065
rect 35529 16065 35541 16068
rect 35575 16065 35587 16099
rect 39390 16096 39396 16108
rect 39351 16068 39396 16096
rect 35529 16059 35587 16065
rect 39390 16056 39396 16068
rect 39448 16056 39454 16108
rect 42797 16099 42855 16105
rect 42797 16065 42809 16099
rect 42843 16096 42855 16099
rect 43990 16096 43996 16108
rect 42843 16068 43996 16096
rect 42843 16065 42855 16068
rect 42797 16059 42855 16065
rect 43990 16056 43996 16068
rect 44048 16056 44054 16108
rect 45005 16099 45063 16105
rect 45005 16065 45017 16099
rect 45051 16096 45063 16099
rect 45278 16096 45284 16108
rect 45051 16068 45284 16096
rect 45051 16065 45063 16068
rect 45005 16059 45063 16065
rect 45278 16056 45284 16068
rect 45336 16056 45342 16108
rect 33183 16000 33916 16028
rect 38013 16031 38071 16037
rect 33183 15997 33195 16000
rect 33137 15991 33195 15997
rect 29641 15963 29699 15969
rect 29641 15960 29653 15963
rect 29604 15932 29653 15960
rect 29604 15920 29610 15932
rect 29641 15929 29653 15932
rect 29687 15929 29699 15963
rect 29641 15923 29699 15929
rect 29917 15963 29975 15969
rect 29917 15929 29929 15963
rect 29963 15960 29975 15963
rect 30282 15960 30288 15972
rect 29963 15932 30288 15960
rect 29963 15929 29975 15932
rect 29917 15923 29975 15929
rect 30282 15920 30288 15932
rect 30340 15920 30346 15972
rect 33796 15969 33824 16000
rect 38013 15997 38025 16031
rect 38059 16028 38071 16031
rect 40589 16031 40647 16037
rect 38059 16000 39528 16028
rect 38059 15997 38071 16000
rect 38013 15991 38071 15997
rect 33781 15963 33839 15969
rect 33781 15929 33793 15963
rect 33827 15929 33839 15963
rect 33781 15923 33839 15929
rect 33873 15963 33931 15969
rect 33873 15929 33885 15963
rect 33919 15960 33931 15963
rect 33962 15960 33968 15972
rect 33919 15932 33968 15960
rect 33919 15929 33931 15932
rect 33873 15923 33931 15929
rect 33962 15920 33968 15932
rect 34020 15960 34026 15972
rect 34330 15960 34336 15972
rect 34020 15932 34336 15960
rect 34020 15920 34026 15932
rect 34330 15920 34336 15932
rect 34388 15920 34394 15972
rect 35710 15920 35716 15972
rect 35768 15969 35774 15972
rect 35768 15963 35832 15969
rect 35768 15929 35786 15963
rect 35820 15929 35832 15963
rect 35768 15923 35832 15929
rect 35768 15920 35774 15923
rect 38654 15920 38660 15972
rect 38712 15960 38718 15972
rect 39500 15969 39528 16000
rect 40589 15997 40601 16031
rect 40635 16028 40647 16031
rect 40681 16031 40739 16037
rect 40681 16028 40693 16031
rect 40635 16000 40693 16028
rect 40635 15997 40647 16000
rect 40589 15991 40647 15997
rect 40681 15997 40693 16000
rect 40727 16028 40739 16031
rect 40770 16028 40776 16040
rect 40727 16000 40776 16028
rect 40727 15997 40739 16000
rect 40681 15991 40739 15997
rect 40770 15988 40776 16000
rect 40828 15988 40834 16040
rect 40948 16031 41006 16037
rect 40948 15997 40960 16031
rect 40994 16028 41006 16031
rect 41230 16028 41236 16040
rect 40994 16000 41236 16028
rect 40994 15997 41006 16000
rect 40948 15991 41006 15997
rect 41230 15988 41236 16000
rect 41288 16028 41294 16040
rect 41414 16028 41420 16040
rect 41288 16000 41420 16028
rect 41288 15988 41294 16000
rect 41414 15988 41420 16000
rect 41472 15988 41478 16040
rect 43257 16031 43315 16037
rect 43257 16028 43269 16031
rect 43180 16000 43269 16028
rect 39393 15963 39451 15969
rect 39393 15960 39405 15963
rect 38712 15932 39405 15960
rect 38712 15920 38718 15932
rect 39393 15929 39405 15932
rect 39439 15929 39451 15963
rect 39393 15923 39451 15929
rect 39485 15963 39543 15969
rect 39485 15929 39497 15963
rect 39531 15960 39543 15963
rect 40862 15960 40868 15972
rect 39531 15932 40868 15960
rect 39531 15929 39543 15932
rect 39485 15923 39543 15929
rect 40862 15920 40868 15932
rect 40920 15920 40926 15972
rect 43180 15904 43208 16000
rect 43257 15997 43269 16000
rect 43303 15997 43315 16031
rect 46216 16028 46244 16127
rect 47121 16031 47179 16037
rect 47121 16028 47133 16031
rect 43257 15991 43315 15997
rect 45020 16000 46244 16028
rect 46492 16000 47133 16028
rect 44542 15920 44548 15972
rect 44600 15960 44606 15972
rect 45020 15969 45048 16000
rect 45005 15963 45063 15969
rect 45005 15960 45017 15963
rect 44600 15932 45017 15960
rect 44600 15920 44606 15932
rect 45005 15929 45017 15932
rect 45051 15929 45063 15963
rect 45005 15923 45063 15929
rect 45097 15963 45155 15969
rect 45097 15929 45109 15963
rect 45143 15929 45155 15963
rect 45097 15923 45155 15929
rect 26602 15892 26608 15904
rect 25516 15864 26608 15892
rect 26602 15852 26608 15864
rect 26660 15892 26666 15904
rect 26878 15892 26884 15904
rect 26660 15864 26884 15892
rect 26660 15852 26666 15864
rect 26878 15852 26884 15864
rect 26936 15892 26942 15904
rect 27433 15895 27491 15901
rect 27433 15892 27445 15895
rect 26936 15864 27445 15892
rect 26936 15852 26942 15864
rect 27433 15861 27445 15864
rect 27479 15892 27491 15895
rect 28166 15892 28172 15904
rect 27479 15864 28172 15892
rect 27479 15861 27491 15864
rect 27433 15855 27491 15861
rect 28166 15852 28172 15864
rect 28224 15852 28230 15904
rect 28350 15892 28356 15904
rect 28311 15864 28356 15892
rect 28350 15852 28356 15864
rect 28408 15852 28414 15904
rect 28994 15852 29000 15904
rect 29052 15892 29058 15904
rect 29825 15895 29883 15901
rect 29825 15892 29837 15895
rect 29052 15864 29837 15892
rect 29052 15852 29058 15864
rect 29825 15861 29837 15864
rect 29871 15861 29883 15895
rect 29825 15855 29883 15861
rect 30374 15852 30380 15904
rect 30432 15892 30438 15904
rect 30558 15892 30564 15904
rect 30432 15864 30564 15892
rect 30432 15852 30438 15864
rect 30558 15852 30564 15864
rect 30616 15892 30622 15904
rect 30653 15895 30711 15901
rect 30653 15892 30665 15895
rect 30616 15864 30665 15892
rect 30616 15852 30622 15864
rect 30653 15861 30665 15864
rect 30699 15892 30711 15895
rect 31389 15895 31447 15901
rect 31389 15892 31401 15895
rect 30699 15864 31401 15892
rect 30699 15861 30711 15864
rect 30653 15855 30711 15861
rect 31389 15861 31401 15864
rect 31435 15861 31447 15895
rect 31389 15855 31447 15861
rect 32122 15852 32128 15904
rect 32180 15892 32186 15904
rect 32217 15895 32275 15901
rect 32217 15892 32229 15895
rect 32180 15864 32229 15892
rect 32180 15852 32186 15864
rect 32217 15861 32229 15864
rect 32263 15892 32275 15895
rect 32950 15892 32956 15904
rect 32263 15864 32956 15892
rect 32263 15861 32275 15864
rect 32217 15855 32275 15861
rect 32950 15852 32956 15864
rect 33008 15852 33014 15904
rect 37918 15852 37924 15904
rect 37976 15892 37982 15904
rect 38286 15892 38292 15904
rect 37976 15864 38292 15892
rect 37976 15852 37982 15864
rect 38286 15852 38292 15864
rect 38344 15892 38350 15904
rect 39853 15895 39911 15901
rect 39853 15892 39865 15895
rect 38344 15864 39865 15892
rect 38344 15852 38350 15864
rect 39853 15861 39865 15864
rect 39899 15892 39911 15895
rect 40221 15895 40279 15901
rect 40221 15892 40233 15895
rect 39899 15864 40233 15892
rect 39899 15861 39911 15864
rect 39853 15855 39911 15861
rect 40221 15861 40233 15864
rect 40267 15892 40279 15895
rect 40589 15895 40647 15901
rect 40589 15892 40601 15895
rect 40267 15864 40601 15892
rect 40267 15861 40279 15864
rect 40221 15855 40279 15861
rect 40589 15861 40601 15864
rect 40635 15861 40647 15895
rect 42058 15892 42064 15904
rect 42019 15864 42064 15892
rect 40589 15855 40647 15861
rect 42058 15852 42064 15864
rect 42116 15852 42122 15904
rect 43162 15892 43168 15904
rect 43123 15864 43168 15892
rect 43162 15852 43168 15864
rect 43220 15852 43226 15904
rect 43438 15892 43444 15904
rect 43399 15864 43444 15892
rect 43438 15852 43444 15864
rect 43496 15852 43502 15904
rect 44266 15892 44272 15904
rect 44227 15864 44272 15892
rect 44266 15852 44272 15864
rect 44324 15852 44330 15904
rect 44818 15852 44824 15904
rect 44876 15892 44882 15904
rect 45112 15892 45140 15923
rect 45554 15920 45560 15972
rect 45612 15960 45618 15972
rect 46492 15969 46520 16000
rect 47121 15997 47133 16000
rect 47167 16028 47179 16031
rect 47486 16028 47492 16040
rect 47167 16000 47492 16028
rect 47167 15997 47179 16000
rect 47121 15991 47179 15997
rect 47486 15988 47492 16000
rect 47544 15988 47550 16040
rect 46477 15963 46535 15969
rect 46477 15960 46489 15963
rect 45612 15932 46489 15960
rect 45612 15920 45618 15932
rect 46477 15929 46489 15932
rect 46523 15929 46535 15963
rect 46477 15923 46535 15929
rect 46566 15920 46572 15972
rect 46624 15960 46630 15972
rect 46753 15963 46811 15969
rect 46753 15960 46765 15963
rect 46624 15932 46765 15960
rect 46624 15920 46630 15932
rect 46753 15929 46765 15932
rect 46799 15960 46811 15963
rect 47581 15963 47639 15969
rect 47581 15960 47593 15963
rect 46799 15932 47593 15960
rect 46799 15929 46811 15932
rect 46753 15923 46811 15929
rect 47581 15929 47593 15932
rect 47627 15929 47639 15963
rect 47581 15923 47639 15929
rect 44876 15864 45140 15892
rect 45925 15895 45983 15901
rect 44876 15852 44882 15864
rect 45925 15861 45937 15895
rect 45971 15892 45983 15895
rect 46382 15892 46388 15904
rect 45971 15864 46388 15892
rect 45971 15861 45983 15864
rect 45925 15855 45983 15861
rect 46382 15852 46388 15864
rect 46440 15892 46446 15904
rect 46661 15895 46719 15901
rect 46661 15892 46673 15895
rect 46440 15864 46673 15892
rect 46440 15852 46446 15864
rect 46661 15861 46673 15864
rect 46707 15861 46719 15895
rect 46661 15855 46719 15861
rect 1104 15802 48852 15824
rect 1104 15750 19606 15802
rect 19658 15750 19670 15802
rect 19722 15750 19734 15802
rect 19786 15750 19798 15802
rect 19850 15750 48852 15802
rect 1104 15728 48852 15750
rect 25593 15691 25651 15697
rect 25593 15657 25605 15691
rect 25639 15688 25651 15691
rect 25774 15688 25780 15700
rect 25639 15660 25780 15688
rect 25639 15657 25651 15660
rect 25593 15651 25651 15657
rect 25774 15648 25780 15660
rect 25832 15648 25838 15700
rect 26786 15648 26792 15700
rect 26844 15688 26850 15700
rect 26881 15691 26939 15697
rect 26881 15688 26893 15691
rect 26844 15660 26893 15688
rect 26844 15648 26850 15660
rect 26881 15657 26893 15660
rect 26927 15657 26939 15691
rect 29546 15688 29552 15700
rect 29507 15660 29552 15688
rect 26881 15651 26939 15657
rect 29546 15648 29552 15660
rect 29604 15648 29610 15700
rect 31294 15688 31300 15700
rect 31255 15660 31300 15688
rect 31294 15648 31300 15660
rect 31352 15648 31358 15700
rect 38654 15648 38660 15700
rect 38712 15688 38718 15700
rect 38841 15691 38899 15697
rect 38841 15688 38853 15691
rect 38712 15660 38853 15688
rect 38712 15648 38718 15660
rect 38841 15657 38853 15660
rect 38887 15657 38899 15691
rect 38841 15651 38899 15657
rect 39301 15691 39359 15697
rect 39301 15657 39313 15691
rect 39347 15688 39359 15691
rect 39390 15688 39396 15700
rect 39347 15660 39396 15688
rect 39347 15657 39359 15660
rect 39301 15651 39359 15657
rect 39390 15648 39396 15660
rect 39448 15648 39454 15700
rect 40589 15691 40647 15697
rect 40589 15657 40601 15691
rect 40635 15688 40647 15691
rect 40770 15688 40776 15700
rect 40635 15660 40776 15688
rect 40635 15657 40647 15660
rect 40589 15651 40647 15657
rect 40770 15648 40776 15660
rect 40828 15688 40834 15700
rect 41230 15688 41236 15700
rect 40828 15660 41236 15688
rect 40828 15648 40834 15660
rect 41230 15648 41236 15660
rect 41288 15648 41294 15700
rect 43438 15648 43444 15700
rect 43496 15688 43502 15700
rect 43901 15691 43959 15697
rect 43901 15688 43913 15691
rect 43496 15660 43913 15688
rect 43496 15648 43502 15660
rect 43901 15657 43913 15660
rect 43947 15688 43959 15691
rect 44174 15688 44180 15700
rect 43947 15660 44180 15688
rect 43947 15657 43959 15660
rect 43901 15651 43959 15657
rect 44174 15648 44180 15660
rect 44232 15648 44238 15700
rect 44542 15688 44548 15700
rect 44503 15660 44548 15688
rect 44542 15648 44548 15660
rect 44600 15648 44606 15700
rect 45281 15691 45339 15697
rect 45281 15657 45293 15691
rect 45327 15688 45339 15691
rect 45462 15688 45468 15700
rect 45327 15660 45468 15688
rect 45327 15657 45339 15660
rect 45281 15651 45339 15657
rect 45462 15648 45468 15660
rect 45520 15648 45526 15700
rect 47486 15688 47492 15700
rect 47447 15660 47492 15688
rect 47486 15648 47492 15660
rect 47544 15648 47550 15700
rect 28436 15623 28494 15629
rect 28436 15589 28448 15623
rect 28482 15620 28494 15623
rect 28626 15620 28632 15632
rect 28482 15592 28632 15620
rect 28482 15589 28494 15592
rect 28436 15583 28494 15589
rect 28626 15580 28632 15592
rect 28684 15620 28690 15632
rect 28994 15620 29000 15632
rect 28684 15592 29000 15620
rect 28684 15580 28690 15592
rect 28994 15580 29000 15592
rect 29052 15580 29058 15632
rect 33042 15580 33048 15632
rect 33100 15620 33106 15632
rect 33505 15623 33563 15629
rect 33505 15620 33517 15623
rect 33100 15592 33517 15620
rect 33100 15580 33106 15592
rect 33505 15589 33517 15592
rect 33551 15620 33563 15623
rect 34591 15623 34649 15629
rect 34591 15620 34603 15623
rect 33551 15592 34603 15620
rect 33551 15589 33563 15592
rect 33505 15583 33563 15589
rect 34591 15589 34603 15592
rect 34637 15589 34649 15623
rect 34591 15583 34649 15589
rect 35069 15623 35127 15629
rect 35069 15589 35081 15623
rect 35115 15620 35127 15623
rect 35250 15620 35256 15632
rect 35115 15592 35256 15620
rect 35115 15589 35127 15592
rect 35069 15583 35127 15589
rect 35250 15580 35256 15592
rect 35308 15580 35314 15632
rect 38013 15623 38071 15629
rect 38013 15589 38025 15623
rect 38059 15620 38071 15623
rect 38194 15620 38200 15632
rect 38059 15592 38200 15620
rect 38059 15589 38071 15592
rect 38013 15583 38071 15589
rect 38194 15580 38200 15592
rect 38252 15620 38258 15632
rect 41049 15623 41107 15629
rect 41049 15620 41061 15623
rect 38252 15592 41061 15620
rect 38252 15580 38258 15592
rect 41049 15589 41061 15592
rect 41095 15620 41107 15623
rect 41138 15620 41144 15632
rect 41095 15592 41144 15620
rect 41095 15589 41107 15592
rect 41049 15583 41107 15589
rect 41138 15580 41144 15592
rect 41196 15620 41202 15632
rect 42058 15620 42064 15632
rect 41196 15592 42064 15620
rect 41196 15580 41202 15592
rect 42058 15580 42064 15592
rect 42116 15580 42122 15632
rect 43070 15580 43076 15632
rect 43128 15620 43134 15632
rect 43717 15623 43775 15629
rect 43717 15620 43729 15623
rect 43128 15592 43729 15620
rect 43128 15580 43134 15592
rect 43717 15589 43729 15592
rect 43763 15620 43775 15623
rect 44082 15620 44088 15632
rect 43763 15592 44088 15620
rect 43763 15589 43775 15592
rect 43717 15583 43775 15589
rect 44082 15580 44088 15592
rect 44140 15580 44146 15632
rect 28166 15552 28172 15564
rect 28127 15524 28172 15552
rect 28166 15512 28172 15524
rect 28224 15512 28230 15564
rect 30650 15552 30656 15564
rect 30563 15524 30656 15552
rect 30650 15512 30656 15524
rect 30708 15552 30714 15564
rect 31294 15552 31300 15564
rect 30708 15524 31300 15552
rect 30708 15512 30714 15524
rect 31294 15512 31300 15524
rect 31352 15512 31358 15564
rect 34790 15512 34796 15564
rect 34848 15552 34854 15564
rect 34885 15555 34943 15561
rect 34885 15552 34897 15555
rect 34848 15524 34897 15552
rect 34848 15512 34854 15524
rect 34885 15521 34897 15524
rect 34931 15552 34943 15555
rect 35529 15555 35587 15561
rect 35529 15552 35541 15555
rect 34931 15524 35541 15552
rect 34931 15521 34943 15524
rect 34885 15515 34943 15521
rect 35529 15521 35541 15524
rect 35575 15552 35587 15555
rect 35710 15552 35716 15564
rect 35575 15524 35716 15552
rect 35575 15521 35587 15524
rect 35529 15515 35587 15521
rect 35710 15512 35716 15524
rect 35768 15512 35774 15564
rect 46106 15552 46112 15564
rect 46067 15524 46112 15552
rect 46106 15512 46112 15524
rect 46164 15512 46170 15564
rect 46382 15561 46388 15564
rect 46376 15552 46388 15561
rect 46343 15524 46388 15552
rect 46376 15515 46388 15524
rect 46382 15512 46388 15515
rect 46440 15512 46446 15564
rect 33502 15484 33508 15496
rect 33463 15456 33508 15484
rect 33502 15444 33508 15456
rect 33560 15444 33566 15496
rect 33597 15487 33655 15493
rect 33597 15453 33609 15487
rect 33643 15484 33655 15487
rect 34422 15484 34428 15496
rect 33643 15456 34428 15484
rect 33643 15453 33655 15456
rect 33597 15447 33655 15453
rect 31757 15419 31815 15425
rect 31757 15385 31769 15419
rect 31803 15416 31815 15419
rect 33612 15416 33640 15447
rect 34422 15444 34428 15456
rect 34480 15444 34486 15496
rect 35161 15487 35219 15493
rect 35161 15453 35173 15487
rect 35207 15453 35219 15487
rect 35161 15447 35219 15453
rect 35176 15416 35204 15447
rect 40862 15444 40868 15496
rect 40920 15484 40926 15496
rect 41325 15487 41383 15493
rect 41325 15484 41337 15487
rect 40920 15456 41337 15484
rect 40920 15444 40926 15456
rect 41325 15453 41337 15456
rect 41371 15484 41383 15487
rect 43990 15484 43996 15496
rect 41371 15456 41828 15484
rect 43951 15456 43996 15484
rect 41371 15453 41383 15456
rect 41325 15447 41383 15453
rect 31803 15388 33640 15416
rect 34440 15388 35204 15416
rect 31803 15385 31815 15388
rect 31757 15379 31815 15385
rect 34440 15360 34468 15388
rect 30377 15351 30435 15357
rect 30377 15317 30389 15351
rect 30423 15348 30435 15351
rect 30650 15348 30656 15360
rect 30423 15320 30656 15348
rect 30423 15317 30435 15320
rect 30377 15311 30435 15317
rect 30650 15308 30656 15320
rect 30708 15308 30714 15360
rect 30834 15348 30840 15360
rect 30795 15320 30840 15348
rect 30834 15308 30840 15320
rect 30892 15308 30898 15360
rect 32306 15348 32312 15360
rect 32267 15320 32312 15348
rect 32306 15308 32312 15320
rect 32364 15308 32370 15360
rect 33045 15351 33103 15357
rect 33045 15317 33057 15351
rect 33091 15348 33103 15351
rect 33134 15348 33140 15360
rect 33091 15320 33140 15348
rect 33091 15317 33103 15320
rect 33045 15311 33103 15317
rect 33134 15308 33140 15320
rect 33192 15308 33198 15360
rect 34422 15348 34428 15360
rect 34383 15320 34428 15348
rect 34422 15308 34428 15320
rect 34480 15308 34486 15360
rect 40773 15351 40831 15357
rect 40773 15317 40785 15351
rect 40819 15348 40831 15351
rect 41322 15348 41328 15360
rect 40819 15320 41328 15348
rect 40819 15317 40831 15320
rect 40773 15311 40831 15317
rect 41322 15308 41328 15320
rect 41380 15308 41386 15360
rect 41800 15357 41828 15456
rect 43990 15444 43996 15456
rect 44048 15444 44054 15496
rect 43254 15376 43260 15428
rect 43312 15416 43318 15428
rect 43441 15419 43499 15425
rect 43441 15416 43453 15419
rect 43312 15388 43453 15416
rect 43312 15376 43318 15388
rect 43441 15385 43453 15388
rect 43487 15385 43499 15419
rect 43441 15379 43499 15385
rect 41785 15351 41843 15357
rect 41785 15317 41797 15351
rect 41831 15348 41843 15351
rect 42334 15348 42340 15360
rect 41831 15320 42340 15348
rect 41831 15317 41843 15320
rect 41785 15311 41843 15317
rect 42334 15308 42340 15320
rect 42392 15308 42398 15360
rect 44818 15348 44824 15360
rect 44779 15320 44824 15348
rect 44818 15308 44824 15320
rect 44876 15308 44882 15360
rect 1104 15258 48852 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 34966 15258
rect 35018 15206 35030 15258
rect 35082 15206 35094 15258
rect 35146 15206 35158 15258
rect 35210 15206 48852 15258
rect 1104 15184 48852 15206
rect 28166 15144 28172 15156
rect 28127 15116 28172 15144
rect 28166 15104 28172 15116
rect 28224 15104 28230 15156
rect 28626 15144 28632 15156
rect 28587 15116 28632 15144
rect 28626 15104 28632 15116
rect 28684 15104 28690 15156
rect 30374 15144 30380 15156
rect 30335 15116 30380 15144
rect 30374 15104 30380 15116
rect 30432 15104 30438 15156
rect 31294 15144 31300 15156
rect 31255 15116 31300 15144
rect 31294 15104 31300 15116
rect 31352 15104 31358 15156
rect 31754 15104 31760 15156
rect 31812 15144 31818 15156
rect 31941 15147 31999 15153
rect 31941 15144 31953 15147
rect 31812 15116 31953 15144
rect 31812 15104 31818 15116
rect 31941 15113 31953 15116
rect 31987 15113 31999 15147
rect 31941 15107 31999 15113
rect 32953 15147 33011 15153
rect 32953 15113 32965 15147
rect 32999 15144 33011 15147
rect 33042 15144 33048 15156
rect 32999 15116 33048 15144
rect 32999 15113 33011 15116
rect 32953 15107 33011 15113
rect 33042 15104 33048 15116
rect 33100 15104 33106 15156
rect 33134 15104 33140 15156
rect 33192 15144 33198 15156
rect 33229 15147 33287 15153
rect 33229 15144 33241 15147
rect 33192 15116 33241 15144
rect 33192 15104 33198 15116
rect 33229 15113 33241 15116
rect 33275 15113 33287 15147
rect 33229 15107 33287 15113
rect 29089 15011 29147 15017
rect 29089 14977 29101 15011
rect 29135 15008 29147 15011
rect 30929 15011 30987 15017
rect 30929 15008 30941 15011
rect 29135 14980 30941 15008
rect 29135 14977 29147 14980
rect 29089 14971 29147 14977
rect 30929 14977 30941 14980
rect 30975 15008 30987 15011
rect 32306 15008 32312 15020
rect 30975 14980 32312 15008
rect 30975 14977 30987 14980
rect 30929 14971 30987 14977
rect 32306 14968 32312 14980
rect 32364 15008 32370 15020
rect 32493 15011 32551 15017
rect 32493 15008 32505 15011
rect 32364 14980 32505 15008
rect 32364 14968 32370 14980
rect 32493 14977 32505 14980
rect 32539 14977 32551 15011
rect 32493 14971 32551 14977
rect 30650 14940 30656 14952
rect 30611 14912 30656 14940
rect 30650 14900 30656 14912
rect 30708 14900 30714 14952
rect 31938 14900 31944 14952
rect 31996 14940 32002 14952
rect 32217 14943 32275 14949
rect 32217 14940 32229 14943
rect 31996 14912 32229 14940
rect 31996 14900 32002 14912
rect 32217 14909 32229 14912
rect 32263 14940 32275 14943
rect 33244 14940 33272 15107
rect 34790 15104 34796 15156
rect 34848 15144 34854 15156
rect 36541 15147 36599 15153
rect 36541 15144 36553 15147
rect 34848 15116 36553 15144
rect 34848 15104 34854 15116
rect 36541 15113 36553 15116
rect 36587 15113 36599 15147
rect 40770 15144 40776 15156
rect 40731 15116 40776 15144
rect 36541 15107 36599 15113
rect 40770 15104 40776 15116
rect 40828 15104 40834 15156
rect 41138 15144 41144 15156
rect 41099 15116 41144 15144
rect 41138 15104 41144 15116
rect 41196 15104 41202 15156
rect 43070 15144 43076 15156
rect 43031 15116 43076 15144
rect 43070 15104 43076 15116
rect 43128 15104 43134 15156
rect 44174 15144 44180 15156
rect 44135 15116 44180 15144
rect 44174 15104 44180 15116
rect 44232 15104 44238 15156
rect 46106 15104 46112 15156
rect 46164 15144 46170 15156
rect 46293 15147 46351 15153
rect 46293 15144 46305 15147
rect 46164 15116 46305 15144
rect 46164 15104 46170 15116
rect 46293 15113 46305 15116
rect 46339 15113 46351 15147
rect 46293 15107 46351 15113
rect 46842 15104 46848 15156
rect 46900 15144 46906 15156
rect 47305 15147 47363 15153
rect 47305 15144 47317 15147
rect 46900 15116 47317 15144
rect 46900 15104 46906 15116
rect 47305 15113 47317 15116
rect 47351 15113 47363 15147
rect 47305 15107 47363 15113
rect 40313 15079 40371 15085
rect 40313 15045 40325 15079
rect 40359 15076 40371 15079
rect 40862 15076 40868 15088
rect 40359 15048 40868 15076
rect 40359 15045 40371 15048
rect 40313 15039 40371 15045
rect 40862 15036 40868 15048
rect 40920 15036 40926 15088
rect 41693 15079 41751 15085
rect 41693 15045 41705 15079
rect 41739 15045 41751 15079
rect 41693 15039 41751 15045
rect 41708 15008 41736 15039
rect 42518 15036 42524 15088
rect 42576 15076 42582 15088
rect 43257 15079 43315 15085
rect 43257 15076 43269 15079
rect 42576 15048 43269 15076
rect 42576 15036 42582 15048
rect 43257 15045 43269 15048
rect 43303 15045 43315 15079
rect 46934 15076 46940 15088
rect 46895 15048 46940 15076
rect 43257 15039 43315 15045
rect 46934 15036 46940 15048
rect 46992 15036 46998 15088
rect 43625 15011 43683 15017
rect 43625 15008 43637 15011
rect 41708 14980 43637 15008
rect 43625 14977 43637 14980
rect 43671 15008 43683 15011
rect 44545 15011 44603 15017
rect 44545 15008 44557 15011
rect 43671 14980 44557 15008
rect 43671 14977 43683 14980
rect 43625 14971 43683 14977
rect 44545 14977 44557 14980
rect 44591 14977 44603 15011
rect 44545 14971 44603 14977
rect 33413 14943 33471 14949
rect 33413 14940 33425 14943
rect 32263 14912 32628 14940
rect 33244 14912 33425 14940
rect 32263 14909 32275 14912
rect 32217 14903 32275 14909
rect 30193 14875 30251 14881
rect 30193 14841 30205 14875
rect 30239 14872 30251 14875
rect 30834 14872 30840 14884
rect 30239 14844 30840 14872
rect 30239 14841 30251 14844
rect 30193 14835 30251 14841
rect 30834 14832 30840 14844
rect 30892 14832 30898 14884
rect 32600 14872 32628 14912
rect 33413 14909 33425 14912
rect 33459 14909 33471 14943
rect 35158 14940 35164 14952
rect 35119 14912 35164 14940
rect 33413 14903 33471 14909
rect 35158 14900 35164 14912
rect 35216 14900 35222 14952
rect 37918 14940 37924 14952
rect 37752 14912 37924 14940
rect 34333 14875 34391 14881
rect 32600 14844 33640 14872
rect 27614 14804 27620 14816
rect 27575 14776 27620 14804
rect 27614 14764 27620 14776
rect 27672 14764 27678 14816
rect 29733 14807 29791 14813
rect 29733 14773 29745 14807
rect 29779 14804 29791 14807
rect 30282 14804 30288 14816
rect 29779 14776 30288 14804
rect 29779 14773 29791 14776
rect 29733 14767 29791 14773
rect 30282 14764 30288 14776
rect 30340 14764 30346 14816
rect 31662 14804 31668 14816
rect 31623 14776 31668 14804
rect 31662 14764 31668 14776
rect 31720 14804 31726 14816
rect 33612 14813 33640 14844
rect 34333 14841 34345 14875
rect 34379 14872 34391 14875
rect 34701 14875 34759 14881
rect 34701 14872 34713 14875
rect 34379 14844 34713 14872
rect 34379 14841 34391 14844
rect 34333 14835 34391 14841
rect 34701 14841 34713 14844
rect 34747 14872 34759 14875
rect 35250 14872 35256 14884
rect 34747 14844 35256 14872
rect 34747 14841 34759 14844
rect 34701 14835 34759 14841
rect 35250 14832 35256 14844
rect 35308 14872 35314 14884
rect 35428 14875 35486 14881
rect 35428 14872 35440 14875
rect 35308 14844 35440 14872
rect 35308 14832 35314 14844
rect 35428 14841 35440 14844
rect 35474 14872 35486 14875
rect 36262 14872 36268 14884
rect 35474 14844 36268 14872
rect 35474 14841 35486 14844
rect 35428 14835 35486 14841
rect 36262 14832 36268 14844
rect 36320 14832 36326 14884
rect 32401 14807 32459 14813
rect 32401 14804 32413 14807
rect 31720 14776 32413 14804
rect 31720 14764 31726 14776
rect 32401 14773 32413 14776
rect 32447 14773 32459 14807
rect 32401 14767 32459 14773
rect 33597 14807 33655 14813
rect 33597 14773 33609 14807
rect 33643 14773 33655 14807
rect 33597 14767 33655 14773
rect 37642 14764 37648 14816
rect 37700 14804 37706 14816
rect 37752 14813 37780 14912
rect 37918 14900 37924 14912
rect 37976 14900 37982 14952
rect 38194 14949 38200 14952
rect 38188 14940 38200 14949
rect 38155 14912 38200 14940
rect 38188 14903 38200 14912
rect 38194 14900 38200 14903
rect 38252 14900 38258 14952
rect 41414 14900 41420 14952
rect 41472 14940 41478 14952
rect 41782 14940 41788 14952
rect 41472 14912 41788 14940
rect 41472 14900 41478 14912
rect 41782 14900 41788 14912
rect 41840 14900 41846 14952
rect 42245 14943 42303 14949
rect 42245 14909 42257 14943
rect 42291 14940 42303 14943
rect 42334 14940 42340 14952
rect 42291 14912 42340 14940
rect 42291 14909 42303 14912
rect 42245 14903 42303 14909
rect 42334 14900 42340 14912
rect 42392 14900 42398 14952
rect 42794 14900 42800 14952
rect 42852 14940 42858 14952
rect 43254 14940 43260 14952
rect 42852 14912 43260 14940
rect 42852 14900 42858 14912
rect 43254 14900 43260 14912
rect 43312 14940 43318 14952
rect 43809 14943 43867 14949
rect 43809 14940 43821 14943
rect 43312 14912 43821 14940
rect 43312 14900 43318 14912
rect 43809 14909 43821 14912
rect 43855 14940 43867 14943
rect 44450 14940 44456 14952
rect 43855 14912 44456 14940
rect 43855 14909 43867 14912
rect 43809 14903 43867 14909
rect 44450 14900 44456 14912
rect 44508 14940 44514 14952
rect 44818 14940 44824 14952
rect 44508 14912 44824 14940
rect 44508 14900 44514 14912
rect 44818 14900 44824 14912
rect 44876 14940 44882 14952
rect 44913 14943 44971 14949
rect 44913 14940 44925 14943
rect 44876 14912 44925 14940
rect 44876 14900 44882 14912
rect 44913 14909 44925 14912
rect 44959 14909 44971 14943
rect 44913 14903 44971 14909
rect 46753 14943 46811 14949
rect 46753 14909 46765 14943
rect 46799 14940 46811 14943
rect 46842 14940 46848 14952
rect 46799 14912 46848 14940
rect 46799 14909 46811 14912
rect 46753 14903 46811 14909
rect 46842 14900 46848 14912
rect 46900 14900 46906 14952
rect 41966 14872 41972 14884
rect 41927 14844 41972 14872
rect 41966 14832 41972 14844
rect 42024 14832 42030 14884
rect 45925 14875 45983 14881
rect 42628 14844 43116 14872
rect 42628 14816 42656 14844
rect 37737 14807 37795 14813
rect 37737 14804 37749 14807
rect 37700 14776 37749 14804
rect 37700 14764 37706 14776
rect 37737 14773 37749 14776
rect 37783 14773 37795 14807
rect 39298 14804 39304 14816
rect 39259 14776 39304 14804
rect 37737 14767 37795 14773
rect 39298 14764 39304 14776
rect 39356 14764 39362 14816
rect 41509 14807 41567 14813
rect 41509 14773 41521 14807
rect 41555 14804 41567 14807
rect 41782 14804 41788 14816
rect 41555 14776 41788 14804
rect 41555 14773 41567 14776
rect 41509 14767 41567 14773
rect 41782 14764 41788 14776
rect 41840 14804 41846 14816
rect 42153 14807 42211 14813
rect 42153 14804 42165 14807
rect 41840 14776 42165 14804
rect 41840 14764 41846 14776
rect 42153 14773 42165 14776
rect 42199 14773 42211 14807
rect 42610 14804 42616 14816
rect 42571 14776 42616 14804
rect 42153 14767 42211 14773
rect 42610 14764 42616 14776
rect 42668 14764 42674 14816
rect 43088 14804 43116 14844
rect 45925 14841 45937 14875
rect 45971 14872 45983 14875
rect 46382 14872 46388 14884
rect 45971 14844 46388 14872
rect 45971 14841 45983 14844
rect 45925 14835 45983 14841
rect 46382 14832 46388 14844
rect 46440 14872 46446 14884
rect 46440 14844 46888 14872
rect 46440 14832 46446 14844
rect 46860 14816 46888 14844
rect 43717 14807 43775 14813
rect 43717 14804 43729 14807
rect 43088 14776 43729 14804
rect 43717 14773 43729 14776
rect 43763 14773 43775 14807
rect 43717 14767 43775 14773
rect 46842 14764 46848 14816
rect 46900 14764 46906 14816
rect 1104 14714 48852 14736
rect 1104 14662 19606 14714
rect 19658 14662 19670 14714
rect 19722 14662 19734 14714
rect 19786 14662 19798 14714
rect 19850 14662 48852 14714
rect 1104 14640 48852 14662
rect 28350 14560 28356 14612
rect 28408 14600 28414 14612
rect 28813 14603 28871 14609
rect 28813 14600 28825 14603
rect 28408 14572 28825 14600
rect 28408 14560 28414 14572
rect 28813 14569 28825 14572
rect 28859 14600 28871 14603
rect 30285 14603 30343 14609
rect 28859 14572 29960 14600
rect 28859 14569 28871 14572
rect 28813 14563 28871 14569
rect 27522 14532 27528 14544
rect 26896 14504 27528 14532
rect 26896 14476 26924 14504
rect 27522 14492 27528 14504
rect 27580 14492 27586 14544
rect 29362 14492 29368 14544
rect 29420 14532 29426 14544
rect 29932 14541 29960 14572
rect 30285 14569 30297 14603
rect 30331 14600 30343 14603
rect 30650 14600 30656 14612
rect 30331 14572 30656 14600
rect 30331 14569 30343 14572
rect 30285 14563 30343 14569
rect 30650 14560 30656 14572
rect 30708 14560 30714 14612
rect 31113 14603 31171 14609
rect 31113 14569 31125 14603
rect 31159 14600 31171 14603
rect 31662 14600 31668 14612
rect 31159 14572 31668 14600
rect 31159 14569 31171 14572
rect 31113 14563 31171 14569
rect 31662 14560 31668 14572
rect 31720 14560 31726 14612
rect 31938 14600 31944 14612
rect 31899 14572 31944 14600
rect 31938 14560 31944 14572
rect 31996 14560 32002 14612
rect 32306 14560 32312 14612
rect 32364 14600 32370 14612
rect 32401 14603 32459 14609
rect 32401 14600 32413 14603
rect 32364 14572 32413 14600
rect 32364 14560 32370 14572
rect 32401 14569 32413 14572
rect 32447 14569 32459 14603
rect 32401 14563 32459 14569
rect 33502 14560 33508 14612
rect 33560 14600 33566 14612
rect 33597 14603 33655 14609
rect 33597 14600 33609 14603
rect 33560 14572 33609 14600
rect 33560 14560 33566 14572
rect 33597 14569 33609 14572
rect 33643 14569 33655 14603
rect 33597 14563 33655 14569
rect 34609 14603 34667 14609
rect 34609 14569 34621 14603
rect 34655 14600 34667 14603
rect 34790 14600 34796 14612
rect 34655 14572 34796 14600
rect 34655 14569 34667 14572
rect 34609 14563 34667 14569
rect 34790 14560 34796 14572
rect 34848 14560 34854 14612
rect 39114 14600 39120 14612
rect 39075 14572 39120 14600
rect 39114 14560 39120 14572
rect 39172 14560 39178 14612
rect 40129 14603 40187 14609
rect 40129 14569 40141 14603
rect 40175 14600 40187 14603
rect 41693 14603 41751 14609
rect 40175 14572 40908 14600
rect 40175 14569 40187 14572
rect 40129 14563 40187 14569
rect 40880 14544 40908 14572
rect 41693 14569 41705 14603
rect 41739 14600 41751 14603
rect 41966 14600 41972 14612
rect 41739 14572 41972 14600
rect 41739 14569 41751 14572
rect 41693 14563 41751 14569
rect 41966 14560 41972 14572
rect 42024 14560 42030 14612
rect 42242 14600 42248 14612
rect 42203 14572 42248 14600
rect 42242 14560 42248 14572
rect 42300 14560 42306 14612
rect 43165 14603 43223 14609
rect 43165 14569 43177 14603
rect 43211 14600 43223 14603
rect 43990 14600 43996 14612
rect 43211 14572 43996 14600
rect 43211 14569 43223 14572
rect 43165 14563 43223 14569
rect 43990 14560 43996 14572
rect 44048 14560 44054 14612
rect 46937 14603 46995 14609
rect 46937 14569 46949 14603
rect 46983 14569 46995 14603
rect 46937 14563 46995 14569
rect 29825 14535 29883 14541
rect 29825 14532 29837 14535
rect 29420 14504 29837 14532
rect 29420 14492 29426 14504
rect 29825 14501 29837 14504
rect 29871 14501 29883 14535
rect 29825 14495 29883 14501
rect 29917 14535 29975 14541
rect 29917 14501 29929 14535
rect 29963 14532 29975 14535
rect 30006 14532 30012 14544
rect 29963 14504 30012 14532
rect 29963 14501 29975 14504
rect 29917 14495 29975 14501
rect 30006 14492 30012 14504
rect 30064 14532 30070 14544
rect 30064 14504 32352 14532
rect 30064 14492 30070 14504
rect 26602 14464 26608 14476
rect 26563 14436 26608 14464
rect 26602 14424 26608 14436
rect 26660 14424 26666 14476
rect 26878 14473 26884 14476
rect 26872 14464 26884 14473
rect 26839 14436 26884 14464
rect 26872 14427 26884 14436
rect 26878 14424 26884 14427
rect 26936 14424 26942 14476
rect 29181 14467 29239 14473
rect 29181 14433 29193 14467
rect 29227 14464 29239 14467
rect 29641 14467 29699 14473
rect 29641 14464 29653 14467
rect 29227 14436 29653 14464
rect 29227 14433 29239 14436
rect 29181 14427 29239 14433
rect 29641 14433 29653 14436
rect 29687 14464 29699 14467
rect 29730 14464 29736 14476
rect 29687 14436 29736 14464
rect 29687 14433 29699 14436
rect 29641 14427 29699 14433
rect 29730 14424 29736 14436
rect 29788 14424 29794 14476
rect 30101 14467 30159 14473
rect 30101 14433 30113 14467
rect 30147 14464 30159 14467
rect 30653 14467 30711 14473
rect 30653 14464 30665 14467
rect 30147 14436 30665 14464
rect 30147 14433 30159 14436
rect 30101 14427 30159 14433
rect 30653 14433 30665 14436
rect 30699 14433 30711 14467
rect 30926 14464 30932 14476
rect 30887 14436 30932 14464
rect 30653 14427 30711 14433
rect 8386 14328 8392 14340
rect 8347 14300 8392 14328
rect 8386 14288 8392 14300
rect 8444 14288 8450 14340
rect 29365 14331 29423 14337
rect 29365 14297 29377 14331
rect 29411 14328 29423 14331
rect 30116 14328 30144 14427
rect 30926 14424 30932 14436
rect 30984 14424 30990 14476
rect 32122 14424 32128 14476
rect 32180 14464 32186 14476
rect 32217 14467 32275 14473
rect 32217 14464 32229 14467
rect 32180 14436 32229 14464
rect 32180 14424 32186 14436
rect 32217 14433 32229 14436
rect 32263 14433 32275 14467
rect 32217 14427 32275 14433
rect 32324 14340 32352 14504
rect 39298 14492 39304 14544
rect 39356 14532 39362 14544
rect 40727 14535 40785 14541
rect 40727 14532 40739 14535
rect 39356 14504 40739 14532
rect 39356 14492 39362 14504
rect 40727 14501 40739 14504
rect 40773 14501 40785 14535
rect 40862 14532 40868 14544
rect 40823 14504 40868 14532
rect 40727 14495 40785 14501
rect 40862 14492 40868 14504
rect 40920 14492 40926 14544
rect 41984 14532 42012 14560
rect 42794 14532 42800 14544
rect 41984 14504 42800 14532
rect 42794 14492 42800 14504
rect 42852 14492 42858 14544
rect 43070 14492 43076 14544
rect 43128 14532 43134 14544
rect 44082 14532 44088 14544
rect 43128 14504 44088 14532
rect 43128 14492 43134 14504
rect 44082 14492 44088 14504
rect 44140 14532 44146 14544
rect 44361 14535 44419 14541
rect 44361 14532 44373 14535
rect 44140 14504 44373 14532
rect 44140 14492 44146 14504
rect 44361 14501 44373 14504
rect 44407 14501 44419 14535
rect 44361 14495 44419 14501
rect 44450 14492 44456 14544
rect 44508 14532 44514 14544
rect 46952 14532 46980 14563
rect 44508 14504 46980 14532
rect 44508 14492 44514 14504
rect 38004 14467 38062 14473
rect 38004 14433 38016 14467
rect 38050 14464 38062 14467
rect 38286 14464 38292 14476
rect 38050 14436 38292 14464
rect 38050 14433 38062 14436
rect 38004 14427 38062 14433
rect 38286 14424 38292 14436
rect 38344 14424 38350 14476
rect 42061 14467 42119 14473
rect 42061 14433 42073 14467
rect 42107 14464 42119 14467
rect 42518 14464 42524 14476
rect 42107 14436 42524 14464
rect 42107 14433 42119 14436
rect 42061 14427 42119 14433
rect 42518 14424 42524 14436
rect 42576 14424 42582 14476
rect 46753 14467 46811 14473
rect 46753 14433 46765 14467
rect 46799 14464 46811 14467
rect 47210 14464 47216 14476
rect 46799 14436 47216 14464
rect 46799 14433 46811 14436
rect 46753 14427 46811 14433
rect 47210 14424 47216 14436
rect 47268 14424 47274 14476
rect 37642 14356 37648 14408
rect 37700 14396 37706 14408
rect 37737 14399 37795 14405
rect 37737 14396 37749 14399
rect 37700 14368 37749 14396
rect 37700 14356 37706 14368
rect 37737 14365 37749 14368
rect 37783 14365 37795 14399
rect 40678 14396 40684 14408
rect 40639 14368 40684 14396
rect 37737 14359 37795 14365
rect 40678 14356 40684 14368
rect 40736 14356 40742 14408
rect 44266 14396 44272 14408
rect 44227 14368 44272 14396
rect 44266 14356 44272 14368
rect 44324 14356 44330 14408
rect 29411 14300 30144 14328
rect 29411 14297 29423 14300
rect 29365 14291 29423 14297
rect 32306 14288 32312 14340
rect 32364 14328 32370 14340
rect 32953 14331 33011 14337
rect 32953 14328 32965 14331
rect 32364 14300 32965 14328
rect 32364 14288 32370 14300
rect 32953 14297 32965 14300
rect 32999 14328 33011 14331
rect 34514 14328 34520 14340
rect 32999 14300 34520 14328
rect 32999 14297 33011 14300
rect 32953 14291 33011 14297
rect 34514 14288 34520 14300
rect 34572 14288 34578 14340
rect 40313 14331 40371 14337
rect 40313 14297 40325 14331
rect 40359 14328 40371 14331
rect 42610 14328 42616 14340
rect 40359 14300 42616 14328
rect 40359 14297 40371 14300
rect 40313 14291 40371 14297
rect 42610 14288 42616 14300
rect 42668 14288 42674 14340
rect 43162 14288 43168 14340
rect 43220 14328 43226 14340
rect 43901 14331 43959 14337
rect 43901 14328 43913 14331
rect 43220 14300 43913 14328
rect 43220 14288 43226 14300
rect 43901 14297 43913 14300
rect 43947 14297 43959 14331
rect 43901 14291 43959 14297
rect 46201 14331 46259 14337
rect 46201 14297 46213 14331
rect 46247 14328 46259 14331
rect 46750 14328 46756 14340
rect 46247 14300 46756 14328
rect 46247 14297 46259 14300
rect 46201 14291 46259 14297
rect 46750 14288 46756 14300
rect 46808 14288 46814 14340
rect 19794 14260 19800 14272
rect 19755 14232 19800 14260
rect 19794 14220 19800 14232
rect 19852 14220 19858 14272
rect 27982 14260 27988 14272
rect 27943 14232 27988 14260
rect 27982 14220 27988 14232
rect 28040 14220 28046 14272
rect 31570 14260 31576 14272
rect 31531 14232 31576 14260
rect 31570 14220 31576 14232
rect 31628 14220 31634 14272
rect 33321 14263 33379 14269
rect 33321 14229 33333 14263
rect 33367 14260 33379 14263
rect 33594 14260 33600 14272
rect 33367 14232 33600 14260
rect 33367 14229 33379 14232
rect 33321 14223 33379 14229
rect 33594 14220 33600 14232
rect 33652 14220 33658 14272
rect 33962 14260 33968 14272
rect 33923 14232 33968 14260
rect 33962 14220 33968 14232
rect 34020 14220 34026 14272
rect 35250 14260 35256 14272
rect 35211 14232 35256 14260
rect 35250 14220 35256 14232
rect 35308 14220 35314 14272
rect 43622 14260 43628 14272
rect 43583 14232 43628 14260
rect 43622 14220 43628 14232
rect 43680 14220 43686 14272
rect 46566 14260 46572 14272
rect 46527 14232 46572 14260
rect 46566 14220 46572 14232
rect 46624 14220 46630 14272
rect 1104 14170 48852 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 34966 14170
rect 35018 14118 35030 14170
rect 35082 14118 35094 14170
rect 35146 14118 35158 14170
rect 35210 14118 48852 14170
rect 1104 14096 48852 14118
rect 26602 14056 26608 14068
rect 26563 14028 26608 14056
rect 26602 14016 26608 14028
rect 26660 14016 26666 14068
rect 26878 14016 26884 14068
rect 26936 14056 26942 14068
rect 26973 14059 27031 14065
rect 26973 14056 26985 14059
rect 26936 14028 26985 14056
rect 26936 14016 26942 14028
rect 26973 14025 26985 14028
rect 27019 14025 27031 14059
rect 29730 14056 29736 14068
rect 29691 14028 29736 14056
rect 26973 14019 27031 14025
rect 29730 14016 29736 14028
rect 29788 14016 29794 14068
rect 30926 14016 30932 14068
rect 30984 14056 30990 14068
rect 31021 14059 31079 14065
rect 31021 14056 31033 14059
rect 30984 14028 31033 14056
rect 30984 14016 30990 14028
rect 31021 14025 31033 14028
rect 31067 14056 31079 14059
rect 31757 14059 31815 14065
rect 31757 14056 31769 14059
rect 31067 14028 31769 14056
rect 31067 14025 31079 14028
rect 31021 14019 31079 14025
rect 31757 14025 31769 14028
rect 31803 14025 31815 14059
rect 36262 14056 36268 14068
rect 36223 14028 36268 14056
rect 31757 14019 31815 14025
rect 36262 14016 36268 14028
rect 36320 14016 36326 14068
rect 39298 14016 39304 14068
rect 39356 14056 39362 14068
rect 39853 14059 39911 14065
rect 39853 14056 39865 14059
rect 39356 14028 39865 14056
rect 39356 14016 39362 14028
rect 39853 14025 39865 14028
rect 39899 14025 39911 14059
rect 39853 14019 39911 14025
rect 41782 14016 41788 14068
rect 41840 14056 41846 14068
rect 41877 14059 41935 14065
rect 41877 14056 41889 14059
rect 41840 14028 41889 14056
rect 41840 14016 41846 14028
rect 41877 14025 41889 14028
rect 41923 14025 41935 14059
rect 42518 14056 42524 14068
rect 42479 14028 42524 14056
rect 41877 14019 41935 14025
rect 42518 14016 42524 14028
rect 42576 14016 42582 14068
rect 43070 14056 43076 14068
rect 43031 14028 43076 14056
rect 43070 14016 43076 14028
rect 43128 14016 43134 14068
rect 44266 14016 44272 14068
rect 44324 14056 44330 14068
rect 45465 14059 45523 14065
rect 45465 14056 45477 14059
rect 44324 14028 45477 14056
rect 44324 14016 44330 14028
rect 45465 14025 45477 14028
rect 45511 14056 45523 14059
rect 46201 14059 46259 14065
rect 46201 14056 46213 14059
rect 45511 14028 46213 14056
rect 45511 14025 45523 14028
rect 45465 14019 45523 14025
rect 46201 14025 46213 14028
rect 46247 14025 46259 14059
rect 47210 14056 47216 14068
rect 47171 14028 47216 14056
rect 46201 14019 46259 14025
rect 47210 14016 47216 14028
rect 47268 14016 47274 14068
rect 19334 13948 19340 14000
rect 19392 13988 19398 14000
rect 19797 13991 19855 13997
rect 19797 13988 19809 13991
rect 19392 13960 19809 13988
rect 19392 13948 19398 13960
rect 19797 13957 19809 13960
rect 19843 13957 19855 13991
rect 19797 13951 19855 13957
rect 27617 13991 27675 13997
rect 27617 13957 27629 13991
rect 27663 13988 27675 13991
rect 29362 13988 29368 14000
rect 27663 13960 29368 13988
rect 27663 13957 27675 13960
rect 27617 13951 27675 13957
rect 29362 13948 29368 13960
rect 29420 13948 29426 14000
rect 33321 13991 33379 13997
rect 33321 13988 33333 13991
rect 32048 13960 33333 13988
rect 19613 13923 19671 13929
rect 19613 13889 19625 13923
rect 19659 13920 19671 13923
rect 20254 13920 20260 13932
rect 19659 13892 20260 13920
rect 19659 13889 19671 13892
rect 19613 13883 19671 13889
rect 20254 13880 20260 13892
rect 20312 13880 20318 13932
rect 28077 13923 28135 13929
rect 28077 13889 28089 13923
rect 28123 13920 28135 13923
rect 28626 13920 28632 13932
rect 28123 13892 28632 13920
rect 28123 13889 28135 13892
rect 28077 13883 28135 13889
rect 28626 13880 28632 13892
rect 28684 13880 28690 13932
rect 30282 13920 30288 13932
rect 29012 13892 30288 13920
rect 8205 13855 8263 13861
rect 8205 13821 8217 13855
rect 8251 13852 8263 13855
rect 8294 13852 8300 13864
rect 8251 13824 8300 13852
rect 8251 13821 8263 13824
rect 8205 13815 8263 13821
rect 8294 13812 8300 13824
rect 8352 13812 8358 13864
rect 8386 13812 8392 13864
rect 8444 13852 8450 13864
rect 8553 13855 8611 13861
rect 8553 13852 8565 13855
rect 8444 13824 8565 13852
rect 8444 13812 8450 13824
rect 8553 13821 8565 13824
rect 8599 13821 8611 13855
rect 8553 13815 8611 13821
rect 19245 13855 19303 13861
rect 19245 13821 19257 13855
rect 19291 13852 19303 13855
rect 20349 13855 20407 13861
rect 20349 13852 20361 13855
rect 19291 13824 20361 13852
rect 19291 13821 19303 13824
rect 19245 13815 19303 13821
rect 20349 13821 20361 13824
rect 20395 13852 20407 13855
rect 20622 13852 20628 13864
rect 20395 13824 20628 13852
rect 20395 13821 20407 13824
rect 20349 13815 20407 13821
rect 20622 13812 20628 13824
rect 20680 13812 20686 13864
rect 27614 13812 27620 13864
rect 27672 13852 27678 13864
rect 28169 13855 28227 13861
rect 28169 13852 28181 13855
rect 27672 13824 28181 13852
rect 27672 13812 27678 13824
rect 28169 13821 28181 13824
rect 28215 13852 28227 13855
rect 29012 13852 29040 13892
rect 30282 13880 30288 13892
rect 30340 13880 30346 13932
rect 28215 13824 29040 13852
rect 29089 13855 29147 13861
rect 28215 13821 28227 13824
rect 28169 13815 28227 13821
rect 29089 13821 29101 13855
rect 29135 13852 29147 13855
rect 30009 13855 30067 13861
rect 30009 13852 30021 13855
rect 29135 13824 30021 13852
rect 29135 13821 29147 13824
rect 29089 13815 29147 13821
rect 30009 13821 30021 13824
rect 30055 13852 30067 13855
rect 30055 13824 30420 13852
rect 30055 13821 30067 13824
rect 30009 13815 30067 13821
rect 19794 13744 19800 13796
rect 19852 13784 19858 13796
rect 20257 13787 20315 13793
rect 20257 13784 20269 13787
rect 19852 13756 20269 13784
rect 19852 13744 19858 13756
rect 20257 13753 20269 13756
rect 20303 13753 20315 13787
rect 20257 13747 20315 13753
rect 27982 13744 27988 13796
rect 28040 13784 28046 13796
rect 28077 13787 28135 13793
rect 28077 13784 28089 13787
rect 28040 13756 28089 13784
rect 28040 13744 28046 13756
rect 28077 13753 28089 13756
rect 28123 13753 28135 13787
rect 30392 13784 30420 13824
rect 31570 13812 31576 13864
rect 31628 13852 31634 13864
rect 32048 13861 32076 13960
rect 33321 13957 33333 13960
rect 33367 13957 33379 13991
rect 33962 13988 33968 14000
rect 33875 13960 33968 13988
rect 33321 13951 33379 13957
rect 32306 13920 32312 13932
rect 32267 13892 32312 13920
rect 32306 13880 32312 13892
rect 32364 13880 32370 13932
rect 32858 13880 32864 13932
rect 32916 13920 32922 13932
rect 33888 13929 33916 13960
rect 33962 13948 33968 13960
rect 34020 13988 34026 14000
rect 34422 13988 34428 14000
rect 34020 13960 34428 13988
rect 34020 13948 34026 13960
rect 34422 13948 34428 13960
rect 34480 13948 34486 14000
rect 33873 13923 33931 13929
rect 33873 13920 33885 13923
rect 32916 13892 33885 13920
rect 32916 13880 32922 13892
rect 33873 13889 33885 13892
rect 33919 13889 33931 13923
rect 33873 13883 33931 13889
rect 40034 13880 40040 13932
rect 40092 13920 40098 13932
rect 40313 13923 40371 13929
rect 40313 13920 40325 13923
rect 40092 13892 40325 13920
rect 40092 13880 40098 13892
rect 40313 13889 40325 13892
rect 40359 13920 40371 13923
rect 46661 13923 46719 13929
rect 40359 13892 40540 13920
rect 40359 13889 40371 13892
rect 40313 13883 40371 13889
rect 32033 13855 32091 13861
rect 32033 13852 32045 13855
rect 31628 13824 32045 13852
rect 31628 13812 31634 13824
rect 32033 13821 32045 13824
rect 32079 13821 32091 13855
rect 32033 13815 32091 13821
rect 32122 13812 32128 13864
rect 32180 13852 32186 13864
rect 32677 13855 32735 13861
rect 32677 13852 32689 13855
rect 32180 13824 32689 13852
rect 32180 13812 32186 13824
rect 32677 13821 32689 13824
rect 32723 13821 32735 13855
rect 33594 13852 33600 13864
rect 33555 13824 33600 13852
rect 32677 13815 32735 13821
rect 33594 13812 33600 13824
rect 33652 13852 33658 13864
rect 34241 13855 34299 13861
rect 34241 13852 34253 13855
rect 33652 13824 34253 13852
rect 33652 13812 33658 13824
rect 34241 13821 34253 13824
rect 34287 13852 34299 13855
rect 34790 13852 34796 13864
rect 34287 13824 34796 13852
rect 34287 13821 34299 13824
rect 34241 13815 34299 13821
rect 34790 13812 34796 13824
rect 34848 13812 34854 13864
rect 35158 13861 35164 13864
rect 34885 13855 34943 13861
rect 34885 13821 34897 13855
rect 34931 13821 34943 13855
rect 34885 13815 34943 13821
rect 35152 13815 35164 13861
rect 35216 13852 35222 13864
rect 35216 13824 35252 13852
rect 31018 13784 31024 13796
rect 30392 13756 31024 13784
rect 28077 13747 28135 13753
rect 31018 13744 31024 13756
rect 31076 13744 31082 13796
rect 33870 13744 33876 13796
rect 33928 13784 33934 13796
rect 34609 13787 34667 13793
rect 34609 13784 34621 13787
rect 33928 13756 34621 13784
rect 33928 13744 33934 13756
rect 34609 13753 34621 13756
rect 34655 13784 34667 13787
rect 34900 13784 34928 13815
rect 35158 13812 35164 13815
rect 35216 13812 35222 13824
rect 35710 13812 35716 13864
rect 35768 13812 35774 13864
rect 37642 13812 37648 13864
rect 37700 13852 37706 13864
rect 40512 13861 40540 13892
rect 46661 13889 46673 13923
rect 46707 13920 46719 13923
rect 46750 13920 46756 13932
rect 46707 13892 46756 13920
rect 46707 13889 46719 13892
rect 46661 13883 46719 13889
rect 46750 13880 46756 13892
rect 46808 13880 46814 13932
rect 37921 13855 37979 13861
rect 37921 13852 37933 13855
rect 37700 13824 37933 13852
rect 37700 13812 37706 13824
rect 37921 13821 37933 13824
rect 37967 13852 37979 13855
rect 39577 13855 39635 13861
rect 37967 13824 38608 13852
rect 37967 13821 37979 13824
rect 37921 13815 37979 13821
rect 35250 13784 35256 13796
rect 34655 13756 35256 13784
rect 34655 13753 34667 13756
rect 34609 13747 34667 13753
rect 35250 13744 35256 13756
rect 35308 13744 35314 13796
rect 35728 13784 35756 13812
rect 36262 13784 36268 13796
rect 35728 13756 36268 13784
rect 36262 13744 36268 13756
rect 36320 13744 36326 13796
rect 38580 13784 38608 13824
rect 39577 13821 39589 13855
rect 39623 13852 39635 13855
rect 40497 13855 40555 13861
rect 39623 13824 40448 13852
rect 39623 13821 39635 13824
rect 39577 13815 39635 13821
rect 39206 13784 39212 13796
rect 38580 13756 39212 13784
rect 39206 13744 39212 13756
rect 39264 13744 39270 13796
rect 40420 13784 40448 13824
rect 40497 13821 40509 13855
rect 40543 13852 40555 13855
rect 41322 13852 41328 13864
rect 40543 13824 41328 13852
rect 40543 13821 40555 13824
rect 40497 13815 40555 13821
rect 41322 13812 41328 13824
rect 41380 13812 41386 13864
rect 43533 13855 43591 13861
rect 43533 13852 43545 13855
rect 43364 13824 43545 13852
rect 40678 13784 40684 13796
rect 40420 13756 40684 13784
rect 40678 13744 40684 13756
rect 40736 13793 40742 13796
rect 40736 13787 40800 13793
rect 40736 13753 40754 13787
rect 40788 13753 40800 13787
rect 40736 13747 40800 13753
rect 40736 13744 40742 13747
rect 4157 13719 4215 13725
rect 4157 13685 4169 13719
rect 4203 13716 4215 13719
rect 4706 13716 4712 13728
rect 4203 13688 4712 13716
rect 4203 13685 4215 13688
rect 4157 13679 4215 13685
rect 4706 13676 4712 13688
rect 4764 13676 4770 13728
rect 8754 13676 8760 13728
rect 8812 13716 8818 13728
rect 9677 13719 9735 13725
rect 9677 13716 9689 13719
rect 8812 13688 9689 13716
rect 8812 13676 8818 13688
rect 9677 13685 9689 13688
rect 9723 13685 9735 13719
rect 27430 13716 27436 13728
rect 27343 13688 27436 13716
rect 9677 13679 9735 13685
rect 27430 13676 27436 13688
rect 27488 13716 27494 13728
rect 28000 13716 28028 13744
rect 43364 13728 43392 13824
rect 43533 13821 43545 13824
rect 43579 13821 43591 13855
rect 43533 13815 43591 13821
rect 43622 13812 43628 13864
rect 43680 13852 43686 13864
rect 43789 13855 43847 13861
rect 43789 13852 43801 13855
rect 43680 13824 43801 13852
rect 43680 13812 43686 13824
rect 43789 13821 43801 13824
rect 43835 13852 43847 13855
rect 43835 13824 44128 13852
rect 43835 13821 43847 13824
rect 43789 13815 43847 13821
rect 44100 13784 44128 13824
rect 45462 13812 45468 13864
rect 45520 13852 45526 13864
rect 46566 13852 46572 13864
rect 45520 13824 46572 13852
rect 45520 13812 45526 13824
rect 46566 13812 46572 13824
rect 46624 13852 46630 13864
rect 46624 13824 46796 13852
rect 46624 13812 46630 13824
rect 44726 13784 44732 13796
rect 44100 13756 44732 13784
rect 44726 13744 44732 13756
rect 44784 13744 44790 13796
rect 46768 13793 46796 13824
rect 46753 13787 46811 13793
rect 46753 13753 46765 13787
rect 46799 13784 46811 13787
rect 47026 13784 47032 13796
rect 46799 13756 47032 13784
rect 46799 13753 46811 13756
rect 46753 13747 46811 13753
rect 47026 13744 47032 13756
rect 47084 13744 47090 13796
rect 28626 13716 28632 13728
rect 27488 13688 28028 13716
rect 28587 13688 28632 13716
rect 27488 13676 27494 13688
rect 28626 13676 28632 13688
rect 28684 13676 28690 13728
rect 29549 13719 29607 13725
rect 29549 13685 29561 13719
rect 29595 13716 29607 13719
rect 29914 13716 29920 13728
rect 29595 13688 29920 13716
rect 29595 13685 29607 13688
rect 29549 13679 29607 13685
rect 29914 13676 29920 13688
rect 29972 13716 29978 13728
rect 30193 13719 30251 13725
rect 30193 13716 30205 13719
rect 29972 13688 30205 13716
rect 29972 13676 29978 13688
rect 30193 13685 30205 13688
rect 30239 13685 30251 13719
rect 30193 13679 30251 13685
rect 31573 13719 31631 13725
rect 31573 13685 31585 13719
rect 31619 13716 31631 13719
rect 32214 13716 32220 13728
rect 31619 13688 32220 13716
rect 31619 13685 31631 13688
rect 31573 13679 31631 13685
rect 32214 13676 32220 13688
rect 32272 13676 32278 13728
rect 33137 13719 33195 13725
rect 33137 13685 33149 13719
rect 33183 13716 33195 13719
rect 33778 13716 33784 13728
rect 33183 13688 33784 13716
rect 33183 13685 33195 13688
rect 33137 13679 33195 13685
rect 33778 13676 33784 13688
rect 33836 13676 33842 13728
rect 37366 13716 37372 13728
rect 37327 13688 37372 13716
rect 37366 13676 37372 13688
rect 37424 13676 37430 13728
rect 38286 13716 38292 13728
rect 38247 13688 38292 13716
rect 38286 13676 38292 13688
rect 38344 13676 38350 13728
rect 43346 13716 43352 13728
rect 43307 13688 43352 13716
rect 43346 13676 43352 13688
rect 43404 13676 43410 13728
rect 44910 13716 44916 13728
rect 44871 13688 44916 13716
rect 44910 13676 44916 13688
rect 44968 13676 44974 13728
rect 45925 13719 45983 13725
rect 45925 13685 45937 13719
rect 45971 13716 45983 13719
rect 46382 13716 46388 13728
rect 45971 13688 46388 13716
rect 45971 13685 45983 13688
rect 45925 13679 45983 13685
rect 46382 13676 46388 13688
rect 46440 13716 46446 13728
rect 46661 13719 46719 13725
rect 46661 13716 46673 13719
rect 46440 13688 46673 13716
rect 46440 13676 46446 13688
rect 46661 13685 46673 13688
rect 46707 13685 46719 13719
rect 46661 13679 46719 13685
rect 1104 13626 48852 13648
rect 1104 13574 19606 13626
rect 19658 13574 19670 13626
rect 19722 13574 19734 13626
rect 19786 13574 19798 13626
rect 19850 13574 48852 13626
rect 1104 13552 48852 13574
rect 4617 13515 4675 13521
rect 4617 13481 4629 13515
rect 4663 13512 4675 13515
rect 4798 13512 4804 13524
rect 4663 13484 4804 13512
rect 4663 13481 4675 13484
rect 4617 13475 4675 13481
rect 4798 13472 4804 13484
rect 4856 13512 4862 13524
rect 5626 13512 5632 13524
rect 4856 13484 5632 13512
rect 4856 13472 4862 13484
rect 5626 13472 5632 13484
rect 5684 13472 5690 13524
rect 29362 13512 29368 13524
rect 29323 13484 29368 13512
rect 29362 13472 29368 13484
rect 29420 13472 29426 13524
rect 31018 13512 31024 13524
rect 30979 13484 31024 13512
rect 31018 13472 31024 13484
rect 31076 13512 31082 13524
rect 33226 13512 33232 13524
rect 31076 13484 33232 13512
rect 31076 13472 31082 13484
rect 33226 13472 33232 13484
rect 33284 13512 33290 13524
rect 33505 13515 33563 13521
rect 33505 13512 33517 13515
rect 33284 13484 33517 13512
rect 33284 13472 33290 13484
rect 33505 13481 33517 13484
rect 33551 13481 33563 13515
rect 33505 13475 33563 13481
rect 34514 13472 34520 13524
rect 34572 13512 34578 13524
rect 35805 13515 35863 13521
rect 35805 13512 35817 13515
rect 34572 13484 35817 13512
rect 34572 13472 34578 13484
rect 35805 13481 35817 13484
rect 35851 13481 35863 13515
rect 40678 13512 40684 13524
rect 40639 13484 40684 13512
rect 35805 13475 35863 13481
rect 40678 13472 40684 13484
rect 40736 13512 40742 13524
rect 41233 13515 41291 13521
rect 41233 13512 41245 13515
rect 40736 13484 41245 13512
rect 40736 13472 40742 13484
rect 41233 13481 41245 13484
rect 41279 13481 41291 13515
rect 41233 13475 41291 13481
rect 43165 13515 43223 13521
rect 43165 13481 43177 13515
rect 43211 13512 43223 13515
rect 43254 13512 43260 13524
rect 43211 13484 43260 13512
rect 43211 13481 43223 13484
rect 43165 13475 43223 13481
rect 43254 13472 43260 13484
rect 43312 13472 43318 13524
rect 44726 13512 44732 13524
rect 44687 13484 44732 13512
rect 44726 13472 44732 13484
rect 44784 13472 44790 13524
rect 46934 13472 46940 13524
rect 46992 13512 46998 13524
rect 47489 13515 47547 13521
rect 47489 13512 47501 13515
rect 46992 13484 47501 13512
rect 46992 13472 46998 13484
rect 47489 13481 47501 13484
rect 47535 13481 47547 13515
rect 47489 13475 47547 13481
rect 4706 13444 4712 13456
rect 4667 13416 4712 13444
rect 4706 13404 4712 13416
rect 4764 13444 4770 13456
rect 6273 13447 6331 13453
rect 6273 13444 6285 13447
rect 4764 13416 6285 13444
rect 4764 13404 4770 13416
rect 6273 13413 6285 13416
rect 6319 13413 6331 13447
rect 6273 13407 6331 13413
rect 2038 13308 2044 13320
rect 1951 13280 2044 13308
rect 2038 13268 2044 13280
rect 2096 13308 2102 13320
rect 3881 13311 3939 13317
rect 3881 13308 3893 13311
rect 2096 13280 3893 13308
rect 2096 13268 2102 13280
rect 3881 13277 3893 13280
rect 3927 13308 3939 13311
rect 4614 13308 4620 13320
rect 3927 13280 4620 13308
rect 3927 13277 3939 13280
rect 3881 13271 3939 13277
rect 4614 13268 4620 13280
rect 4672 13268 4678 13320
rect 1486 13132 1492 13184
rect 1544 13172 1550 13184
rect 1581 13175 1639 13181
rect 1581 13172 1593 13175
rect 1544 13144 1593 13172
rect 1544 13132 1550 13144
rect 1581 13141 1593 13144
rect 1627 13141 1639 13175
rect 1581 13135 1639 13141
rect 4062 13132 4068 13184
rect 4120 13172 4126 13184
rect 4157 13175 4215 13181
rect 4157 13172 4169 13175
rect 4120 13144 4169 13172
rect 4120 13132 4126 13144
rect 4157 13141 4169 13144
rect 4203 13141 4215 13175
rect 6288 13172 6316 13407
rect 19334 13404 19340 13456
rect 19392 13444 19398 13456
rect 27430 13453 27436 13456
rect 19797 13447 19855 13453
rect 19797 13444 19809 13447
rect 19392 13416 19809 13444
rect 19392 13404 19398 13416
rect 19797 13413 19809 13416
rect 19843 13413 19855 13447
rect 27424 13444 27436 13453
rect 27391 13416 27436 13444
rect 19797 13407 19855 13413
rect 27424 13407 27436 13416
rect 27430 13404 27436 13407
rect 27488 13404 27494 13456
rect 29914 13453 29920 13456
rect 29908 13444 29920 13453
rect 29875 13416 29920 13444
rect 29908 13407 29920 13416
rect 29914 13404 29920 13407
rect 29972 13404 29978 13456
rect 32674 13444 32680 13456
rect 32635 13416 32680 13444
rect 32674 13404 32680 13416
rect 32732 13404 32738 13456
rect 32769 13447 32827 13453
rect 32769 13413 32781 13447
rect 32815 13444 32827 13447
rect 32858 13444 32864 13456
rect 32815 13416 32864 13444
rect 32815 13413 32827 13416
rect 32769 13407 32827 13413
rect 32858 13404 32864 13416
rect 32916 13404 32922 13456
rect 35342 13444 35348 13456
rect 35303 13416 35348 13444
rect 35342 13404 35348 13416
rect 35400 13404 35406 13456
rect 37553 13447 37611 13453
rect 37553 13413 37565 13447
rect 37599 13444 37611 13447
rect 38102 13444 38108 13456
rect 37599 13416 38108 13444
rect 37599 13413 37611 13416
rect 37553 13407 37611 13413
rect 38102 13404 38108 13416
rect 38160 13444 38166 13456
rect 38289 13447 38347 13453
rect 38289 13444 38301 13447
rect 38160 13416 38301 13444
rect 38160 13404 38166 13416
rect 38289 13413 38301 13416
rect 38335 13413 38347 13447
rect 38289 13407 38347 13413
rect 39298 13404 39304 13456
rect 39356 13444 39362 13456
rect 39546 13447 39604 13453
rect 39546 13444 39558 13447
rect 39356 13416 39558 13444
rect 39356 13404 39362 13416
rect 39546 13413 39558 13416
rect 39592 13413 39604 13447
rect 39546 13407 39604 13413
rect 42794 13404 42800 13456
rect 42852 13444 42858 13456
rect 43594 13447 43652 13453
rect 43594 13444 43606 13447
rect 42852 13416 43606 13444
rect 42852 13404 42858 13416
rect 43594 13413 43606 13416
rect 43640 13413 43652 13447
rect 43594 13407 43652 13413
rect 6730 13385 6736 13388
rect 6724 13339 6736 13385
rect 6788 13376 6794 13388
rect 19610 13376 19616 13388
rect 6788 13348 6824 13376
rect 19571 13348 19616 13376
rect 6730 13336 6736 13339
rect 6788 13336 6794 13348
rect 19610 13336 19616 13348
rect 19668 13336 19674 13388
rect 26602 13336 26608 13388
rect 26660 13376 26666 13388
rect 27154 13376 27160 13388
rect 26660 13348 27160 13376
rect 26660 13336 26666 13348
rect 27154 13336 27160 13348
rect 27212 13336 27218 13388
rect 31941 13379 31999 13385
rect 31941 13345 31953 13379
rect 31987 13376 31999 13379
rect 32493 13379 32551 13385
rect 32493 13376 32505 13379
rect 31987 13348 32505 13376
rect 31987 13345 31999 13348
rect 31941 13339 31999 13345
rect 32493 13345 32505 13348
rect 32539 13376 32551 13379
rect 33042 13376 33048 13388
rect 32539 13348 33048 13376
rect 32539 13345 32551 13348
rect 32493 13339 32551 13345
rect 33042 13336 33048 13348
rect 33100 13336 33106 13388
rect 33318 13336 33324 13388
rect 33376 13376 33382 13388
rect 33781 13379 33839 13385
rect 33781 13376 33793 13379
rect 33376 13348 33793 13376
rect 33376 13336 33382 13348
rect 33781 13345 33793 13348
rect 33827 13345 33839 13379
rect 33781 13339 33839 13345
rect 6454 13308 6460 13320
rect 6415 13280 6460 13308
rect 6454 13268 6460 13280
rect 6512 13268 6518 13320
rect 18874 13268 18880 13320
rect 18932 13308 18938 13320
rect 19889 13311 19947 13317
rect 19889 13308 19901 13311
rect 18932 13280 19901 13308
rect 18932 13268 18938 13280
rect 19889 13277 19901 13280
rect 19935 13277 19947 13311
rect 29638 13308 29644 13320
rect 29599 13280 29644 13308
rect 19889 13271 19947 13277
rect 29638 13268 29644 13280
rect 29696 13268 29702 13320
rect 35360 13308 35388 13404
rect 35621 13379 35679 13385
rect 35621 13345 35633 13379
rect 35667 13376 35679 13379
rect 36170 13376 36176 13388
rect 35667 13348 36176 13376
rect 35667 13345 35679 13348
rect 35621 13339 35679 13345
rect 36170 13336 36176 13348
rect 36228 13336 36234 13388
rect 46017 13379 46075 13385
rect 46017 13345 46029 13379
rect 46063 13376 46075 13379
rect 46376 13379 46434 13385
rect 46376 13376 46388 13379
rect 46063 13348 46388 13376
rect 46063 13345 46075 13348
rect 46017 13339 46075 13345
rect 46376 13345 46388 13348
rect 46422 13376 46434 13379
rect 46750 13376 46756 13388
rect 46422 13348 46756 13376
rect 46422 13345 46434 13348
rect 46376 13339 46434 13345
rect 46750 13336 46756 13348
rect 46808 13336 46814 13388
rect 36630 13308 36636 13320
rect 35360 13280 36636 13308
rect 36630 13268 36636 13280
rect 36688 13268 36694 13320
rect 37366 13268 37372 13320
rect 37424 13308 37430 13320
rect 38194 13308 38200 13320
rect 37424 13280 38200 13308
rect 37424 13268 37430 13280
rect 38194 13268 38200 13280
rect 38252 13268 38258 13320
rect 38286 13268 38292 13320
rect 38344 13308 38350 13320
rect 38381 13311 38439 13317
rect 38381 13308 38393 13311
rect 38344 13280 38393 13308
rect 38344 13268 38350 13280
rect 38381 13277 38393 13280
rect 38427 13277 38439 13311
rect 38381 13271 38439 13277
rect 39206 13268 39212 13320
rect 39264 13308 39270 13320
rect 39301 13311 39359 13317
rect 39301 13308 39313 13311
rect 39264 13280 39313 13308
rect 39264 13268 39270 13280
rect 39301 13277 39313 13280
rect 39347 13277 39359 13311
rect 43346 13308 43352 13320
rect 43307 13280 43352 13308
rect 39301 13271 39359 13277
rect 43346 13268 43352 13280
rect 43404 13268 43410 13320
rect 46106 13308 46112 13320
rect 46067 13280 46112 13308
rect 46106 13268 46112 13280
rect 46164 13268 46170 13320
rect 32214 13240 32220 13252
rect 32175 13212 32220 13240
rect 32214 13200 32220 13212
rect 32272 13200 32278 13252
rect 37826 13240 37832 13252
rect 37787 13212 37832 13240
rect 37826 13200 37832 13212
rect 37884 13200 37890 13252
rect 7190 13172 7196 13184
rect 6288 13144 7196 13172
rect 4157 13135 4215 13141
rect 7190 13132 7196 13144
rect 7248 13132 7254 13184
rect 7374 13132 7380 13184
rect 7432 13172 7438 13184
rect 7837 13175 7895 13181
rect 7837 13172 7849 13175
rect 7432 13144 7849 13172
rect 7432 13132 7438 13144
rect 7837 13141 7849 13144
rect 7883 13141 7895 13175
rect 7837 13135 7895 13141
rect 19337 13175 19395 13181
rect 19337 13141 19349 13175
rect 19383 13172 19395 13175
rect 20257 13175 20315 13181
rect 20257 13172 20269 13175
rect 19383 13144 20269 13172
rect 19383 13141 19395 13144
rect 19337 13135 19395 13141
rect 20257 13141 20269 13144
rect 20303 13172 20315 13175
rect 20346 13172 20352 13184
rect 20303 13144 20352 13172
rect 20303 13141 20315 13144
rect 20257 13135 20315 13141
rect 20346 13132 20352 13144
rect 20404 13132 20410 13184
rect 28537 13175 28595 13181
rect 28537 13141 28549 13175
rect 28583 13172 28595 13175
rect 28626 13172 28632 13184
rect 28583 13144 28632 13172
rect 28583 13141 28595 13144
rect 28537 13135 28595 13141
rect 28626 13132 28632 13144
rect 28684 13132 28690 13184
rect 32766 13132 32772 13184
rect 32824 13172 32830 13184
rect 33137 13175 33195 13181
rect 33137 13172 33149 13175
rect 32824 13144 33149 13172
rect 32824 13132 32830 13144
rect 33137 13141 33149 13144
rect 33183 13172 33195 13175
rect 33870 13172 33876 13184
rect 33183 13144 33876 13172
rect 33183 13141 33195 13144
rect 33137 13135 33195 13141
rect 33870 13132 33876 13144
rect 33928 13132 33934 13184
rect 36170 13172 36176 13184
rect 36131 13144 36176 13172
rect 36170 13132 36176 13144
rect 36228 13132 36234 13184
rect 36906 13172 36912 13184
rect 36867 13144 36912 13172
rect 36906 13132 36912 13144
rect 36964 13132 36970 13184
rect 1104 13082 48852 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 34966 13082
rect 35018 13030 35030 13082
rect 35082 13030 35094 13082
rect 35146 13030 35158 13082
rect 35210 13030 48852 13082
rect 1104 13008 48852 13030
rect 5626 12968 5632 12980
rect 5587 12940 5632 12968
rect 5626 12928 5632 12940
rect 5684 12928 5690 12980
rect 6454 12968 6460 12980
rect 6415 12940 6460 12968
rect 6454 12928 6460 12940
rect 6512 12928 6518 12980
rect 7650 12928 7656 12980
rect 7708 12968 7714 12980
rect 7929 12971 7987 12977
rect 7929 12968 7941 12971
rect 7708 12940 7941 12968
rect 7708 12928 7714 12940
rect 7929 12937 7941 12940
rect 7975 12968 7987 12971
rect 9861 12971 9919 12977
rect 9861 12968 9873 12971
rect 7975 12940 9873 12968
rect 7975 12937 7987 12940
rect 7929 12931 7987 12937
rect 9861 12937 9873 12940
rect 9907 12937 9919 12971
rect 9861 12931 9919 12937
rect 19337 12971 19395 12977
rect 19337 12937 19349 12971
rect 19383 12968 19395 12971
rect 19426 12968 19432 12980
rect 19383 12940 19432 12968
rect 19383 12937 19395 12940
rect 19337 12931 19395 12937
rect 19426 12928 19432 12940
rect 19484 12968 19490 12980
rect 19610 12968 19616 12980
rect 19484 12940 19616 12968
rect 19484 12928 19490 12940
rect 19610 12928 19616 12940
rect 19668 12928 19674 12980
rect 27154 12968 27160 12980
rect 27115 12940 27160 12968
rect 27154 12928 27160 12940
rect 27212 12928 27218 12980
rect 27430 12928 27436 12980
rect 27488 12968 27494 12980
rect 27525 12971 27583 12977
rect 27525 12968 27537 12971
rect 27488 12940 27537 12968
rect 27488 12928 27494 12940
rect 27525 12937 27537 12940
rect 27571 12937 27583 12971
rect 27525 12931 27583 12937
rect 29914 12928 29920 12980
rect 29972 12968 29978 12980
rect 30009 12971 30067 12977
rect 30009 12968 30021 12971
rect 29972 12940 30021 12968
rect 29972 12928 29978 12940
rect 30009 12937 30021 12940
rect 30055 12937 30067 12971
rect 30009 12931 30067 12937
rect 32674 12928 32680 12980
rect 32732 12968 32738 12980
rect 34333 12971 34391 12977
rect 34333 12968 34345 12971
rect 32732 12940 34345 12968
rect 32732 12928 32738 12940
rect 34333 12937 34345 12940
rect 34379 12937 34391 12971
rect 36262 12968 36268 12980
rect 36223 12940 36268 12968
rect 34333 12931 34391 12937
rect 36262 12928 36268 12940
rect 36320 12928 36326 12980
rect 38194 12928 38200 12980
rect 38252 12968 38258 12980
rect 38749 12971 38807 12977
rect 38749 12968 38761 12971
rect 38252 12940 38761 12968
rect 38252 12928 38258 12940
rect 38749 12937 38761 12940
rect 38795 12937 38807 12971
rect 38749 12931 38807 12937
rect 39298 12928 39304 12980
rect 39356 12968 39362 12980
rect 39669 12971 39727 12977
rect 39669 12968 39681 12971
rect 39356 12940 39681 12968
rect 39356 12928 39362 12940
rect 39669 12937 39681 12940
rect 39715 12937 39727 12971
rect 39669 12931 39727 12937
rect 41417 12971 41475 12977
rect 41417 12937 41429 12971
rect 41463 12968 41475 12971
rect 43346 12968 43352 12980
rect 41463 12940 43352 12968
rect 41463 12937 41475 12940
rect 41417 12931 41475 12937
rect 6914 12860 6920 12912
rect 6972 12900 6978 12912
rect 6972 12872 7017 12900
rect 6972 12860 6978 12872
rect 31754 12860 31760 12912
rect 31812 12900 31818 12912
rect 32858 12900 32864 12912
rect 31812 12872 32864 12900
rect 31812 12860 31818 12872
rect 32858 12860 32864 12872
rect 32916 12860 32922 12912
rect 39206 12860 39212 12912
rect 39264 12900 39270 12912
rect 39393 12903 39451 12909
rect 39393 12900 39405 12903
rect 39264 12872 39405 12900
rect 39264 12860 39270 12872
rect 39393 12869 39405 12872
rect 39439 12900 39451 12903
rect 39942 12900 39948 12912
rect 39439 12872 39948 12900
rect 39439 12869 39451 12872
rect 39393 12863 39451 12869
rect 39942 12860 39948 12872
rect 40000 12860 40006 12912
rect 41524 12844 41552 12940
rect 43346 12928 43352 12940
rect 43404 12928 43410 12980
rect 44082 12968 44088 12980
rect 44043 12940 44088 12968
rect 44082 12928 44088 12940
rect 44140 12928 44146 12980
rect 45097 12971 45155 12977
rect 45097 12937 45109 12971
rect 45143 12968 45155 12971
rect 45462 12968 45468 12980
rect 45143 12940 45468 12968
rect 45143 12937 45155 12940
rect 45097 12931 45155 12937
rect 42794 12860 42800 12912
rect 42852 12900 42858 12912
rect 42889 12903 42947 12909
rect 42889 12900 42901 12903
rect 42852 12872 42901 12900
rect 42852 12860 42858 12872
rect 42889 12869 42901 12872
rect 42935 12900 42947 12903
rect 43809 12903 43867 12909
rect 43809 12900 43821 12903
rect 42935 12872 43821 12900
rect 42935 12869 42947 12872
rect 42889 12863 42947 12869
rect 43809 12869 43821 12872
rect 43855 12869 43867 12903
rect 43809 12863 43867 12869
rect 6822 12792 6828 12844
rect 6880 12832 6886 12844
rect 7374 12832 7380 12844
rect 6880 12804 7380 12832
rect 6880 12792 6886 12804
rect 7374 12792 7380 12804
rect 7432 12792 7438 12844
rect 20346 12832 20352 12844
rect 20307 12804 20352 12832
rect 20346 12792 20352 12804
rect 20404 12792 20410 12844
rect 41506 12832 41512 12844
rect 41419 12804 41512 12832
rect 41506 12792 41512 12804
rect 41564 12792 41570 12844
rect 44542 12832 44548 12844
rect 44455 12804 44548 12832
rect 44542 12792 44548 12804
rect 44600 12832 44606 12844
rect 44910 12832 44916 12844
rect 44600 12804 44916 12832
rect 44600 12792 44606 12804
rect 44910 12792 44916 12804
rect 44968 12792 44974 12844
rect 1486 12764 1492 12776
rect 1447 12736 1492 12764
rect 1486 12724 1492 12736
rect 1544 12724 1550 12776
rect 1756 12767 1814 12773
rect 1756 12733 1768 12767
rect 1802 12764 1814 12767
rect 2038 12764 2044 12776
rect 1802 12736 2044 12764
rect 1802 12733 1814 12736
rect 1756 12727 1814 12733
rect 2038 12724 2044 12736
rect 2096 12724 2102 12776
rect 4154 12764 4160 12776
rect 4067 12736 4160 12764
rect 4154 12724 4160 12736
rect 4212 12764 4218 12776
rect 4249 12767 4307 12773
rect 4249 12764 4261 12767
rect 4212 12736 4261 12764
rect 4212 12724 4218 12736
rect 4249 12733 4261 12736
rect 4295 12764 4307 12767
rect 6454 12764 6460 12776
rect 4295 12736 6460 12764
rect 4295 12733 4307 12736
rect 4249 12727 4307 12733
rect 6454 12724 6460 12736
rect 6512 12764 6518 12776
rect 7006 12764 7012 12776
rect 6512 12736 7012 12764
rect 6512 12724 6518 12736
rect 7006 12724 7012 12736
rect 7064 12724 7070 12776
rect 7190 12724 7196 12776
rect 7248 12764 7254 12776
rect 7469 12767 7527 12773
rect 7469 12764 7481 12767
rect 7248 12736 7481 12764
rect 7248 12724 7254 12736
rect 7469 12733 7481 12736
rect 7515 12733 7527 12767
rect 7469 12727 7527 12733
rect 8294 12724 8300 12776
rect 8352 12764 8358 12776
rect 8754 12773 8760 12776
rect 8481 12767 8539 12773
rect 8481 12764 8493 12767
rect 8352 12736 8493 12764
rect 8352 12724 8358 12736
rect 8481 12733 8493 12736
rect 8527 12764 8539 12767
rect 8748 12764 8760 12773
rect 8527 12736 8616 12764
rect 8715 12736 8760 12764
rect 8527 12733 8539 12736
rect 8481 12727 8539 12733
rect 3789 12699 3847 12705
rect 3789 12665 3801 12699
rect 3835 12696 3847 12699
rect 4494 12699 4552 12705
rect 4494 12696 4506 12699
rect 3835 12668 4506 12696
rect 3835 12665 3847 12668
rect 3789 12659 3847 12665
rect 4494 12665 4506 12668
rect 4540 12696 4552 12699
rect 5534 12696 5540 12708
rect 4540 12668 5540 12696
rect 4540 12665 4552 12668
rect 4494 12659 4552 12665
rect 5534 12656 5540 12668
rect 5592 12656 5598 12708
rect 2682 12588 2688 12640
rect 2740 12628 2746 12640
rect 2869 12631 2927 12637
rect 2869 12628 2881 12631
rect 2740 12600 2881 12628
rect 2740 12588 2746 12600
rect 2869 12597 2881 12600
rect 2915 12597 2927 12631
rect 2869 12591 2927 12597
rect 6730 12588 6736 12640
rect 6788 12628 6794 12640
rect 7377 12631 7435 12637
rect 7377 12628 7389 12631
rect 6788 12600 7389 12628
rect 6788 12588 6794 12600
rect 7377 12597 7389 12600
rect 7423 12628 7435 12631
rect 7650 12628 7656 12640
rect 7423 12600 7656 12628
rect 7423 12597 7435 12600
rect 7377 12591 7435 12597
rect 7650 12588 7656 12600
rect 7708 12588 7714 12640
rect 8389 12631 8447 12637
rect 8389 12597 8401 12631
rect 8435 12628 8447 12631
rect 8588 12628 8616 12736
rect 8748 12727 8760 12736
rect 8754 12724 8760 12727
rect 8812 12724 8818 12776
rect 19889 12767 19947 12773
rect 19889 12733 19901 12767
rect 19935 12764 19947 12767
rect 19978 12764 19984 12776
rect 19935 12736 19984 12764
rect 19935 12733 19947 12736
rect 19889 12727 19947 12733
rect 19978 12724 19984 12736
rect 20036 12724 20042 12776
rect 20254 12724 20260 12776
rect 20312 12764 20318 12776
rect 20625 12767 20683 12773
rect 20625 12764 20637 12767
rect 20312 12736 20637 12764
rect 20312 12724 20318 12736
rect 20625 12733 20637 12736
rect 20671 12733 20683 12767
rect 20625 12727 20683 12733
rect 32122 12724 32128 12776
rect 32180 12764 32186 12776
rect 32766 12764 32772 12776
rect 32180 12736 32772 12764
rect 32180 12724 32186 12736
rect 32766 12724 32772 12736
rect 32824 12764 32830 12776
rect 33226 12773 33232 12776
rect 32953 12767 33011 12773
rect 32953 12764 32965 12767
rect 32824 12736 32965 12764
rect 32824 12724 32830 12736
rect 32953 12733 32965 12736
rect 32999 12733 33011 12767
rect 33220 12764 33232 12773
rect 33187 12736 33232 12764
rect 32953 12727 33011 12733
rect 33220 12727 33232 12736
rect 33226 12724 33232 12727
rect 33284 12724 33290 12776
rect 34606 12724 34612 12776
rect 34664 12764 34670 12776
rect 34885 12767 34943 12773
rect 34885 12764 34897 12767
rect 34664 12736 34897 12764
rect 34664 12724 34670 12736
rect 34885 12733 34897 12736
rect 34931 12733 34943 12767
rect 36814 12764 36820 12776
rect 36775 12736 36820 12764
rect 34885 12727 34943 12733
rect 36814 12724 36820 12736
rect 36872 12724 36878 12776
rect 36906 12724 36912 12776
rect 36964 12764 36970 12776
rect 41782 12773 41788 12776
rect 37073 12767 37131 12773
rect 37073 12764 37085 12767
rect 36964 12736 37085 12764
rect 36964 12724 36970 12736
rect 37073 12733 37085 12736
rect 37119 12764 37131 12767
rect 41776 12764 41788 12773
rect 37119 12736 37228 12764
rect 37119 12733 37131 12736
rect 37073 12727 37131 12733
rect 37200 12708 37228 12736
rect 41708 12736 41788 12764
rect 31113 12699 31171 12705
rect 31113 12665 31125 12699
rect 31159 12665 31171 12699
rect 31113 12659 31171 12665
rect 32861 12699 32919 12705
rect 32861 12665 32873 12699
rect 32907 12665 32919 12699
rect 32861 12659 32919 12665
rect 9582 12628 9588 12640
rect 8435 12600 9588 12628
rect 8435 12597 8447 12600
rect 8389 12591 8447 12597
rect 9582 12588 9588 12600
rect 9640 12588 9646 12640
rect 18874 12628 18880 12640
rect 18835 12600 18880 12628
rect 18874 12588 18880 12600
rect 18932 12588 18938 12640
rect 19797 12631 19855 12637
rect 19797 12597 19809 12631
rect 19843 12628 19855 12631
rect 20351 12631 20409 12637
rect 20351 12628 20363 12631
rect 19843 12600 20363 12628
rect 19843 12597 19855 12600
rect 19797 12591 19855 12597
rect 20351 12597 20363 12600
rect 20397 12628 20409 12631
rect 20438 12628 20444 12640
rect 20397 12600 20444 12628
rect 20397 12597 20409 12600
rect 20351 12591 20409 12597
rect 20438 12588 20444 12600
rect 20496 12588 20502 12640
rect 20714 12588 20720 12640
rect 20772 12628 20778 12640
rect 21729 12631 21787 12637
rect 21729 12628 21741 12631
rect 20772 12600 21741 12628
rect 20772 12588 20778 12600
rect 21729 12597 21741 12600
rect 21775 12597 21787 12631
rect 29638 12628 29644 12640
rect 29599 12600 29644 12628
rect 21729 12591 21787 12597
rect 29638 12588 29644 12600
rect 29696 12588 29702 12640
rect 31018 12628 31024 12640
rect 30979 12600 31024 12628
rect 31018 12588 31024 12600
rect 31076 12628 31082 12640
rect 31128 12628 31156 12659
rect 31076 12600 31156 12628
rect 32876 12628 32904 12659
rect 33778 12656 33784 12708
rect 33836 12696 33842 12708
rect 35130 12699 35188 12705
rect 35130 12696 35142 12699
rect 33836 12668 35142 12696
rect 33836 12656 33842 12668
rect 35130 12665 35142 12668
rect 35176 12696 35188 12699
rect 35250 12696 35256 12708
rect 35176 12668 35256 12696
rect 35176 12665 35188 12668
rect 35130 12659 35188 12665
rect 35250 12656 35256 12668
rect 35308 12656 35314 12708
rect 37182 12656 37188 12708
rect 37240 12656 37246 12708
rect 41049 12699 41107 12705
rect 41049 12665 41061 12699
rect 41095 12696 41107 12699
rect 41708 12696 41736 12736
rect 41776 12727 41788 12736
rect 41782 12724 41788 12727
rect 41840 12724 41846 12776
rect 43346 12724 43352 12776
rect 43404 12764 43410 12776
rect 43533 12767 43591 12773
rect 43533 12764 43545 12767
rect 43404 12736 43545 12764
rect 43404 12724 43410 12736
rect 43533 12733 43545 12736
rect 43579 12764 43591 12767
rect 44082 12764 44088 12776
rect 43579 12736 44088 12764
rect 43579 12733 43591 12736
rect 43533 12727 43591 12733
rect 44082 12724 44088 12736
rect 44140 12724 44146 12776
rect 44637 12767 44695 12773
rect 44637 12733 44649 12767
rect 44683 12764 44695 12767
rect 45112 12764 45140 12931
rect 45462 12928 45468 12940
rect 45520 12928 45526 12980
rect 46750 12928 46756 12980
rect 46808 12968 46814 12980
rect 47489 12971 47547 12977
rect 47489 12968 47501 12971
rect 46808 12940 47501 12968
rect 46808 12928 46814 12940
rect 47489 12937 47501 12940
rect 47535 12937 47547 12971
rect 47489 12931 47547 12937
rect 46106 12764 46112 12776
rect 44683 12736 45140 12764
rect 45848 12736 46112 12764
rect 44683 12733 44695 12736
rect 44637 12727 44695 12733
rect 41095 12668 41736 12696
rect 41095 12665 41107 12668
rect 41049 12659 41107 12665
rect 33226 12628 33232 12640
rect 32876 12600 33232 12628
rect 31076 12588 31082 12600
rect 33226 12588 33232 12600
rect 33284 12588 33290 12640
rect 38194 12628 38200 12640
rect 38155 12600 38200 12628
rect 38194 12588 38200 12600
rect 38252 12588 38258 12640
rect 41322 12588 41328 12640
rect 41380 12628 41386 12640
rect 41506 12628 41512 12640
rect 41380 12600 41512 12628
rect 41380 12588 41386 12600
rect 41506 12588 41512 12600
rect 41564 12588 41570 12640
rect 44082 12588 44088 12640
rect 44140 12628 44146 12640
rect 44545 12631 44603 12637
rect 44545 12628 44557 12631
rect 44140 12600 44557 12628
rect 44140 12588 44146 12600
rect 44545 12597 44557 12600
rect 44591 12628 44603 12631
rect 44726 12628 44732 12640
rect 44591 12600 44732 12628
rect 44591 12597 44603 12600
rect 44545 12591 44603 12597
rect 44726 12588 44732 12600
rect 44784 12588 44790 12640
rect 45554 12628 45560 12640
rect 45515 12600 45560 12628
rect 45554 12588 45560 12600
rect 45612 12628 45618 12640
rect 45848 12637 45876 12736
rect 46106 12724 46112 12736
rect 46164 12724 46170 12776
rect 46382 12773 46388 12776
rect 46376 12764 46388 12773
rect 46343 12736 46388 12764
rect 46376 12727 46388 12736
rect 46382 12724 46388 12727
rect 46440 12724 46446 12776
rect 45833 12631 45891 12637
rect 45833 12628 45845 12631
rect 45612 12600 45845 12628
rect 45612 12588 45618 12600
rect 45833 12597 45845 12600
rect 45879 12597 45891 12631
rect 45833 12591 45891 12597
rect 1104 12538 48852 12560
rect 1104 12486 19606 12538
rect 19658 12486 19670 12538
rect 19722 12486 19734 12538
rect 19786 12486 19798 12538
rect 19850 12486 48852 12538
rect 1104 12464 48852 12486
rect 4614 12384 4620 12436
rect 4672 12424 4678 12436
rect 5445 12427 5503 12433
rect 5445 12424 5457 12427
rect 4672 12396 5457 12424
rect 4672 12384 4678 12396
rect 5445 12393 5457 12396
rect 5491 12393 5503 12427
rect 5445 12387 5503 12393
rect 5534 12384 5540 12436
rect 5592 12424 5598 12436
rect 6365 12427 6423 12433
rect 6365 12424 6377 12427
rect 5592 12396 6377 12424
rect 5592 12384 5598 12396
rect 6365 12393 6377 12396
rect 6411 12424 6423 12427
rect 6822 12424 6828 12436
rect 6411 12396 6828 12424
rect 6411 12393 6423 12396
rect 6365 12387 6423 12393
rect 6822 12384 6828 12396
rect 6880 12384 6886 12436
rect 7650 12424 7656 12436
rect 7611 12396 7656 12424
rect 7650 12384 7656 12396
rect 7708 12384 7714 12436
rect 8573 12427 8631 12433
rect 8573 12393 8585 12427
rect 8619 12424 8631 12427
rect 8754 12424 8760 12436
rect 8619 12396 8760 12424
rect 8619 12393 8631 12396
rect 8573 12387 8631 12393
rect 8754 12384 8760 12396
rect 8812 12384 8818 12436
rect 19334 12424 19340 12436
rect 19295 12396 19340 12424
rect 19334 12384 19340 12396
rect 19392 12384 19398 12436
rect 19426 12384 19432 12436
rect 19484 12424 19490 12436
rect 19521 12427 19579 12433
rect 19521 12424 19533 12427
rect 19484 12396 19533 12424
rect 19484 12384 19490 12396
rect 19521 12393 19533 12396
rect 19567 12393 19579 12427
rect 19521 12387 19579 12393
rect 20073 12427 20131 12433
rect 20073 12393 20085 12427
rect 20119 12424 20131 12427
rect 20254 12424 20260 12436
rect 20119 12396 20260 12424
rect 20119 12393 20131 12396
rect 20073 12387 20131 12393
rect 20254 12384 20260 12396
rect 20312 12384 20318 12436
rect 22278 12424 22284 12436
rect 22239 12396 22284 12424
rect 22278 12384 22284 12396
rect 22336 12384 22342 12436
rect 29733 12427 29791 12433
rect 29733 12393 29745 12427
rect 29779 12424 29791 12427
rect 29914 12424 29920 12436
rect 29779 12396 29920 12424
rect 29779 12393 29791 12396
rect 29733 12387 29791 12393
rect 29914 12384 29920 12396
rect 29972 12384 29978 12436
rect 31573 12427 31631 12433
rect 31573 12393 31585 12427
rect 31619 12424 31631 12427
rect 31662 12424 31668 12436
rect 31619 12396 31668 12424
rect 31619 12393 31631 12396
rect 31573 12387 31631 12393
rect 31662 12384 31668 12396
rect 31720 12384 31726 12436
rect 33134 12384 33140 12436
rect 33192 12424 33198 12436
rect 33505 12427 33563 12433
rect 33505 12424 33517 12427
rect 33192 12396 33517 12424
rect 33192 12384 33198 12396
rect 33505 12393 33517 12396
rect 33551 12424 33563 12427
rect 34238 12424 34244 12436
rect 33551 12396 34244 12424
rect 33551 12393 33563 12396
rect 33505 12387 33563 12393
rect 34238 12384 34244 12396
rect 34296 12384 34302 12436
rect 35250 12384 35256 12436
rect 35308 12424 35314 12436
rect 35989 12427 36047 12433
rect 35989 12424 36001 12427
rect 35308 12396 36001 12424
rect 35308 12384 35314 12396
rect 35989 12393 36001 12396
rect 36035 12393 36047 12427
rect 35989 12387 36047 12393
rect 37553 12427 37611 12433
rect 37553 12393 37565 12427
rect 37599 12424 37611 12427
rect 38194 12424 38200 12436
rect 37599 12396 38200 12424
rect 37599 12393 37611 12396
rect 37553 12387 37611 12393
rect 38194 12384 38200 12396
rect 38252 12384 38258 12436
rect 41046 12384 41052 12436
rect 41104 12424 41110 12436
rect 41325 12427 41383 12433
rect 41325 12424 41337 12427
rect 41104 12396 41337 12424
rect 41104 12384 41110 12396
rect 41325 12393 41337 12396
rect 41371 12393 41383 12427
rect 44082 12424 44088 12436
rect 44043 12396 44088 12424
rect 41325 12387 41383 12393
rect 44082 12384 44088 12396
rect 44140 12384 44146 12436
rect 47026 12384 47032 12436
rect 47084 12424 47090 12436
rect 47673 12427 47731 12433
rect 47673 12424 47685 12427
rect 47084 12396 47685 12424
rect 47084 12384 47090 12396
rect 47673 12393 47685 12396
rect 47719 12393 47731 12427
rect 47673 12387 47731 12393
rect 1756 12359 1814 12365
rect 1756 12325 1768 12359
rect 1802 12356 1814 12359
rect 2314 12356 2320 12368
rect 1802 12328 2320 12356
rect 1802 12325 1814 12328
rect 1756 12319 1814 12325
rect 2314 12316 2320 12328
rect 2372 12356 2378 12368
rect 2682 12356 2688 12368
rect 2372 12328 2688 12356
rect 2372 12316 2378 12328
rect 2682 12316 2688 12328
rect 2740 12316 2746 12368
rect 3881 12359 3939 12365
rect 3881 12325 3893 12359
rect 3927 12356 3939 12359
rect 4332 12359 4390 12365
rect 4332 12356 4344 12359
rect 3927 12328 4344 12356
rect 3927 12325 3939 12328
rect 3881 12319 3939 12325
rect 4332 12325 4344 12328
rect 4378 12356 4390 12359
rect 4798 12356 4804 12368
rect 4378 12328 4804 12356
rect 4378 12325 4390 12328
rect 4332 12319 4390 12325
rect 4798 12316 4804 12328
rect 4856 12316 4862 12368
rect 7098 12356 7104 12368
rect 7059 12328 7104 12356
rect 7098 12316 7104 12328
rect 7156 12316 7162 12368
rect 18230 12316 18236 12368
rect 18288 12356 18294 12368
rect 18509 12359 18567 12365
rect 18509 12356 18521 12359
rect 18288 12328 18521 12356
rect 18288 12316 18294 12328
rect 18509 12325 18521 12328
rect 18555 12356 18567 12359
rect 20622 12356 20628 12368
rect 18555 12328 20628 12356
rect 18555 12325 18567 12328
rect 18509 12319 18567 12325
rect 20622 12316 20628 12328
rect 20680 12316 20686 12368
rect 20806 12316 20812 12368
rect 20864 12356 20870 12368
rect 21168 12359 21226 12365
rect 21168 12356 21180 12359
rect 20864 12328 21180 12356
rect 20864 12316 20870 12328
rect 21168 12325 21180 12328
rect 21214 12356 21226 12359
rect 21358 12356 21364 12368
rect 21214 12328 21364 12356
rect 21214 12325 21226 12328
rect 21168 12319 21226 12325
rect 21358 12316 21364 12328
rect 21416 12316 21422 12368
rect 29638 12356 29644 12368
rect 28368 12328 29644 12356
rect 28368 12300 28396 12328
rect 29638 12316 29644 12328
rect 29696 12316 29702 12368
rect 31941 12359 31999 12365
rect 31941 12325 31953 12359
rect 31987 12356 31999 12359
rect 32392 12359 32450 12365
rect 32392 12356 32404 12359
rect 31987 12328 32404 12356
rect 31987 12325 31999 12328
rect 31941 12319 31999 12325
rect 32392 12325 32404 12328
rect 32438 12356 32450 12359
rect 32674 12356 32680 12368
rect 32438 12328 32680 12356
rect 32438 12325 32450 12328
rect 32392 12319 32450 12325
rect 32674 12316 32680 12328
rect 32732 12316 32738 12368
rect 34256 12356 34284 12384
rect 34854 12359 34912 12365
rect 34854 12356 34866 12359
rect 34256 12328 34866 12356
rect 34854 12325 34866 12328
rect 34900 12325 34912 12359
rect 34854 12319 34912 12325
rect 36814 12316 36820 12368
rect 36872 12356 36878 12368
rect 36909 12359 36967 12365
rect 36909 12356 36921 12359
rect 36872 12328 36921 12356
rect 36872 12316 36878 12328
rect 36909 12325 36921 12328
rect 36955 12356 36967 12359
rect 37642 12356 37648 12368
rect 36955 12328 37648 12356
rect 36955 12325 36967 12328
rect 36909 12319 36967 12325
rect 37642 12316 37648 12328
rect 37700 12316 37706 12368
rect 38562 12356 38568 12368
rect 38523 12328 38568 12356
rect 38562 12316 38568 12328
rect 38620 12316 38626 12368
rect 39758 12316 39764 12368
rect 39816 12356 39822 12368
rect 40129 12359 40187 12365
rect 40129 12356 40141 12359
rect 39816 12328 40141 12356
rect 39816 12316 39822 12328
rect 40129 12325 40141 12328
rect 40175 12325 40187 12359
rect 40129 12319 40187 12325
rect 45002 12316 45008 12368
rect 45060 12356 45066 12368
rect 45462 12356 45468 12368
rect 45060 12328 45468 12356
rect 45060 12316 45066 12328
rect 45462 12316 45468 12328
rect 45520 12316 45526 12368
rect 1486 12288 1492 12300
rect 1399 12260 1492 12288
rect 1486 12248 1492 12260
rect 1544 12288 1550 12300
rect 4154 12288 4160 12300
rect 1544 12260 4160 12288
rect 1544 12248 1550 12260
rect 4154 12248 4160 12260
rect 4212 12248 4218 12300
rect 6914 12288 6920 12300
rect 6875 12260 6920 12288
rect 6914 12248 6920 12260
rect 6972 12248 6978 12300
rect 9950 12297 9956 12300
rect 9944 12288 9956 12297
rect 9911 12260 9956 12288
rect 9944 12251 9956 12260
rect 9950 12248 9956 12251
rect 10008 12248 10014 12300
rect 17862 12248 17868 12300
rect 17920 12288 17926 12300
rect 18325 12291 18383 12297
rect 18325 12288 18337 12291
rect 17920 12260 18337 12288
rect 17920 12248 17926 12260
rect 18325 12257 18337 12260
rect 18371 12288 18383 12291
rect 19886 12288 19892 12300
rect 18371 12260 19892 12288
rect 18371 12257 18383 12260
rect 18325 12251 18383 12257
rect 19886 12248 19892 12260
rect 19944 12248 19950 12300
rect 27154 12248 27160 12300
rect 27212 12288 27218 12300
rect 28350 12288 28356 12300
rect 27212 12260 28356 12288
rect 27212 12248 27218 12260
rect 28350 12248 28356 12260
rect 28408 12248 28414 12300
rect 28626 12297 28632 12300
rect 28620 12288 28632 12297
rect 28587 12260 28632 12288
rect 28620 12251 28632 12260
rect 28626 12248 28632 12251
rect 28684 12248 28690 12300
rect 36832 12288 36860 12316
rect 38378 12288 38384 12300
rect 34624 12260 36860 12288
rect 38339 12260 38384 12288
rect 3970 12180 3976 12232
rect 4028 12220 4034 12232
rect 4065 12223 4123 12229
rect 4065 12220 4077 12223
rect 4028 12192 4077 12220
rect 4028 12180 4034 12192
rect 4065 12189 4077 12192
rect 4111 12220 4123 12223
rect 4172 12220 4200 12248
rect 34624 12232 34652 12260
rect 38378 12248 38384 12260
rect 38436 12248 38442 12300
rect 41141 12291 41199 12297
rect 41141 12288 41153 12291
rect 40052 12260 41153 12288
rect 40052 12232 40080 12260
rect 41141 12257 41153 12260
rect 41187 12288 41199 12291
rect 41506 12288 41512 12300
rect 41187 12260 41512 12288
rect 41187 12257 41199 12260
rect 41141 12251 41199 12257
rect 41506 12248 41512 12260
rect 41564 12248 41570 12300
rect 44453 12291 44511 12297
rect 44453 12257 44465 12291
rect 44499 12288 44511 12291
rect 44542 12288 44548 12300
rect 44499 12260 44548 12288
rect 44499 12257 44511 12260
rect 44453 12251 44511 12257
rect 44542 12248 44548 12260
rect 44600 12288 44606 12300
rect 45278 12297 45284 12300
rect 45272 12288 45284 12297
rect 44600 12260 45284 12288
rect 44600 12248 44606 12260
rect 45272 12251 45284 12260
rect 45278 12248 45284 12251
rect 45336 12248 45342 12300
rect 47486 12288 47492 12300
rect 47447 12260 47492 12288
rect 47486 12248 47492 12260
rect 47544 12248 47550 12300
rect 4111 12192 4200 12220
rect 4111 12189 4123 12192
rect 4065 12183 4123 12189
rect 6454 12180 6460 12232
rect 6512 12220 6518 12232
rect 7193 12223 7251 12229
rect 7193 12220 7205 12223
rect 6512 12192 7205 12220
rect 6512 12180 6518 12192
rect 7193 12189 7205 12192
rect 7239 12189 7251 12223
rect 9674 12220 9680 12232
rect 9635 12192 9680 12220
rect 7193 12183 7251 12189
rect 9674 12180 9680 12192
rect 9732 12180 9738 12232
rect 18506 12180 18512 12232
rect 18564 12220 18570 12232
rect 18601 12223 18659 12229
rect 18601 12220 18613 12223
rect 18564 12192 18613 12220
rect 18564 12180 18570 12192
rect 18601 12189 18613 12192
rect 18647 12189 18659 12223
rect 20898 12220 20904 12232
rect 20859 12192 20904 12220
rect 18601 12183 18659 12189
rect 20898 12180 20904 12192
rect 20956 12180 20962 12232
rect 32122 12220 32128 12232
rect 32083 12192 32128 12220
rect 32122 12180 32128 12192
rect 32180 12180 32186 12232
rect 33870 12180 33876 12232
rect 33928 12220 33934 12232
rect 34425 12223 34483 12229
rect 34425 12220 34437 12223
rect 33928 12192 34437 12220
rect 33928 12180 33934 12192
rect 34425 12189 34437 12192
rect 34471 12220 34483 12223
rect 34606 12220 34612 12232
rect 34471 12192 34612 12220
rect 34471 12189 34483 12192
rect 34425 12183 34483 12189
rect 34606 12180 34612 12192
rect 34664 12180 34670 12232
rect 37274 12180 37280 12232
rect 37332 12220 37338 12232
rect 38657 12223 38715 12229
rect 38657 12220 38669 12223
rect 37332 12192 38669 12220
rect 37332 12180 37338 12192
rect 38657 12189 38669 12192
rect 38703 12220 38715 12223
rect 39022 12220 39028 12232
rect 38703 12192 39028 12220
rect 38703 12189 38715 12192
rect 38657 12183 38715 12189
rect 39022 12180 39028 12192
rect 39080 12180 39086 12232
rect 40034 12220 40040 12232
rect 39947 12192 40040 12220
rect 40034 12180 40040 12192
rect 40092 12180 40098 12232
rect 40218 12220 40224 12232
rect 40179 12192 40224 12220
rect 40218 12180 40224 12192
rect 40276 12180 40282 12232
rect 45002 12220 45008 12232
rect 44963 12192 45008 12220
rect 45002 12180 45008 12192
rect 45060 12180 45066 12232
rect 38102 12152 38108 12164
rect 38063 12124 38108 12152
rect 38102 12112 38108 12124
rect 38160 12112 38166 12164
rect 46382 12152 46388 12164
rect 46295 12124 46388 12152
rect 46382 12112 46388 12124
rect 46440 12152 46446 12164
rect 46937 12155 46995 12161
rect 46937 12152 46949 12155
rect 46440 12124 46949 12152
rect 46440 12112 46446 12124
rect 46937 12121 46949 12124
rect 46983 12121 46995 12155
rect 46937 12115 46995 12121
rect 2866 12084 2872 12096
rect 2827 12056 2872 12084
rect 2866 12044 2872 12056
rect 2924 12044 2930 12096
rect 3513 12087 3571 12093
rect 3513 12053 3525 12087
rect 3559 12084 3571 12087
rect 3878 12084 3884 12096
rect 3559 12056 3884 12084
rect 3559 12053 3571 12056
rect 3513 12047 3571 12053
rect 3878 12044 3884 12056
rect 3936 12044 3942 12096
rect 5534 12044 5540 12096
rect 5592 12084 5598 12096
rect 6641 12087 6699 12093
rect 6641 12084 6653 12087
rect 5592 12056 6653 12084
rect 5592 12044 5598 12056
rect 6641 12053 6653 12056
rect 6687 12053 6699 12087
rect 6641 12047 6699 12053
rect 11057 12087 11115 12093
rect 11057 12053 11069 12087
rect 11103 12084 11115 12087
rect 11238 12084 11244 12096
rect 11103 12056 11244 12084
rect 11103 12053 11115 12056
rect 11057 12047 11115 12053
rect 11238 12044 11244 12056
rect 11296 12044 11302 12096
rect 13630 12084 13636 12096
rect 13591 12056 13636 12084
rect 13630 12044 13636 12056
rect 13688 12044 13694 12096
rect 16022 12084 16028 12096
rect 15983 12056 16028 12084
rect 16022 12044 16028 12056
rect 16080 12044 16086 12096
rect 18049 12087 18107 12093
rect 18049 12053 18061 12087
rect 18095 12084 18107 12087
rect 18598 12084 18604 12096
rect 18095 12056 18604 12084
rect 18095 12053 18107 12056
rect 18049 12047 18107 12053
rect 18598 12044 18604 12056
rect 18656 12044 18662 12096
rect 19061 12087 19119 12093
rect 19061 12053 19073 12087
rect 19107 12084 19119 12087
rect 19242 12084 19248 12096
rect 19107 12056 19248 12084
rect 19107 12053 19119 12056
rect 19061 12047 19119 12053
rect 19242 12044 19248 12056
rect 19300 12044 19306 12096
rect 19978 12044 19984 12096
rect 20036 12084 20042 12096
rect 20438 12084 20444 12096
rect 20036 12056 20444 12084
rect 20036 12044 20042 12056
rect 20438 12044 20444 12056
rect 20496 12044 20502 12096
rect 23566 12044 23572 12096
rect 23624 12084 23630 12096
rect 23661 12087 23719 12093
rect 23661 12084 23673 12087
rect 23624 12056 23673 12084
rect 23624 12044 23630 12056
rect 23661 12053 23673 12056
rect 23707 12053 23719 12087
rect 23661 12047 23719 12053
rect 33226 12044 33232 12096
rect 33284 12084 33290 12096
rect 34057 12087 34115 12093
rect 34057 12084 34069 12087
rect 33284 12056 34069 12084
rect 33284 12044 33290 12056
rect 34057 12053 34069 12056
rect 34103 12053 34115 12087
rect 39666 12084 39672 12096
rect 39627 12056 39672 12084
rect 34057 12047 34115 12053
rect 39666 12044 39672 12056
rect 39724 12044 39730 12096
rect 40862 12084 40868 12096
rect 40823 12056 40868 12084
rect 40862 12044 40868 12056
rect 40920 12044 40926 12096
rect 1104 11994 48852 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 34966 11994
rect 35018 11942 35030 11994
rect 35082 11942 35094 11994
rect 35146 11942 35158 11994
rect 35210 11942 48852 11994
rect 1104 11920 48852 11942
rect 1486 11840 1492 11892
rect 1544 11880 1550 11892
rect 1581 11883 1639 11889
rect 1581 11880 1593 11883
rect 1544 11852 1593 11880
rect 1544 11840 1550 11852
rect 1581 11849 1593 11852
rect 1627 11849 1639 11883
rect 2866 11880 2872 11892
rect 2827 11852 2872 11880
rect 1581 11843 1639 11849
rect 2866 11840 2872 11852
rect 2924 11840 2930 11892
rect 3970 11840 3976 11892
rect 4028 11880 4034 11892
rect 4341 11883 4399 11889
rect 4341 11880 4353 11883
rect 4028 11852 4353 11880
rect 4028 11840 4034 11852
rect 4341 11849 4353 11852
rect 4387 11849 4399 11883
rect 4798 11880 4804 11892
rect 4759 11852 4804 11880
rect 4341 11843 4399 11849
rect 4798 11840 4804 11852
rect 4856 11840 4862 11892
rect 5534 11880 5540 11892
rect 5495 11852 5540 11880
rect 5534 11840 5540 11852
rect 5592 11840 5598 11892
rect 6273 11883 6331 11889
rect 6273 11849 6285 11883
rect 6319 11880 6331 11883
rect 6914 11880 6920 11892
rect 6319 11852 6920 11880
rect 6319 11849 6331 11852
rect 6273 11843 6331 11849
rect 6914 11840 6920 11852
rect 6972 11840 6978 11892
rect 9950 11840 9956 11892
rect 10008 11880 10014 11892
rect 10045 11883 10103 11889
rect 10045 11880 10057 11883
rect 10008 11852 10057 11880
rect 10008 11840 10014 11852
rect 10045 11849 10057 11852
rect 10091 11849 10103 11883
rect 10045 11843 10103 11849
rect 16117 11883 16175 11889
rect 16117 11849 16129 11883
rect 16163 11880 16175 11883
rect 17862 11880 17868 11892
rect 16163 11852 17868 11880
rect 16163 11849 16175 11852
rect 16117 11843 16175 11849
rect 17862 11840 17868 11852
rect 17920 11840 17926 11892
rect 18230 11880 18236 11892
rect 18191 11852 18236 11880
rect 18230 11840 18236 11852
rect 18288 11840 18294 11892
rect 21358 11880 21364 11892
rect 21319 11852 21364 11880
rect 21358 11840 21364 11852
rect 21416 11840 21422 11892
rect 25038 11880 25044 11892
rect 24999 11852 25044 11880
rect 25038 11840 25044 11852
rect 25096 11840 25102 11892
rect 28350 11880 28356 11892
rect 28311 11852 28356 11880
rect 28350 11840 28356 11852
rect 28408 11840 28414 11892
rect 28626 11840 28632 11892
rect 28684 11880 28690 11892
rect 28721 11883 28779 11889
rect 28721 11880 28733 11883
rect 28684 11852 28733 11880
rect 28684 11840 28690 11852
rect 28721 11849 28733 11852
rect 28767 11849 28779 11883
rect 32122 11880 32128 11892
rect 32083 11852 32128 11880
rect 28721 11843 28779 11849
rect 32122 11840 32128 11852
rect 32180 11840 32186 11892
rect 32585 11883 32643 11889
rect 32585 11849 32597 11883
rect 32631 11880 32643 11883
rect 32674 11880 32680 11892
rect 32631 11852 32680 11880
rect 32631 11849 32643 11852
rect 32585 11843 32643 11849
rect 32674 11840 32680 11852
rect 32732 11840 32738 11892
rect 34238 11880 34244 11892
rect 34199 11852 34244 11880
rect 34238 11840 34244 11852
rect 34296 11840 34302 11892
rect 34606 11880 34612 11892
rect 34567 11852 34612 11880
rect 34606 11840 34612 11852
rect 34664 11840 34670 11892
rect 35161 11883 35219 11889
rect 35161 11849 35173 11883
rect 35207 11880 35219 11883
rect 35250 11880 35256 11892
rect 35207 11852 35256 11880
rect 35207 11849 35219 11852
rect 35161 11843 35219 11849
rect 35250 11840 35256 11852
rect 35308 11840 35314 11892
rect 39022 11880 39028 11892
rect 38983 11852 39028 11880
rect 39022 11840 39028 11852
rect 39080 11840 39086 11892
rect 39669 11883 39727 11889
rect 39669 11849 39681 11883
rect 39715 11880 39727 11883
rect 39758 11880 39764 11892
rect 39715 11852 39764 11880
rect 39715 11849 39727 11852
rect 39669 11843 39727 11849
rect 39758 11840 39764 11852
rect 39816 11840 39822 11892
rect 40034 11880 40040 11892
rect 39995 11852 40040 11880
rect 40034 11840 40040 11852
rect 40092 11840 40098 11892
rect 45278 11840 45284 11892
rect 45336 11880 45342 11892
rect 45373 11883 45431 11889
rect 45373 11880 45385 11883
rect 45336 11852 45385 11880
rect 45336 11840 45342 11852
rect 45373 11849 45385 11852
rect 45419 11849 45431 11883
rect 47486 11880 47492 11892
rect 47447 11852 47492 11880
rect 45373 11843 45431 11849
rect 47486 11840 47492 11852
rect 47544 11840 47550 11892
rect 1857 11815 1915 11821
rect 1857 11781 1869 11815
rect 1903 11812 1915 11815
rect 2774 11812 2780 11824
rect 1903 11784 2780 11812
rect 1903 11781 1915 11784
rect 1857 11775 1915 11781
rect 2774 11772 2780 11784
rect 2832 11772 2838 11824
rect 2317 11747 2375 11753
rect 2317 11713 2329 11747
rect 2363 11744 2375 11747
rect 2406 11744 2412 11756
rect 2363 11716 2412 11744
rect 2363 11713 2375 11716
rect 2317 11707 2375 11713
rect 2406 11704 2412 11716
rect 2464 11744 2470 11756
rect 2884 11744 2912 11840
rect 3418 11812 3424 11824
rect 3379 11784 3424 11812
rect 3418 11772 3424 11784
rect 3476 11772 3482 11824
rect 2464 11716 2912 11744
rect 2464 11704 2470 11716
rect 5552 11676 5580 11840
rect 6641 11815 6699 11821
rect 6641 11781 6653 11815
rect 6687 11812 6699 11815
rect 7098 11812 7104 11824
rect 6687 11784 7104 11812
rect 6687 11781 6699 11784
rect 6641 11775 6699 11781
rect 7098 11772 7104 11784
rect 7156 11812 7162 11824
rect 7561 11815 7619 11821
rect 7561 11812 7573 11815
rect 7156 11784 7573 11812
rect 7156 11772 7162 11784
rect 7561 11781 7573 11784
rect 7607 11781 7619 11815
rect 7561 11775 7619 11781
rect 11425 11815 11483 11821
rect 11425 11781 11437 11815
rect 11471 11812 11483 11815
rect 12434 11812 12440 11824
rect 11471 11784 12440 11812
rect 11471 11781 11483 11784
rect 11425 11775 11483 11781
rect 12434 11772 12440 11784
rect 12492 11772 12498 11824
rect 20898 11772 20904 11824
rect 20956 11812 20962 11824
rect 20993 11815 21051 11821
rect 20993 11812 21005 11815
rect 20956 11784 21005 11812
rect 20956 11772 20962 11784
rect 20993 11781 21005 11784
rect 21039 11812 21051 11815
rect 22186 11812 22192 11824
rect 21039 11784 22192 11812
rect 21039 11781 21051 11784
rect 20993 11775 21051 11781
rect 22186 11772 22192 11784
rect 22244 11812 22250 11824
rect 23385 11815 23443 11821
rect 23385 11812 23397 11815
rect 22244 11784 23397 11812
rect 22244 11772 22250 11784
rect 23385 11781 23397 11784
rect 23431 11812 23443 11815
rect 23431 11784 23704 11812
rect 23431 11781 23443 11784
rect 23385 11775 23443 11781
rect 23676 11756 23704 11784
rect 34514 11772 34520 11824
rect 34572 11812 34578 11824
rect 35621 11815 35679 11821
rect 35621 11812 35633 11815
rect 34572 11784 35633 11812
rect 34572 11772 34578 11784
rect 35621 11781 35633 11784
rect 35667 11781 35679 11815
rect 35621 11775 35679 11781
rect 7650 11704 7656 11756
rect 7708 11744 7714 11756
rect 8021 11747 8079 11753
rect 8021 11744 8033 11747
rect 7708 11716 8033 11744
rect 7708 11704 7714 11716
rect 8021 11713 8033 11716
rect 8067 11744 8079 11747
rect 8754 11744 8760 11756
rect 8067 11716 8760 11744
rect 8067 11713 8079 11716
rect 8021 11707 8079 11713
rect 8754 11704 8760 11716
rect 8812 11704 8818 11756
rect 9674 11704 9680 11756
rect 9732 11744 9738 11756
rect 9769 11747 9827 11753
rect 9769 11744 9781 11747
rect 9732 11716 9781 11744
rect 9732 11704 9738 11716
rect 9769 11713 9781 11716
rect 9815 11744 9827 11747
rect 11882 11744 11888 11756
rect 9815 11716 11888 11744
rect 9815 11713 9827 11716
rect 9769 11707 9827 11713
rect 11882 11704 11888 11716
rect 11940 11744 11946 11756
rect 13357 11747 13415 11753
rect 13357 11744 13369 11747
rect 11940 11716 13369 11744
rect 11940 11704 11946 11716
rect 13357 11713 13369 11716
rect 13403 11744 13415 11747
rect 13538 11744 13544 11756
rect 13403 11716 13544 11744
rect 13403 11713 13415 11716
rect 13357 11707 13415 11713
rect 13538 11704 13544 11716
rect 13596 11704 13602 11756
rect 16022 11704 16028 11756
rect 16080 11744 16086 11756
rect 16669 11747 16727 11753
rect 16669 11744 16681 11747
rect 16080 11716 16681 11744
rect 16080 11704 16086 11716
rect 16669 11713 16681 11716
rect 16715 11713 16727 11747
rect 23658 11744 23664 11756
rect 23571 11716 23664 11744
rect 16669 11707 16727 11713
rect 23658 11704 23664 11716
rect 23716 11704 23722 11756
rect 37553 11747 37611 11753
rect 37553 11713 37565 11747
rect 37599 11744 37611 11747
rect 37642 11744 37648 11756
rect 37599 11716 37648 11744
rect 37599 11713 37611 11716
rect 37553 11707 37611 11713
rect 37642 11704 37648 11716
rect 37700 11704 37706 11756
rect 5629 11679 5687 11685
rect 5629 11676 5641 11679
rect 5552 11648 5641 11676
rect 5629 11645 5641 11648
rect 5675 11645 5687 11679
rect 5629 11639 5687 11645
rect 11146 11636 11152 11688
rect 11204 11676 11210 11688
rect 11241 11679 11299 11685
rect 11241 11676 11253 11679
rect 11204 11648 11253 11676
rect 11204 11636 11210 11648
rect 11241 11645 11253 11648
rect 11287 11676 11299 11679
rect 11793 11679 11851 11685
rect 11793 11676 11805 11679
rect 11287 11648 11805 11676
rect 11287 11645 11299 11648
rect 11241 11639 11299 11645
rect 11793 11645 11805 11648
rect 11839 11676 11851 11679
rect 12342 11676 12348 11688
rect 11839 11648 12348 11676
rect 11839 11645 11851 11648
rect 11793 11639 11851 11645
rect 12342 11636 12348 11648
rect 12400 11636 12406 11688
rect 13630 11636 13636 11688
rect 13688 11676 13694 11688
rect 13797 11679 13855 11685
rect 13797 11676 13809 11679
rect 13688 11648 13809 11676
rect 13688 11636 13694 11648
rect 13797 11645 13809 11648
rect 13843 11645 13855 11679
rect 18969 11679 19027 11685
rect 18969 11676 18981 11679
rect 13797 11639 13855 11645
rect 15488 11648 16620 11676
rect 2314 11608 2320 11620
rect 2275 11580 2320 11608
rect 2314 11568 2320 11580
rect 2372 11568 2378 11620
rect 2409 11611 2467 11617
rect 2409 11577 2421 11611
rect 2455 11608 2467 11611
rect 2682 11608 2688 11620
rect 2455 11580 2688 11608
rect 2455 11577 2467 11580
rect 2409 11571 2467 11577
rect 2682 11568 2688 11580
rect 2740 11568 2746 11620
rect 2774 11568 2780 11620
rect 2832 11608 2838 11620
rect 3697 11611 3755 11617
rect 3697 11608 3709 11611
rect 2832 11580 3709 11608
rect 2832 11568 2838 11580
rect 3697 11577 3709 11580
rect 3743 11577 3755 11611
rect 3970 11608 3976 11620
rect 3931 11580 3976 11608
rect 3697 11571 3755 11577
rect 3970 11568 3976 11580
rect 4028 11568 4034 11620
rect 7190 11568 7196 11620
rect 7248 11608 7254 11620
rect 7834 11608 7840 11620
rect 7248 11580 7840 11608
rect 7248 11568 7254 11580
rect 7834 11568 7840 11580
rect 7892 11608 7898 11620
rect 8113 11611 8171 11617
rect 8113 11608 8125 11611
rect 7892 11580 8125 11608
rect 7892 11568 7898 11580
rect 8113 11577 8125 11580
rect 8159 11577 8171 11611
rect 8113 11571 8171 11577
rect 15488 11552 15516 11648
rect 16592 11617 16620 11648
rect 18800 11648 18981 11676
rect 16393 11611 16451 11617
rect 16393 11577 16405 11611
rect 16439 11577 16451 11611
rect 16393 11571 16451 11577
rect 16577 11611 16635 11617
rect 16577 11577 16589 11611
rect 16623 11577 16635 11611
rect 16577 11571 16635 11577
rect 3237 11543 3295 11549
rect 3237 11509 3249 11543
rect 3283 11540 3295 11543
rect 3881 11543 3939 11549
rect 3881 11540 3893 11543
rect 3283 11512 3893 11540
rect 3283 11509 3295 11512
rect 3237 11503 3295 11509
rect 3881 11509 3893 11512
rect 3927 11540 3939 11543
rect 4062 11540 4068 11552
rect 3927 11512 4068 11540
rect 3927 11509 3939 11512
rect 3881 11503 3939 11509
rect 4062 11500 4068 11512
rect 4120 11500 4126 11552
rect 5810 11540 5816 11552
rect 5771 11512 5816 11540
rect 5810 11500 5816 11512
rect 5868 11500 5874 11552
rect 7377 11543 7435 11549
rect 7377 11509 7389 11543
rect 7423 11540 7435 11543
rect 8021 11543 8079 11549
rect 8021 11540 8033 11543
rect 7423 11512 8033 11540
rect 7423 11509 7435 11512
rect 7377 11503 7435 11509
rect 8021 11509 8033 11512
rect 8067 11540 8079 11543
rect 8386 11540 8392 11552
rect 8067 11512 8392 11540
rect 8067 11509 8079 11512
rect 8021 11503 8079 11509
rect 8386 11500 8392 11512
rect 8444 11500 8450 11552
rect 14918 11540 14924 11552
rect 14879 11512 14924 11540
rect 14918 11500 14924 11512
rect 14976 11500 14982 11552
rect 15470 11540 15476 11552
rect 15431 11512 15476 11540
rect 15470 11500 15476 11512
rect 15528 11500 15534 11552
rect 15838 11540 15844 11552
rect 15799 11512 15844 11540
rect 15838 11500 15844 11512
rect 15896 11540 15902 11552
rect 16408 11540 16436 11571
rect 15896 11512 16436 11540
rect 15896 11500 15902 11512
rect 18138 11500 18144 11552
rect 18196 11540 18202 11552
rect 18800 11549 18828 11648
rect 18969 11645 18981 11648
rect 19015 11645 19027 11679
rect 18969 11639 19027 11645
rect 35437 11679 35495 11685
rect 35437 11645 35449 11679
rect 35483 11676 35495 11679
rect 40773 11679 40831 11685
rect 35483 11648 36032 11676
rect 35483 11645 35495 11648
rect 35437 11639 35495 11645
rect 19242 11617 19248 11620
rect 19236 11608 19248 11617
rect 19203 11580 19248 11608
rect 19236 11571 19248 11580
rect 19242 11568 19248 11571
rect 19300 11568 19306 11620
rect 23566 11568 23572 11620
rect 23624 11608 23630 11620
rect 23906 11611 23964 11617
rect 23906 11608 23918 11611
rect 23624 11580 23918 11608
rect 23624 11568 23630 11580
rect 23906 11577 23918 11580
rect 23952 11577 23964 11611
rect 23906 11571 23964 11577
rect 18785 11543 18843 11549
rect 18785 11540 18797 11543
rect 18196 11512 18797 11540
rect 18196 11500 18202 11512
rect 18785 11509 18797 11512
rect 18831 11509 18843 11543
rect 18785 11503 18843 11509
rect 20349 11543 20407 11549
rect 20349 11509 20361 11543
rect 20395 11540 20407 11543
rect 20622 11540 20628 11552
rect 20395 11512 20628 11540
rect 20395 11509 20407 11512
rect 20349 11503 20407 11509
rect 20622 11500 20628 11512
rect 20680 11500 20686 11552
rect 36004 11549 36032 11648
rect 40773 11645 40785 11679
rect 40819 11676 40831 11679
rect 41509 11679 41567 11685
rect 41509 11676 41521 11679
rect 40819 11648 41521 11676
rect 40819 11645 40831 11648
rect 40773 11639 40831 11645
rect 41509 11645 41521 11648
rect 41555 11676 41567 11679
rect 42702 11676 42708 11688
rect 41555 11648 42708 11676
rect 41555 11645 41567 11648
rect 41509 11639 41567 11645
rect 42702 11636 42708 11648
rect 42760 11636 42766 11688
rect 37185 11611 37243 11617
rect 37185 11577 37197 11611
rect 37231 11608 37243 11611
rect 37890 11611 37948 11617
rect 37890 11608 37902 11611
rect 37231 11580 37902 11608
rect 37231 11577 37243 11580
rect 37185 11571 37243 11577
rect 37890 11577 37902 11580
rect 37936 11608 37948 11611
rect 40862 11608 40868 11620
rect 37936 11580 40868 11608
rect 37936 11577 37948 11580
rect 37890 11571 37948 11577
rect 40862 11568 40868 11580
rect 40920 11608 40926 11620
rect 40957 11611 41015 11617
rect 40957 11608 40969 11611
rect 40920 11580 40969 11608
rect 40920 11568 40926 11580
rect 40957 11577 40969 11580
rect 41003 11577 41015 11611
rect 40957 11571 41015 11577
rect 35989 11543 36047 11549
rect 35989 11509 36001 11543
rect 36035 11540 36047 11543
rect 36078 11540 36084 11552
rect 36035 11512 36084 11540
rect 36035 11509 36047 11512
rect 35989 11503 36047 11509
rect 36078 11500 36084 11512
rect 36136 11500 36142 11552
rect 41138 11540 41144 11552
rect 41099 11512 41144 11540
rect 41138 11500 41144 11512
rect 41196 11500 41202 11552
rect 41506 11500 41512 11552
rect 41564 11540 41570 11552
rect 41785 11543 41843 11549
rect 41785 11540 41797 11543
rect 41564 11512 41797 11540
rect 41564 11500 41570 11512
rect 41785 11509 41797 11512
rect 41831 11509 41843 11543
rect 41785 11503 41843 11509
rect 44174 11500 44180 11552
rect 44232 11540 44238 11552
rect 45002 11540 45008 11552
rect 44232 11512 45008 11540
rect 44232 11500 44238 11512
rect 45002 11500 45008 11512
rect 45060 11500 45066 11552
rect 1104 11450 48852 11472
rect 1104 11398 19606 11450
rect 19658 11398 19670 11450
rect 19722 11398 19734 11450
rect 19786 11398 19798 11450
rect 19850 11398 48852 11450
rect 1104 11376 48852 11398
rect 2406 11336 2412 11348
rect 2367 11308 2412 11336
rect 2406 11296 2412 11308
rect 2464 11296 2470 11348
rect 2682 11336 2688 11348
rect 2643 11308 2688 11336
rect 2682 11296 2688 11308
rect 2740 11296 2746 11348
rect 2774 11296 2780 11348
rect 2832 11336 2838 11348
rect 5442 11345 5448 11348
rect 3329 11339 3387 11345
rect 3329 11336 3341 11339
rect 2832 11308 3341 11336
rect 2832 11296 2838 11308
rect 3329 11305 3341 11308
rect 3375 11305 3387 11339
rect 3329 11299 3387 11305
rect 5435 11339 5448 11345
rect 5435 11305 5447 11339
rect 5500 11336 5506 11348
rect 5500 11308 5535 11336
rect 5435 11299 5448 11305
rect 5442 11296 5448 11299
rect 5500 11296 5506 11308
rect 5810 11296 5816 11348
rect 5868 11336 5874 11348
rect 5905 11339 5963 11345
rect 5905 11336 5917 11339
rect 5868 11308 5917 11336
rect 5868 11296 5874 11308
rect 5905 11305 5917 11308
rect 5951 11305 5963 11339
rect 5905 11299 5963 11305
rect 7561 11339 7619 11345
rect 7561 11305 7573 11339
rect 7607 11336 7619 11339
rect 7650 11336 7656 11348
rect 7607 11308 7656 11336
rect 7607 11305 7619 11308
rect 7561 11299 7619 11305
rect 7650 11296 7656 11308
rect 7708 11296 7714 11348
rect 12713 11339 12771 11345
rect 12713 11305 12725 11339
rect 12759 11336 12771 11339
rect 13078 11336 13084 11348
rect 12759 11308 13084 11336
rect 12759 11305 12771 11308
rect 12713 11299 12771 11305
rect 13078 11296 13084 11308
rect 13136 11336 13142 11348
rect 13357 11339 13415 11345
rect 13357 11336 13369 11339
rect 13136 11308 13369 11336
rect 13136 11296 13142 11308
rect 13357 11305 13369 11308
rect 13403 11336 13415 11339
rect 13630 11336 13636 11348
rect 13403 11308 13636 11336
rect 13403 11305 13415 11308
rect 13357 11299 13415 11305
rect 13630 11296 13636 11308
rect 13688 11296 13694 11348
rect 14185 11339 14243 11345
rect 14185 11305 14197 11339
rect 14231 11336 14243 11339
rect 15838 11336 15844 11348
rect 14231 11308 15844 11336
rect 14231 11305 14243 11308
rect 14185 11299 14243 11305
rect 15838 11296 15844 11308
rect 15896 11296 15902 11348
rect 37274 11296 37280 11348
rect 37332 11336 37338 11348
rect 37461 11339 37519 11345
rect 37461 11336 37473 11339
rect 37332 11308 37473 11336
rect 37332 11296 37338 11308
rect 37461 11305 37473 11308
rect 37507 11305 37519 11339
rect 37461 11299 37519 11305
rect 37921 11339 37979 11345
rect 37921 11305 37933 11339
rect 37967 11336 37979 11339
rect 38378 11336 38384 11348
rect 37967 11308 38384 11336
rect 37967 11305 37979 11308
rect 37921 11299 37979 11305
rect 38378 11296 38384 11308
rect 38436 11296 38442 11348
rect 38562 11296 38568 11348
rect 38620 11336 38626 11348
rect 38657 11339 38715 11345
rect 38657 11336 38669 11339
rect 38620 11308 38669 11336
rect 38620 11296 38626 11308
rect 38657 11305 38669 11308
rect 38703 11336 38715 11339
rect 39025 11339 39083 11345
rect 39025 11336 39037 11339
rect 38703 11308 39037 11336
rect 38703 11305 38715 11308
rect 38657 11299 38715 11305
rect 39025 11305 39037 11308
rect 39071 11305 39083 11339
rect 39025 11299 39083 11305
rect 40862 11296 40868 11348
rect 40920 11336 40926 11348
rect 42061 11339 42119 11345
rect 42061 11336 42073 11339
rect 40920 11308 42073 11336
rect 40920 11296 40926 11308
rect 42061 11305 42073 11308
rect 42107 11305 42119 11339
rect 42061 11299 42119 11305
rect 1673 11271 1731 11277
rect 1673 11237 1685 11271
rect 1719 11268 1731 11271
rect 2041 11271 2099 11277
rect 2041 11268 2053 11271
rect 1719 11240 2053 11268
rect 1719 11237 1731 11240
rect 1673 11231 1731 11237
rect 2041 11237 2053 11240
rect 2087 11268 2099 11271
rect 2314 11268 2320 11280
rect 2087 11240 2320 11268
rect 2087 11237 2099 11240
rect 2041 11231 2099 11237
rect 2314 11228 2320 11240
rect 2372 11228 2378 11280
rect 11882 11268 11888 11280
rect 11348 11240 11888 11268
rect 3418 11160 3424 11212
rect 3476 11200 3482 11212
rect 4249 11203 4307 11209
rect 4249 11200 4261 11203
rect 3476 11172 4261 11200
rect 3476 11160 3482 11172
rect 4249 11169 4261 11172
rect 4295 11200 4307 11203
rect 4614 11200 4620 11212
rect 4295 11172 4620 11200
rect 4295 11169 4307 11172
rect 4249 11163 4307 11169
rect 4614 11160 4620 11172
rect 4672 11160 4678 11212
rect 10229 11203 10287 11209
rect 10229 11169 10241 11203
rect 10275 11200 10287 11203
rect 10686 11200 10692 11212
rect 10275 11172 10692 11200
rect 10275 11169 10287 11172
rect 10229 11163 10287 11169
rect 10686 11160 10692 11172
rect 10744 11160 10750 11212
rect 11348 11209 11376 11240
rect 11882 11228 11888 11240
rect 11940 11228 11946 11280
rect 14918 11228 14924 11280
rect 14976 11268 14982 11280
rect 15924 11271 15982 11277
rect 15924 11268 15936 11271
rect 14976 11240 15936 11268
rect 14976 11228 14982 11240
rect 15924 11237 15936 11240
rect 15970 11268 15982 11271
rect 16022 11268 16028 11280
rect 15970 11240 16028 11268
rect 15970 11237 15982 11240
rect 15924 11231 15982 11237
rect 16022 11228 16028 11240
rect 16080 11228 16086 11280
rect 26234 11228 26240 11280
rect 26292 11268 26298 11280
rect 26872 11271 26930 11277
rect 26872 11268 26884 11271
rect 26292 11240 26884 11268
rect 26292 11228 26298 11240
rect 26872 11237 26884 11240
rect 26918 11268 26930 11271
rect 27522 11268 27528 11280
rect 26918 11240 27528 11268
rect 26918 11237 26930 11240
rect 26872 11231 26930 11237
rect 27522 11228 27528 11240
rect 27580 11228 27586 11280
rect 33686 11228 33692 11280
rect 33744 11268 33750 11280
rect 34118 11271 34176 11277
rect 34118 11268 34130 11271
rect 33744 11240 34130 11268
rect 33744 11228 33750 11240
rect 34118 11237 34130 11240
rect 34164 11268 34176 11271
rect 34238 11268 34244 11280
rect 34164 11240 34244 11268
rect 34164 11237 34176 11240
rect 34118 11231 34176 11237
rect 34238 11228 34244 11240
rect 34296 11228 34302 11280
rect 41322 11268 41328 11280
rect 40696 11240 41328 11268
rect 11606 11209 11612 11212
rect 11333 11203 11391 11209
rect 11333 11169 11345 11203
rect 11379 11169 11391 11203
rect 11600 11200 11612 11209
rect 11567 11172 11612 11200
rect 11333 11163 11391 11169
rect 11600 11163 11612 11172
rect 11606 11160 11612 11163
rect 11664 11160 11670 11212
rect 13538 11160 13544 11212
rect 13596 11200 13602 11212
rect 15654 11200 15660 11212
rect 13596 11172 15660 11200
rect 13596 11160 13602 11172
rect 15654 11160 15660 11172
rect 15712 11160 15718 11212
rect 18414 11209 18420 11212
rect 18049 11203 18107 11209
rect 18049 11169 18061 11203
rect 18095 11200 18107 11203
rect 18408 11200 18420 11209
rect 18095 11172 18420 11200
rect 18095 11169 18107 11172
rect 18049 11163 18107 11169
rect 18408 11163 18420 11172
rect 5813 11135 5871 11141
rect 5813 11132 5825 11135
rect 5000 11104 5825 11132
rect 5000 11008 5028 11104
rect 5813 11101 5825 11104
rect 5859 11101 5871 11135
rect 5813 11095 5871 11101
rect 5902 11092 5908 11144
rect 5960 11132 5966 11144
rect 5997 11135 6055 11141
rect 5997 11132 6009 11135
rect 5960 11104 6009 11132
rect 5960 11092 5966 11104
rect 5997 11101 6009 11104
rect 6043 11101 6055 11135
rect 5997 11095 6055 11101
rect 5261 11067 5319 11073
rect 5261 11033 5273 11067
rect 5307 11064 5319 11067
rect 5534 11064 5540 11076
rect 5307 11036 5540 11064
rect 5307 11033 5319 11036
rect 5261 11027 5319 11033
rect 5534 11024 5540 11036
rect 5592 11024 5598 11076
rect 6454 11064 6460 11076
rect 5644 11036 6460 11064
rect 4433 10999 4491 11005
rect 4433 10965 4445 10999
rect 4479 10996 4491 10999
rect 4982 10996 4988 11008
rect 4479 10968 4988 10996
rect 4479 10965 4491 10968
rect 4433 10959 4491 10965
rect 4982 10956 4988 10968
rect 5040 10956 5046 11008
rect 5442 10956 5448 11008
rect 5500 10996 5506 11008
rect 5644 10996 5672 11036
rect 6454 11024 6460 11036
rect 6512 11064 6518 11076
rect 7466 11064 7472 11076
rect 6512 11036 7472 11064
rect 6512 11024 6518 11036
rect 7466 11024 7472 11036
rect 7524 11024 7530 11076
rect 10410 11064 10416 11076
rect 10371 11036 10416 11064
rect 10410 11024 10416 11036
rect 10468 11024 10474 11076
rect 17037 11067 17095 11073
rect 17037 11033 17049 11067
rect 17083 11064 17095 11067
rect 18064 11064 18092 11163
rect 18414 11160 18420 11163
rect 18472 11160 18478 11212
rect 22445 11203 22503 11209
rect 22445 11200 22457 11203
rect 22112 11172 22457 11200
rect 18138 11092 18144 11144
rect 18196 11132 18202 11144
rect 18196 11104 18289 11132
rect 18196 11092 18202 11104
rect 17083 11036 18092 11064
rect 17083 11033 17095 11036
rect 17037 11027 17095 11033
rect 5500 10968 5672 10996
rect 6917 10999 6975 11005
rect 5500 10956 5506 10968
rect 6917 10965 6929 10999
rect 6963 10996 6975 10999
rect 7190 10996 7196 11008
rect 6963 10968 7196 10996
rect 6963 10965 6975 10968
rect 6917 10959 6975 10965
rect 7190 10956 7196 10968
rect 7248 10956 7254 11008
rect 7834 10996 7840 11008
rect 7795 10968 7840 10996
rect 7834 10956 7840 10968
rect 7892 10956 7898 11008
rect 8478 10996 8484 11008
rect 8439 10968 8484 10996
rect 8478 10956 8484 10968
rect 8536 10956 8542 11008
rect 17770 10956 17776 11008
rect 17828 10996 17834 11008
rect 18156 10996 18184 11092
rect 19242 11064 19248 11076
rect 19076 11036 19248 11064
rect 17828 10968 18184 10996
rect 17828 10956 17834 10968
rect 18506 10956 18512 11008
rect 18564 10996 18570 11008
rect 19076 10996 19104 11036
rect 19242 11024 19248 11036
rect 19300 11064 19306 11076
rect 19521 11067 19579 11073
rect 19521 11064 19533 11067
rect 19300 11036 19533 11064
rect 19300 11024 19306 11036
rect 19521 11033 19533 11036
rect 19567 11033 19579 11067
rect 19521 11027 19579 11033
rect 20441 11067 20499 11073
rect 20441 11033 20453 11067
rect 20487 11064 20499 11067
rect 20898 11064 20904 11076
rect 20487 11036 20904 11064
rect 20487 11033 20499 11036
rect 20441 11027 20499 11033
rect 20898 11024 20904 11036
rect 20956 11024 20962 11076
rect 18564 10968 19104 10996
rect 18564 10956 18570 10968
rect 20714 10956 20720 11008
rect 20772 10996 20778 11008
rect 22112 10996 22140 11172
rect 22445 11169 22457 11172
rect 22491 11169 22503 11203
rect 26602 11200 26608 11212
rect 26515 11172 26608 11200
rect 22445 11163 22503 11169
rect 26602 11160 26608 11172
rect 26660 11200 26666 11212
rect 27154 11200 27160 11212
rect 26660 11172 27160 11200
rect 26660 11160 26666 11172
rect 27154 11160 27160 11172
rect 27212 11160 27218 11212
rect 28350 11160 28356 11212
rect 28408 11200 28414 11212
rect 29089 11203 29147 11209
rect 29089 11200 29101 11203
rect 28408 11172 29101 11200
rect 28408 11160 28414 11172
rect 29089 11169 29101 11172
rect 29135 11169 29147 11203
rect 29089 11163 29147 11169
rect 29356 11203 29414 11209
rect 29356 11169 29368 11203
rect 29402 11200 29414 11203
rect 29638 11200 29644 11212
rect 29402 11172 29644 11200
rect 29402 11169 29414 11172
rect 29356 11163 29414 11169
rect 29638 11160 29644 11172
rect 29696 11160 29702 11212
rect 33873 11203 33931 11209
rect 33873 11169 33885 11203
rect 33919 11200 33931 11203
rect 33962 11200 33968 11212
rect 33919 11172 33968 11200
rect 33919 11169 33931 11172
rect 33873 11163 33931 11169
rect 33962 11160 33968 11172
rect 34020 11160 34026 11212
rect 37734 11200 37740 11212
rect 37695 11172 37740 11200
rect 37734 11160 37740 11172
rect 37792 11160 37798 11212
rect 38841 11203 38899 11209
rect 38841 11169 38853 11203
rect 38887 11200 38899 11203
rect 39666 11200 39672 11212
rect 38887 11172 39672 11200
rect 38887 11169 38899 11172
rect 38841 11163 38899 11169
rect 39666 11160 39672 11172
rect 39724 11160 39730 11212
rect 40696 11209 40724 11240
rect 41322 11228 41328 11240
rect 41380 11228 41386 11280
rect 43622 11228 43628 11280
rect 43680 11268 43686 11280
rect 43901 11271 43959 11277
rect 43901 11268 43913 11271
rect 43680 11240 43913 11268
rect 43680 11228 43686 11240
rect 43901 11237 43913 11240
rect 43947 11237 43959 11271
rect 43901 11231 43959 11237
rect 40954 11209 40960 11212
rect 40681 11203 40739 11209
rect 40681 11169 40693 11203
rect 40727 11169 40739 11203
rect 40681 11163 40739 11169
rect 40948 11163 40960 11209
rect 41012 11200 41018 11212
rect 41012 11172 41048 11200
rect 40954 11160 40960 11163
rect 41012 11160 41018 11172
rect 43070 11160 43076 11212
rect 43128 11200 43134 11212
rect 43717 11203 43775 11209
rect 43717 11200 43729 11203
rect 43128 11172 43729 11200
rect 43128 11160 43134 11172
rect 43717 11169 43729 11172
rect 43763 11169 43775 11203
rect 43717 11163 43775 11169
rect 22186 11092 22192 11144
rect 22244 11132 22250 11144
rect 43993 11135 44051 11141
rect 22244 11104 22289 11132
rect 22244 11092 22250 11104
rect 43993 11101 44005 11135
rect 44039 11101 44051 11135
rect 43993 11095 44051 11101
rect 23566 11064 23572 11076
rect 23400 11036 23572 11064
rect 22186 10996 22192 11008
rect 20772 10968 22192 10996
rect 20772 10956 20778 10968
rect 22186 10956 22192 10968
rect 22244 10956 22250 11008
rect 23106 10956 23112 11008
rect 23164 10996 23170 11008
rect 23400 10996 23428 11036
rect 23566 11024 23572 11036
rect 23624 11024 23630 11076
rect 27982 11064 27988 11076
rect 27943 11036 27988 11064
rect 27982 11024 27988 11036
rect 28040 11024 28046 11076
rect 30466 11064 30472 11076
rect 30427 11036 30472 11064
rect 30466 11024 30472 11036
rect 30524 11024 30530 11076
rect 39853 11067 39911 11073
rect 39853 11033 39865 11067
rect 39899 11064 39911 11067
rect 40218 11064 40224 11076
rect 39899 11036 40224 11064
rect 39899 11033 39911 11036
rect 39853 11027 39911 11033
rect 40218 11024 40224 11036
rect 40276 11064 40282 11076
rect 40586 11064 40592 11076
rect 40276 11036 40592 11064
rect 40276 11024 40282 11036
rect 40586 11024 40592 11036
rect 40644 11024 40650 11076
rect 43162 11064 43168 11076
rect 43123 11036 43168 11064
rect 43162 11024 43168 11036
rect 43220 11064 43226 11076
rect 44008 11064 44036 11095
rect 43220 11036 44036 11064
rect 43220 11024 43226 11036
rect 23164 10968 23428 10996
rect 35253 10999 35311 11005
rect 23164 10956 23170 10968
rect 35253 10965 35265 10999
rect 35299 10996 35311 10999
rect 35342 10996 35348 11008
rect 35299 10968 35348 10996
rect 35299 10965 35311 10968
rect 35253 10959 35311 10965
rect 35342 10956 35348 10968
rect 35400 10996 35406 11008
rect 35805 10999 35863 11005
rect 35805 10996 35817 10999
rect 35400 10968 35817 10996
rect 35400 10956 35406 10968
rect 35805 10965 35817 10968
rect 35851 10965 35863 10999
rect 35805 10959 35863 10965
rect 39485 10999 39543 11005
rect 39485 10965 39497 10999
rect 39531 10996 39543 10999
rect 39574 10996 39580 11008
rect 39531 10968 39580 10996
rect 39531 10965 39543 10968
rect 39485 10959 39543 10965
rect 39574 10956 39580 10968
rect 39632 10956 39638 11008
rect 43438 10996 43444 11008
rect 43399 10968 43444 10996
rect 43438 10956 43444 10968
rect 43496 10956 43502 11008
rect 1104 10906 48852 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 34966 10906
rect 35018 10854 35030 10906
rect 35082 10854 35094 10906
rect 35146 10854 35158 10906
rect 35210 10854 48852 10906
rect 1104 10832 48852 10854
rect 4341 10795 4399 10801
rect 4341 10761 4353 10795
rect 4387 10792 4399 10795
rect 4614 10792 4620 10804
rect 4387 10764 4620 10792
rect 4387 10761 4399 10764
rect 4341 10755 4399 10761
rect 4614 10752 4620 10764
rect 4672 10752 4678 10804
rect 4982 10792 4988 10804
rect 4943 10764 4988 10792
rect 4982 10752 4988 10764
rect 5040 10752 5046 10804
rect 5258 10792 5264 10804
rect 5219 10764 5264 10792
rect 5258 10752 5264 10764
rect 5316 10752 5322 10804
rect 5810 10752 5816 10804
rect 5868 10792 5874 10804
rect 6181 10795 6239 10801
rect 6181 10792 6193 10795
rect 5868 10764 6193 10792
rect 5868 10752 5874 10764
rect 6181 10761 6193 10764
rect 6227 10761 6239 10795
rect 11054 10792 11060 10804
rect 11015 10764 11060 10792
rect 6181 10755 6239 10761
rect 11054 10752 11060 10764
rect 11112 10752 11118 10804
rect 11882 10792 11888 10804
rect 11843 10764 11888 10792
rect 11882 10752 11888 10764
rect 11940 10752 11946 10804
rect 12526 10792 12532 10804
rect 12487 10764 12532 10792
rect 12526 10752 12532 10764
rect 12584 10752 12590 10804
rect 15654 10792 15660 10804
rect 15615 10764 15660 10792
rect 15654 10752 15660 10764
rect 15712 10752 15718 10804
rect 16022 10792 16028 10804
rect 15983 10764 16028 10792
rect 16022 10752 16028 10764
rect 16080 10752 16086 10804
rect 18414 10752 18420 10804
rect 18472 10792 18478 10804
rect 19061 10795 19119 10801
rect 19061 10792 19073 10795
rect 18472 10764 19073 10792
rect 18472 10752 18478 10764
rect 19061 10761 19073 10764
rect 19107 10761 19119 10795
rect 19061 10755 19119 10761
rect 22278 10752 22284 10804
rect 22336 10792 22342 10804
rect 22741 10795 22799 10801
rect 22741 10792 22753 10795
rect 22336 10764 22753 10792
rect 22336 10752 22342 10764
rect 22741 10761 22753 10764
rect 22787 10761 22799 10795
rect 22741 10755 22799 10761
rect 25869 10795 25927 10801
rect 25869 10761 25881 10795
rect 25915 10792 25927 10795
rect 26142 10792 26148 10804
rect 25915 10764 26148 10792
rect 25915 10761 25927 10764
rect 25869 10755 25927 10761
rect 26142 10752 26148 10764
rect 26200 10752 26206 10804
rect 27246 10792 27252 10804
rect 27207 10764 27252 10792
rect 27246 10752 27252 10764
rect 27304 10752 27310 10804
rect 28353 10795 28411 10801
rect 28353 10761 28365 10795
rect 28399 10792 28411 10795
rect 29638 10792 29644 10804
rect 28399 10764 29644 10792
rect 28399 10761 28411 10764
rect 28353 10755 28411 10761
rect 29638 10752 29644 10764
rect 29696 10792 29702 10804
rect 30653 10795 30711 10801
rect 30653 10792 30665 10795
rect 29696 10764 30665 10792
rect 29696 10752 29702 10764
rect 30653 10761 30665 10764
rect 30699 10761 30711 10795
rect 33870 10792 33876 10804
rect 33831 10764 33876 10792
rect 30653 10755 30711 10761
rect 33870 10752 33876 10764
rect 33928 10752 33934 10804
rect 34238 10792 34244 10804
rect 34199 10764 34244 10792
rect 34238 10752 34244 10764
rect 34296 10752 34302 10804
rect 37734 10752 37740 10804
rect 37792 10792 37798 10804
rect 38381 10795 38439 10801
rect 38381 10792 38393 10795
rect 37792 10764 38393 10792
rect 37792 10752 37798 10764
rect 38381 10761 38393 10764
rect 38427 10792 38439 10795
rect 38427 10764 38976 10792
rect 38427 10761 38439 10764
rect 38381 10755 38439 10761
rect 6914 10724 6920 10736
rect 6875 10696 6920 10724
rect 6914 10684 6920 10696
rect 6972 10684 6978 10736
rect 11422 10724 11428 10736
rect 11383 10696 11428 10724
rect 11422 10684 11428 10696
rect 11480 10684 11486 10736
rect 18141 10727 18199 10733
rect 18141 10693 18153 10727
rect 18187 10724 18199 10727
rect 19242 10724 19248 10736
rect 18187 10696 19248 10724
rect 18187 10693 18199 10696
rect 18141 10687 18199 10693
rect 19242 10684 19248 10696
rect 19300 10684 19306 10736
rect 33888 10724 33916 10752
rect 34609 10727 34667 10733
rect 34609 10724 34621 10727
rect 33888 10696 34621 10724
rect 34609 10693 34621 10696
rect 34655 10724 34667 10727
rect 34790 10724 34796 10736
rect 34655 10696 34796 10724
rect 34655 10693 34667 10696
rect 34609 10687 34667 10693
rect 34790 10684 34796 10696
rect 34848 10724 34854 10736
rect 38948 10733 38976 10764
rect 39666 10752 39672 10804
rect 39724 10792 39730 10804
rect 39853 10795 39911 10801
rect 39853 10792 39865 10795
rect 39724 10764 39865 10792
rect 39724 10752 39730 10764
rect 39853 10761 39865 10764
rect 39899 10761 39911 10795
rect 39853 10755 39911 10761
rect 40954 10752 40960 10804
rect 41012 10792 41018 10804
rect 41049 10795 41107 10801
rect 41049 10792 41061 10795
rect 41012 10764 41061 10792
rect 41012 10752 41018 10764
rect 41049 10761 41061 10764
rect 41095 10761 41107 10795
rect 41506 10792 41512 10804
rect 41467 10764 41512 10792
rect 41049 10755 41107 10761
rect 41506 10752 41512 10764
rect 41564 10752 41570 10804
rect 43070 10752 43076 10804
rect 43128 10792 43134 10804
rect 44729 10795 44787 10801
rect 44729 10792 44741 10795
rect 43128 10764 44741 10792
rect 43128 10752 43134 10764
rect 44729 10761 44741 10764
rect 44775 10761 44787 10795
rect 44729 10755 44787 10761
rect 37921 10727 37979 10733
rect 34848 10696 35020 10724
rect 34848 10684 34854 10696
rect 1486 10616 1492 10668
rect 1544 10656 1550 10668
rect 1581 10659 1639 10665
rect 1581 10656 1593 10659
rect 1544 10628 1593 10656
rect 1544 10616 1550 10628
rect 1581 10625 1593 10628
rect 1627 10625 1639 10659
rect 7466 10656 7472 10668
rect 7427 10628 7472 10656
rect 1581 10619 1639 10625
rect 7466 10616 7472 10628
rect 7524 10656 7530 10668
rect 7837 10659 7895 10665
rect 7837 10656 7849 10659
rect 7524 10628 7849 10656
rect 7524 10616 7530 10628
rect 7837 10625 7849 10628
rect 7883 10625 7895 10659
rect 7837 10619 7895 10625
rect 11054 10616 11060 10668
rect 11112 10656 11118 10668
rect 11606 10656 11612 10668
rect 11112 10628 11612 10656
rect 11112 10616 11118 10628
rect 11606 10616 11612 10628
rect 11664 10656 11670 10668
rect 12161 10659 12219 10665
rect 12161 10656 12173 10659
rect 11664 10628 12173 10656
rect 11664 10616 11670 10628
rect 12161 10625 12173 10628
rect 12207 10625 12219 10659
rect 13078 10656 13084 10668
rect 13039 10628 13084 10656
rect 12161 10619 12219 10625
rect 13078 10616 13084 10628
rect 13136 10616 13142 10668
rect 20254 10616 20260 10668
rect 20312 10656 20318 10668
rect 20809 10659 20867 10665
rect 20809 10656 20821 10659
rect 20312 10628 20821 10656
rect 20312 10616 20318 10628
rect 20809 10625 20821 10628
rect 20855 10625 20867 10659
rect 20809 10619 20867 10625
rect 20898 10616 20904 10668
rect 20956 10656 20962 10668
rect 21085 10659 21143 10665
rect 21085 10656 21097 10659
rect 20956 10628 21097 10656
rect 20956 10616 20962 10628
rect 21085 10625 21097 10628
rect 21131 10625 21143 10659
rect 21085 10619 21143 10625
rect 28350 10616 28356 10668
rect 28408 10656 28414 10668
rect 28629 10659 28687 10665
rect 28629 10656 28641 10659
rect 28408 10628 28641 10656
rect 28408 10616 28414 10628
rect 28629 10625 28641 10628
rect 28675 10656 28687 10659
rect 28997 10659 29055 10665
rect 28997 10656 29009 10659
rect 28675 10628 29009 10656
rect 28675 10625 28687 10628
rect 28629 10619 28687 10625
rect 28997 10625 29009 10628
rect 29043 10656 29055 10659
rect 29270 10656 29276 10668
rect 29043 10628 29276 10656
rect 29043 10625 29055 10628
rect 28997 10619 29055 10625
rect 29270 10616 29276 10628
rect 29328 10616 29334 10668
rect 34992 10665 35020 10696
rect 37921 10693 37933 10727
rect 37967 10724 37979 10727
rect 38657 10727 38715 10733
rect 38657 10724 38669 10727
rect 37967 10696 38669 10724
rect 37967 10693 37979 10696
rect 37921 10687 37979 10693
rect 38657 10693 38669 10696
rect 38703 10693 38715 10727
rect 38657 10687 38715 10693
rect 38933 10727 38991 10733
rect 38933 10693 38945 10727
rect 38979 10724 38991 10727
rect 39758 10724 39764 10736
rect 38979 10696 39764 10724
rect 38979 10693 38991 10696
rect 38933 10687 38991 10693
rect 34977 10659 35035 10665
rect 34977 10625 34989 10659
rect 35023 10625 35035 10659
rect 38672 10656 38700 10687
rect 39758 10684 39764 10696
rect 39816 10684 39822 10736
rect 40773 10727 40831 10733
rect 40773 10693 40785 10727
rect 40819 10724 40831 10727
rect 41322 10724 41328 10736
rect 40819 10696 41328 10724
rect 40819 10693 40831 10696
rect 40773 10687 40831 10693
rect 41322 10684 41328 10696
rect 41380 10684 41386 10736
rect 38672 10628 39436 10656
rect 34977 10619 35035 10625
rect 1848 10591 1906 10597
rect 1848 10557 1860 10591
rect 1894 10588 1906 10591
rect 2406 10588 2412 10600
rect 1894 10560 2412 10588
rect 1894 10557 1906 10560
rect 1848 10551 1906 10557
rect 2406 10548 2412 10560
rect 2464 10548 2470 10600
rect 5534 10588 5540 10600
rect 5495 10560 5540 10588
rect 5534 10548 5540 10560
rect 5592 10548 5598 10600
rect 7190 10588 7196 10600
rect 7151 10560 7196 10588
rect 7190 10548 7196 10560
rect 7248 10548 7254 10600
rect 8297 10591 8355 10597
rect 8297 10557 8309 10591
rect 8343 10588 8355 10591
rect 8389 10591 8447 10597
rect 8389 10588 8401 10591
rect 8343 10560 8401 10588
rect 8343 10557 8355 10560
rect 8297 10551 8355 10557
rect 8389 10557 8401 10560
rect 8435 10557 8447 10591
rect 8389 10551 8447 10557
rect 4709 10523 4767 10529
rect 4709 10489 4721 10523
rect 4755 10520 4767 10523
rect 5813 10523 5871 10529
rect 5813 10520 5825 10523
rect 4755 10492 5825 10520
rect 4755 10489 4767 10492
rect 4709 10483 4767 10489
rect 5813 10489 5825 10492
rect 5859 10520 5871 10523
rect 5902 10520 5908 10532
rect 5859 10492 5908 10520
rect 5859 10489 5871 10492
rect 5813 10483 5871 10489
rect 5902 10480 5908 10492
rect 5960 10480 5966 10532
rect 8404 10520 8432 10551
rect 8478 10548 8484 10600
rect 8536 10588 8542 10600
rect 8645 10591 8703 10597
rect 8645 10588 8657 10591
rect 8536 10560 8657 10588
rect 8536 10548 8542 10560
rect 8645 10557 8657 10560
rect 8691 10557 8703 10591
rect 8645 10551 8703 10557
rect 11146 10548 11152 10600
rect 11204 10588 11210 10600
rect 11241 10591 11299 10597
rect 11241 10588 11253 10591
rect 11204 10560 11253 10588
rect 11204 10548 11210 10560
rect 11241 10557 11253 10560
rect 11287 10557 11299 10591
rect 11241 10551 11299 10557
rect 12434 10548 12440 10600
rect 12492 10588 12498 10600
rect 12805 10591 12863 10597
rect 12805 10588 12817 10591
rect 12492 10560 12817 10588
rect 12492 10548 12498 10560
rect 12805 10557 12817 10560
rect 12851 10588 12863 10591
rect 13449 10591 13507 10597
rect 13449 10588 13461 10591
rect 12851 10560 13461 10588
rect 12851 10557 12863 10560
rect 12805 10551 12863 10557
rect 13449 10557 13461 10560
rect 13495 10557 13507 10591
rect 13449 10551 13507 10557
rect 18506 10548 18512 10600
rect 18564 10588 18570 10600
rect 18693 10591 18751 10597
rect 18693 10588 18705 10591
rect 18564 10560 18705 10588
rect 18564 10548 18570 10560
rect 18693 10557 18705 10560
rect 18739 10557 18751 10591
rect 18693 10551 18751 10557
rect 19889 10591 19947 10597
rect 19889 10557 19901 10591
rect 19935 10588 19947 10591
rect 20349 10591 20407 10597
rect 20349 10588 20361 10591
rect 19935 10560 20361 10588
rect 19935 10557 19947 10560
rect 19889 10551 19947 10557
rect 20349 10557 20361 10560
rect 20395 10588 20407 10591
rect 20438 10588 20444 10600
rect 20395 10560 20444 10588
rect 20395 10557 20407 10560
rect 20349 10551 20407 10557
rect 20438 10548 20444 10560
rect 20496 10548 20502 10600
rect 37645 10591 37703 10597
rect 37645 10557 37657 10591
rect 37691 10588 37703 10591
rect 37737 10591 37795 10597
rect 37737 10588 37749 10591
rect 37691 10560 37749 10588
rect 37691 10557 37703 10560
rect 37645 10551 37703 10557
rect 37737 10557 37749 10560
rect 37783 10588 37795 10591
rect 37826 10588 37832 10600
rect 37783 10560 37832 10588
rect 37783 10557 37795 10560
rect 37737 10551 37795 10557
rect 37826 10548 37832 10560
rect 37884 10548 37890 10600
rect 9674 10520 9680 10532
rect 8404 10492 9680 10520
rect 9674 10480 9680 10492
rect 9732 10480 9738 10532
rect 12986 10520 12992 10532
rect 12947 10492 12992 10520
rect 12986 10480 12992 10492
rect 13044 10480 13050 10532
rect 17497 10523 17555 10529
rect 17497 10489 17509 10523
rect 17543 10520 17555 10523
rect 17862 10520 17868 10532
rect 17543 10492 17868 10520
rect 17543 10489 17555 10492
rect 17497 10483 17555 10489
rect 17862 10480 17868 10492
rect 17920 10520 17926 10532
rect 18417 10523 18475 10529
rect 18417 10520 18429 10523
rect 17920 10492 18429 10520
rect 17920 10480 17926 10492
rect 18417 10489 18429 10492
rect 18463 10489 18475 10523
rect 18598 10520 18604 10532
rect 18559 10492 18604 10520
rect 18417 10483 18475 10489
rect 18598 10480 18604 10492
rect 18656 10480 18662 10532
rect 25961 10523 26019 10529
rect 25961 10489 25973 10523
rect 26007 10520 26019 10523
rect 26050 10520 26056 10532
rect 26007 10492 26056 10520
rect 26007 10489 26019 10492
rect 25961 10483 26019 10489
rect 26050 10480 26056 10492
rect 26108 10480 26114 10532
rect 29546 10529 29552 10532
rect 29540 10520 29552 10529
rect 29507 10492 29552 10520
rect 29540 10483 29552 10492
rect 29546 10480 29552 10483
rect 29604 10480 29610 10532
rect 35244 10523 35302 10529
rect 35244 10489 35256 10523
rect 35290 10520 35302 10523
rect 35342 10520 35348 10532
rect 35290 10492 35348 10520
rect 35290 10489 35302 10492
rect 35244 10483 35302 10489
rect 35342 10480 35348 10492
rect 35400 10480 35406 10532
rect 39206 10520 39212 10532
rect 39167 10492 39212 10520
rect 39206 10480 39212 10492
rect 39264 10480 39270 10532
rect 39408 10529 39436 10628
rect 43349 10591 43407 10597
rect 43349 10557 43361 10591
rect 43395 10588 43407 10591
rect 43395 10560 43760 10588
rect 43395 10557 43407 10560
rect 43349 10551 43407 10557
rect 39393 10523 39451 10529
rect 39393 10489 39405 10523
rect 39439 10489 39451 10523
rect 39393 10483 39451 10489
rect 39485 10523 39543 10529
rect 39485 10489 39497 10523
rect 39531 10520 39543 10523
rect 39574 10520 39580 10532
rect 39531 10492 39580 10520
rect 39531 10489 39543 10492
rect 39485 10483 39543 10489
rect 39574 10480 39580 10492
rect 39632 10480 39638 10532
rect 41782 10520 41788 10532
rect 41743 10492 41788 10520
rect 41782 10480 41788 10492
rect 41840 10480 41846 10532
rect 42058 10520 42064 10532
rect 42019 10492 42064 10520
rect 42058 10480 42064 10492
rect 42116 10480 42122 10532
rect 43622 10529 43628 10532
rect 42521 10523 42579 10529
rect 42521 10489 42533 10523
rect 42567 10520 42579 10523
rect 42889 10523 42947 10529
rect 42889 10520 42901 10523
rect 42567 10492 42901 10520
rect 42567 10489 42579 10492
rect 42521 10483 42579 10489
rect 42889 10489 42901 10492
rect 42935 10520 42947 10523
rect 43616 10520 43628 10529
rect 42935 10492 43628 10520
rect 42935 10489 42947 10492
rect 42889 10483 42947 10489
rect 43616 10483 43628 10492
rect 43622 10480 43628 10483
rect 43680 10480 43686 10532
rect 2498 10412 2504 10464
rect 2556 10452 2562 10464
rect 2961 10455 3019 10461
rect 2961 10452 2973 10455
rect 2556 10424 2973 10452
rect 2556 10412 2562 10424
rect 2961 10421 2973 10424
rect 3007 10421 3019 10455
rect 2961 10415 3019 10421
rect 5258 10412 5264 10464
rect 5316 10452 5322 10464
rect 5721 10455 5779 10461
rect 5721 10452 5733 10455
rect 5316 10424 5733 10452
rect 5316 10412 5322 10424
rect 5721 10421 5733 10424
rect 5767 10421 5779 10455
rect 5721 10415 5779 10421
rect 6546 10412 6552 10464
rect 6604 10452 6610 10464
rect 6641 10455 6699 10461
rect 6641 10452 6653 10455
rect 6604 10424 6653 10452
rect 6604 10412 6610 10424
rect 6641 10421 6653 10424
rect 6687 10452 6699 10455
rect 7377 10455 7435 10461
rect 7377 10452 7389 10455
rect 6687 10424 7389 10452
rect 6687 10421 6699 10424
rect 6641 10415 6699 10421
rect 7377 10421 7389 10424
rect 7423 10421 7435 10455
rect 9766 10452 9772 10464
rect 9727 10424 9772 10452
rect 7377 10415 7435 10421
rect 9766 10412 9772 10424
rect 9824 10412 9830 10464
rect 10413 10455 10471 10461
rect 10413 10421 10425 10455
rect 10459 10452 10471 10455
rect 10686 10452 10692 10464
rect 10459 10424 10692 10452
rect 10459 10421 10471 10424
rect 10413 10415 10471 10421
rect 10686 10412 10692 10424
rect 10744 10412 10750 10464
rect 17770 10452 17776 10464
rect 17731 10424 17776 10452
rect 17770 10412 17776 10424
rect 17828 10412 17834 10464
rect 20257 10455 20315 10461
rect 20257 10421 20269 10455
rect 20303 10452 20315 10455
rect 20811 10455 20869 10461
rect 20811 10452 20823 10455
rect 20303 10424 20823 10452
rect 20303 10421 20315 10424
rect 20257 10415 20315 10421
rect 20811 10421 20823 10424
rect 20857 10452 20869 10455
rect 20990 10452 20996 10464
rect 20857 10424 20996 10452
rect 20857 10421 20869 10424
rect 20811 10415 20869 10421
rect 20990 10412 20996 10424
rect 21048 10412 21054 10464
rect 21450 10412 21456 10464
rect 21508 10452 21514 10464
rect 22189 10455 22247 10461
rect 22189 10452 22201 10455
rect 21508 10424 22201 10452
rect 21508 10412 21514 10424
rect 22189 10421 22201 10424
rect 22235 10421 22247 10455
rect 22189 10415 22247 10421
rect 23014 10412 23020 10464
rect 23072 10452 23078 10464
rect 23661 10455 23719 10461
rect 23661 10452 23673 10455
rect 23072 10424 23673 10452
rect 23072 10412 23078 10424
rect 23661 10421 23673 10424
rect 23707 10421 23719 10455
rect 36354 10452 36360 10464
rect 36315 10424 36360 10452
rect 23661 10415 23719 10421
rect 36354 10412 36360 10424
rect 36412 10412 36418 10464
rect 41966 10452 41972 10464
rect 41927 10424 41972 10452
rect 41966 10412 41972 10424
rect 42024 10412 42030 10464
rect 43257 10455 43315 10461
rect 43257 10421 43269 10455
rect 43303 10452 43315 10455
rect 43732 10452 43760 10560
rect 44082 10452 44088 10464
rect 43303 10424 44088 10452
rect 43303 10421 43315 10424
rect 43257 10415 43315 10421
rect 44082 10412 44088 10424
rect 44140 10412 44146 10464
rect 1104 10362 48852 10384
rect 1104 10310 19606 10362
rect 19658 10310 19670 10362
rect 19722 10310 19734 10362
rect 19786 10310 19798 10362
rect 19850 10310 48852 10362
rect 1104 10288 48852 10310
rect 1486 10208 1492 10260
rect 1544 10248 1550 10260
rect 1581 10251 1639 10257
rect 1581 10248 1593 10251
rect 1544 10220 1593 10248
rect 1544 10208 1550 10220
rect 1581 10217 1593 10220
rect 1627 10217 1639 10251
rect 2498 10248 2504 10260
rect 2459 10220 2504 10248
rect 1581 10211 1639 10217
rect 2498 10208 2504 10220
rect 2556 10208 2562 10260
rect 4341 10251 4399 10257
rect 4341 10217 4353 10251
rect 4387 10248 4399 10251
rect 5258 10248 5264 10260
rect 4387 10220 5264 10248
rect 4387 10217 4399 10220
rect 4341 10211 4399 10217
rect 5258 10208 5264 10220
rect 5316 10208 5322 10260
rect 5534 10248 5540 10260
rect 5495 10220 5540 10248
rect 5534 10208 5540 10220
rect 5592 10208 5598 10260
rect 5902 10248 5908 10260
rect 5863 10220 5908 10248
rect 5902 10208 5908 10220
rect 5960 10208 5966 10260
rect 8478 10208 8484 10260
rect 8536 10248 8542 10260
rect 8573 10251 8631 10257
rect 8573 10248 8585 10251
rect 8536 10220 8585 10248
rect 8536 10208 8542 10220
rect 8573 10217 8585 10220
rect 8619 10217 8631 10251
rect 8573 10211 8631 10217
rect 12342 10208 12348 10260
rect 12400 10248 12406 10260
rect 12713 10251 12771 10257
rect 12713 10248 12725 10251
rect 12400 10220 12725 10248
rect 12400 10208 12406 10220
rect 12713 10217 12725 10220
rect 12759 10217 12771 10251
rect 12713 10211 12771 10217
rect 12986 10208 12992 10260
rect 13044 10248 13050 10260
rect 13173 10251 13231 10257
rect 13173 10248 13185 10251
rect 13044 10220 13185 10248
rect 13044 10208 13050 10220
rect 13173 10217 13185 10220
rect 13219 10217 13231 10251
rect 17862 10248 17868 10260
rect 17823 10220 17868 10248
rect 13173 10211 13231 10217
rect 17862 10208 17868 10220
rect 17920 10208 17926 10260
rect 18417 10251 18475 10257
rect 18417 10217 18429 10251
rect 18463 10248 18475 10251
rect 18506 10248 18512 10260
rect 18463 10220 18512 10248
rect 18463 10217 18475 10220
rect 18417 10211 18475 10217
rect 18506 10208 18512 10220
rect 18564 10208 18570 10260
rect 18598 10208 18604 10260
rect 18656 10248 18662 10260
rect 18693 10251 18751 10257
rect 18693 10248 18705 10251
rect 18656 10220 18705 10248
rect 18656 10208 18662 10220
rect 18693 10217 18705 10220
rect 18739 10217 18751 10251
rect 18693 10211 18751 10217
rect 20254 10208 20260 10260
rect 20312 10248 20318 10260
rect 20349 10251 20407 10257
rect 20349 10248 20361 10251
rect 20312 10220 20361 10248
rect 20312 10208 20318 10220
rect 20349 10217 20361 10220
rect 20395 10217 20407 10251
rect 20349 10211 20407 10217
rect 20983 10251 21041 10257
rect 20983 10217 20995 10251
rect 21029 10248 21041 10251
rect 23017 10251 23075 10257
rect 23017 10248 23029 10251
rect 21029 10220 23029 10248
rect 21029 10217 21041 10220
rect 20983 10211 21041 10217
rect 23017 10217 23029 10220
rect 23063 10248 23075 10251
rect 23198 10248 23204 10260
rect 23063 10220 23204 10248
rect 23063 10217 23075 10220
rect 23017 10211 23075 10217
rect 2038 10140 2044 10192
rect 2096 10180 2102 10192
rect 2593 10183 2651 10189
rect 2593 10180 2605 10183
rect 2096 10152 2605 10180
rect 2096 10140 2102 10152
rect 2593 10149 2605 10152
rect 2639 10180 2651 10183
rect 2682 10180 2688 10192
rect 2639 10152 2688 10180
rect 2639 10149 2651 10152
rect 2593 10143 2651 10149
rect 2682 10140 2688 10152
rect 2740 10140 2746 10192
rect 7009 10183 7067 10189
rect 7009 10149 7021 10183
rect 7055 10180 7067 10183
rect 7098 10180 7104 10192
rect 7055 10152 7104 10180
rect 7055 10149 7067 10152
rect 7009 10143 7067 10149
rect 7098 10140 7104 10152
rect 7156 10140 7162 10192
rect 11146 10140 11152 10192
rect 11204 10180 11210 10192
rect 12526 10180 12532 10192
rect 11204 10152 12532 10180
rect 11204 10140 11210 10152
rect 12526 10140 12532 10152
rect 12584 10140 12590 10192
rect 15841 10183 15899 10189
rect 15841 10149 15853 10183
rect 15887 10180 15899 10183
rect 15930 10180 15936 10192
rect 15887 10152 15936 10180
rect 15887 10149 15899 10152
rect 15841 10143 15899 10149
rect 15930 10140 15936 10152
rect 15988 10140 15994 10192
rect 20364 10180 20392 10211
rect 23198 10208 23204 10220
rect 23256 10208 23262 10260
rect 25406 10248 25412 10260
rect 25367 10220 25412 10248
rect 25406 10208 25412 10220
rect 25464 10208 25470 10260
rect 26602 10208 26608 10260
rect 26660 10248 26666 10260
rect 26697 10251 26755 10257
rect 26697 10248 26709 10251
rect 26660 10220 26709 10248
rect 26660 10208 26666 10220
rect 26697 10217 26709 10220
rect 26743 10217 26755 10251
rect 26697 10211 26755 10217
rect 28718 10208 28724 10260
rect 28776 10248 28782 10260
rect 28997 10251 29055 10257
rect 28997 10248 29009 10251
rect 28776 10220 29009 10248
rect 28776 10208 28782 10220
rect 28997 10217 29009 10220
rect 29043 10248 29055 10251
rect 29638 10248 29644 10260
rect 29043 10220 29644 10248
rect 29043 10217 29055 10220
rect 28997 10211 29055 10217
rect 29638 10208 29644 10220
rect 29696 10208 29702 10260
rect 34238 10208 34244 10260
rect 34296 10248 34302 10260
rect 35437 10251 35495 10257
rect 35437 10248 35449 10251
rect 34296 10220 35449 10248
rect 34296 10208 34302 10220
rect 35437 10217 35449 10220
rect 35483 10217 35495 10251
rect 35437 10211 35495 10217
rect 38933 10251 38991 10257
rect 38933 10217 38945 10251
rect 38979 10248 38991 10251
rect 39206 10248 39212 10260
rect 38979 10220 39212 10248
rect 38979 10217 38991 10220
rect 38933 10211 38991 10217
rect 39206 10208 39212 10220
rect 39264 10248 39270 10260
rect 39485 10251 39543 10257
rect 39485 10248 39497 10251
rect 39264 10220 39497 10248
rect 39264 10208 39270 10220
rect 39485 10217 39497 10220
rect 39531 10217 39543 10251
rect 40586 10248 40592 10260
rect 40547 10220 40592 10248
rect 39485 10211 39543 10217
rect 40586 10208 40592 10220
rect 40644 10208 40650 10260
rect 41782 10248 41788 10260
rect 41743 10220 41788 10248
rect 41782 10208 41788 10220
rect 41840 10248 41846 10260
rect 42337 10251 42395 10257
rect 42337 10248 42349 10251
rect 41840 10220 42349 10248
rect 41840 10208 41846 10220
rect 42337 10217 42349 10220
rect 42383 10217 42395 10251
rect 43070 10248 43076 10260
rect 43031 10220 43076 10248
rect 42337 10211 42395 10217
rect 43070 10208 43076 10220
rect 43128 10208 43134 10260
rect 46934 10248 46940 10260
rect 46895 10220 46940 10248
rect 46934 10208 46940 10220
rect 46992 10208 46998 10260
rect 21266 10180 21272 10192
rect 20364 10152 21272 10180
rect 21266 10140 21272 10152
rect 21324 10140 21330 10192
rect 21450 10180 21456 10192
rect 21411 10152 21456 10180
rect 21450 10140 21456 10152
rect 21508 10140 21514 10192
rect 21545 10183 21603 10189
rect 21545 10149 21557 10183
rect 21591 10180 21603 10183
rect 21726 10180 21732 10192
rect 21591 10152 21732 10180
rect 21591 10149 21603 10152
rect 21545 10143 21603 10149
rect 21726 10140 21732 10152
rect 21784 10180 21790 10192
rect 22186 10180 22192 10192
rect 21784 10152 22192 10180
rect 21784 10140 21790 10152
rect 22186 10140 22192 10152
rect 22244 10140 22250 10192
rect 26050 10180 26056 10192
rect 26011 10152 26056 10180
rect 26050 10140 26056 10152
rect 26108 10140 26114 10192
rect 27522 10140 27528 10192
rect 27580 10180 27586 10192
rect 28810 10180 28816 10192
rect 27580 10152 28816 10180
rect 27580 10140 27586 10152
rect 28810 10140 28816 10152
rect 28868 10140 28874 10192
rect 37734 10140 37740 10192
rect 37792 10180 37798 10192
rect 38289 10183 38347 10189
rect 38289 10180 38301 10183
rect 37792 10152 38301 10180
rect 37792 10140 37798 10152
rect 38289 10149 38301 10152
rect 38335 10149 38347 10183
rect 38289 10143 38347 10149
rect 39574 10140 39580 10192
rect 39632 10180 39638 10192
rect 41049 10183 41107 10189
rect 41049 10180 41061 10183
rect 39632 10152 41061 10180
rect 39632 10140 39638 10152
rect 41049 10149 41061 10152
rect 41095 10180 41107 10183
rect 42058 10180 42064 10192
rect 41095 10152 42064 10180
rect 41095 10149 41107 10152
rect 41049 10143 41107 10149
rect 42058 10140 42064 10152
rect 42116 10140 42122 10192
rect 43438 10140 43444 10192
rect 43496 10180 43502 10192
rect 43717 10183 43775 10189
rect 43717 10180 43729 10183
rect 43496 10152 43729 10180
rect 43496 10140 43502 10152
rect 43717 10149 43729 10152
rect 43763 10149 43775 10183
rect 43898 10180 43904 10192
rect 43859 10152 43904 10180
rect 43717 10143 43775 10149
rect 43898 10140 43904 10152
rect 43956 10140 43962 10192
rect 4157 10115 4215 10121
rect 4157 10081 4169 10115
rect 4203 10112 4215 10115
rect 4614 10112 4620 10124
rect 4203 10084 4620 10112
rect 4203 10081 4215 10084
rect 4157 10075 4215 10081
rect 4614 10072 4620 10084
rect 4672 10072 4678 10124
rect 5350 10112 5356 10124
rect 5311 10084 5356 10112
rect 5350 10072 5356 10084
rect 5408 10072 5414 10124
rect 8389 10115 8447 10121
rect 8389 10081 8401 10115
rect 8435 10112 8447 10115
rect 9766 10112 9772 10124
rect 8435 10084 9772 10112
rect 8435 10081 8447 10084
rect 8389 10075 8447 10081
rect 9766 10072 9772 10084
rect 9824 10112 9830 10124
rect 9944 10115 10002 10121
rect 9944 10112 9956 10115
rect 9824 10084 9956 10112
rect 9824 10072 9830 10084
rect 9944 10081 9956 10084
rect 9990 10112 10002 10115
rect 10410 10112 10416 10124
rect 9990 10084 10416 10112
rect 9990 10081 10002 10084
rect 9944 10075 10002 10081
rect 10410 10072 10416 10084
rect 10468 10072 10474 10124
rect 15654 10112 15660 10124
rect 15615 10084 15660 10112
rect 15654 10072 15660 10084
rect 15712 10072 15718 10124
rect 34514 10072 34520 10124
rect 34572 10112 34578 10124
rect 35529 10115 35587 10121
rect 35529 10112 35541 10115
rect 34572 10084 35541 10112
rect 34572 10072 34578 10084
rect 35529 10081 35541 10084
rect 35575 10112 35587 10115
rect 35802 10112 35808 10124
rect 35575 10084 35808 10112
rect 35575 10081 35587 10084
rect 35529 10075 35587 10081
rect 35802 10072 35808 10084
rect 35860 10072 35866 10124
rect 38102 10112 38108 10124
rect 38063 10084 38108 10112
rect 38102 10072 38108 10084
rect 38160 10072 38166 10124
rect 39298 10112 39304 10124
rect 39259 10084 39304 10112
rect 39298 10072 39304 10084
rect 39356 10072 39362 10124
rect 40405 10115 40463 10121
rect 40405 10081 40417 10115
rect 40451 10112 40463 10115
rect 40770 10112 40776 10124
rect 40451 10084 40776 10112
rect 40451 10081 40463 10084
rect 40405 10075 40463 10081
rect 40770 10072 40776 10084
rect 40828 10112 40834 10124
rect 41138 10112 41144 10124
rect 40828 10084 41144 10112
rect 40828 10072 40834 10084
rect 41138 10072 41144 10084
rect 41196 10072 41202 10124
rect 42153 10115 42211 10121
rect 42153 10081 42165 10115
rect 42199 10112 42211 10115
rect 42426 10112 42432 10124
rect 42199 10084 42432 10112
rect 42199 10081 42211 10084
rect 42153 10075 42211 10081
rect 42426 10072 42432 10084
rect 42484 10112 42490 10124
rect 45830 10121 45836 10124
rect 45824 10112 45836 10121
rect 42484 10084 43484 10112
rect 45791 10084 45836 10112
rect 42484 10072 42490 10084
rect 2498 10044 2504 10056
rect 2459 10016 2504 10044
rect 2498 10004 2504 10016
rect 2556 10004 2562 10056
rect 7006 10044 7012 10056
rect 6967 10016 7012 10044
rect 7006 10004 7012 10016
rect 7064 10004 7070 10056
rect 7101 10047 7159 10053
rect 7101 10013 7113 10047
rect 7147 10044 7159 10047
rect 7282 10044 7288 10056
rect 7147 10016 7288 10044
rect 7147 10013 7159 10016
rect 7101 10007 7159 10013
rect 7282 10004 7288 10016
rect 7340 10044 7346 10056
rect 7834 10044 7840 10056
rect 7340 10016 7840 10044
rect 7340 10004 7346 10016
rect 7834 10004 7840 10016
rect 7892 10044 7898 10056
rect 8665 10047 8723 10053
rect 8665 10044 8677 10047
rect 7892 10016 8677 10044
rect 7892 10004 7898 10016
rect 8665 10013 8677 10016
rect 8711 10044 8723 10047
rect 9033 10047 9091 10053
rect 9033 10044 9045 10047
rect 8711 10016 9045 10044
rect 8711 10013 8723 10016
rect 8665 10007 8723 10013
rect 9033 10013 9045 10016
rect 9079 10013 9091 10047
rect 9674 10044 9680 10056
rect 9635 10016 9680 10044
rect 9033 10007 9091 10013
rect 9674 10004 9680 10016
rect 9732 10004 9738 10056
rect 12802 10044 12808 10056
rect 12763 10016 12808 10044
rect 12802 10004 12808 10016
rect 12860 10004 12866 10056
rect 15194 10004 15200 10056
rect 15252 10044 15258 10056
rect 15933 10047 15991 10053
rect 15933 10044 15945 10047
rect 15252 10016 15945 10044
rect 15252 10004 15258 10016
rect 15933 10013 15945 10016
rect 15979 10013 15991 10047
rect 23014 10044 23020 10056
rect 22975 10016 23020 10044
rect 15933 10007 15991 10013
rect 23014 10004 23020 10016
rect 23072 10004 23078 10056
rect 23106 10004 23112 10056
rect 23164 10044 23170 10056
rect 25314 10044 25320 10056
rect 23164 10016 23209 10044
rect 25275 10016 25320 10044
rect 23164 10004 23170 10016
rect 25314 10004 25320 10016
rect 25372 10004 25378 10056
rect 25498 10044 25504 10056
rect 25459 10016 25504 10044
rect 25498 10004 25504 10016
rect 25556 10004 25562 10056
rect 28994 10004 29000 10056
rect 29052 10044 29058 10056
rect 29089 10047 29147 10053
rect 29089 10044 29101 10047
rect 29052 10016 29101 10044
rect 29052 10004 29058 10016
rect 29089 10013 29101 10016
rect 29135 10013 29147 10047
rect 35342 10044 35348 10056
rect 35303 10016 35348 10044
rect 29089 10007 29147 10013
rect 35342 10004 35348 10016
rect 35400 10004 35406 10056
rect 38381 10047 38439 10053
rect 38381 10013 38393 10047
rect 38427 10044 38439 10047
rect 38562 10044 38568 10056
rect 38427 10016 38568 10044
rect 38427 10013 38439 10016
rect 38381 10007 38439 10013
rect 38562 10004 38568 10016
rect 38620 10004 38626 10056
rect 6546 9976 6552 9988
rect 6507 9948 6552 9976
rect 6546 9936 6552 9948
rect 6604 9936 6610 9988
rect 7024 9976 7052 10004
rect 7561 9979 7619 9985
rect 7561 9976 7573 9979
rect 7024 9948 7573 9976
rect 7561 9945 7573 9948
rect 7607 9945 7619 9979
rect 7561 9939 7619 9945
rect 10686 9936 10692 9988
rect 10744 9976 10750 9988
rect 12253 9979 12311 9985
rect 12253 9976 12265 9979
rect 10744 9948 12265 9976
rect 10744 9936 10750 9948
rect 12253 9945 12265 9948
rect 12299 9945 12311 9979
rect 12253 9939 12311 9945
rect 24765 9979 24823 9985
rect 24765 9945 24777 9979
rect 24811 9976 24823 9979
rect 25516 9976 25544 10004
rect 37826 9976 37832 9988
rect 24811 9948 25544 9976
rect 37787 9948 37832 9976
rect 24811 9945 24823 9948
rect 24765 9939 24823 9945
rect 37826 9936 37832 9948
rect 37884 9936 37890 9988
rect 43456 9985 43484 10084
rect 45824 10075 45836 10084
rect 45830 10072 45836 10075
rect 45888 10072 45894 10124
rect 43622 10004 43628 10056
rect 43680 10044 43686 10056
rect 43993 10047 44051 10053
rect 43993 10044 44005 10047
rect 43680 10016 44005 10044
rect 43680 10004 43686 10016
rect 43993 10013 44005 10016
rect 44039 10013 44051 10047
rect 45554 10044 45560 10056
rect 45515 10016 45560 10044
rect 43993 10007 44051 10013
rect 45554 10004 45560 10016
rect 45612 10004 45618 10056
rect 43441 9979 43499 9985
rect 43441 9945 43453 9979
rect 43487 9945 43499 9979
rect 43441 9939 43499 9945
rect 2041 9911 2099 9917
rect 2041 9877 2053 9911
rect 2087 9908 2099 9911
rect 2682 9908 2688 9920
rect 2087 9880 2688 9908
rect 2087 9877 2099 9880
rect 2041 9871 2099 9877
rect 2682 9868 2688 9880
rect 2740 9868 2746 9920
rect 4706 9908 4712 9920
rect 4667 9880 4712 9908
rect 4706 9868 4712 9880
rect 4764 9908 4770 9920
rect 5442 9908 5448 9920
rect 4764 9880 5448 9908
rect 4764 9868 4770 9880
rect 5442 9868 5448 9880
rect 5500 9868 5506 9920
rect 7190 9868 7196 9920
rect 7248 9908 7254 9920
rect 8113 9911 8171 9917
rect 8113 9908 8125 9911
rect 7248 9880 8125 9908
rect 7248 9868 7254 9880
rect 8113 9877 8125 9880
rect 8159 9877 8171 9911
rect 11054 9908 11060 9920
rect 11015 9880 11060 9908
rect 8113 9871 8171 9877
rect 11054 9868 11060 9880
rect 11112 9868 11118 9920
rect 15378 9908 15384 9920
rect 15339 9880 15384 9908
rect 15378 9868 15384 9880
rect 15436 9868 15442 9920
rect 22557 9911 22615 9917
rect 22557 9877 22569 9911
rect 22603 9908 22615 9911
rect 23566 9908 23572 9920
rect 22603 9880 23572 9908
rect 22603 9877 22615 9880
rect 22557 9871 22615 9877
rect 23566 9868 23572 9880
rect 23624 9868 23630 9920
rect 24946 9908 24952 9920
rect 24907 9880 24952 9908
rect 24946 9868 24952 9880
rect 25004 9868 25010 9920
rect 28534 9908 28540 9920
rect 28495 9880 28540 9908
rect 28534 9868 28540 9880
rect 28592 9868 28598 9920
rect 29546 9908 29552 9920
rect 29459 9880 29552 9908
rect 29546 9868 29552 9880
rect 29604 9908 29610 9920
rect 30006 9908 30012 9920
rect 29604 9880 30012 9908
rect 29604 9868 29610 9880
rect 30006 9868 30012 9880
rect 30064 9868 30070 9920
rect 34977 9911 35035 9917
rect 34977 9877 34989 9911
rect 35023 9908 35035 9911
rect 35434 9908 35440 9920
rect 35023 9880 35440 9908
rect 35023 9877 35035 9880
rect 34977 9871 35035 9877
rect 35434 9868 35440 9880
rect 35492 9868 35498 9920
rect 41509 9911 41567 9917
rect 41509 9877 41521 9911
rect 41555 9908 41567 9911
rect 41966 9908 41972 9920
rect 41555 9880 41972 9908
rect 41555 9877 41567 9880
rect 41509 9871 41567 9877
rect 41966 9868 41972 9880
rect 42024 9868 42030 9920
rect 44266 9868 44272 9920
rect 44324 9908 44330 9920
rect 44545 9911 44603 9917
rect 44545 9908 44557 9911
rect 44324 9880 44557 9908
rect 44324 9868 44330 9880
rect 44545 9877 44557 9880
rect 44591 9908 44603 9911
rect 45094 9908 45100 9920
rect 44591 9880 45100 9908
rect 44591 9877 44603 9880
rect 44545 9871 44603 9877
rect 45094 9868 45100 9880
rect 45152 9868 45158 9920
rect 1104 9818 48852 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 34966 9818
rect 35018 9766 35030 9818
rect 35082 9766 35094 9818
rect 35146 9766 35158 9818
rect 35210 9766 48852 9818
rect 1104 9744 48852 9766
rect 2498 9664 2504 9716
rect 2556 9704 2562 9716
rect 5350 9704 5356 9716
rect 2556 9676 2728 9704
rect 5311 9676 5356 9704
rect 2556 9664 2562 9676
rect 2700 9636 2728 9676
rect 5350 9664 5356 9676
rect 5408 9664 5414 9716
rect 5629 9707 5687 9713
rect 5629 9673 5641 9707
rect 5675 9704 5687 9707
rect 5902 9704 5908 9716
rect 5675 9676 5908 9704
rect 5675 9673 5687 9676
rect 5629 9667 5687 9673
rect 5902 9664 5908 9676
rect 5960 9664 5966 9716
rect 7006 9704 7012 9716
rect 6967 9676 7012 9704
rect 7006 9664 7012 9676
rect 7064 9664 7070 9716
rect 8478 9664 8484 9716
rect 8536 9704 8542 9716
rect 8941 9707 8999 9713
rect 8941 9704 8953 9707
rect 8536 9676 8953 9704
rect 8536 9664 8542 9676
rect 8941 9673 8953 9676
rect 8987 9673 8999 9707
rect 8941 9667 8999 9673
rect 12526 9664 12532 9716
rect 12584 9704 12590 9716
rect 12621 9707 12679 9713
rect 12621 9704 12633 9707
rect 12584 9676 12633 9704
rect 12584 9664 12590 9676
rect 12621 9673 12633 9676
rect 12667 9673 12679 9707
rect 12621 9667 12679 9673
rect 12802 9664 12808 9716
rect 12860 9704 12866 9716
rect 12989 9707 13047 9713
rect 12989 9704 13001 9707
rect 12860 9676 13001 9704
rect 12860 9664 12866 9676
rect 12989 9673 13001 9676
rect 13035 9673 13047 9707
rect 12989 9667 13047 9673
rect 15654 9664 15660 9716
rect 15712 9704 15718 9716
rect 20993 9707 21051 9713
rect 15712 9676 16528 9704
rect 15712 9664 15718 9676
rect 2774 9636 2780 9648
rect 2700 9608 2780 9636
rect 2774 9596 2780 9608
rect 2832 9636 2838 9648
rect 3973 9639 4031 9645
rect 2832 9608 2925 9636
rect 2832 9596 2838 9608
rect 3973 9605 3985 9639
rect 4019 9636 4031 9639
rect 4614 9636 4620 9648
rect 4019 9608 4620 9636
rect 4019 9605 4031 9608
rect 3973 9599 4031 9605
rect 4614 9596 4620 9608
rect 4672 9636 4678 9648
rect 4893 9639 4951 9645
rect 4893 9636 4905 9639
rect 4672 9608 4905 9636
rect 4672 9596 4678 9608
rect 4893 9605 4905 9608
rect 4939 9605 4951 9639
rect 4893 9599 4951 9605
rect 2682 9528 2688 9580
rect 2740 9568 2746 9580
rect 3697 9571 3755 9577
rect 3697 9568 3709 9571
rect 2740 9540 3709 9568
rect 2740 9528 2746 9540
rect 3697 9537 3709 9540
rect 3743 9568 3755 9571
rect 7024 9568 7052 9664
rect 11425 9639 11483 9645
rect 11425 9605 11437 9639
rect 11471 9636 11483 9639
rect 12820 9636 12848 9664
rect 11471 9608 12848 9636
rect 16500 9636 16528 9676
rect 20993 9673 21005 9707
rect 21039 9704 21051 9707
rect 21450 9704 21456 9716
rect 21039 9676 21456 9704
rect 21039 9673 21051 9676
rect 20993 9667 21051 9673
rect 21450 9664 21456 9676
rect 21508 9664 21514 9716
rect 21726 9704 21732 9716
rect 21687 9676 21732 9704
rect 21726 9664 21732 9676
rect 21784 9664 21790 9716
rect 22557 9707 22615 9713
rect 22557 9673 22569 9707
rect 22603 9704 22615 9707
rect 23014 9704 23020 9716
rect 22603 9676 23020 9704
rect 22603 9673 22615 9676
rect 22557 9667 22615 9673
rect 23014 9664 23020 9676
rect 23072 9664 23078 9716
rect 23198 9704 23204 9716
rect 23159 9676 23204 9704
rect 23198 9664 23204 9676
rect 23256 9664 23262 9716
rect 25406 9704 25412 9716
rect 25148 9676 25412 9704
rect 16666 9636 16672 9648
rect 16500 9608 16672 9636
rect 11471 9605 11483 9608
rect 11425 9599 11483 9605
rect 16666 9596 16672 9608
rect 16724 9636 16730 9648
rect 16853 9639 16911 9645
rect 16853 9636 16865 9639
rect 16724 9608 16865 9636
rect 16724 9596 16730 9608
rect 16853 9605 16865 9608
rect 16899 9605 16911 9639
rect 21266 9636 21272 9648
rect 21227 9608 21272 9636
rect 16853 9599 16911 9605
rect 21266 9596 21272 9608
rect 21324 9596 21330 9648
rect 21468 9636 21496 9664
rect 21910 9636 21916 9648
rect 21468 9608 21916 9636
rect 21910 9596 21916 9608
rect 21968 9596 21974 9648
rect 22925 9639 22983 9645
rect 22925 9605 22937 9639
rect 22971 9636 22983 9639
rect 23106 9636 23112 9648
rect 22971 9608 23112 9636
rect 22971 9605 22983 9608
rect 22925 9599 22983 9605
rect 23106 9596 23112 9608
rect 23164 9596 23170 9648
rect 24578 9596 24584 9648
rect 24636 9636 24642 9648
rect 24765 9639 24823 9645
rect 24765 9636 24777 9639
rect 24636 9608 24777 9636
rect 24636 9596 24642 9608
rect 24765 9605 24777 9608
rect 24811 9636 24823 9639
rect 25148 9636 25176 9676
rect 25406 9664 25412 9676
rect 25464 9664 25470 9716
rect 27617 9707 27675 9713
rect 27617 9673 27629 9707
rect 27663 9704 27675 9707
rect 27798 9704 27804 9716
rect 27663 9676 27804 9704
rect 27663 9673 27675 9676
rect 27617 9667 27675 9673
rect 27798 9664 27804 9676
rect 27856 9704 27862 9716
rect 28534 9704 28540 9716
rect 27856 9676 28540 9704
rect 27856 9664 27862 9676
rect 28534 9664 28540 9676
rect 28592 9664 28598 9716
rect 28718 9704 28724 9716
rect 28679 9676 28724 9704
rect 28718 9664 28724 9676
rect 28776 9664 28782 9716
rect 28810 9664 28816 9716
rect 28868 9704 28874 9716
rect 28868 9676 28948 9704
rect 28868 9664 28874 9676
rect 27154 9636 27160 9648
rect 24811 9608 25176 9636
rect 27115 9608 27160 9636
rect 24811 9605 24823 9608
rect 24765 9599 24823 9605
rect 27154 9596 27160 9608
rect 27212 9596 27218 9648
rect 28920 9636 28948 9676
rect 29270 9664 29276 9716
rect 29328 9704 29334 9716
rect 29917 9707 29975 9713
rect 29917 9704 29929 9707
rect 29328 9676 29929 9704
rect 29328 9664 29334 9676
rect 29917 9673 29929 9676
rect 29963 9673 29975 9707
rect 29917 9667 29975 9673
rect 28997 9639 29055 9645
rect 28997 9636 29009 9639
rect 28920 9608 29009 9636
rect 28997 9605 29009 9608
rect 29043 9605 29055 9639
rect 28997 9599 29055 9605
rect 12253 9571 12311 9577
rect 3743 9540 4476 9568
rect 7024 9540 7696 9568
rect 3743 9537 3755 9540
rect 3697 9531 3755 9537
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9500 1455 9503
rect 1486 9500 1492 9512
rect 1443 9472 1492 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 1486 9460 1492 9472
rect 1544 9460 1550 9512
rect 1664 9503 1722 9509
rect 1664 9469 1676 9503
rect 1710 9500 1722 9503
rect 2406 9500 2412 9512
rect 1710 9472 2412 9500
rect 1710 9469 1722 9472
rect 1664 9463 1722 9469
rect 2406 9460 2412 9472
rect 2464 9460 2470 9512
rect 3421 9435 3479 9441
rect 3421 9401 3433 9435
rect 3467 9432 3479 9435
rect 4154 9432 4160 9444
rect 3467 9404 4160 9432
rect 3467 9401 3479 9404
rect 3421 9395 3479 9401
rect 4154 9392 4160 9404
rect 4212 9432 4218 9444
rect 4448 9441 4476 9540
rect 4982 9460 4988 9512
rect 5040 9500 5046 9512
rect 5445 9503 5503 9509
rect 5445 9500 5457 9503
rect 5040 9472 5457 9500
rect 5040 9460 5046 9472
rect 5445 9469 5457 9472
rect 5491 9500 5503 9503
rect 5997 9503 6055 9509
rect 5997 9500 6009 9503
rect 5491 9472 6009 9500
rect 5491 9469 5503 9472
rect 5445 9463 5503 9469
rect 5997 9469 6009 9472
rect 6043 9469 6055 9503
rect 5997 9463 6055 9469
rect 7561 9503 7619 9509
rect 7561 9469 7573 9503
rect 7607 9469 7619 9503
rect 7668 9500 7696 9540
rect 12253 9537 12265 9571
rect 12299 9568 12311 9571
rect 12342 9568 12348 9580
rect 12299 9540 12348 9568
rect 12299 9537 12311 9540
rect 12253 9531 12311 9537
rect 12342 9528 12348 9540
rect 12400 9528 12406 9580
rect 29932 9568 29960 9667
rect 34238 9664 34244 9716
rect 34296 9704 34302 9716
rect 34609 9707 34667 9713
rect 34609 9704 34621 9707
rect 34296 9676 34621 9704
rect 34296 9664 34302 9676
rect 34609 9673 34621 9676
rect 34655 9673 34667 9707
rect 34609 9667 34667 9673
rect 34790 9664 34796 9716
rect 34848 9704 34854 9716
rect 35345 9707 35403 9713
rect 35345 9704 35357 9707
rect 34848 9676 35357 9704
rect 34848 9664 34854 9676
rect 35345 9673 35357 9676
rect 35391 9673 35403 9707
rect 37734 9704 37740 9716
rect 37695 9676 37740 9704
rect 35345 9667 35403 9673
rect 34333 9639 34391 9645
rect 34333 9605 34345 9639
rect 34379 9636 34391 9639
rect 34514 9636 34520 9648
rect 34379 9608 34520 9636
rect 34379 9605 34391 9608
rect 34333 9599 34391 9605
rect 34514 9596 34520 9608
rect 34572 9596 34578 9648
rect 30098 9568 30104 9580
rect 29932 9540 30104 9568
rect 30098 9528 30104 9540
rect 30156 9528 30162 9580
rect 35360 9568 35388 9667
rect 37734 9664 37740 9676
rect 37792 9664 37798 9716
rect 40770 9704 40776 9716
rect 40731 9676 40776 9704
rect 40770 9664 40776 9676
rect 40828 9664 40834 9716
rect 41414 9664 41420 9716
rect 41472 9704 41478 9716
rect 41690 9704 41696 9716
rect 41472 9676 41696 9704
rect 41472 9664 41478 9676
rect 41690 9664 41696 9676
rect 41748 9664 41754 9716
rect 43438 9664 43444 9716
rect 43496 9704 43502 9716
rect 43717 9707 43775 9713
rect 43717 9704 43729 9707
rect 43496 9676 43729 9704
rect 43496 9664 43502 9676
rect 43717 9673 43729 9676
rect 43763 9673 43775 9707
rect 43717 9667 43775 9673
rect 42337 9639 42395 9645
rect 42337 9605 42349 9639
rect 42383 9636 42395 9639
rect 42794 9636 42800 9648
rect 42383 9608 42800 9636
rect 42383 9605 42395 9608
rect 42337 9599 42395 9605
rect 42794 9596 42800 9608
rect 42852 9596 42858 9648
rect 43349 9639 43407 9645
rect 43349 9605 43361 9639
rect 43395 9636 43407 9639
rect 43898 9636 43904 9648
rect 43395 9608 43904 9636
rect 43395 9605 43407 9608
rect 43349 9599 43407 9605
rect 43898 9596 43904 9608
rect 43956 9636 43962 9648
rect 44545 9639 44603 9645
rect 44545 9636 44557 9639
rect 43956 9608 44557 9636
rect 43956 9596 43962 9608
rect 44545 9605 44557 9608
rect 44591 9605 44603 9639
rect 46934 9636 46940 9648
rect 46895 9608 46940 9636
rect 44545 9599 44603 9605
rect 46934 9596 46940 9608
rect 46992 9596 46998 9648
rect 47394 9636 47400 9648
rect 47355 9608 47400 9636
rect 47394 9596 47400 9608
rect 47452 9596 47458 9648
rect 35526 9568 35532 9580
rect 35360 9540 35532 9568
rect 35526 9528 35532 9540
rect 35584 9528 35590 9580
rect 41690 9528 41696 9580
rect 41748 9568 41754 9580
rect 42058 9568 42064 9580
rect 41748 9540 42064 9568
rect 41748 9528 41754 9540
rect 42058 9528 42064 9540
rect 42116 9528 42122 9580
rect 7834 9509 7840 9512
rect 7817 9503 7840 9509
rect 7817 9500 7829 9503
rect 7668 9472 7829 9500
rect 7561 9463 7619 9469
rect 7817 9469 7829 9472
rect 7892 9500 7898 9512
rect 10413 9503 10471 9509
rect 7892 9472 7965 9500
rect 7817 9463 7840 9469
rect 4249 9435 4307 9441
rect 4249 9432 4261 9435
rect 4212 9404 4261 9432
rect 4212 9392 4218 9404
rect 4249 9401 4261 9404
rect 4295 9401 4307 9435
rect 4249 9395 4307 9401
rect 4433 9435 4491 9441
rect 4433 9401 4445 9435
rect 4479 9401 4491 9435
rect 4433 9395 4491 9401
rect 4525 9435 4583 9441
rect 4525 9401 4537 9435
rect 4571 9432 4583 9435
rect 4706 9432 4712 9444
rect 4571 9404 4712 9432
rect 4571 9401 4583 9404
rect 4525 9395 4583 9401
rect 3970 9324 3976 9376
rect 4028 9364 4034 9376
rect 4540 9364 4568 9395
rect 4706 9392 4712 9404
rect 4764 9392 4770 9444
rect 6454 9392 6460 9444
rect 6512 9432 6518 9444
rect 7377 9435 7435 9441
rect 7377 9432 7389 9435
rect 6512 9404 7389 9432
rect 6512 9392 6518 9404
rect 7377 9401 7389 9404
rect 7423 9432 7435 9435
rect 7576 9432 7604 9463
rect 7834 9460 7840 9463
rect 7892 9460 7898 9472
rect 10413 9469 10425 9503
rect 10459 9500 10471 9503
rect 11241 9503 11299 9509
rect 11241 9500 11253 9503
rect 10459 9472 11253 9500
rect 10459 9469 10471 9472
rect 10413 9463 10471 9469
rect 11241 9469 11253 9472
rect 11287 9500 11299 9503
rect 11793 9503 11851 9509
rect 11793 9500 11805 9503
rect 11287 9472 11805 9500
rect 11287 9469 11299 9472
rect 11241 9463 11299 9469
rect 11793 9469 11805 9472
rect 11839 9469 11851 9503
rect 11793 9463 11851 9469
rect 14461 9503 14519 9509
rect 14461 9469 14473 9503
rect 14507 9500 14519 9503
rect 14553 9503 14611 9509
rect 14553 9500 14565 9503
rect 14507 9472 14565 9500
rect 14507 9469 14519 9472
rect 14461 9463 14519 9469
rect 14553 9469 14565 9472
rect 14599 9500 14611 9503
rect 15286 9500 15292 9512
rect 14599 9472 15292 9500
rect 14599 9469 14611 9472
rect 14553 9463 14611 9469
rect 15286 9460 15292 9472
rect 15344 9500 15350 9512
rect 15562 9500 15568 9512
rect 15344 9472 15568 9500
rect 15344 9460 15350 9472
rect 15562 9460 15568 9472
rect 15620 9460 15626 9512
rect 24949 9503 25007 9509
rect 24949 9469 24961 9503
rect 24995 9500 25007 9503
rect 25225 9503 25283 9509
rect 25225 9500 25237 9503
rect 24995 9472 25237 9500
rect 24995 9469 25007 9472
rect 24949 9463 25007 9469
rect 25225 9469 25237 9472
rect 25271 9469 25283 9503
rect 28077 9503 28135 9509
rect 28077 9500 28089 9503
rect 25225 9463 25283 9469
rect 27908 9472 28089 9500
rect 7423 9404 7604 9432
rect 7423 9401 7435 9404
rect 7377 9395 7435 9401
rect 9950 9392 9956 9444
rect 10008 9432 10014 9444
rect 10045 9435 10103 9441
rect 10045 9432 10057 9435
rect 10008 9404 10057 9432
rect 10008 9392 10014 9404
rect 10045 9401 10057 9404
rect 10091 9401 10103 9435
rect 10045 9395 10103 9401
rect 6546 9364 6552 9376
rect 4028 9336 4568 9364
rect 6507 9336 6552 9364
rect 4028 9324 4034 9336
rect 6546 9324 6552 9336
rect 6604 9364 6610 9376
rect 7098 9364 7104 9376
rect 6604 9336 7104 9364
rect 6604 9324 6610 9336
rect 7098 9324 7104 9336
rect 7156 9324 7162 9376
rect 9674 9364 9680 9376
rect 9635 9336 9680 9364
rect 9674 9324 9680 9336
rect 9732 9324 9738 9376
rect 10060 9364 10088 9395
rect 10134 9392 10140 9444
rect 10192 9432 10198 9444
rect 10229 9435 10287 9441
rect 10229 9432 10241 9435
rect 10192 9404 10241 9432
rect 10192 9392 10198 9404
rect 10229 9401 10241 9404
rect 10275 9432 10287 9435
rect 10962 9432 10968 9444
rect 10275 9404 10968 9432
rect 10275 9401 10287 9404
rect 10229 9395 10287 9401
rect 10962 9392 10968 9404
rect 11020 9392 11026 9444
rect 14642 9392 14648 9444
rect 14700 9432 14706 9444
rect 14798 9435 14856 9441
rect 14798 9432 14810 9435
rect 14700 9404 14810 9432
rect 14700 9392 14706 9404
rect 14798 9401 14810 9404
rect 14844 9401 14856 9435
rect 14798 9395 14856 9401
rect 24029 9435 24087 9441
rect 24029 9401 24041 9435
rect 24075 9432 24087 9435
rect 24397 9435 24455 9441
rect 24397 9432 24409 9435
rect 24075 9404 24409 9432
rect 24075 9401 24087 9404
rect 24029 9395 24087 9401
rect 24397 9401 24409 9404
rect 24443 9432 24455 9435
rect 25314 9432 25320 9444
rect 24443 9404 25320 9432
rect 24443 9401 24455 9404
rect 24397 9395 24455 9401
rect 25314 9392 25320 9404
rect 25372 9432 25378 9444
rect 25492 9435 25550 9441
rect 25492 9432 25504 9435
rect 25372 9404 25504 9432
rect 25372 9392 25378 9404
rect 25492 9401 25504 9404
rect 25538 9432 25550 9435
rect 26050 9432 26056 9444
rect 25538 9404 26056 9432
rect 25538 9401 25550 9404
rect 25492 9395 25550 9401
rect 26050 9392 26056 9404
rect 26108 9392 26114 9444
rect 27908 9376 27936 9472
rect 28077 9469 28089 9472
rect 28123 9469 28135 9503
rect 28077 9463 28135 9469
rect 40770 9460 40776 9512
rect 40828 9500 40834 9512
rect 41417 9503 41475 9509
rect 41417 9500 41429 9503
rect 40828 9472 41429 9500
rect 40828 9460 40834 9472
rect 41417 9469 41429 9472
rect 41463 9500 41475 9503
rect 42889 9503 42947 9509
rect 42889 9500 42901 9503
rect 41463 9472 42901 9500
rect 41463 9469 41475 9472
rect 41417 9463 41475 9469
rect 42889 9469 42901 9472
rect 42935 9500 42947 9503
rect 43162 9500 43168 9512
rect 42935 9472 43168 9500
rect 42935 9469 42947 9472
rect 42889 9463 42947 9469
rect 43162 9460 43168 9472
rect 43220 9500 43226 9512
rect 44266 9500 44272 9512
rect 43220 9472 44272 9500
rect 43220 9460 43226 9472
rect 44266 9460 44272 9472
rect 44324 9460 44330 9512
rect 45830 9500 45836 9512
rect 44836 9472 45836 9500
rect 44836 9444 44864 9472
rect 45830 9460 45836 9472
rect 45888 9500 45894 9512
rect 46293 9503 46351 9509
rect 46293 9500 46305 9503
rect 45888 9472 46305 9500
rect 45888 9460 45894 9472
rect 46293 9469 46305 9472
rect 46339 9500 46351 9503
rect 46474 9500 46480 9512
rect 46339 9472 46480 9500
rect 46339 9469 46351 9472
rect 46293 9463 46351 9469
rect 46474 9460 46480 9472
rect 46532 9460 46538 9512
rect 46753 9503 46811 9509
rect 46753 9469 46765 9503
rect 46799 9500 46811 9503
rect 47412 9500 47440 9596
rect 46799 9472 47440 9500
rect 46799 9469 46811 9472
rect 46753 9463 46811 9469
rect 30374 9441 30380 9444
rect 30368 9432 30380 9441
rect 30335 9404 30380 9432
rect 30368 9395 30380 9404
rect 30374 9392 30380 9395
rect 30432 9392 30438 9444
rect 35796 9435 35854 9441
rect 35796 9401 35808 9435
rect 35842 9432 35854 9435
rect 36354 9432 36360 9444
rect 35842 9404 36360 9432
rect 35842 9401 35854 9404
rect 35796 9395 35854 9401
rect 36354 9392 36360 9404
rect 36412 9392 36418 9444
rect 41785 9435 41843 9441
rect 41785 9401 41797 9435
rect 41831 9432 41843 9435
rect 42610 9432 42616 9444
rect 41831 9404 42616 9432
rect 41831 9401 41843 9404
rect 41785 9395 41843 9401
rect 42610 9392 42616 9404
rect 42668 9392 42674 9444
rect 44818 9432 44824 9444
rect 44779 9404 44824 9432
rect 44818 9392 44824 9404
rect 44876 9392 44882 9444
rect 45094 9432 45100 9444
rect 45055 9404 45100 9432
rect 45094 9392 45100 9404
rect 45152 9392 45158 9444
rect 10689 9367 10747 9373
rect 10689 9364 10701 9367
rect 10060 9336 10701 9364
rect 10689 9333 10701 9336
rect 10735 9333 10747 9367
rect 15930 9364 15936 9376
rect 15891 9336 15936 9364
rect 10689 9327 10747 9333
rect 15930 9324 15936 9336
rect 15988 9364 15994 9376
rect 16485 9367 16543 9373
rect 16485 9364 16497 9367
rect 15988 9336 16497 9364
rect 15988 9324 15994 9336
rect 16485 9333 16497 9336
rect 16531 9333 16543 9367
rect 16485 9327 16543 9333
rect 24670 9324 24676 9376
rect 24728 9364 24734 9376
rect 24949 9367 25007 9373
rect 24949 9364 24961 9367
rect 24728 9336 24961 9364
rect 24728 9324 24734 9336
rect 24949 9333 24961 9336
rect 24995 9364 25007 9367
rect 25041 9367 25099 9373
rect 25041 9364 25053 9367
rect 24995 9336 25053 9364
rect 24995 9333 25007 9336
rect 24949 9327 25007 9333
rect 25041 9333 25053 9336
rect 25087 9333 25099 9367
rect 26602 9364 26608 9376
rect 26563 9336 26608 9364
rect 25041 9327 25099 9333
rect 26602 9324 26608 9336
rect 26660 9324 26666 9376
rect 27890 9364 27896 9376
rect 27851 9336 27896 9364
rect 27890 9324 27896 9336
rect 27948 9324 27954 9376
rect 28258 9364 28264 9376
rect 28219 9336 28264 9364
rect 28258 9324 28264 9336
rect 28316 9324 28322 9376
rect 30006 9324 30012 9376
rect 30064 9364 30070 9376
rect 31481 9367 31539 9373
rect 31481 9364 31493 9367
rect 30064 9336 31493 9364
rect 30064 9324 30070 9336
rect 31481 9333 31493 9336
rect 31527 9333 31539 9367
rect 31481 9327 31539 9333
rect 36446 9324 36452 9376
rect 36504 9364 36510 9376
rect 36909 9367 36967 9373
rect 36909 9364 36921 9367
rect 36504 9336 36921 9364
rect 36504 9324 36510 9336
rect 36909 9333 36921 9336
rect 36955 9333 36967 9367
rect 38102 9364 38108 9376
rect 38063 9336 38108 9364
rect 36909 9327 36967 9333
rect 38102 9324 38108 9336
rect 38160 9324 38166 9376
rect 38562 9364 38568 9376
rect 38523 9336 38568 9364
rect 38562 9324 38568 9336
rect 38620 9324 38626 9376
rect 38654 9324 38660 9376
rect 38712 9364 38718 9376
rect 39298 9364 39304 9376
rect 38712 9336 39304 9364
rect 38712 9324 38718 9336
rect 39298 9324 39304 9336
rect 39356 9324 39362 9376
rect 42153 9367 42211 9373
rect 42153 9333 42165 9367
rect 42199 9364 42211 9367
rect 42518 9364 42524 9376
rect 42199 9336 42524 9364
rect 42199 9333 42211 9336
rect 42153 9327 42211 9333
rect 42518 9324 42524 9336
rect 42576 9364 42582 9376
rect 42797 9367 42855 9373
rect 42797 9364 42809 9367
rect 42576 9336 42809 9364
rect 42576 9324 42582 9336
rect 42797 9333 42809 9336
rect 42843 9333 42855 9367
rect 42797 9327 42855 9333
rect 44361 9367 44419 9373
rect 44361 9333 44373 9367
rect 44407 9364 44419 9367
rect 45002 9364 45008 9376
rect 44407 9336 45008 9364
rect 44407 9333 44419 9336
rect 44361 9327 44419 9333
rect 45002 9324 45008 9336
rect 45060 9324 45066 9376
rect 45186 9324 45192 9376
rect 45244 9364 45250 9376
rect 45554 9364 45560 9376
rect 45244 9336 45560 9364
rect 45244 9324 45250 9336
rect 45554 9324 45560 9336
rect 45612 9324 45618 9376
rect 1104 9274 48852 9296
rect 1104 9222 19606 9274
rect 19658 9222 19670 9274
rect 19722 9222 19734 9274
rect 19786 9222 19798 9274
rect 19850 9222 48852 9274
rect 1104 9200 48852 9222
rect 1486 9120 1492 9172
rect 1544 9160 1550 9172
rect 1581 9163 1639 9169
rect 1581 9160 1593 9163
rect 1544 9132 1593 9160
rect 1544 9120 1550 9132
rect 1581 9129 1593 9132
rect 1627 9129 1639 9163
rect 1581 9123 1639 9129
rect 2041 9163 2099 9169
rect 2041 9129 2053 9163
rect 2087 9160 2099 9163
rect 2406 9160 2412 9172
rect 2087 9132 2412 9160
rect 2087 9129 2099 9132
rect 2041 9123 2099 9129
rect 2406 9120 2412 9132
rect 2464 9120 2470 9172
rect 2774 9120 2780 9172
rect 2832 9160 2838 9172
rect 7834 9160 7840 9172
rect 2832 9132 2877 9160
rect 7795 9132 7840 9160
rect 2832 9120 2838 9132
rect 7834 9120 7840 9132
rect 7892 9120 7898 9172
rect 8478 9160 8484 9172
rect 8439 9132 8484 9160
rect 8478 9120 8484 9132
rect 8536 9120 8542 9172
rect 8849 9163 8907 9169
rect 8849 9129 8861 9163
rect 8895 9160 8907 9163
rect 10410 9160 10416 9172
rect 8895 9132 10416 9160
rect 8895 9129 8907 9132
rect 8849 9123 8907 9129
rect 10410 9120 10416 9132
rect 10468 9120 10474 9172
rect 16666 9160 16672 9172
rect 16627 9132 16672 9160
rect 16666 9120 16672 9132
rect 16724 9120 16730 9172
rect 26050 9160 26056 9172
rect 26011 9132 26056 9160
rect 26050 9120 26056 9132
rect 26108 9120 26114 9172
rect 26602 9120 26608 9172
rect 26660 9160 26666 9172
rect 27065 9163 27123 9169
rect 27065 9160 27077 9163
rect 26660 9132 27077 9160
rect 26660 9120 26666 9132
rect 27065 9129 27077 9132
rect 27111 9129 27123 9163
rect 27065 9123 27123 9129
rect 29546 9120 29552 9172
rect 29604 9160 29610 9172
rect 29641 9163 29699 9169
rect 29641 9160 29653 9163
rect 29604 9132 29653 9160
rect 29604 9120 29610 9132
rect 29641 9129 29653 9132
rect 29687 9160 29699 9163
rect 30193 9163 30251 9169
rect 30193 9160 30205 9163
rect 29687 9132 30205 9160
rect 29687 9129 29699 9132
rect 29641 9123 29699 9129
rect 30193 9129 30205 9132
rect 30239 9160 30251 9163
rect 30374 9160 30380 9172
rect 30239 9132 30380 9160
rect 30239 9129 30251 9132
rect 30193 9123 30251 9129
rect 30374 9120 30380 9132
rect 30432 9160 30438 9172
rect 33505 9163 33563 9169
rect 33505 9160 33517 9163
rect 30432 9132 33517 9160
rect 30432 9120 30438 9132
rect 33505 9129 33517 9132
rect 33551 9129 33563 9163
rect 33505 9123 33563 9129
rect 34977 9163 35035 9169
rect 34977 9129 34989 9163
rect 35023 9160 35035 9163
rect 35342 9160 35348 9172
rect 35023 9132 35348 9160
rect 35023 9129 35035 9132
rect 34977 9123 35035 9129
rect 35342 9120 35348 9132
rect 35400 9120 35406 9172
rect 35621 9163 35679 9169
rect 35621 9129 35633 9163
rect 35667 9160 35679 9163
rect 35986 9160 35992 9172
rect 35667 9132 35992 9160
rect 35667 9129 35679 9132
rect 35621 9123 35679 9129
rect 35986 9120 35992 9132
rect 36044 9160 36050 9172
rect 36354 9160 36360 9172
rect 36044 9132 36360 9160
rect 36044 9120 36050 9132
rect 36354 9120 36360 9132
rect 36412 9160 36418 9172
rect 36449 9163 36507 9169
rect 36449 9160 36461 9163
rect 36412 9132 36461 9160
rect 36412 9120 36418 9132
rect 36449 9129 36461 9132
rect 36495 9129 36507 9163
rect 40034 9160 40040 9172
rect 36449 9123 36507 9129
rect 38948 9132 39436 9160
rect 39947 9132 40040 9160
rect 38948 9104 38976 9132
rect 4614 9092 4620 9104
rect 4575 9064 4620 9092
rect 4614 9052 4620 9064
rect 4672 9052 4678 9104
rect 7282 9092 7288 9104
rect 6288 9064 7288 9092
rect 2038 8984 2044 9036
rect 2096 9024 2102 9036
rect 4709 9027 4767 9033
rect 4709 9024 4721 9027
rect 2096 8996 4721 9024
rect 2096 8984 2102 8996
rect 4709 8993 4721 8996
rect 4755 9024 4767 9027
rect 5166 9024 5172 9036
rect 4755 8996 5172 9024
rect 4755 8993 4767 8996
rect 4709 8987 4767 8993
rect 5166 8984 5172 8996
rect 5224 9024 5230 9036
rect 6288 9033 6316 9064
rect 7282 9052 7288 9064
rect 7340 9052 7346 9104
rect 10134 9092 10140 9104
rect 10095 9064 10140 9092
rect 10134 9052 10140 9064
rect 10192 9052 10198 9104
rect 12250 9101 12256 9104
rect 12244 9092 12256 9101
rect 12211 9064 12256 9092
rect 12244 9055 12256 9064
rect 12250 9052 12256 9055
rect 12308 9052 12314 9104
rect 24578 9092 24584 9104
rect 24539 9064 24584 9092
rect 24578 9052 24584 9064
rect 24636 9092 24642 9104
rect 24918 9095 24976 9101
rect 24918 9092 24930 9095
rect 24636 9064 24930 9092
rect 24636 9052 24642 9064
rect 24918 9061 24930 9064
rect 24964 9061 24976 9095
rect 27154 9092 27160 9104
rect 27115 9064 27160 9092
rect 24918 9055 24976 9061
rect 27154 9052 27160 9064
rect 27212 9052 27218 9104
rect 27798 9052 27804 9104
rect 27856 9092 27862 9104
rect 27893 9095 27951 9101
rect 27893 9092 27905 9095
rect 27856 9064 27905 9092
rect 27856 9052 27862 9064
rect 27893 9061 27905 9064
rect 27939 9061 27951 9095
rect 28074 9092 28080 9104
rect 28035 9064 28080 9092
rect 27893 9055 27951 9061
rect 28074 9052 28080 9064
rect 28132 9052 28138 9104
rect 29086 9052 29092 9104
rect 29144 9092 29150 9104
rect 29457 9095 29515 9101
rect 29457 9092 29469 9095
rect 29144 9064 29469 9092
rect 29144 9052 29150 9064
rect 29457 9061 29469 9064
rect 29503 9092 29515 9095
rect 30006 9092 30012 9104
rect 29503 9064 30012 9092
rect 29503 9061 29515 9064
rect 29457 9055 29515 9061
rect 30006 9052 30012 9064
rect 30064 9052 30070 9104
rect 35802 9052 35808 9104
rect 35860 9092 35866 9104
rect 38930 9092 38936 9104
rect 35860 9064 36584 9092
rect 38843 9064 38936 9092
rect 35860 9052 35866 9064
rect 6273 9027 6331 9033
rect 6273 9024 6285 9027
rect 5224 8996 6285 9024
rect 5224 8984 5230 8996
rect 6273 8993 6285 8996
rect 6319 8993 6331 9027
rect 6273 8987 6331 8993
rect 6546 8984 6552 9036
rect 6604 9024 6610 9036
rect 6713 9027 6771 9033
rect 6713 9024 6725 9027
rect 6604 8996 6725 9024
rect 6604 8984 6610 8996
rect 6713 8993 6725 8996
rect 6759 8993 6771 9027
rect 6713 8987 6771 8993
rect 15010 8984 15016 9036
rect 15068 9024 15074 9036
rect 15545 9027 15603 9033
rect 15545 9024 15557 9027
rect 15068 8996 15557 9024
rect 15068 8984 15074 8996
rect 15545 8993 15557 8996
rect 15591 9024 15603 9027
rect 15930 9024 15936 9036
rect 15591 8996 15936 9024
rect 15591 8993 15603 8996
rect 15545 8987 15603 8993
rect 15930 8984 15936 8996
rect 15988 8984 15994 9036
rect 18046 9033 18052 9036
rect 18040 9024 18052 9033
rect 18007 8996 18052 9024
rect 18040 8987 18052 8996
rect 18046 8984 18052 8987
rect 18104 8984 18110 9036
rect 22278 9024 22284 9036
rect 22239 8996 22284 9024
rect 22278 8984 22284 8996
rect 22336 8984 22342 9036
rect 22548 9027 22606 9033
rect 22548 8993 22560 9027
rect 22594 9024 22606 9027
rect 22922 9024 22928 9036
rect 22594 8996 22928 9024
rect 22594 8993 22606 8996
rect 22548 8987 22606 8993
rect 22922 8984 22928 8996
rect 22980 8984 22986 9036
rect 27172 9024 27200 9052
rect 28537 9027 28595 9033
rect 28537 9024 28549 9027
rect 27172 8996 28549 9024
rect 28537 8993 28549 8996
rect 28583 9024 28595 9027
rect 28905 9027 28963 9033
rect 28905 9024 28917 9027
rect 28583 8996 28917 9024
rect 28583 8993 28595 8996
rect 28537 8987 28595 8993
rect 28905 8993 28917 8996
rect 28951 9024 28963 9027
rect 28994 9024 29000 9036
rect 28951 8996 29000 9024
rect 28951 8993 28963 8996
rect 28905 8987 28963 8993
rect 28994 8984 29000 8996
rect 29052 9024 29058 9036
rect 29733 9027 29791 9033
rect 29733 9024 29745 9027
rect 29052 8996 29745 9024
rect 29052 8984 29058 8996
rect 29733 8993 29745 8996
rect 29779 9024 29791 9027
rect 30190 9024 30196 9036
rect 29779 8996 30196 9024
rect 29779 8993 29791 8996
rect 29733 8987 29791 8993
rect 30190 8984 30196 8996
rect 30248 9024 30254 9036
rect 30469 9027 30527 9033
rect 30469 9024 30481 9027
rect 30248 8996 30481 9024
rect 30248 8984 30254 8996
rect 30469 8993 30481 8996
rect 30515 9024 30527 9027
rect 30834 9024 30840 9036
rect 30515 8996 30840 9024
rect 30515 8993 30527 8996
rect 30469 8987 30527 8993
rect 30834 8984 30840 8996
rect 30892 8984 30898 9036
rect 31846 8984 31852 9036
rect 31904 9024 31910 9036
rect 32381 9027 32439 9033
rect 32381 9024 32393 9027
rect 31904 8996 32393 9024
rect 31904 8984 31910 8996
rect 32381 8993 32393 8996
rect 32427 8993 32439 9027
rect 32381 8987 32439 8993
rect 4617 8959 4675 8965
rect 4617 8925 4629 8959
rect 4663 8925 4675 8959
rect 6454 8956 6460 8968
rect 6415 8928 6460 8956
rect 4617 8919 4675 8925
rect 4154 8888 4160 8900
rect 4115 8860 4160 8888
rect 4154 8848 4160 8860
rect 4212 8848 4218 8900
rect 4632 8888 4660 8919
rect 6454 8916 6460 8928
rect 6512 8916 6518 8968
rect 11974 8956 11980 8968
rect 11935 8928 11980 8956
rect 11974 8916 11980 8928
rect 12032 8916 12038 8968
rect 15286 8956 15292 8968
rect 15247 8928 15292 8956
rect 15286 8916 15292 8928
rect 15344 8916 15350 8968
rect 17770 8956 17776 8968
rect 17731 8928 17776 8956
rect 17770 8916 17776 8928
rect 17828 8916 17834 8968
rect 20898 8956 20904 8968
rect 20859 8928 20904 8956
rect 20898 8916 20904 8928
rect 20956 8916 20962 8968
rect 24670 8956 24676 8968
rect 24631 8928 24676 8956
rect 24670 8916 24676 8928
rect 24728 8916 24734 8968
rect 27062 8956 27068 8968
rect 27023 8928 27068 8956
rect 27062 8916 27068 8928
rect 27120 8916 27126 8968
rect 28166 8956 28172 8968
rect 28127 8928 28172 8956
rect 28166 8916 28172 8928
rect 28224 8916 28230 8968
rect 30098 8916 30104 8968
rect 30156 8956 30162 8968
rect 31570 8956 31576 8968
rect 30156 8928 31576 8956
rect 30156 8916 30162 8928
rect 31570 8916 31576 8928
rect 31628 8956 31634 8968
rect 32125 8959 32183 8965
rect 32125 8956 32137 8959
rect 31628 8928 32137 8956
rect 31628 8916 31634 8928
rect 32125 8925 32137 8928
rect 32171 8925 32183 8959
rect 36446 8956 36452 8968
rect 36407 8928 36452 8956
rect 32125 8919 32183 8925
rect 36446 8916 36452 8928
rect 36504 8916 36510 8968
rect 36556 8965 36584 9064
rect 38930 9052 38936 9064
rect 38988 9052 38994 9104
rect 39114 9092 39120 9104
rect 39075 9064 39120 9092
rect 39114 9052 39120 9064
rect 39172 9052 39178 9104
rect 39408 9092 39436 9132
rect 40034 9120 40040 9132
rect 40092 9160 40098 9172
rect 41966 9160 41972 9172
rect 40092 9132 40816 9160
rect 41927 9132 41972 9160
rect 40092 9120 40098 9132
rect 40788 9104 40816 9132
rect 41966 9120 41972 9132
rect 42024 9120 42030 9172
rect 42426 9160 42432 9172
rect 42387 9132 42432 9160
rect 42426 9120 42432 9132
rect 42484 9120 42490 9172
rect 44545 9163 44603 9169
rect 44545 9129 44557 9163
rect 44591 9160 44603 9163
rect 44818 9160 44824 9172
rect 44591 9132 44824 9160
rect 44591 9129 44603 9132
rect 44545 9123 44603 9129
rect 44818 9120 44824 9132
rect 44876 9120 44882 9172
rect 46474 9160 46480 9172
rect 46435 9132 46480 9160
rect 46474 9120 46480 9132
rect 46532 9120 46538 9172
rect 40203 9095 40261 9101
rect 40203 9092 40215 9095
rect 39408 9064 40215 9092
rect 40203 9061 40215 9064
rect 40249 9061 40261 9095
rect 40678 9092 40684 9104
rect 40639 9064 40684 9092
rect 40203 9055 40261 9061
rect 40678 9052 40684 9064
rect 40736 9052 40742 9104
rect 40770 9052 40776 9104
rect 40828 9092 40834 9104
rect 40828 9064 40873 9092
rect 40828 9052 40834 9064
rect 45002 9052 45008 9104
rect 45060 9092 45066 9104
rect 45364 9095 45422 9101
rect 45364 9092 45376 9095
rect 45060 9064 45376 9092
rect 45060 9052 45066 9064
rect 45364 9061 45376 9064
rect 45410 9092 45422 9095
rect 45554 9092 45560 9104
rect 45410 9064 45560 9092
rect 45410 9061 45422 9064
rect 45364 9055 45422 9061
rect 45554 9052 45560 9064
rect 45612 9052 45618 9104
rect 38473 9027 38531 9033
rect 38473 8993 38485 9027
rect 38519 9024 38531 9027
rect 38562 9024 38568 9036
rect 38519 8996 38568 9024
rect 38519 8993 38531 8996
rect 38473 8987 38531 8993
rect 38562 8984 38568 8996
rect 38620 9024 38626 9036
rect 40494 9024 40500 9036
rect 38620 8996 39252 9024
rect 40455 8996 40500 9024
rect 38620 8984 38626 8996
rect 39224 8968 39252 8996
rect 40494 8984 40500 8996
rect 40552 8984 40558 9036
rect 41785 9027 41843 9033
rect 41785 8993 41797 9027
rect 41831 9024 41843 9027
rect 42426 9024 42432 9036
rect 41831 8996 42432 9024
rect 41831 8993 41843 8996
rect 41785 8987 41843 8993
rect 42426 8984 42432 8996
rect 42484 8984 42490 9036
rect 45186 9024 45192 9036
rect 45112 8996 45192 9024
rect 36541 8959 36599 8965
rect 36541 8925 36553 8959
rect 36587 8956 36599 8959
rect 36722 8956 36728 8968
rect 36587 8928 36728 8956
rect 36587 8925 36599 8928
rect 36541 8919 36599 8925
rect 36722 8916 36728 8928
rect 36780 8916 36786 8968
rect 39206 8956 39212 8968
rect 39167 8928 39212 8956
rect 39206 8916 39212 8928
rect 39264 8916 39270 8968
rect 44174 8916 44180 8968
rect 44232 8956 44238 8968
rect 44818 8956 44824 8968
rect 44232 8928 44824 8956
rect 44232 8916 44238 8928
rect 44818 8916 44824 8928
rect 44876 8956 44882 8968
rect 45112 8965 45140 8996
rect 45186 8984 45192 8996
rect 45244 8984 45250 9036
rect 45097 8959 45155 8965
rect 45097 8956 45109 8959
rect 44876 8928 45109 8956
rect 44876 8916 44882 8928
rect 45097 8925 45109 8928
rect 45143 8925 45155 8959
rect 45097 8919 45155 8925
rect 4798 8888 4804 8900
rect 4632 8860 4804 8888
rect 4798 8848 4804 8860
rect 4856 8848 4862 8900
rect 13814 8848 13820 8900
rect 13872 8888 13878 8900
rect 15013 8891 15071 8897
rect 15013 8888 15025 8891
rect 13872 8860 15025 8888
rect 13872 8848 13878 8860
rect 15013 8857 15025 8860
rect 15059 8888 15071 8891
rect 15102 8888 15108 8900
rect 15059 8860 15108 8888
rect 15059 8857 15071 8860
rect 15013 8851 15071 8857
rect 15102 8848 15108 8860
rect 15160 8848 15166 8900
rect 27617 8891 27675 8897
rect 27617 8857 27629 8891
rect 27663 8888 27675 8891
rect 27890 8888 27896 8900
rect 27663 8860 27896 8888
rect 27663 8857 27675 8860
rect 27617 8851 27675 8857
rect 27890 8848 27896 8860
rect 27948 8848 27954 8900
rect 35989 8891 36047 8897
rect 35989 8857 36001 8891
rect 36035 8888 36047 8891
rect 38102 8888 38108 8900
rect 36035 8860 38108 8888
rect 36035 8857 36047 8860
rect 35989 8851 36047 8857
rect 38102 8848 38108 8860
rect 38160 8848 38166 8900
rect 38654 8888 38660 8900
rect 38615 8860 38660 8888
rect 38654 8848 38660 8860
rect 38712 8848 38718 8900
rect 12618 8780 12624 8832
rect 12676 8820 12682 8832
rect 13357 8823 13415 8829
rect 13357 8820 13369 8823
rect 12676 8792 13369 8820
rect 12676 8780 12682 8792
rect 13357 8789 13369 8792
rect 13403 8789 13415 8823
rect 14642 8820 14648 8832
rect 14603 8792 14648 8820
rect 13357 8783 13415 8789
rect 14642 8780 14648 8792
rect 14700 8780 14706 8832
rect 17586 8820 17592 8832
rect 17547 8792 17592 8820
rect 17586 8780 17592 8792
rect 17644 8780 17650 8832
rect 17678 8780 17684 8832
rect 17736 8820 17742 8832
rect 19153 8823 19211 8829
rect 19153 8820 19165 8823
rect 17736 8792 19165 8820
rect 17736 8780 17742 8792
rect 19153 8789 19165 8792
rect 19199 8789 19211 8823
rect 19153 8783 19211 8789
rect 20806 8780 20812 8832
rect 20864 8820 20870 8832
rect 23661 8823 23719 8829
rect 23661 8820 23673 8823
rect 20864 8792 23673 8820
rect 20864 8780 20870 8792
rect 23661 8789 23673 8792
rect 23707 8789 23719 8823
rect 23661 8783 23719 8789
rect 26234 8780 26240 8832
rect 26292 8820 26298 8832
rect 26605 8823 26663 8829
rect 26605 8820 26617 8823
rect 26292 8792 26617 8820
rect 26292 8780 26298 8792
rect 26605 8789 26617 8792
rect 26651 8789 26663 8823
rect 29178 8820 29184 8832
rect 29139 8792 29184 8820
rect 26605 8783 26663 8789
rect 29178 8780 29184 8792
rect 29236 8780 29242 8832
rect 30742 8780 30748 8832
rect 30800 8820 30806 8832
rect 31849 8823 31907 8829
rect 31849 8820 31861 8823
rect 30800 8792 31861 8820
rect 30800 8780 30806 8792
rect 31849 8789 31861 8792
rect 31895 8820 31907 8823
rect 32490 8820 32496 8832
rect 31895 8792 32496 8820
rect 31895 8789 31907 8792
rect 31849 8783 31907 8789
rect 32490 8780 32496 8792
rect 32548 8780 32554 8832
rect 43073 8823 43131 8829
rect 43073 8789 43085 8823
rect 43119 8820 43131 8823
rect 43622 8820 43628 8832
rect 43119 8792 43628 8820
rect 43119 8789 43131 8792
rect 43073 8783 43131 8789
rect 43622 8780 43628 8792
rect 43680 8780 43686 8832
rect 1104 8730 48852 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 34966 8730
rect 35018 8678 35030 8730
rect 35082 8678 35094 8730
rect 35146 8678 35158 8730
rect 35210 8678 48852 8730
rect 1104 8656 48852 8678
rect 2038 8616 2044 8628
rect 1999 8588 2044 8616
rect 2038 8576 2044 8588
rect 2096 8576 2102 8628
rect 3881 8619 3939 8625
rect 3881 8585 3893 8619
rect 3927 8616 3939 8619
rect 4525 8619 4583 8625
rect 4525 8616 4537 8619
rect 3927 8588 4537 8616
rect 3927 8585 3939 8588
rect 3881 8579 3939 8585
rect 4525 8585 4537 8588
rect 4571 8616 4583 8619
rect 4614 8616 4620 8628
rect 4571 8588 4620 8616
rect 4571 8585 4583 8588
rect 4525 8579 4583 8585
rect 4614 8576 4620 8588
rect 4672 8576 4678 8628
rect 4798 8616 4804 8628
rect 4759 8588 4804 8616
rect 4798 8576 4804 8588
rect 4856 8616 4862 8628
rect 6089 8619 6147 8625
rect 6089 8616 6101 8619
rect 4856 8588 6101 8616
rect 4856 8576 4862 8588
rect 6089 8585 6101 8588
rect 6135 8585 6147 8619
rect 6089 8579 6147 8585
rect 1486 8508 1492 8560
rect 1544 8548 1550 8560
rect 2317 8551 2375 8557
rect 2317 8548 2329 8551
rect 1544 8520 2329 8548
rect 1544 8508 1550 8520
rect 2317 8517 2329 8520
rect 2363 8548 2375 8551
rect 5166 8548 5172 8560
rect 2363 8520 2544 8548
rect 5127 8520 5172 8548
rect 2363 8517 2375 8520
rect 2317 8511 2375 8517
rect 2516 8489 2544 8520
rect 5166 8508 5172 8520
rect 5224 8508 5230 8560
rect 2501 8483 2559 8489
rect 2501 8449 2513 8483
rect 2547 8449 2559 8483
rect 6104 8480 6132 8579
rect 6546 8576 6552 8628
rect 6604 8616 6610 8628
rect 8205 8619 8263 8625
rect 8205 8616 8217 8619
rect 6604 8588 8217 8616
rect 6604 8576 6610 8588
rect 8205 8585 8217 8588
rect 8251 8585 8263 8619
rect 15010 8616 15016 8628
rect 14971 8588 15016 8616
rect 8205 8579 8263 8585
rect 15010 8576 15016 8588
rect 15068 8576 15074 8628
rect 15286 8616 15292 8628
rect 15247 8588 15292 8616
rect 15286 8576 15292 8588
rect 15344 8616 15350 8628
rect 17405 8619 17463 8625
rect 17405 8616 17417 8619
rect 15344 8588 17417 8616
rect 15344 8576 15350 8588
rect 17405 8585 17417 8588
rect 17451 8616 17463 8619
rect 17770 8616 17776 8628
rect 17451 8588 17776 8616
rect 17451 8585 17463 8588
rect 17405 8579 17463 8585
rect 17770 8576 17776 8588
rect 17828 8576 17834 8628
rect 22278 8576 22284 8628
rect 22336 8616 22342 8628
rect 22465 8619 22523 8625
rect 22465 8616 22477 8619
rect 22336 8588 22477 8616
rect 22336 8576 22342 8588
rect 22465 8585 22477 8588
rect 22511 8585 22523 8619
rect 22922 8616 22928 8628
rect 22835 8588 22928 8616
rect 22465 8579 22523 8585
rect 16390 8548 16396 8560
rect 16351 8520 16396 8548
rect 16390 8508 16396 8520
rect 16448 8508 16454 8560
rect 6104 8452 6960 8480
rect 2501 8443 2559 8449
rect 2516 8344 2544 8443
rect 2774 8421 2780 8424
rect 2768 8375 2780 8421
rect 2832 8412 2838 8424
rect 6825 8415 6883 8421
rect 2832 8384 2868 8412
rect 2774 8372 2780 8375
rect 2832 8372 2838 8384
rect 6825 8381 6837 8415
rect 6871 8381 6883 8415
rect 6932 8412 6960 8452
rect 14642 8440 14648 8492
rect 14700 8480 14706 8492
rect 15841 8483 15899 8489
rect 15841 8480 15853 8483
rect 14700 8452 15853 8480
rect 14700 8440 14706 8452
rect 15841 8449 15853 8452
rect 15887 8480 15899 8483
rect 16853 8483 16911 8489
rect 16853 8480 16865 8483
rect 15887 8452 16865 8480
rect 15887 8449 15899 8452
rect 15841 8443 15899 8449
rect 16853 8449 16865 8452
rect 16899 8480 16911 8483
rect 17678 8480 17684 8492
rect 16899 8452 17684 8480
rect 16899 8449 16911 8452
rect 16853 8443 16911 8449
rect 17678 8440 17684 8452
rect 17736 8440 17742 8492
rect 17788 8480 17816 8576
rect 22480 8548 22508 8579
rect 22922 8576 22928 8588
rect 22980 8616 22986 8628
rect 25041 8619 25099 8625
rect 25041 8616 25053 8619
rect 22980 8588 25053 8616
rect 22980 8576 22986 8588
rect 25041 8585 25053 8588
rect 25087 8585 25099 8619
rect 25041 8579 25099 8585
rect 27062 8576 27068 8628
rect 27120 8616 27126 8628
rect 27120 8588 27568 8616
rect 27120 8576 27126 8588
rect 27540 8557 27568 8588
rect 28074 8576 28080 8628
rect 28132 8616 28138 8628
rect 28537 8619 28595 8625
rect 28537 8616 28549 8619
rect 28132 8588 28549 8616
rect 28132 8576 28138 8588
rect 28537 8585 28549 8588
rect 28583 8616 28595 8619
rect 29178 8616 29184 8628
rect 28583 8588 29184 8616
rect 28583 8585 28595 8588
rect 28537 8579 28595 8585
rect 29178 8576 29184 8588
rect 29236 8576 29242 8628
rect 29546 8616 29552 8628
rect 29507 8588 29552 8616
rect 29546 8576 29552 8588
rect 29604 8576 29610 8628
rect 31570 8616 31576 8628
rect 31531 8588 31576 8616
rect 31570 8576 31576 8588
rect 31628 8576 31634 8628
rect 31938 8576 31944 8628
rect 31996 8616 32002 8628
rect 33137 8619 33195 8625
rect 33137 8616 33149 8619
rect 31996 8588 33149 8616
rect 31996 8576 32002 8588
rect 33137 8585 33149 8588
rect 33183 8585 33195 8619
rect 35986 8616 35992 8628
rect 35947 8588 35992 8616
rect 33137 8579 33195 8585
rect 35986 8576 35992 8588
rect 36044 8576 36050 8628
rect 38930 8616 38936 8628
rect 38891 8588 38936 8616
rect 38930 8576 38936 8588
rect 38988 8576 38994 8628
rect 40494 8576 40500 8628
rect 40552 8616 40558 8628
rect 41877 8619 41935 8625
rect 41877 8616 41889 8619
rect 40552 8588 41889 8616
rect 40552 8576 40558 8588
rect 41877 8585 41889 8588
rect 41923 8585 41935 8619
rect 42426 8616 42432 8628
rect 42387 8588 42432 8616
rect 41877 8579 41935 8585
rect 42426 8576 42432 8588
rect 42484 8616 42490 8628
rect 43073 8619 43131 8625
rect 43073 8616 43085 8619
rect 42484 8588 43085 8616
rect 42484 8576 42490 8588
rect 43073 8585 43085 8588
rect 43119 8585 43131 8619
rect 43073 8579 43131 8585
rect 23385 8551 23443 8557
rect 23385 8548 23397 8551
rect 22480 8520 23397 8548
rect 23385 8517 23397 8520
rect 23431 8517 23443 8551
rect 23385 8511 23443 8517
rect 27525 8551 27583 8557
rect 27525 8517 27537 8551
rect 27571 8548 27583 8551
rect 28169 8551 28227 8557
rect 28169 8548 28181 8551
rect 27571 8520 28181 8548
rect 27571 8517 27583 8520
rect 27525 8511 27583 8517
rect 28169 8517 28181 8520
rect 28215 8517 28227 8551
rect 29086 8548 29092 8560
rect 29047 8520 29092 8548
rect 28169 8511 28227 8517
rect 18049 8483 18107 8489
rect 18049 8480 18061 8483
rect 17788 8452 18061 8480
rect 18049 8449 18061 8452
rect 18095 8449 18107 8483
rect 18049 8443 18107 8449
rect 7081 8415 7139 8421
rect 7081 8412 7093 8415
rect 6932 8384 7093 8412
rect 6825 8375 6883 8381
rect 7081 8381 7093 8384
rect 7127 8381 7139 8415
rect 7081 8375 7139 8381
rect 2516 8316 2728 8344
rect 2700 8276 2728 8316
rect 6454 8304 6460 8356
rect 6512 8344 6518 8356
rect 6549 8347 6607 8353
rect 6549 8344 6561 8347
rect 6512 8316 6561 8344
rect 6512 8304 6518 8316
rect 6549 8313 6561 8316
rect 6595 8344 6607 8347
rect 6840 8344 6868 8375
rect 11974 8372 11980 8424
rect 12032 8412 12038 8424
rect 12437 8415 12495 8421
rect 12437 8412 12449 8415
rect 12032 8384 12449 8412
rect 12032 8372 12038 8384
rect 12437 8381 12449 8384
rect 12483 8381 12495 8415
rect 18064 8412 18092 8443
rect 20806 8421 20812 8424
rect 20349 8415 20407 8421
rect 20349 8412 20361 8415
rect 18064 8384 20361 8412
rect 12437 8375 12495 8381
rect 20349 8381 20361 8384
rect 20395 8412 20407 8415
rect 20533 8415 20591 8421
rect 20533 8412 20545 8415
rect 20395 8384 20545 8412
rect 20395 8381 20407 8384
rect 20349 8375 20407 8381
rect 20533 8381 20545 8384
rect 20579 8381 20591 8415
rect 20800 8412 20812 8421
rect 20767 8384 20812 8412
rect 20533 8375 20591 8381
rect 20800 8375 20812 8384
rect 20806 8372 20812 8375
rect 20864 8372 20870 8424
rect 23400 8412 23428 8511
rect 29086 8508 29092 8520
rect 29144 8508 29150 8560
rect 29362 8508 29368 8560
rect 29420 8548 29426 8560
rect 30285 8551 30343 8557
rect 30285 8548 30297 8551
rect 29420 8520 30297 8548
rect 29420 8508 29426 8520
rect 30285 8517 30297 8520
rect 30331 8517 30343 8551
rect 30285 8511 30343 8517
rect 25685 8483 25743 8489
rect 25685 8449 25697 8483
rect 25731 8480 25743 8483
rect 30101 8483 30159 8489
rect 25731 8452 26280 8480
rect 25731 8449 25743 8452
rect 25685 8443 25743 8449
rect 23661 8415 23719 8421
rect 23661 8412 23673 8415
rect 23400 8384 23673 8412
rect 23661 8381 23673 8384
rect 23707 8412 23719 8415
rect 24670 8412 24676 8424
rect 23707 8384 24676 8412
rect 23707 8381 23719 8384
rect 23661 8375 23719 8381
rect 6914 8344 6920 8356
rect 6595 8316 6920 8344
rect 6595 8313 6607 8316
rect 6549 8307 6607 8313
rect 6914 8304 6920 8316
rect 6972 8304 6978 8356
rect 11517 8347 11575 8353
rect 11517 8313 11529 8347
rect 11563 8344 11575 8347
rect 12526 8344 12532 8356
rect 11563 8316 12532 8344
rect 11563 8313 11575 8316
rect 11517 8307 11575 8313
rect 12526 8304 12532 8316
rect 12584 8344 12590 8356
rect 12682 8347 12740 8353
rect 12682 8344 12694 8347
rect 12584 8316 12694 8344
rect 12584 8304 12590 8316
rect 12682 8313 12694 8316
rect 12728 8313 12740 8347
rect 12682 8307 12740 8313
rect 16209 8347 16267 8353
rect 16209 8313 16221 8347
rect 16255 8344 16267 8347
rect 16942 8344 16948 8356
rect 16255 8316 16620 8344
rect 16903 8316 16948 8344
rect 16255 8313 16267 8316
rect 16209 8307 16267 8313
rect 4062 8276 4068 8288
rect 2700 8248 4068 8276
rect 4062 8236 4068 8248
rect 4120 8236 4126 8288
rect 9674 8236 9680 8288
rect 9732 8276 9738 8288
rect 11793 8279 11851 8285
rect 11793 8276 11805 8279
rect 9732 8248 11805 8276
rect 9732 8236 9738 8248
rect 11793 8245 11805 8248
rect 11839 8276 11851 8279
rect 11974 8276 11980 8288
rect 11839 8248 11980 8276
rect 11839 8245 11851 8248
rect 11793 8239 11851 8245
rect 11974 8236 11980 8248
rect 12032 8276 12038 8288
rect 12161 8279 12219 8285
rect 12161 8276 12173 8279
rect 12032 8248 12173 8276
rect 12032 8236 12038 8248
rect 12161 8245 12173 8248
rect 12207 8245 12219 8279
rect 12161 8239 12219 8245
rect 12894 8236 12900 8288
rect 12952 8276 12958 8288
rect 13817 8279 13875 8285
rect 13817 8276 13829 8279
rect 12952 8248 13829 8276
rect 12952 8236 12958 8248
rect 13817 8245 13829 8248
rect 13863 8245 13875 8279
rect 16592 8276 16620 8316
rect 16942 8304 16948 8316
rect 17000 8304 17006 8356
rect 17586 8304 17592 8356
rect 17644 8344 17650 8356
rect 18316 8347 18374 8353
rect 18316 8344 18328 8347
rect 17644 8316 18328 8344
rect 17644 8304 17650 8316
rect 18316 8313 18328 8316
rect 18362 8344 18374 8347
rect 18506 8344 18512 8356
rect 18362 8316 18512 8344
rect 18362 8313 18374 8316
rect 18316 8307 18374 8313
rect 18506 8304 18512 8316
rect 18564 8344 18570 8356
rect 18564 8316 21956 8344
rect 18564 8304 18570 8316
rect 16850 8276 16856 8288
rect 16592 8248 16856 8276
rect 13817 8239 13875 8245
rect 16850 8236 16856 8248
rect 16908 8236 16914 8288
rect 18598 8236 18604 8288
rect 18656 8276 18662 8288
rect 21928 8285 21956 8316
rect 19429 8279 19487 8285
rect 19429 8276 19441 8279
rect 18656 8248 19441 8276
rect 18656 8236 18662 8248
rect 19429 8245 19441 8248
rect 19475 8245 19487 8279
rect 19429 8239 19487 8245
rect 21913 8279 21971 8285
rect 21913 8245 21925 8279
rect 21959 8245 21971 8279
rect 23768 8276 23796 8384
rect 24670 8372 24676 8384
rect 24728 8412 24734 8424
rect 25961 8415 26019 8421
rect 25961 8412 25973 8415
rect 24728 8384 25973 8412
rect 24728 8372 24734 8384
rect 25961 8381 25973 8384
rect 26007 8412 26019 8415
rect 26145 8415 26203 8421
rect 26145 8412 26157 8415
rect 26007 8384 26157 8412
rect 26007 8381 26019 8384
rect 25961 8375 26019 8381
rect 23934 8353 23940 8356
rect 23928 8344 23940 8353
rect 23895 8316 23940 8344
rect 23928 8307 23940 8316
rect 23934 8304 23940 8307
rect 23992 8304 23998 8356
rect 23842 8276 23848 8288
rect 23768 8248 23848 8276
rect 21913 8239 21971 8245
rect 23842 8236 23848 8248
rect 23900 8236 23906 8288
rect 26068 8276 26096 8384
rect 26145 8381 26157 8384
rect 26191 8381 26203 8415
rect 26145 8375 26203 8381
rect 26252 8344 26280 8452
rect 30101 8449 30113 8483
rect 30147 8480 30159 8483
rect 30742 8480 30748 8492
rect 30147 8452 30748 8480
rect 30147 8449 30159 8452
rect 30101 8443 30159 8449
rect 30742 8440 30748 8452
rect 30800 8440 30806 8492
rect 30834 8440 30840 8492
rect 30892 8480 30898 8492
rect 31588 8480 31616 8576
rect 42794 8548 42800 8560
rect 42755 8520 42800 8548
rect 42794 8508 42800 8520
rect 42852 8508 42858 8560
rect 46934 8548 46940 8560
rect 46895 8520 46940 8548
rect 46934 8508 46940 8520
rect 46992 8508 46998 8560
rect 31757 8483 31815 8489
rect 31757 8480 31769 8483
rect 30892 8452 30937 8480
rect 31588 8452 31769 8480
rect 30892 8440 30898 8452
rect 31757 8449 31769 8452
rect 31803 8449 31815 8483
rect 31757 8443 31815 8449
rect 30576 8384 31708 8412
rect 26412 8347 26470 8353
rect 26412 8344 26424 8347
rect 26252 8316 26424 8344
rect 26412 8313 26424 8316
rect 26458 8344 26470 8347
rect 26510 8344 26516 8356
rect 26458 8316 26516 8344
rect 26458 8313 26470 8316
rect 26412 8307 26470 8313
rect 26510 8304 26516 8316
rect 26568 8304 26574 8356
rect 30576 8353 30604 8384
rect 30561 8347 30619 8353
rect 30561 8344 30573 8347
rect 30300 8316 30573 8344
rect 30300 8288 30328 8316
rect 30561 8313 30573 8316
rect 30607 8313 30619 8347
rect 30742 8344 30748 8356
rect 30703 8316 30748 8344
rect 30561 8307 30619 8313
rect 30742 8304 30748 8316
rect 30800 8304 30806 8356
rect 31680 8344 31708 8384
rect 35526 8372 35532 8424
rect 35584 8412 35590 8424
rect 36265 8415 36323 8421
rect 36265 8412 36277 8415
rect 35584 8384 36277 8412
rect 35584 8372 35590 8384
rect 36265 8381 36277 8384
rect 36311 8412 36323 8415
rect 36449 8415 36507 8421
rect 36449 8412 36461 8415
rect 36311 8384 36461 8412
rect 36311 8381 36323 8384
rect 36265 8375 36323 8381
rect 36449 8381 36461 8384
rect 36495 8381 36507 8415
rect 36449 8375 36507 8381
rect 36538 8372 36544 8424
rect 36596 8412 36602 8424
rect 36705 8415 36763 8421
rect 36705 8412 36717 8415
rect 36596 8384 36717 8412
rect 36596 8372 36602 8384
rect 36705 8381 36717 8384
rect 36751 8381 36763 8415
rect 36705 8375 36763 8381
rect 40310 8372 40316 8424
rect 40368 8412 40374 8424
rect 40497 8415 40555 8421
rect 40497 8412 40509 8415
rect 40368 8384 40509 8412
rect 40368 8372 40374 8384
rect 40497 8381 40509 8384
rect 40543 8381 40555 8415
rect 42812 8412 42840 8508
rect 43622 8480 43628 8492
rect 43583 8452 43628 8480
rect 43622 8440 43628 8452
rect 43680 8440 43686 8492
rect 47394 8480 47400 8492
rect 47355 8452 47400 8480
rect 47394 8440 47400 8452
rect 47452 8440 47458 8492
rect 46753 8415 46811 8421
rect 42812 8384 43576 8412
rect 40497 8375 40555 8381
rect 31846 8344 31852 8356
rect 31680 8316 31852 8344
rect 31846 8304 31852 8316
rect 31904 8304 31910 8356
rect 32024 8347 32082 8353
rect 32024 8313 32036 8347
rect 32070 8344 32082 8347
rect 32490 8344 32496 8356
rect 32070 8316 32496 8344
rect 32070 8313 32082 8316
rect 32024 8307 32082 8313
rect 32490 8304 32496 8316
rect 32548 8304 32554 8356
rect 35621 8347 35679 8353
rect 35621 8313 35633 8347
rect 35667 8344 35679 8347
rect 36556 8344 36584 8372
rect 39114 8344 39120 8356
rect 35667 8316 36584 8344
rect 38580 8316 39120 8344
rect 35667 8313 35679 8316
rect 35621 8307 35679 8313
rect 26602 8276 26608 8288
rect 26068 8248 26608 8276
rect 26602 8236 26608 8248
rect 26660 8236 26666 8288
rect 30282 8236 30288 8288
rect 30340 8236 30346 8288
rect 37826 8276 37832 8288
rect 37787 8248 37832 8276
rect 37826 8236 37832 8248
rect 37884 8236 37890 8288
rect 37918 8236 37924 8288
rect 37976 8276 37982 8288
rect 38580 8285 38608 8316
rect 39114 8304 39120 8316
rect 39172 8304 39178 8356
rect 39577 8347 39635 8353
rect 39577 8313 39589 8347
rect 39623 8344 39635 8347
rect 39945 8347 40003 8353
rect 39945 8344 39957 8347
rect 39623 8316 39957 8344
rect 39623 8313 39635 8316
rect 39577 8307 39635 8313
rect 39945 8313 39957 8316
rect 39991 8344 40003 8347
rect 40764 8347 40822 8353
rect 39991 8316 40520 8344
rect 39991 8313 40003 8316
rect 39945 8307 40003 8313
rect 38565 8279 38623 8285
rect 38565 8276 38577 8279
rect 37976 8248 38577 8276
rect 37976 8236 37982 8248
rect 38565 8245 38577 8248
rect 38611 8245 38623 8279
rect 40310 8276 40316 8288
rect 40271 8248 40316 8276
rect 38565 8239 38623 8245
rect 40310 8236 40316 8248
rect 40368 8236 40374 8288
rect 40492 8276 40520 8316
rect 40764 8313 40776 8347
rect 40810 8344 40822 8347
rect 41598 8344 41604 8356
rect 40810 8316 41604 8344
rect 40810 8313 40822 8316
rect 40764 8307 40822 8313
rect 40678 8276 40684 8288
rect 40492 8248 40684 8276
rect 40678 8236 40684 8248
rect 40736 8276 40742 8288
rect 40779 8276 40807 8307
rect 41598 8304 41604 8316
rect 41656 8304 41662 8356
rect 43070 8304 43076 8356
rect 43128 8344 43134 8356
rect 43548 8353 43576 8384
rect 46753 8381 46765 8415
rect 46799 8412 46811 8415
rect 47412 8412 47440 8440
rect 46799 8384 47440 8412
rect 46799 8381 46811 8384
rect 46753 8375 46811 8381
rect 43349 8347 43407 8353
rect 43349 8344 43361 8347
rect 43128 8316 43361 8344
rect 43128 8304 43134 8316
rect 43349 8313 43361 8316
rect 43395 8313 43407 8347
rect 43349 8307 43407 8313
rect 43533 8347 43591 8353
rect 43533 8313 43545 8347
rect 43579 8313 43591 8347
rect 43533 8307 43591 8313
rect 40736 8248 40807 8276
rect 40736 8236 40742 8248
rect 44818 8236 44824 8288
rect 44876 8276 44882 8288
rect 45097 8279 45155 8285
rect 45097 8276 45109 8279
rect 44876 8248 45109 8276
rect 44876 8236 44882 8248
rect 45097 8245 45109 8248
rect 45143 8245 45155 8279
rect 45554 8276 45560 8288
rect 45515 8248 45560 8276
rect 45097 8239 45155 8245
rect 45554 8236 45560 8248
rect 45612 8236 45618 8288
rect 1104 8186 48852 8208
rect 1104 8134 19606 8186
rect 19658 8134 19670 8186
rect 19722 8134 19734 8186
rect 19786 8134 19798 8186
rect 19850 8134 48852 8186
rect 1104 8112 48852 8134
rect 1673 8075 1731 8081
rect 1673 8041 1685 8075
rect 1719 8072 1731 8075
rect 2038 8072 2044 8084
rect 1719 8044 2044 8072
rect 1719 8041 1731 8044
rect 1673 8035 1731 8041
rect 2038 8032 2044 8044
rect 2096 8032 2102 8084
rect 2593 8075 2651 8081
rect 2593 8041 2605 8075
rect 2639 8072 2651 8075
rect 2682 8072 2688 8084
rect 2639 8044 2688 8072
rect 2639 8041 2651 8044
rect 2593 8035 2651 8041
rect 2682 8032 2688 8044
rect 2740 8032 2746 8084
rect 4798 8032 4804 8084
rect 4856 8072 4862 8084
rect 5445 8075 5503 8081
rect 5445 8072 5457 8075
rect 4856 8044 5457 8072
rect 4856 8032 4862 8044
rect 5445 8041 5457 8044
rect 5491 8041 5503 8075
rect 6546 8072 6552 8084
rect 6507 8044 6552 8072
rect 5445 8035 5503 8041
rect 6546 8032 6552 8044
rect 6604 8032 6610 8084
rect 12069 8075 12127 8081
rect 12069 8041 12081 8075
rect 12115 8072 12127 8075
rect 12250 8072 12256 8084
rect 12115 8044 12256 8072
rect 12115 8041 12127 8044
rect 12069 8035 12127 8041
rect 12250 8032 12256 8044
rect 12308 8032 12314 8084
rect 16850 8032 16856 8084
rect 16908 8072 16914 8084
rect 17589 8075 17647 8081
rect 17589 8072 17601 8075
rect 16908 8044 17601 8072
rect 16908 8032 16914 8044
rect 17589 8041 17601 8044
rect 17635 8072 17647 8075
rect 18046 8072 18052 8084
rect 17635 8044 18052 8072
rect 17635 8041 17647 8044
rect 17589 8035 17647 8041
rect 18046 8032 18052 8044
rect 18104 8072 18110 8084
rect 19061 8075 19119 8081
rect 19061 8072 19073 8075
rect 18104 8044 19073 8072
rect 18104 8032 18110 8044
rect 19061 8041 19073 8044
rect 19107 8041 19119 8075
rect 19061 8035 19119 8041
rect 20254 8032 20260 8084
rect 20312 8072 20318 8084
rect 20625 8075 20683 8081
rect 20625 8072 20637 8075
rect 20312 8044 20637 8072
rect 20312 8032 20318 8044
rect 20625 8041 20637 8044
rect 20671 8072 20683 8075
rect 20806 8072 20812 8084
rect 20671 8044 20812 8072
rect 20671 8041 20683 8044
rect 20625 8035 20683 8041
rect 20806 8032 20812 8044
rect 20864 8072 20870 8084
rect 21174 8072 21180 8084
rect 20864 8044 21180 8072
rect 20864 8032 20870 8044
rect 21174 8032 21180 8044
rect 21232 8032 21238 8084
rect 22002 8072 22008 8084
rect 21284 8044 22008 8072
rect 4332 8007 4390 8013
rect 4332 7973 4344 8007
rect 4378 8004 4390 8007
rect 4614 8004 4620 8016
rect 4378 7976 4620 8004
rect 4378 7973 4390 7976
rect 4332 7967 4390 7973
rect 4614 7964 4620 7976
rect 4672 7964 4678 8016
rect 9944 8007 10002 8013
rect 9944 7973 9956 8007
rect 9990 8004 10002 8007
rect 11238 8004 11244 8016
rect 9990 7976 11244 8004
rect 9990 7973 10002 7976
rect 9944 7967 10002 7973
rect 11238 7964 11244 7976
rect 11296 7964 11302 8016
rect 12526 7964 12532 8016
rect 12584 8004 12590 8016
rect 12989 8007 13047 8013
rect 12989 8004 13001 8007
rect 12584 7976 13001 8004
rect 12584 7964 12590 7976
rect 12989 7973 13001 7976
rect 13035 7973 13047 8007
rect 12989 7967 13047 7973
rect 16301 8007 16359 8013
rect 16301 7973 16313 8007
rect 16347 8004 16359 8007
rect 16390 8004 16396 8016
rect 16347 7976 16396 8004
rect 16347 7973 16359 7976
rect 16301 7967 16359 7973
rect 16390 7964 16396 7976
rect 16448 7964 16454 8016
rect 16482 7964 16488 8016
rect 16540 8004 16546 8016
rect 16942 8004 16948 8016
rect 16540 7976 16585 8004
rect 16903 7976 16948 8004
rect 16540 7964 16546 7976
rect 16942 7964 16948 7976
rect 17000 7964 17006 8016
rect 17948 8007 18006 8013
rect 17948 7973 17960 8007
rect 17994 8004 18006 8007
rect 18598 8004 18604 8016
rect 17994 7976 18604 8004
rect 17994 7973 18006 7976
rect 17948 7967 18006 7973
rect 18598 7964 18604 7976
rect 18656 7964 18662 8016
rect 21284 8004 21312 8044
rect 22002 8032 22008 8044
rect 22060 8032 22066 8084
rect 24670 8072 24676 8084
rect 24631 8044 24676 8072
rect 24670 8032 24676 8044
rect 24728 8032 24734 8084
rect 24946 8032 24952 8084
rect 25004 8072 25010 8084
rect 25409 8075 25467 8081
rect 25409 8072 25421 8075
rect 25004 8044 25421 8072
rect 25004 8032 25010 8044
rect 25409 8041 25421 8044
rect 25455 8041 25467 8075
rect 25409 8035 25467 8041
rect 26237 8075 26295 8081
rect 26237 8041 26249 8075
rect 26283 8072 26295 8075
rect 26510 8072 26516 8084
rect 26283 8044 26516 8072
rect 26283 8041 26295 8044
rect 26237 8035 26295 8041
rect 26510 8032 26516 8044
rect 26568 8032 26574 8084
rect 28166 8032 28172 8084
rect 28224 8072 28230 8084
rect 28442 8072 28448 8084
rect 28224 8044 28448 8072
rect 28224 8032 28230 8044
rect 28442 8032 28448 8044
rect 28500 8072 28506 8084
rect 30282 8072 30288 8084
rect 28500 8044 29684 8072
rect 30243 8044 30288 8072
rect 28500 8032 28506 8044
rect 21192 7976 21312 8004
rect 26780 8007 26838 8013
rect 1489 7939 1547 7945
rect 1489 7905 1501 7939
rect 1535 7936 1547 7939
rect 1946 7936 1952 7948
rect 1535 7908 1952 7936
rect 1535 7905 1547 7908
rect 1489 7899 1547 7905
rect 1946 7896 1952 7908
rect 2004 7896 2010 7948
rect 11701 7939 11759 7945
rect 11701 7905 11713 7939
rect 11747 7936 11759 7939
rect 13814 7936 13820 7948
rect 11747 7908 13820 7936
rect 11747 7905 11759 7908
rect 11701 7899 11759 7905
rect 13096 7880 13124 7908
rect 13814 7896 13820 7908
rect 13872 7896 13878 7948
rect 17681 7939 17739 7945
rect 17681 7905 17693 7939
rect 17727 7936 17739 7939
rect 17770 7936 17776 7948
rect 17727 7908 17776 7936
rect 17727 7905 17739 7908
rect 17681 7899 17739 7905
rect 17770 7896 17776 7908
rect 17828 7896 17834 7948
rect 21192 7945 21220 7976
rect 26780 7973 26792 8007
rect 26826 8004 26838 8007
rect 27062 8004 27068 8016
rect 26826 7976 27068 8004
rect 26826 7973 26838 7976
rect 26780 7967 26838 7973
rect 27062 7964 27068 7976
rect 27120 7964 27126 8016
rect 28905 8007 28963 8013
rect 28905 7973 28917 8007
rect 28951 8004 28963 8007
rect 29362 8004 29368 8016
rect 28951 7976 29368 8004
rect 28951 7973 28963 7976
rect 28905 7967 28963 7973
rect 29362 7964 29368 7976
rect 29420 7964 29426 8016
rect 29546 8004 29552 8016
rect 29507 7976 29552 8004
rect 29546 7964 29552 7976
rect 29604 7964 29610 8016
rect 29656 8013 29684 8044
rect 30282 8032 30288 8044
rect 30340 8032 30346 8084
rect 31570 8032 31576 8084
rect 31628 8072 31634 8084
rect 31757 8075 31815 8081
rect 31757 8072 31769 8075
rect 31628 8044 31769 8072
rect 31628 8032 31634 8044
rect 31757 8041 31769 8044
rect 31803 8041 31815 8075
rect 31757 8035 31815 8041
rect 31846 8032 31852 8084
rect 31904 8072 31910 8084
rect 32309 8075 32367 8081
rect 32309 8072 32321 8075
rect 31904 8044 32321 8072
rect 31904 8032 31910 8044
rect 32309 8041 32321 8044
rect 32355 8041 32367 8075
rect 36446 8072 36452 8084
rect 36407 8044 36452 8072
rect 32309 8035 32367 8041
rect 36446 8032 36452 8044
rect 36504 8032 36510 8084
rect 40129 8075 40187 8081
rect 40129 8041 40141 8075
rect 40175 8072 40187 8075
rect 40494 8072 40500 8084
rect 40175 8044 40500 8072
rect 40175 8041 40187 8044
rect 40129 8035 40187 8041
rect 40494 8032 40500 8044
rect 40552 8032 40558 8084
rect 41598 8072 41604 8084
rect 41559 8044 41604 8072
rect 41598 8032 41604 8044
rect 41656 8032 41662 8084
rect 42518 8032 42524 8084
rect 42576 8072 42582 8084
rect 43533 8075 43591 8081
rect 43533 8072 43545 8075
rect 42576 8044 43545 8072
rect 42576 8032 42582 8044
rect 43533 8041 43545 8044
rect 43579 8072 43591 8075
rect 43622 8072 43628 8084
rect 43579 8044 43628 8072
rect 43579 8041 43591 8044
rect 43533 8035 43591 8041
rect 43622 8032 43628 8044
rect 43680 8032 43686 8084
rect 45554 8032 45560 8084
rect 45612 8072 45618 8084
rect 46201 8075 46259 8081
rect 46201 8072 46213 8075
rect 45612 8044 46213 8072
rect 45612 8032 45618 8044
rect 46201 8041 46213 8044
rect 46247 8041 46259 8075
rect 46201 8035 46259 8041
rect 29641 8007 29699 8013
rect 29641 7973 29653 8007
rect 29687 7973 29699 8007
rect 29641 7967 29699 7973
rect 35989 8007 36047 8013
rect 35989 7973 36001 8007
rect 36035 8004 36047 8007
rect 36722 8004 36728 8016
rect 36035 7976 36728 8004
rect 36035 7973 36047 7976
rect 35989 7967 36047 7973
rect 36722 7964 36728 7976
rect 36780 7964 36786 8016
rect 37826 7964 37832 8016
rect 37884 8004 37890 8016
rect 37982 8007 38040 8013
rect 37982 8004 37994 8007
rect 37884 7976 37994 8004
rect 37884 7964 37890 7976
rect 37982 7973 37994 7976
rect 38028 7973 38040 8007
rect 37982 7967 38040 7973
rect 21177 7939 21235 7945
rect 21177 7905 21189 7939
rect 21223 7905 21235 7939
rect 21177 7899 21235 7905
rect 24946 7896 24952 7948
rect 25004 7936 25010 7948
rect 25501 7939 25559 7945
rect 25501 7936 25513 7939
rect 25004 7908 25513 7936
rect 25004 7896 25010 7908
rect 25501 7905 25513 7908
rect 25547 7905 25559 7939
rect 25501 7899 25559 7905
rect 26513 7939 26571 7945
rect 26513 7905 26525 7939
rect 26559 7936 26571 7939
rect 26602 7936 26608 7948
rect 26559 7908 26608 7936
rect 26559 7905 26571 7908
rect 26513 7899 26571 7905
rect 26602 7896 26608 7908
rect 26660 7896 26666 7948
rect 30561 7939 30619 7945
rect 30561 7905 30573 7939
rect 30607 7905 30619 7939
rect 30561 7899 30619 7905
rect 4062 7868 4068 7880
rect 4023 7840 4068 7868
rect 4062 7828 4068 7840
rect 4120 7828 4126 7880
rect 9306 7828 9312 7880
rect 9364 7868 9370 7880
rect 9674 7868 9680 7880
rect 9364 7840 9680 7868
rect 9364 7828 9370 7840
rect 9674 7828 9680 7840
rect 9732 7828 9738 7880
rect 12894 7868 12900 7880
rect 12855 7840 12900 7868
rect 12894 7828 12900 7840
rect 12952 7828 12958 7880
rect 13078 7868 13084 7880
rect 13039 7840 13084 7868
rect 13078 7828 13084 7840
rect 13136 7828 13142 7880
rect 16574 7868 16580 7880
rect 16535 7840 16580 7868
rect 16574 7828 16580 7840
rect 16632 7828 16638 7880
rect 20990 7828 20996 7880
rect 21048 7868 21054 7880
rect 21450 7868 21456 7880
rect 21048 7840 21456 7868
rect 21048 7828 21054 7840
rect 21450 7828 21456 7840
rect 21508 7877 21514 7880
rect 21508 7871 21558 7877
rect 21508 7837 21512 7871
rect 21546 7837 21558 7871
rect 21634 7868 21640 7880
rect 21595 7840 21640 7868
rect 21508 7831 21558 7837
rect 21508 7828 21514 7831
rect 21634 7828 21640 7840
rect 21692 7828 21698 7880
rect 21910 7868 21916 7880
rect 21871 7840 21916 7868
rect 21910 7828 21916 7840
rect 21968 7828 21974 7880
rect 22002 7828 22008 7880
rect 22060 7868 22066 7880
rect 22094 7868 22100 7880
rect 22060 7840 22100 7868
rect 22060 7828 22066 7840
rect 22094 7828 22100 7840
rect 22152 7828 22158 7880
rect 24578 7828 24584 7880
rect 24636 7868 24642 7880
rect 25409 7871 25467 7877
rect 25409 7868 25421 7871
rect 24636 7840 25421 7868
rect 24636 7828 24642 7840
rect 25409 7837 25421 7840
rect 25455 7868 25467 7871
rect 26142 7868 26148 7880
rect 25455 7840 26148 7868
rect 25455 7837 25467 7840
rect 25409 7831 25467 7837
rect 26142 7828 26148 7840
rect 26200 7828 26206 7880
rect 23753 7803 23811 7809
rect 23753 7769 23765 7803
rect 23799 7800 23811 7803
rect 23934 7800 23940 7812
rect 23799 7772 23940 7800
rect 23799 7769 23811 7772
rect 23753 7763 23811 7769
rect 23934 7760 23940 7772
rect 23992 7800 23998 7812
rect 24762 7800 24768 7812
rect 23992 7772 24768 7800
rect 23992 7760 23998 7772
rect 24762 7760 24768 7772
rect 24820 7760 24826 7812
rect 29089 7803 29147 7809
rect 29089 7769 29101 7803
rect 29135 7800 29147 7803
rect 30576 7800 30604 7899
rect 39942 7896 39948 7948
rect 40000 7936 40006 7948
rect 40477 7939 40535 7945
rect 40477 7936 40489 7939
rect 40000 7908 40489 7936
rect 40000 7896 40006 7908
rect 40477 7905 40489 7908
rect 40523 7905 40535 7939
rect 40477 7899 40535 7905
rect 45088 7939 45146 7945
rect 45088 7905 45100 7939
rect 45134 7936 45146 7939
rect 45370 7936 45376 7948
rect 45134 7908 45376 7936
rect 45134 7905 45146 7908
rect 45088 7899 45146 7905
rect 45370 7896 45376 7908
rect 45428 7896 45434 7948
rect 37734 7868 37740 7880
rect 37695 7840 37740 7868
rect 37734 7828 37740 7840
rect 37792 7828 37798 7880
rect 40218 7868 40224 7880
rect 40179 7840 40224 7868
rect 40218 7828 40224 7840
rect 40276 7828 40282 7880
rect 44818 7868 44824 7880
rect 44779 7840 44824 7868
rect 44818 7828 44824 7840
rect 44876 7828 44882 7880
rect 30650 7800 30656 7812
rect 29135 7772 30656 7800
rect 29135 7769 29147 7772
rect 29089 7763 29147 7769
rect 30650 7760 30656 7772
rect 30708 7760 30714 7812
rect 6914 7732 6920 7744
rect 6875 7704 6920 7732
rect 6914 7692 6920 7704
rect 6972 7692 6978 7744
rect 11057 7735 11115 7741
rect 11057 7701 11069 7735
rect 11103 7732 11115 7735
rect 11790 7732 11796 7744
rect 11103 7704 11796 7732
rect 11103 7701 11115 7704
rect 11057 7695 11115 7701
rect 11790 7692 11796 7704
rect 11848 7692 11854 7744
rect 12529 7735 12587 7741
rect 12529 7701 12541 7735
rect 12575 7732 12587 7735
rect 13814 7732 13820 7744
rect 12575 7704 13820 7732
rect 12575 7701 12587 7704
rect 12529 7695 12587 7701
rect 13814 7692 13820 7704
rect 13872 7692 13878 7744
rect 15010 7732 15016 7744
rect 14971 7704 15016 7732
rect 15010 7692 15016 7704
rect 15068 7692 15074 7744
rect 16022 7732 16028 7744
rect 15983 7704 16028 7732
rect 16022 7692 16028 7704
rect 16080 7692 16086 7744
rect 20806 7692 20812 7744
rect 20864 7732 20870 7744
rect 21634 7732 21640 7744
rect 20864 7704 21640 7732
rect 20864 7692 20870 7704
rect 21634 7692 21640 7704
rect 21692 7692 21698 7744
rect 23017 7735 23075 7741
rect 23017 7701 23029 7735
rect 23063 7732 23075 7735
rect 23290 7732 23296 7744
rect 23063 7704 23296 7732
rect 23063 7701 23075 7704
rect 23017 7695 23075 7701
rect 23290 7692 23296 7704
rect 23348 7692 23354 7744
rect 24949 7735 25007 7741
rect 24949 7701 24961 7735
rect 24995 7732 25007 7735
rect 25314 7732 25320 7744
rect 24995 7704 25320 7732
rect 24995 7701 25007 7704
rect 24949 7695 25007 7701
rect 25314 7692 25320 7704
rect 25372 7692 25378 7744
rect 27614 7692 27620 7744
rect 27672 7732 27678 7744
rect 27893 7735 27951 7741
rect 27893 7732 27905 7735
rect 27672 7704 27905 7732
rect 27672 7692 27678 7704
rect 27893 7701 27905 7704
rect 27939 7701 27951 7735
rect 30742 7732 30748 7744
rect 30703 7704 30748 7732
rect 27893 7695 27951 7701
rect 30742 7692 30748 7704
rect 30800 7692 30806 7744
rect 38378 7692 38384 7744
rect 38436 7732 38442 7744
rect 39117 7735 39175 7741
rect 39117 7732 39129 7735
rect 38436 7704 39129 7732
rect 38436 7692 38442 7704
rect 39117 7701 39129 7704
rect 39163 7732 39175 7735
rect 39942 7732 39948 7744
rect 39163 7704 39948 7732
rect 39163 7701 39175 7704
rect 39117 7695 39175 7701
rect 39942 7692 39948 7704
rect 40000 7692 40006 7744
rect 43070 7732 43076 7744
rect 43031 7704 43076 7732
rect 43070 7692 43076 7704
rect 43128 7692 43134 7744
rect 1104 7642 48852 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 34966 7642
rect 35018 7590 35030 7642
rect 35082 7590 35094 7642
rect 35146 7590 35158 7642
rect 35210 7590 48852 7642
rect 1104 7568 48852 7590
rect 4525 7531 4583 7537
rect 4525 7497 4537 7531
rect 4571 7528 4583 7531
rect 4614 7528 4620 7540
rect 4571 7500 4620 7528
rect 4571 7497 4583 7500
rect 4525 7491 4583 7497
rect 4614 7488 4620 7500
rect 4672 7488 4678 7540
rect 11238 7528 11244 7540
rect 11199 7500 11244 7528
rect 11238 7488 11244 7500
rect 11296 7488 11302 7540
rect 11974 7488 11980 7540
rect 12032 7528 12038 7540
rect 12161 7531 12219 7537
rect 12161 7528 12173 7531
rect 12032 7500 12173 7528
rect 12032 7488 12038 7500
rect 12161 7497 12173 7500
rect 12207 7497 12219 7531
rect 12802 7528 12808 7540
rect 12161 7491 12219 7497
rect 12452 7500 12808 7528
rect 5261 7463 5319 7469
rect 5261 7429 5273 7463
rect 5307 7460 5319 7463
rect 5442 7460 5448 7472
rect 5307 7432 5448 7460
rect 5307 7429 5319 7432
rect 5261 7423 5319 7429
rect 5442 7420 5448 7432
rect 5500 7420 5506 7472
rect 11885 7395 11943 7401
rect 11885 7361 11897 7395
rect 11931 7392 11943 7395
rect 12452 7392 12480 7500
rect 12802 7488 12808 7500
rect 12860 7488 12866 7540
rect 16390 7528 16396 7540
rect 16351 7500 16396 7528
rect 16390 7488 16396 7500
rect 16448 7488 16454 7540
rect 17770 7528 17776 7540
rect 17731 7500 17776 7528
rect 17770 7488 17776 7500
rect 17828 7488 17834 7540
rect 20254 7528 20260 7540
rect 20215 7500 20260 7528
rect 20254 7488 20260 7500
rect 20312 7488 20318 7540
rect 20625 7531 20683 7537
rect 20625 7497 20637 7531
rect 20671 7528 20683 7531
rect 20898 7528 20904 7540
rect 20671 7500 20904 7528
rect 20671 7497 20683 7500
rect 20625 7491 20683 7497
rect 20898 7488 20904 7500
rect 20956 7488 20962 7540
rect 21634 7488 21640 7540
rect 21692 7528 21698 7540
rect 22465 7531 22523 7537
rect 22465 7528 22477 7531
rect 21692 7500 22477 7528
rect 21692 7488 21698 7500
rect 22465 7497 22477 7500
rect 22511 7497 22523 7531
rect 24578 7528 24584 7540
rect 24539 7500 24584 7528
rect 22465 7491 22523 7497
rect 24578 7488 24584 7500
rect 24636 7488 24642 7540
rect 24854 7528 24860 7540
rect 24815 7500 24860 7528
rect 24854 7488 24860 7500
rect 24912 7488 24918 7540
rect 26973 7531 27031 7537
rect 26973 7497 26985 7531
rect 27019 7528 27031 7531
rect 27062 7528 27068 7540
rect 27019 7500 27068 7528
rect 27019 7497 27031 7500
rect 26973 7491 27031 7497
rect 27062 7488 27068 7500
rect 27120 7488 27126 7540
rect 29546 7488 29552 7540
rect 29604 7528 29610 7540
rect 29641 7531 29699 7537
rect 29641 7528 29653 7531
rect 29604 7500 29653 7528
rect 29604 7488 29610 7500
rect 29641 7497 29653 7500
rect 29687 7528 29699 7531
rect 30561 7531 30619 7537
rect 30561 7528 30573 7531
rect 29687 7500 30573 7528
rect 29687 7497 29699 7500
rect 29641 7491 29699 7497
rect 30561 7497 30573 7500
rect 30607 7497 30619 7531
rect 30561 7491 30619 7497
rect 31021 7531 31079 7537
rect 31021 7497 31033 7531
rect 31067 7528 31079 7531
rect 31478 7528 31484 7540
rect 31067 7500 31484 7528
rect 31067 7497 31079 7500
rect 31021 7491 31079 7497
rect 15013 7463 15071 7469
rect 15013 7429 15025 7463
rect 15059 7460 15071 7463
rect 15102 7460 15108 7472
rect 15059 7432 15108 7460
rect 15059 7429 15071 7432
rect 15013 7423 15071 7429
rect 15102 7420 15108 7432
rect 15160 7420 15166 7472
rect 16025 7463 16083 7469
rect 16025 7429 16037 7463
rect 16071 7460 16083 7463
rect 16482 7460 16488 7472
rect 16071 7432 16488 7460
rect 16071 7429 16083 7432
rect 16025 7423 16083 7429
rect 16482 7420 16488 7432
rect 16540 7460 16546 7472
rect 18141 7463 18199 7469
rect 18141 7460 18153 7463
rect 16540 7432 18153 7460
rect 16540 7420 16546 7432
rect 18141 7429 18153 7432
rect 18187 7429 18199 7463
rect 20806 7460 20812 7472
rect 20767 7432 20812 7460
rect 18141 7423 18199 7429
rect 20806 7420 20812 7432
rect 20864 7420 20870 7472
rect 11931 7364 12480 7392
rect 17405 7395 17463 7401
rect 11931 7361 11943 7364
rect 11885 7355 11943 7361
rect 17405 7361 17417 7395
rect 17451 7392 17463 7395
rect 18598 7392 18604 7404
rect 17451 7364 18604 7392
rect 17451 7361 17463 7364
rect 17405 7355 17463 7361
rect 18598 7352 18604 7364
rect 18656 7352 18662 7404
rect 20916 7392 20944 7488
rect 21174 7420 21180 7472
rect 21232 7460 21238 7472
rect 21232 7432 21404 7460
rect 21232 7420 21238 7432
rect 21376 7401 21404 7432
rect 21450 7420 21456 7472
rect 21508 7460 21514 7472
rect 21729 7463 21787 7469
rect 21729 7460 21741 7463
rect 21508 7432 21741 7460
rect 21508 7420 21514 7432
rect 21729 7429 21741 7432
rect 21775 7429 21787 7463
rect 21729 7423 21787 7429
rect 21269 7395 21327 7401
rect 21269 7392 21281 7395
rect 20916 7364 21281 7392
rect 21269 7361 21281 7364
rect 21315 7361 21327 7395
rect 21269 7355 21327 7361
rect 21361 7395 21419 7401
rect 21361 7361 21373 7395
rect 21407 7361 21419 7395
rect 21744 7392 21772 7423
rect 21910 7420 21916 7472
rect 21968 7460 21974 7472
rect 22097 7463 22155 7469
rect 22097 7460 22109 7463
rect 21968 7432 22109 7460
rect 21968 7420 21974 7432
rect 22097 7429 22109 7432
rect 22143 7429 22155 7463
rect 27706 7460 27712 7472
rect 27667 7432 27712 7460
rect 22097 7423 22155 7429
rect 27706 7420 27712 7432
rect 27764 7420 27770 7472
rect 22002 7392 22008 7404
rect 21744 7364 22008 7392
rect 21361 7355 21419 7361
rect 22002 7352 22008 7364
rect 22060 7352 22066 7404
rect 28169 7395 28227 7401
rect 28169 7361 28181 7395
rect 28215 7392 28227 7395
rect 28258 7392 28264 7404
rect 28215 7364 28264 7392
rect 28215 7361 28227 7364
rect 28169 7355 28227 7361
rect 28258 7352 28264 7364
rect 28316 7392 28322 7404
rect 28629 7395 28687 7401
rect 28629 7392 28641 7395
rect 28316 7364 28641 7392
rect 28316 7352 28322 7364
rect 28629 7361 28641 7364
rect 28675 7361 28687 7395
rect 28629 7355 28687 7361
rect 29638 7352 29644 7404
rect 29696 7392 29702 7404
rect 30190 7392 30196 7404
rect 29696 7364 30196 7392
rect 29696 7352 29702 7364
rect 30190 7352 30196 7364
rect 30248 7352 30254 7404
rect 31128 7401 31156 7500
rect 31478 7488 31484 7500
rect 31536 7488 31542 7540
rect 32490 7528 32496 7540
rect 32451 7500 32496 7528
rect 32490 7488 32496 7500
rect 32548 7488 32554 7540
rect 37001 7531 37059 7537
rect 37001 7497 37013 7531
rect 37047 7528 37059 7531
rect 37369 7531 37427 7537
rect 37369 7528 37381 7531
rect 37047 7500 37381 7528
rect 37047 7497 37059 7500
rect 37001 7491 37059 7497
rect 37369 7497 37381 7500
rect 37415 7528 37427 7531
rect 37826 7528 37832 7540
rect 37415 7500 37832 7528
rect 37415 7497 37427 7500
rect 37369 7491 37427 7497
rect 37826 7488 37832 7500
rect 37884 7488 37890 7540
rect 37918 7488 37924 7540
rect 37976 7528 37982 7540
rect 39942 7528 39948 7540
rect 37976 7500 38021 7528
rect 39903 7500 39948 7528
rect 37976 7488 37982 7500
rect 39942 7488 39948 7500
rect 40000 7488 40006 7540
rect 42429 7531 42487 7537
rect 42429 7497 42441 7531
rect 42475 7528 42487 7531
rect 42518 7528 42524 7540
rect 42475 7500 42524 7528
rect 42475 7497 42487 7500
rect 42429 7491 42487 7497
rect 42518 7488 42524 7500
rect 42576 7488 42582 7540
rect 36722 7420 36728 7472
rect 36780 7460 36786 7472
rect 36780 7432 38516 7460
rect 36780 7420 36786 7432
rect 31113 7395 31171 7401
rect 31113 7361 31125 7395
rect 31159 7361 31171 7395
rect 38378 7392 38384 7404
rect 38339 7364 38384 7392
rect 31113 7355 31171 7361
rect 38378 7352 38384 7364
rect 38436 7352 38442 7404
rect 38488 7401 38516 7432
rect 38473 7395 38531 7401
rect 38473 7361 38485 7395
rect 38519 7392 38531 7395
rect 38933 7395 38991 7401
rect 38933 7392 38945 7395
rect 38519 7364 38945 7392
rect 38519 7361 38531 7364
rect 38473 7355 38531 7361
rect 38933 7361 38945 7364
rect 38979 7392 38991 7395
rect 39942 7392 39948 7404
rect 38979 7364 39948 7392
rect 38979 7361 38991 7364
rect 38933 7355 38991 7361
rect 39942 7352 39948 7364
rect 40000 7352 40006 7404
rect 9306 7324 9312 7336
rect 9140 7296 9312 7324
rect 5534 7256 5540 7268
rect 5495 7228 5540 7256
rect 5534 7216 5540 7228
rect 5592 7216 5598 7268
rect 5626 7216 5632 7268
rect 5684 7256 5690 7268
rect 5813 7259 5871 7265
rect 5813 7256 5825 7259
rect 5684 7228 5825 7256
rect 5684 7216 5690 7228
rect 5813 7225 5825 7228
rect 5859 7225 5871 7259
rect 5813 7219 5871 7225
rect 1673 7191 1731 7197
rect 1673 7157 1685 7191
rect 1719 7188 1731 7191
rect 1946 7188 1952 7200
rect 1719 7160 1952 7188
rect 1719 7157 1731 7160
rect 1673 7151 1731 7157
rect 1946 7148 1952 7160
rect 2004 7148 2010 7200
rect 4154 7188 4160 7200
rect 4115 7160 4160 7188
rect 4154 7148 4160 7160
rect 4212 7148 4218 7200
rect 5077 7191 5135 7197
rect 5077 7157 5089 7191
rect 5123 7188 5135 7191
rect 5718 7188 5724 7200
rect 5123 7160 5724 7188
rect 5123 7157 5135 7160
rect 5077 7151 5135 7157
rect 5718 7148 5724 7160
rect 5776 7148 5782 7200
rect 6914 7148 6920 7200
rect 6972 7188 6978 7200
rect 9140 7197 9168 7296
rect 9306 7284 9312 7296
rect 9364 7284 9370 7336
rect 11974 7284 11980 7336
rect 12032 7324 12038 7336
rect 12342 7324 12348 7336
rect 12032 7296 12348 7324
rect 12032 7284 12038 7296
rect 12342 7284 12348 7296
rect 12400 7324 12406 7336
rect 12437 7327 12495 7333
rect 12437 7324 12449 7327
rect 12400 7296 12449 7324
rect 12400 7284 12406 7296
rect 12437 7293 12449 7296
rect 12483 7293 12495 7327
rect 12437 7287 12495 7293
rect 14829 7327 14887 7333
rect 14829 7293 14841 7327
rect 14875 7324 14887 7327
rect 14875 7296 15424 7324
rect 14875 7293 14887 7296
rect 14829 7287 14887 7293
rect 15396 7268 15424 7296
rect 16942 7284 16948 7336
rect 17000 7324 17006 7336
rect 18693 7327 18751 7333
rect 18693 7324 18705 7327
rect 17000 7296 18705 7324
rect 17000 7284 17006 7296
rect 18693 7293 18705 7296
rect 18739 7324 18751 7327
rect 19061 7327 19119 7333
rect 19061 7324 19073 7327
rect 18739 7296 19073 7324
rect 18739 7293 18751 7296
rect 18693 7287 18751 7293
rect 19061 7293 19073 7296
rect 19107 7293 19119 7327
rect 19061 7287 19119 7293
rect 19889 7327 19947 7333
rect 19889 7293 19901 7327
rect 19935 7324 19947 7327
rect 21174 7324 21180 7336
rect 19935 7296 21180 7324
rect 19935 7293 19947 7296
rect 19889 7287 19947 7293
rect 21174 7284 21180 7296
rect 21232 7324 21238 7336
rect 21232 7296 21312 7324
rect 21232 7284 21238 7296
rect 9582 7265 9588 7268
rect 9576 7256 9588 7265
rect 9543 7228 9588 7256
rect 9576 7219 9588 7228
rect 9582 7216 9588 7219
rect 9640 7216 9646 7268
rect 12704 7259 12762 7265
rect 12704 7225 12716 7259
rect 12750 7256 12762 7259
rect 12894 7256 12900 7268
rect 12750 7228 12900 7256
rect 12750 7225 12762 7228
rect 12704 7219 12762 7225
rect 12894 7216 12900 7228
rect 12952 7216 12958 7268
rect 15286 7256 15292 7268
rect 15247 7228 15292 7256
rect 15286 7216 15292 7228
rect 15344 7216 15350 7268
rect 15378 7216 15384 7268
rect 15436 7256 15442 7268
rect 15473 7259 15531 7265
rect 15473 7256 15485 7259
rect 15436 7228 15485 7256
rect 15436 7216 15442 7228
rect 15473 7225 15485 7228
rect 15519 7225 15531 7259
rect 15473 7219 15531 7225
rect 15565 7259 15623 7265
rect 15565 7225 15577 7259
rect 15611 7256 15623 7259
rect 15611 7228 15645 7256
rect 15611 7225 15623 7228
rect 15565 7219 15623 7225
rect 8757 7191 8815 7197
rect 8757 7188 8769 7191
rect 6972 7160 8769 7188
rect 6972 7148 6978 7160
rect 8757 7157 8769 7160
rect 8803 7188 8815 7191
rect 9125 7191 9183 7197
rect 9125 7188 9137 7191
rect 8803 7160 9137 7188
rect 8803 7157 8815 7160
rect 8757 7151 8815 7157
rect 9125 7157 9137 7160
rect 9171 7157 9183 7191
rect 9125 7151 9183 7157
rect 10226 7148 10232 7200
rect 10284 7188 10290 7200
rect 10689 7191 10747 7197
rect 10689 7188 10701 7191
rect 10284 7160 10701 7188
rect 10284 7148 10290 7160
rect 10689 7157 10701 7160
rect 10735 7157 10747 7191
rect 10689 7151 10747 7157
rect 12342 7148 12348 7200
rect 12400 7188 12406 7200
rect 12434 7188 12440 7200
rect 12400 7160 12440 7188
rect 12400 7148 12406 7160
rect 12434 7148 12440 7160
rect 12492 7148 12498 7200
rect 13817 7191 13875 7197
rect 13817 7157 13829 7191
rect 13863 7188 13875 7191
rect 13906 7188 13912 7200
rect 13863 7160 13912 7188
rect 13863 7157 13875 7160
rect 13817 7151 13875 7157
rect 13906 7148 13912 7160
rect 13964 7148 13970 7200
rect 15010 7148 15016 7200
rect 15068 7188 15074 7200
rect 15580 7188 15608 7219
rect 18506 7216 18512 7268
rect 18564 7256 18570 7268
rect 21284 7265 21312 7296
rect 22094 7284 22100 7336
rect 22152 7324 22158 7336
rect 22554 7324 22560 7336
rect 22152 7296 22560 7324
rect 22152 7284 22158 7296
rect 22554 7284 22560 7296
rect 22612 7324 22618 7336
rect 22833 7327 22891 7333
rect 22833 7324 22845 7327
rect 22612 7296 22845 7324
rect 22612 7284 22618 7296
rect 22833 7293 22845 7296
rect 22879 7293 22891 7327
rect 25314 7324 25320 7336
rect 25275 7296 25320 7324
rect 22833 7287 22891 7293
rect 25314 7284 25320 7296
rect 25372 7324 25378 7336
rect 25869 7327 25927 7333
rect 25869 7324 25881 7327
rect 25372 7296 25881 7324
rect 25372 7284 25378 7296
rect 25869 7293 25881 7296
rect 25915 7293 25927 7327
rect 25869 7287 25927 7293
rect 29730 7284 29736 7336
rect 29788 7324 29794 7336
rect 29917 7327 29975 7333
rect 29917 7324 29929 7327
rect 29788 7296 29929 7324
rect 29788 7284 29794 7296
rect 29917 7293 29929 7296
rect 29963 7324 29975 7327
rect 33594 7324 33600 7336
rect 29963 7296 30512 7324
rect 33555 7296 33600 7324
rect 29963 7293 29975 7296
rect 29917 7287 29975 7293
rect 18601 7259 18659 7265
rect 18601 7256 18613 7259
rect 18564 7228 18613 7256
rect 18564 7216 18570 7228
rect 18601 7225 18613 7228
rect 18647 7225 18659 7259
rect 18601 7219 18659 7225
rect 21269 7259 21327 7265
rect 21269 7225 21281 7259
rect 21315 7225 21327 7259
rect 28258 7256 28264 7268
rect 28219 7228 28264 7256
rect 21269 7219 21327 7225
rect 28258 7216 28264 7228
rect 28316 7216 28322 7268
rect 30484 7256 30512 7296
rect 33594 7284 33600 7296
rect 33652 7324 33658 7336
rect 34149 7327 34207 7333
rect 34149 7324 34161 7327
rect 33652 7296 34161 7324
rect 33652 7284 33658 7296
rect 34149 7293 34161 7296
rect 34195 7293 34207 7327
rect 40310 7324 40316 7336
rect 40223 7296 40316 7324
rect 34149 7287 34207 7293
rect 40310 7284 40316 7296
rect 40368 7324 40374 7336
rect 40678 7324 40684 7336
rect 40368 7296 40684 7324
rect 40368 7284 40374 7296
rect 40678 7284 40684 7296
rect 40736 7324 40742 7336
rect 40957 7327 41015 7333
rect 40957 7324 40969 7327
rect 40736 7296 40969 7324
rect 40736 7284 40742 7296
rect 40957 7293 40969 7296
rect 41003 7324 41015 7327
rect 41049 7327 41107 7333
rect 41049 7324 41061 7327
rect 41003 7296 41061 7324
rect 41003 7293 41015 7296
rect 40957 7287 41015 7293
rect 41049 7293 41061 7296
rect 41095 7324 41107 7327
rect 43533 7327 43591 7333
rect 43533 7324 43545 7327
rect 41095 7296 43545 7324
rect 41095 7293 41107 7296
rect 41049 7287 41107 7293
rect 43533 7293 43545 7296
rect 43579 7293 43591 7327
rect 43533 7287 43591 7293
rect 31202 7256 31208 7268
rect 30484 7228 31208 7256
rect 31202 7216 31208 7228
rect 31260 7256 31266 7268
rect 31358 7259 31416 7265
rect 31358 7256 31370 7259
rect 31260 7228 31370 7256
rect 31260 7216 31266 7228
rect 31358 7225 31370 7228
rect 31404 7225 31416 7259
rect 31358 7219 31416 7225
rect 40494 7216 40500 7268
rect 40552 7256 40558 7268
rect 41138 7256 41144 7268
rect 40552 7228 41144 7256
rect 40552 7216 40558 7228
rect 41138 7216 41144 7228
rect 41196 7256 41202 7268
rect 41294 7259 41352 7265
rect 41294 7256 41306 7259
rect 41196 7228 41306 7256
rect 41196 7216 41202 7228
rect 41294 7225 41306 7228
rect 41340 7225 41352 7259
rect 43438 7256 43444 7268
rect 43351 7228 43444 7256
rect 41294 7219 41352 7225
rect 43438 7216 43444 7228
rect 43496 7256 43502 7268
rect 43548 7256 43576 7287
rect 43622 7284 43628 7336
rect 43680 7324 43686 7336
rect 43789 7327 43847 7333
rect 43789 7324 43801 7327
rect 43680 7296 43801 7324
rect 43680 7284 43686 7296
rect 43789 7293 43801 7296
rect 43835 7293 43847 7327
rect 43789 7287 43847 7293
rect 46753 7327 46811 7333
rect 46753 7293 46765 7327
rect 46799 7324 46811 7327
rect 46799 7296 47440 7324
rect 46799 7293 46811 7296
rect 46753 7287 46811 7293
rect 44818 7256 44824 7268
rect 43496 7228 44824 7256
rect 43496 7216 43502 7228
rect 44818 7216 44824 7228
rect 44876 7256 44882 7268
rect 44876 7228 45600 7256
rect 44876 7216 44882 7228
rect 16574 7188 16580 7200
rect 15068 7160 16580 7188
rect 15068 7148 15074 7160
rect 16574 7148 16580 7160
rect 16632 7188 16638 7200
rect 16669 7191 16727 7197
rect 16669 7188 16681 7191
rect 16632 7160 16681 7188
rect 16632 7148 16638 7160
rect 16669 7157 16681 7160
rect 16715 7157 16727 7191
rect 16669 7151 16727 7157
rect 23474 7148 23480 7200
rect 23532 7188 23538 7200
rect 23661 7191 23719 7197
rect 23661 7188 23673 7191
rect 23532 7160 23673 7188
rect 23532 7148 23538 7160
rect 23661 7157 23673 7160
rect 23707 7157 23719 7191
rect 25498 7188 25504 7200
rect 25459 7160 25504 7188
rect 23661 7151 23719 7157
rect 25498 7148 25504 7160
rect 25556 7148 25562 7200
rect 26602 7188 26608 7200
rect 26563 7160 26608 7188
rect 26602 7148 26608 7160
rect 26660 7148 26666 7200
rect 27525 7191 27583 7197
rect 27525 7157 27537 7191
rect 27571 7188 27583 7191
rect 28166 7188 28172 7200
rect 27571 7160 28172 7188
rect 27571 7157 27583 7160
rect 27525 7151 27583 7157
rect 28166 7148 28172 7160
rect 28224 7148 28230 7200
rect 29089 7191 29147 7197
rect 29089 7157 29101 7191
rect 29135 7188 29147 7191
rect 30101 7191 30159 7197
rect 30101 7188 30113 7191
rect 29135 7160 30113 7188
rect 29135 7157 29147 7160
rect 29089 7151 29147 7157
rect 30101 7157 30113 7160
rect 30147 7188 30159 7191
rect 30466 7188 30472 7200
rect 30147 7160 30472 7188
rect 30147 7157 30159 7160
rect 30101 7151 30159 7157
rect 30466 7148 30472 7160
rect 30524 7148 30530 7200
rect 33778 7188 33784 7200
rect 33739 7160 33784 7188
rect 33778 7148 33784 7160
rect 33836 7148 33842 7200
rect 37274 7148 37280 7200
rect 37332 7188 37338 7200
rect 37645 7191 37703 7197
rect 37645 7188 37657 7191
rect 37332 7160 37657 7188
rect 37332 7148 37338 7160
rect 37645 7157 37657 7160
rect 37691 7188 37703 7191
rect 37734 7188 37740 7200
rect 37691 7160 37740 7188
rect 37691 7157 37703 7160
rect 37645 7151 37703 7157
rect 37734 7148 37740 7160
rect 37792 7148 37798 7200
rect 37826 7148 37832 7200
rect 37884 7188 37890 7200
rect 38381 7191 38439 7197
rect 38381 7188 38393 7191
rect 37884 7160 38393 7188
rect 37884 7148 37890 7160
rect 38381 7157 38393 7160
rect 38427 7157 38439 7191
rect 38381 7151 38439 7157
rect 44174 7148 44180 7200
rect 44232 7188 44238 7200
rect 45572 7197 45600 7228
rect 47412 7200 47440 7296
rect 44913 7191 44971 7197
rect 44913 7188 44925 7191
rect 44232 7160 44925 7188
rect 44232 7148 44238 7160
rect 44913 7157 44925 7160
rect 44959 7157 44971 7191
rect 44913 7151 44971 7157
rect 45557 7191 45615 7197
rect 45557 7157 45569 7191
rect 45603 7188 45615 7191
rect 45830 7188 45836 7200
rect 45603 7160 45836 7188
rect 45603 7157 45615 7160
rect 45557 7151 45615 7157
rect 45830 7148 45836 7160
rect 45888 7148 45894 7200
rect 46934 7188 46940 7200
rect 46895 7160 46940 7188
rect 46934 7148 46940 7160
rect 46992 7148 46998 7200
rect 47394 7188 47400 7200
rect 47355 7160 47400 7188
rect 47394 7148 47400 7160
rect 47452 7148 47458 7200
rect 1104 7098 48852 7120
rect 1104 7046 19606 7098
rect 19658 7046 19670 7098
rect 19722 7046 19734 7098
rect 19786 7046 19798 7098
rect 19850 7046 48852 7098
rect 1104 7024 48852 7046
rect 9401 6987 9459 6993
rect 9401 6953 9413 6987
rect 9447 6984 9459 6987
rect 9582 6984 9588 6996
rect 9447 6956 9588 6984
rect 9447 6953 9459 6956
rect 9401 6947 9459 6953
rect 9582 6944 9588 6956
rect 9640 6944 9646 6996
rect 10226 6984 10232 6996
rect 10187 6956 10232 6984
rect 10226 6944 10232 6956
rect 10284 6944 10290 6996
rect 11238 6944 11244 6996
rect 11296 6984 11302 6996
rect 11606 6984 11612 6996
rect 11296 6956 11612 6984
rect 11296 6944 11302 6956
rect 11606 6944 11612 6956
rect 11664 6984 11670 6996
rect 11793 6987 11851 6993
rect 11793 6984 11805 6987
rect 11664 6956 11805 6984
rect 11664 6944 11670 6956
rect 11793 6953 11805 6956
rect 11839 6953 11851 6987
rect 12526 6984 12532 6996
rect 12487 6956 12532 6984
rect 11793 6947 11851 6953
rect 12526 6944 12532 6956
rect 12584 6944 12590 6996
rect 12894 6984 12900 6996
rect 12855 6956 12900 6984
rect 12894 6944 12900 6956
rect 12952 6944 12958 6996
rect 15286 6944 15292 6996
rect 15344 6944 15350 6996
rect 18509 6987 18567 6993
rect 18509 6953 18521 6987
rect 18555 6984 18567 6987
rect 18598 6984 18604 6996
rect 18555 6956 18604 6984
rect 18555 6953 18567 6956
rect 18509 6947 18567 6953
rect 18598 6944 18604 6956
rect 18656 6944 18662 6996
rect 29730 6984 29736 6996
rect 29691 6956 29736 6984
rect 29730 6944 29736 6956
rect 29788 6944 29794 6996
rect 30650 6984 30656 6996
rect 30611 6956 30656 6984
rect 30650 6944 30656 6956
rect 30708 6944 30714 6996
rect 38378 6984 38384 6996
rect 38339 6956 38384 6984
rect 38378 6944 38384 6956
rect 38436 6944 38442 6996
rect 41138 6984 41144 6996
rect 41099 6956 41144 6984
rect 41138 6944 41144 6956
rect 41196 6944 41202 6996
rect 3326 6876 3332 6928
rect 3384 6916 3390 6928
rect 4154 6916 4160 6928
rect 3384 6888 4160 6916
rect 3384 6876 3390 6888
rect 4154 6876 4160 6888
rect 4212 6916 4218 6928
rect 4212 6888 5488 6916
rect 4212 6876 4218 6888
rect 2869 6851 2927 6857
rect 2869 6817 2881 6851
rect 2915 6848 2927 6851
rect 3234 6848 3240 6860
rect 2915 6820 3240 6848
rect 2915 6817 2927 6820
rect 2869 6811 2927 6817
rect 3234 6808 3240 6820
rect 3292 6808 3298 6860
rect 5460 6848 5488 6888
rect 5534 6876 5540 6928
rect 5592 6916 5598 6928
rect 6822 6916 6828 6928
rect 5592 6888 6828 6916
rect 5592 6876 5598 6888
rect 6822 6876 6828 6888
rect 6880 6876 6886 6928
rect 15304 6916 15332 6944
rect 21637 6919 21695 6925
rect 21637 6916 21649 6919
rect 15120 6888 15332 6916
rect 21376 6888 21649 6916
rect 6178 6857 6184 6860
rect 5460 6820 5948 6848
rect 5920 6792 5948 6820
rect 6172 6811 6184 6857
rect 6236 6848 6242 6860
rect 10042 6848 10048 6860
rect 6236 6820 6272 6848
rect 10003 6820 10048 6848
rect 6178 6808 6184 6811
rect 6236 6808 6242 6820
rect 10042 6808 10048 6820
rect 10100 6808 10106 6860
rect 11885 6851 11943 6857
rect 11885 6848 11897 6851
rect 10336 6820 11897 6848
rect 5534 6780 5540 6792
rect 5184 6752 5540 6780
rect 3053 6715 3111 6721
rect 3053 6681 3065 6715
rect 3099 6712 3111 6715
rect 3970 6712 3976 6724
rect 3099 6684 3976 6712
rect 3099 6681 3111 6684
rect 3053 6675 3111 6681
rect 3970 6672 3976 6684
rect 4028 6672 4034 6724
rect 4154 6672 4160 6724
rect 4212 6712 4218 6724
rect 5184 6721 5212 6752
rect 5534 6740 5540 6752
rect 5592 6740 5598 6792
rect 5902 6780 5908 6792
rect 5863 6752 5908 6780
rect 5902 6740 5908 6752
rect 5960 6740 5966 6792
rect 9490 6740 9496 6792
rect 9548 6780 9554 6792
rect 10336 6789 10364 6820
rect 11885 6817 11897 6820
rect 11931 6848 11943 6851
rect 11974 6848 11980 6860
rect 11931 6820 11980 6848
rect 11931 6817 11943 6820
rect 11885 6811 11943 6817
rect 11974 6808 11980 6820
rect 12032 6808 12038 6860
rect 13814 6808 13820 6860
rect 13872 6848 13878 6860
rect 14921 6851 14979 6857
rect 14921 6848 14933 6851
rect 13872 6820 14933 6848
rect 13872 6808 13878 6820
rect 14921 6817 14933 6820
rect 14967 6848 14979 6851
rect 15120 6848 15148 6888
rect 21376 6860 21404 6888
rect 21637 6885 21649 6888
rect 21683 6885 21695 6919
rect 28258 6916 28264 6928
rect 21637 6879 21695 6885
rect 27540 6888 28264 6916
rect 14967 6820 15148 6848
rect 14967 6817 14979 6820
rect 14921 6811 14979 6817
rect 15194 6808 15200 6860
rect 15252 6848 15258 6860
rect 15289 6851 15347 6857
rect 15289 6848 15301 6851
rect 15252 6820 15301 6848
rect 15252 6808 15258 6820
rect 15289 6817 15301 6820
rect 15335 6848 15347 6851
rect 15470 6848 15476 6860
rect 15335 6820 15476 6848
rect 15335 6817 15347 6820
rect 15289 6811 15347 6817
rect 15470 6808 15476 6820
rect 15528 6808 15534 6860
rect 16022 6808 16028 6860
rect 16080 6848 16086 6860
rect 16390 6848 16396 6860
rect 16080 6820 16396 6848
rect 16080 6808 16086 6820
rect 16390 6808 16396 6820
rect 16448 6808 16454 6860
rect 18141 6851 18199 6857
rect 18141 6817 18153 6851
rect 18187 6848 18199 6851
rect 18506 6848 18512 6860
rect 18187 6820 18512 6848
rect 18187 6817 18199 6820
rect 18141 6811 18199 6817
rect 18506 6808 18512 6820
rect 18564 6808 18570 6860
rect 21358 6808 21364 6860
rect 21416 6808 21422 6860
rect 21453 6851 21511 6857
rect 21453 6817 21465 6851
rect 21499 6848 21511 6851
rect 21910 6848 21916 6860
rect 21499 6820 21916 6848
rect 21499 6817 21511 6820
rect 21453 6811 21511 6817
rect 21910 6808 21916 6820
rect 21968 6808 21974 6860
rect 24946 6848 24952 6860
rect 24907 6820 24952 6848
rect 24946 6808 24952 6820
rect 25004 6808 25010 6860
rect 26513 6851 26571 6857
rect 26513 6817 26525 6851
rect 26559 6848 26571 6851
rect 26878 6848 26884 6860
rect 26559 6820 26884 6848
rect 26559 6817 26571 6820
rect 26513 6811 26571 6817
rect 26878 6808 26884 6820
rect 26936 6808 26942 6860
rect 10321 6783 10379 6789
rect 10321 6780 10333 6783
rect 9548 6752 10333 6780
rect 9548 6740 9554 6752
rect 10321 6749 10333 6752
rect 10367 6749 10379 6783
rect 11790 6780 11796 6792
rect 11751 6752 11796 6780
rect 10321 6743 10379 6749
rect 11790 6740 11796 6752
rect 11848 6740 11854 6792
rect 19797 6783 19855 6789
rect 19797 6749 19809 6783
rect 19843 6780 19855 6783
rect 20530 6780 20536 6792
rect 19843 6752 20536 6780
rect 19843 6749 19855 6752
rect 19797 6743 19855 6749
rect 20530 6740 20536 6752
rect 20588 6740 20594 6792
rect 21729 6783 21787 6789
rect 21729 6749 21741 6783
rect 21775 6780 21787 6783
rect 22922 6780 22928 6792
rect 21775 6752 22928 6780
rect 21775 6749 21787 6752
rect 21729 6743 21787 6749
rect 22922 6740 22928 6752
rect 22980 6740 22986 6792
rect 23934 6780 23940 6792
rect 23895 6752 23940 6780
rect 23934 6740 23940 6752
rect 23992 6740 23998 6792
rect 5169 6715 5227 6721
rect 5169 6712 5181 6715
rect 4212 6684 5181 6712
rect 4212 6672 4218 6684
rect 5169 6681 5181 6684
rect 5215 6681 5227 6715
rect 5169 6675 5227 6681
rect 8205 6715 8263 6721
rect 8205 6681 8217 6715
rect 8251 6712 8263 6715
rect 21174 6712 21180 6724
rect 8251 6684 9444 6712
rect 21135 6684 21180 6712
rect 8251 6681 8263 6684
rect 8205 6675 8263 6681
rect 9416 6656 9444 6684
rect 21174 6672 21180 6684
rect 21232 6672 21238 6724
rect 27540 6721 27568 6888
rect 28258 6876 28264 6888
rect 28316 6876 28322 6928
rect 28442 6876 28448 6928
rect 28500 6916 28506 6928
rect 29178 6916 29184 6928
rect 28500 6888 29184 6916
rect 28500 6876 28506 6888
rect 29178 6876 29184 6888
rect 29236 6876 29242 6928
rect 33778 6876 33784 6928
rect 33836 6916 33842 6928
rect 34149 6919 34207 6925
rect 34149 6916 34161 6919
rect 33836 6888 34161 6916
rect 33836 6876 33842 6888
rect 34149 6885 34161 6888
rect 34195 6885 34207 6919
rect 34149 6879 34207 6885
rect 34330 6876 34336 6928
rect 34388 6916 34394 6928
rect 34388 6888 34433 6916
rect 34388 6876 34394 6888
rect 27614 6808 27620 6860
rect 27672 6848 27678 6860
rect 27965 6851 28023 6857
rect 27965 6848 27977 6851
rect 27672 6820 27977 6848
rect 27672 6808 27678 6820
rect 27965 6817 27977 6820
rect 28011 6817 28023 6851
rect 27965 6811 28023 6817
rect 32490 6808 32496 6860
rect 32548 6848 32554 6860
rect 32677 6851 32735 6857
rect 32677 6848 32689 6851
rect 32548 6820 32689 6848
rect 32548 6808 32554 6820
rect 32677 6817 32689 6820
rect 32723 6817 32735 6851
rect 32677 6811 32735 6817
rect 42610 6808 42616 6860
rect 42668 6848 42674 6860
rect 43605 6851 43663 6857
rect 43605 6848 43617 6851
rect 42668 6820 43617 6848
rect 42668 6808 42674 6820
rect 43605 6817 43617 6820
rect 43651 6848 43663 6851
rect 44174 6848 44180 6860
rect 43651 6820 44180 6848
rect 43651 6817 43663 6820
rect 43605 6811 43663 6817
rect 44174 6808 44180 6820
rect 44232 6808 44238 6860
rect 44726 6808 44732 6860
rect 44784 6848 44790 6860
rect 46106 6857 46112 6860
rect 46089 6851 46112 6857
rect 46089 6848 46101 6851
rect 44784 6820 46101 6848
rect 44784 6808 44790 6820
rect 46089 6817 46101 6820
rect 46164 6848 46170 6860
rect 46164 6820 46237 6848
rect 46089 6811 46112 6817
rect 46106 6808 46112 6811
rect 46164 6808 46170 6820
rect 27706 6780 27712 6792
rect 27667 6752 27712 6780
rect 27706 6740 27712 6752
rect 27764 6740 27770 6792
rect 34425 6783 34483 6789
rect 34425 6780 34437 6783
rect 33704 6752 34437 6780
rect 27525 6715 27583 6721
rect 27525 6712 27537 6715
rect 26252 6684 27537 6712
rect 26252 6656 26280 6684
rect 27525 6681 27537 6684
rect 27571 6681 27583 6715
rect 27525 6675 27583 6681
rect 33704 6656 33732 6752
rect 34425 6749 34437 6752
rect 34471 6749 34483 6783
rect 35345 6783 35403 6789
rect 35345 6780 35357 6783
rect 34425 6743 34483 6749
rect 35268 6752 35357 6780
rect 35268 6656 35296 6752
rect 35345 6749 35357 6752
rect 35391 6749 35403 6783
rect 37826 6780 37832 6792
rect 37787 6752 37832 6780
rect 35345 6743 35403 6749
rect 37826 6740 37832 6752
rect 37884 6740 37890 6792
rect 43346 6780 43352 6792
rect 43307 6752 43352 6780
rect 43346 6740 43352 6752
rect 43404 6740 43410 6792
rect 45830 6780 45836 6792
rect 45791 6752 45836 6780
rect 45830 6740 45836 6752
rect 45888 6740 45894 6792
rect 4706 6604 4712 6656
rect 4764 6644 4770 6656
rect 5537 6647 5595 6653
rect 5537 6644 5549 6647
rect 4764 6616 5549 6644
rect 4764 6604 4770 6616
rect 5537 6613 5549 6616
rect 5583 6644 5595 6647
rect 5626 6644 5632 6656
rect 5583 6616 5632 6644
rect 5583 6613 5595 6616
rect 5537 6607 5595 6613
rect 5626 6604 5632 6616
rect 5684 6604 5690 6656
rect 5718 6604 5724 6656
rect 5776 6644 5782 6656
rect 6178 6644 6184 6656
rect 5776 6616 6184 6644
rect 5776 6604 5782 6616
rect 6178 6604 6184 6616
rect 6236 6644 6242 6656
rect 7285 6647 7343 6653
rect 7285 6644 7297 6647
rect 6236 6616 7297 6644
rect 6236 6604 6242 6616
rect 7285 6613 7297 6616
rect 7331 6613 7343 6647
rect 7285 6607 7343 6613
rect 9398 6604 9404 6656
rect 9456 6644 9462 6656
rect 9769 6647 9827 6653
rect 9769 6644 9781 6647
rect 9456 6616 9781 6644
rect 9456 6604 9462 6616
rect 9769 6613 9781 6616
rect 9815 6613 9827 6647
rect 11330 6644 11336 6656
rect 11291 6616 11336 6644
rect 9769 6607 9827 6613
rect 11330 6604 11336 6616
rect 11388 6604 11394 6656
rect 13265 6647 13323 6653
rect 13265 6613 13277 6647
rect 13311 6644 13323 6647
rect 13354 6644 13360 6656
rect 13311 6616 13360 6644
rect 13311 6613 13323 6616
rect 13265 6607 13323 6613
rect 13354 6604 13360 6616
rect 13412 6604 13418 6656
rect 15473 6647 15531 6653
rect 15473 6613 15485 6647
rect 15519 6644 15531 6647
rect 15746 6644 15752 6656
rect 15519 6616 15752 6644
rect 15519 6613 15531 6616
rect 15473 6607 15531 6613
rect 15746 6604 15752 6616
rect 15804 6604 15810 6656
rect 15930 6604 15936 6656
rect 15988 6644 15994 6656
rect 16577 6647 16635 6653
rect 16577 6644 16589 6647
rect 15988 6616 16589 6644
rect 15988 6604 15994 6616
rect 16577 6613 16589 6616
rect 16623 6613 16635 6647
rect 23750 6644 23756 6656
rect 23711 6616 23756 6644
rect 16577 6607 16635 6613
rect 23750 6604 23756 6616
rect 23808 6604 23814 6656
rect 26234 6604 26240 6656
rect 26292 6644 26298 6656
rect 26292 6616 26337 6644
rect 26292 6604 26298 6616
rect 26510 6604 26516 6656
rect 26568 6644 26574 6656
rect 26697 6647 26755 6653
rect 26697 6644 26709 6647
rect 26568 6616 26709 6644
rect 26568 6604 26574 6616
rect 26697 6613 26709 6616
rect 26743 6613 26755 6647
rect 29086 6644 29092 6656
rect 29047 6616 29092 6644
rect 26697 6607 26755 6613
rect 29086 6604 29092 6616
rect 29144 6604 29150 6656
rect 30377 6647 30435 6653
rect 30377 6613 30389 6647
rect 30423 6644 30435 6647
rect 30558 6644 30564 6656
rect 30423 6616 30564 6644
rect 30423 6613 30435 6616
rect 30377 6607 30435 6613
rect 30558 6604 30564 6616
rect 30616 6604 30622 6656
rect 31202 6644 31208 6656
rect 31163 6616 31208 6644
rect 31202 6604 31208 6616
rect 31260 6604 31266 6656
rect 32490 6644 32496 6656
rect 32451 6616 32496 6644
rect 32490 6604 32496 6616
rect 32548 6604 32554 6656
rect 32861 6647 32919 6653
rect 32861 6613 32873 6647
rect 32907 6644 32919 6647
rect 33318 6644 33324 6656
rect 32907 6616 33324 6644
rect 32907 6613 32919 6616
rect 32861 6607 32919 6613
rect 33318 6604 33324 6616
rect 33376 6604 33382 6656
rect 33686 6644 33692 6656
rect 33647 6616 33692 6644
rect 33686 6604 33692 6616
rect 33744 6604 33750 6656
rect 33870 6644 33876 6656
rect 33831 6616 33876 6644
rect 33870 6604 33876 6616
rect 33928 6604 33934 6656
rect 35250 6644 35256 6656
rect 35211 6616 35256 6644
rect 35250 6604 35256 6616
rect 35308 6604 35314 6656
rect 44726 6644 44732 6656
rect 44687 6616 44732 6644
rect 44726 6604 44732 6616
rect 44784 6604 44790 6656
rect 45370 6644 45376 6656
rect 45283 6616 45376 6644
rect 45370 6604 45376 6616
rect 45428 6644 45434 6656
rect 47213 6647 47271 6653
rect 47213 6644 47225 6647
rect 45428 6616 47225 6644
rect 45428 6604 45434 6616
rect 47213 6613 47225 6616
rect 47259 6613 47271 6647
rect 47213 6607 47271 6613
rect 1104 6554 48852 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 34966 6554
rect 35018 6502 35030 6554
rect 35082 6502 35094 6554
rect 35146 6502 35158 6554
rect 35210 6502 48852 6554
rect 1104 6480 48852 6502
rect 3326 6440 3332 6452
rect 3160 6412 3332 6440
rect 3160 6313 3188 6412
rect 3326 6400 3332 6412
rect 3384 6400 3390 6452
rect 6270 6440 6276 6452
rect 6231 6412 6276 6440
rect 6270 6400 6276 6412
rect 6328 6400 6334 6452
rect 9306 6400 9312 6452
rect 9364 6440 9370 6452
rect 9493 6443 9551 6449
rect 9493 6440 9505 6443
rect 9364 6412 9505 6440
rect 9364 6400 9370 6412
rect 9493 6409 9505 6412
rect 9539 6409 9551 6443
rect 9493 6403 9551 6409
rect 8202 6372 8208 6384
rect 8163 6344 8208 6372
rect 8202 6332 8208 6344
rect 8260 6332 8266 6384
rect 3145 6307 3203 6313
rect 3145 6273 3157 6307
rect 3191 6273 3203 6307
rect 3145 6267 3203 6273
rect 8665 6307 8723 6313
rect 8665 6273 8677 6307
rect 8711 6304 8723 6307
rect 9398 6304 9404 6316
rect 8711 6276 9404 6304
rect 8711 6273 8723 6276
rect 8665 6267 8723 6273
rect 9398 6264 9404 6276
rect 9456 6264 9462 6316
rect 9508 6304 9536 6403
rect 10042 6400 10048 6452
rect 10100 6440 10106 6452
rect 11057 6443 11115 6449
rect 11057 6440 11069 6443
rect 10100 6412 11069 6440
rect 10100 6400 10106 6412
rect 11057 6409 11069 6412
rect 11103 6409 11115 6443
rect 11606 6440 11612 6452
rect 11567 6412 11612 6440
rect 11057 6403 11115 6409
rect 11606 6400 11612 6412
rect 11664 6400 11670 6452
rect 11790 6400 11796 6452
rect 11848 6440 11854 6452
rect 11977 6443 12035 6449
rect 11977 6440 11989 6443
rect 11848 6412 11989 6440
rect 11848 6400 11854 6412
rect 11977 6409 11989 6412
rect 12023 6409 12035 6443
rect 16390 6440 16396 6452
rect 16351 6412 16396 6440
rect 11977 6403 12035 6409
rect 16390 6400 16396 6412
rect 16448 6400 16454 6452
rect 17954 6400 17960 6452
rect 18012 6440 18018 6452
rect 18230 6440 18236 6452
rect 18012 6412 18236 6440
rect 18012 6400 18018 6412
rect 18230 6400 18236 6412
rect 18288 6440 18294 6452
rect 19521 6443 19579 6449
rect 19521 6440 19533 6443
rect 18288 6412 19533 6440
rect 18288 6400 18294 6412
rect 19521 6409 19533 6412
rect 19567 6409 19579 6443
rect 19521 6403 19579 6409
rect 21729 6443 21787 6449
rect 21729 6409 21741 6443
rect 21775 6440 21787 6443
rect 21910 6440 21916 6452
rect 21775 6412 21916 6440
rect 21775 6409 21787 6412
rect 21729 6403 21787 6409
rect 13081 6375 13139 6381
rect 13081 6341 13093 6375
rect 13127 6372 13139 6375
rect 13630 6372 13636 6384
rect 13127 6344 13636 6372
rect 13127 6341 13139 6344
rect 13081 6335 13139 6341
rect 13630 6332 13636 6344
rect 13688 6332 13694 6384
rect 15473 6375 15531 6381
rect 15473 6341 15485 6375
rect 15519 6372 15531 6375
rect 16482 6372 16488 6384
rect 15519 6344 16488 6372
rect 15519 6341 15531 6344
rect 15473 6335 15531 6341
rect 16482 6332 16488 6344
rect 16540 6332 16546 6384
rect 9677 6307 9735 6313
rect 9677 6304 9689 6307
rect 9508 6276 9689 6304
rect 9677 6273 9689 6276
rect 9723 6273 9735 6307
rect 9677 6267 9735 6273
rect 14553 6307 14611 6313
rect 14553 6273 14565 6307
rect 14599 6304 14611 6307
rect 15838 6304 15844 6316
rect 14599 6276 15844 6304
rect 14599 6273 14611 6276
rect 14553 6267 14611 6273
rect 15838 6264 15844 6276
rect 15896 6304 15902 6316
rect 16025 6307 16083 6313
rect 16025 6304 16037 6307
rect 15896 6276 16037 6304
rect 15896 6264 15902 6276
rect 16025 6273 16037 6276
rect 16071 6273 16083 6307
rect 19536 6304 19564 6403
rect 21910 6400 21916 6412
rect 21968 6400 21974 6452
rect 22465 6443 22523 6449
rect 22465 6409 22477 6443
rect 22511 6440 22523 6443
rect 22922 6440 22928 6452
rect 22511 6412 22928 6440
rect 22511 6409 22523 6412
rect 22465 6403 22523 6409
rect 22922 6400 22928 6412
rect 22980 6400 22986 6452
rect 23842 6440 23848 6452
rect 23676 6412 23848 6440
rect 23676 6313 23704 6412
rect 23842 6400 23848 6412
rect 23900 6400 23906 6452
rect 24854 6400 24860 6452
rect 24912 6440 24918 6452
rect 25041 6443 25099 6449
rect 25041 6440 25053 6443
rect 24912 6412 25053 6440
rect 24912 6400 24918 6412
rect 25041 6409 25053 6412
rect 25087 6409 25099 6443
rect 25041 6403 25099 6409
rect 25498 6400 25504 6452
rect 25556 6440 25562 6452
rect 25961 6443 26019 6449
rect 25961 6440 25973 6443
rect 25556 6412 25973 6440
rect 25556 6400 25562 6412
rect 25961 6409 25973 6412
rect 26007 6409 26019 6443
rect 25961 6403 26019 6409
rect 19705 6307 19763 6313
rect 19705 6304 19717 6307
rect 19536 6276 19717 6304
rect 16025 6267 16083 6273
rect 19705 6273 19717 6276
rect 19751 6273 19763 6307
rect 19705 6267 19763 6273
rect 23477 6307 23535 6313
rect 23477 6273 23489 6307
rect 23523 6304 23535 6307
rect 23661 6307 23719 6313
rect 23661 6304 23673 6307
rect 23523 6276 23673 6304
rect 23523 6273 23535 6276
rect 23477 6267 23535 6273
rect 23661 6273 23673 6276
rect 23707 6273 23719 6307
rect 23661 6267 23719 6273
rect 7653 6239 7711 6245
rect 7653 6205 7665 6239
rect 7699 6236 7711 6239
rect 7834 6236 7840 6248
rect 7699 6208 7840 6236
rect 7699 6205 7711 6208
rect 7653 6199 7711 6205
rect 7834 6196 7840 6208
rect 7892 6236 7898 6248
rect 8757 6239 8815 6245
rect 8757 6236 8769 6239
rect 7892 6208 8769 6236
rect 7892 6196 7898 6208
rect 8757 6205 8769 6208
rect 8803 6205 8815 6239
rect 9944 6239 10002 6245
rect 9944 6236 9956 6239
rect 8757 6199 8815 6205
rect 9784 6208 9956 6236
rect 2593 6171 2651 6177
rect 2593 6137 2605 6171
rect 2639 6168 2651 6171
rect 3390 6171 3448 6177
rect 3390 6168 3402 6171
rect 2639 6140 3402 6168
rect 2639 6137 2651 6140
rect 2593 6131 2651 6137
rect 3390 6137 3402 6140
rect 3436 6168 3448 6171
rect 4614 6168 4620 6180
rect 3436 6140 4620 6168
rect 3436 6137 3448 6140
rect 3390 6131 3448 6137
rect 4614 6128 4620 6140
rect 4672 6128 4678 6180
rect 8021 6171 8079 6177
rect 8021 6137 8033 6171
rect 8067 6168 8079 6171
rect 8662 6168 8668 6180
rect 8067 6140 8668 6168
rect 8067 6137 8079 6140
rect 8021 6131 8079 6137
rect 8662 6128 8668 6140
rect 8720 6128 8726 6180
rect 9217 6171 9275 6177
rect 9217 6137 9229 6171
rect 9263 6168 9275 6171
rect 9784 6168 9812 6208
rect 9944 6205 9956 6208
rect 9990 6236 10002 6239
rect 10226 6236 10232 6248
rect 9990 6208 10232 6236
rect 9990 6205 10002 6208
rect 9944 6199 10002 6205
rect 10226 6196 10232 6208
rect 10284 6196 10290 6248
rect 13354 6236 13360 6248
rect 13315 6208 13360 6236
rect 13354 6196 13360 6208
rect 13412 6196 13418 6248
rect 14921 6239 14979 6245
rect 14921 6205 14933 6239
rect 14967 6236 14979 6239
rect 15746 6236 15752 6248
rect 14967 6208 15752 6236
rect 14967 6205 14979 6208
rect 14921 6199 14979 6205
rect 15746 6196 15752 6208
rect 15804 6196 15810 6248
rect 23750 6196 23756 6248
rect 23808 6236 23814 6248
rect 23917 6239 23975 6245
rect 23917 6236 23929 6239
rect 23808 6208 23929 6236
rect 23808 6196 23814 6208
rect 23917 6205 23929 6208
rect 23963 6205 23975 6239
rect 23917 6199 23975 6205
rect 9263 6140 9812 6168
rect 9263 6137 9275 6140
rect 9217 6131 9275 6137
rect 13078 6128 13084 6180
rect 13136 6168 13142 6180
rect 13633 6171 13691 6177
rect 13633 6168 13645 6171
rect 13136 6140 13645 6168
rect 13136 6128 13142 6140
rect 13633 6137 13645 6140
rect 13679 6168 13691 6171
rect 15289 6171 15347 6177
rect 13679 6140 14136 6168
rect 13679 6137 13691 6140
rect 13633 6131 13691 6137
rect 14108 6112 14136 6140
rect 15289 6137 15301 6171
rect 15335 6168 15347 6171
rect 15930 6168 15936 6180
rect 15335 6140 15936 6168
rect 15335 6137 15347 6140
rect 15289 6131 15347 6137
rect 15930 6128 15936 6140
rect 15988 6128 15994 6180
rect 19978 6177 19984 6180
rect 19245 6171 19303 6177
rect 19245 6137 19257 6171
rect 19291 6168 19303 6171
rect 19972 6168 19984 6177
rect 19291 6140 19984 6168
rect 19291 6137 19303 6140
rect 19245 6131 19303 6137
rect 19972 6131 19984 6140
rect 19978 6128 19984 6131
rect 20036 6128 20042 6180
rect 21358 6128 21364 6180
rect 21416 6168 21422 6180
rect 22005 6171 22063 6177
rect 22005 6168 22017 6171
rect 21416 6140 22017 6168
rect 21416 6128 21422 6140
rect 22005 6137 22017 6140
rect 22051 6137 22063 6171
rect 25976 6168 26004 6403
rect 26418 6400 26424 6452
rect 26476 6440 26482 6452
rect 26602 6440 26608 6452
rect 26476 6412 26608 6440
rect 26476 6400 26482 6412
rect 26602 6400 26608 6412
rect 26660 6440 26666 6452
rect 27706 6440 27712 6452
rect 26660 6412 27712 6440
rect 26660 6400 26666 6412
rect 27706 6400 27712 6412
rect 27764 6400 27770 6452
rect 29089 6443 29147 6449
rect 29089 6409 29101 6443
rect 29135 6440 29147 6443
rect 29178 6440 29184 6452
rect 29135 6412 29184 6440
rect 29135 6409 29147 6412
rect 29089 6403 29147 6409
rect 29178 6400 29184 6412
rect 29236 6400 29242 6452
rect 31202 6400 31208 6452
rect 31260 6440 31266 6452
rect 31665 6443 31723 6449
rect 31665 6440 31677 6443
rect 31260 6412 31677 6440
rect 31260 6400 31266 6412
rect 31665 6409 31677 6412
rect 31711 6409 31723 6443
rect 31665 6403 31723 6409
rect 33778 6400 33784 6452
rect 33836 6440 33842 6452
rect 33965 6443 34023 6449
rect 33965 6440 33977 6443
rect 33836 6412 33977 6440
rect 33836 6400 33842 6412
rect 33965 6409 33977 6412
rect 34011 6409 34023 6443
rect 42610 6440 42616 6452
rect 42571 6412 42616 6440
rect 33965 6403 34023 6409
rect 42610 6400 42616 6412
rect 42668 6400 42674 6452
rect 43070 6400 43076 6452
rect 43128 6440 43134 6452
rect 43809 6443 43867 6449
rect 43809 6440 43821 6443
rect 43128 6412 43821 6440
rect 43128 6400 43134 6412
rect 43809 6409 43821 6412
rect 43855 6409 43867 6443
rect 43809 6403 43867 6409
rect 46106 6400 46112 6452
rect 46164 6440 46170 6452
rect 46293 6443 46351 6449
rect 46293 6440 46305 6443
rect 46164 6412 46305 6440
rect 46164 6400 46170 6412
rect 46293 6409 46305 6412
rect 46339 6409 46351 6443
rect 46293 6403 46351 6409
rect 26234 6332 26240 6384
rect 26292 6372 26298 6384
rect 33045 6375 33103 6381
rect 26292 6344 26337 6372
rect 26292 6332 26298 6344
rect 33045 6341 33057 6375
rect 33091 6372 33103 6375
rect 33134 6372 33140 6384
rect 33091 6344 33140 6372
rect 33091 6341 33103 6344
rect 33045 6335 33103 6341
rect 33134 6332 33140 6344
rect 33192 6332 33198 6384
rect 35253 6375 35311 6381
rect 35253 6341 35265 6375
rect 35299 6372 35311 6375
rect 35526 6372 35532 6384
rect 35299 6344 35532 6372
rect 35299 6341 35311 6344
rect 35253 6335 35311 6341
rect 35526 6332 35532 6344
rect 35584 6332 35590 6384
rect 37734 6372 37740 6384
rect 37695 6344 37740 6372
rect 37734 6332 37740 6344
rect 37792 6332 37798 6384
rect 43438 6372 43444 6384
rect 43399 6344 43444 6372
rect 43438 6332 43444 6344
rect 43496 6332 43502 6384
rect 32398 6304 32404 6316
rect 32359 6276 32404 6304
rect 32398 6264 32404 6276
rect 32456 6264 32462 6316
rect 33318 6264 33324 6316
rect 33376 6304 33382 6316
rect 33597 6307 33655 6313
rect 33597 6304 33609 6307
rect 33376 6276 33609 6304
rect 33376 6264 33382 6276
rect 33597 6273 33609 6276
rect 33643 6273 33655 6307
rect 33597 6267 33655 6273
rect 34701 6307 34759 6313
rect 34701 6273 34713 6307
rect 34747 6304 34759 6307
rect 35805 6307 35863 6313
rect 35805 6304 35817 6307
rect 34747 6276 35817 6304
rect 34747 6273 34759 6276
rect 34701 6267 34759 6273
rect 35805 6273 35817 6276
rect 35851 6304 35863 6307
rect 36262 6304 36268 6316
rect 35851 6276 36268 6304
rect 35851 6273 35863 6276
rect 35805 6267 35863 6273
rect 36262 6264 36268 6276
rect 36320 6264 36326 6316
rect 37553 6307 37611 6313
rect 37553 6273 37565 6307
rect 37599 6304 37611 6307
rect 43073 6307 43131 6313
rect 37599 6276 38332 6304
rect 37599 6273 37611 6276
rect 37553 6267 37611 6273
rect 26234 6196 26240 6248
rect 26292 6236 26298 6248
rect 26789 6239 26847 6245
rect 26789 6236 26801 6239
rect 26292 6208 26801 6236
rect 26292 6196 26298 6208
rect 26789 6205 26801 6208
rect 26835 6205 26847 6239
rect 26789 6199 26847 6205
rect 30285 6239 30343 6245
rect 30285 6205 30297 6239
rect 30331 6205 30343 6239
rect 30285 6199 30343 6205
rect 26510 6168 26516 6180
rect 25976 6140 26372 6168
rect 26471 6140 26516 6168
rect 22005 6131 22063 6137
rect 2961 6103 3019 6109
rect 2961 6069 2973 6103
rect 3007 6100 3019 6103
rect 3234 6100 3240 6112
rect 3007 6072 3240 6100
rect 3007 6069 3019 6072
rect 2961 6063 3019 6069
rect 3234 6060 3240 6072
rect 3292 6060 3298 6112
rect 4525 6103 4583 6109
rect 4525 6069 4537 6103
rect 4571 6100 4583 6103
rect 4798 6100 4804 6112
rect 4571 6072 4804 6100
rect 4571 6069 4583 6072
rect 4525 6063 4583 6069
rect 4798 6060 4804 6072
rect 4856 6060 4862 6112
rect 5902 6100 5908 6112
rect 5863 6072 5908 6100
rect 5902 6060 5908 6072
rect 5960 6100 5966 6112
rect 6730 6100 6736 6112
rect 5960 6072 6736 6100
rect 5960 6060 5966 6072
rect 6730 6060 6736 6072
rect 6788 6060 6794 6112
rect 12894 6100 12900 6112
rect 12807 6072 12900 6100
rect 12894 6060 12900 6072
rect 12952 6100 12958 6112
rect 13541 6103 13599 6109
rect 13541 6100 13553 6103
rect 12952 6072 13553 6100
rect 12952 6060 12958 6072
rect 13541 6069 13553 6072
rect 13587 6100 13599 6103
rect 13722 6100 13728 6112
rect 13587 6072 13728 6100
rect 13587 6069 13599 6072
rect 13541 6063 13599 6069
rect 13722 6060 13728 6072
rect 13780 6060 13786 6112
rect 14090 6100 14096 6112
rect 14051 6072 14096 6100
rect 14090 6060 14096 6072
rect 14148 6060 14154 6112
rect 18046 6100 18052 6112
rect 18007 6072 18052 6100
rect 18046 6060 18052 6072
rect 18104 6060 18110 6112
rect 21085 6103 21143 6109
rect 21085 6069 21097 6103
rect 21131 6100 21143 6103
rect 21542 6100 21548 6112
rect 21131 6072 21548 6100
rect 21131 6069 21143 6072
rect 21085 6063 21143 6069
rect 21542 6060 21548 6072
rect 21600 6060 21606 6112
rect 26344 6100 26372 6140
rect 26510 6128 26516 6140
rect 26568 6128 26574 6180
rect 27614 6128 27620 6180
rect 27672 6168 27678 6180
rect 28077 6171 28135 6177
rect 28077 6168 28089 6171
rect 27672 6140 28089 6168
rect 27672 6128 27678 6140
rect 28077 6137 28089 6140
rect 28123 6137 28135 6171
rect 28077 6131 28135 6137
rect 28994 6128 29000 6180
rect 29052 6168 29058 6180
rect 30101 6171 30159 6177
rect 30101 6168 30113 6171
rect 29052 6140 30113 6168
rect 29052 6128 29058 6140
rect 30101 6137 30113 6140
rect 30147 6168 30159 6171
rect 30300 6168 30328 6199
rect 30558 6177 30564 6180
rect 30552 6168 30564 6177
rect 30147 6140 30328 6168
rect 30519 6140 30564 6168
rect 30147 6137 30159 6140
rect 30101 6131 30159 6137
rect 30552 6131 30564 6140
rect 30558 6128 30564 6131
rect 30616 6128 30622 6180
rect 32416 6168 32444 6264
rect 32861 6239 32919 6245
rect 32861 6205 32873 6239
rect 32907 6236 32919 6239
rect 32907 6208 33548 6236
rect 32907 6205 32919 6208
rect 32861 6199 32919 6205
rect 33318 6168 33324 6180
rect 32416 6140 33324 6168
rect 33318 6128 33324 6140
rect 33376 6128 33382 6180
rect 33520 6177 33548 6208
rect 35250 6196 35256 6248
rect 35308 6236 35314 6248
rect 35529 6239 35587 6245
rect 35529 6236 35541 6239
rect 35308 6208 35541 6236
rect 35308 6196 35314 6208
rect 35529 6205 35541 6208
rect 35575 6205 35587 6239
rect 36173 6239 36231 6245
rect 36173 6236 36185 6239
rect 35529 6199 35587 6205
rect 35636 6208 36185 6236
rect 33505 6171 33563 6177
rect 33505 6137 33517 6171
rect 33551 6168 33563 6171
rect 33594 6168 33600 6180
rect 33551 6140 33600 6168
rect 33551 6137 33563 6140
rect 33505 6131 33563 6137
rect 33594 6128 33600 6140
rect 33652 6128 33658 6180
rect 26697 6103 26755 6109
rect 26697 6100 26709 6103
rect 26344 6072 26709 6100
rect 26697 6069 26709 6072
rect 26743 6069 26755 6103
rect 26697 6063 26755 6069
rect 26878 6060 26884 6112
rect 26936 6100 26942 6112
rect 27157 6103 27215 6109
rect 27157 6100 27169 6103
rect 26936 6072 27169 6100
rect 26936 6060 26942 6072
rect 27157 6069 27169 6072
rect 27203 6069 27215 6103
rect 29638 6100 29644 6112
rect 29551 6072 29644 6100
rect 27157 6063 27215 6069
rect 29638 6060 29644 6072
rect 29696 6100 29702 6112
rect 29914 6100 29920 6112
rect 29696 6072 29920 6100
rect 29696 6060 29702 6072
rect 29914 6060 29920 6072
rect 29972 6060 29978 6112
rect 33870 6060 33876 6112
rect 33928 6100 33934 6112
rect 35636 6100 35664 6208
rect 36173 6205 36185 6208
rect 36219 6205 36231 6239
rect 36173 6199 36231 6205
rect 37185 6239 37243 6245
rect 37185 6205 37197 6239
rect 37231 6236 37243 6239
rect 37826 6236 37832 6248
rect 37231 6208 37832 6236
rect 37231 6205 37243 6208
rect 37185 6199 37243 6205
rect 37826 6196 37832 6208
rect 37884 6236 37890 6248
rect 38013 6239 38071 6245
rect 38013 6236 38025 6239
rect 37884 6208 38025 6236
rect 37884 6196 37890 6208
rect 38013 6205 38025 6208
rect 38059 6205 38071 6239
rect 38013 6199 38071 6205
rect 38304 6180 38332 6276
rect 43073 6273 43085 6307
rect 43119 6304 43131 6307
rect 44269 6307 44327 6313
rect 44269 6304 44281 6307
rect 43119 6276 44281 6304
rect 43119 6273 43131 6276
rect 43073 6267 43131 6273
rect 44269 6273 44281 6276
rect 44315 6304 44327 6307
rect 45370 6304 45376 6316
rect 44315 6276 45376 6304
rect 44315 6273 44327 6276
rect 44269 6267 44327 6273
rect 45370 6264 45376 6276
rect 45428 6264 45434 6316
rect 39298 6236 39304 6248
rect 39259 6208 39304 6236
rect 39298 6196 39304 6208
rect 39356 6236 39362 6248
rect 39853 6239 39911 6245
rect 39853 6236 39865 6239
rect 39356 6208 39865 6236
rect 39356 6196 39362 6208
rect 39853 6205 39865 6208
rect 39899 6205 39911 6239
rect 44358 6236 44364 6248
rect 44319 6208 44364 6236
rect 39853 6199 39911 6205
rect 44358 6196 44364 6208
rect 44416 6196 44422 6248
rect 36817 6171 36875 6177
rect 36817 6137 36829 6171
rect 36863 6168 36875 6171
rect 38197 6171 38255 6177
rect 38197 6168 38209 6171
rect 36863 6140 38209 6168
rect 36863 6137 36875 6140
rect 36817 6131 36875 6137
rect 38197 6137 38209 6140
rect 38243 6137 38255 6171
rect 38197 6131 38255 6137
rect 35713 6103 35771 6109
rect 35713 6100 35725 6103
rect 33928 6072 35725 6100
rect 33928 6060 33934 6072
rect 35713 6069 35725 6072
rect 35759 6069 35771 6103
rect 38212 6100 38240 6131
rect 38286 6128 38292 6180
rect 38344 6168 38350 6180
rect 38344 6140 38389 6168
rect 38344 6128 38350 6140
rect 38654 6100 38660 6112
rect 38212 6072 38660 6100
rect 35713 6063 35771 6069
rect 38654 6060 38660 6072
rect 38712 6060 38718 6112
rect 39485 6103 39543 6109
rect 39485 6069 39497 6103
rect 39531 6100 39543 6103
rect 39850 6100 39856 6112
rect 39531 6072 39856 6100
rect 39531 6069 39543 6072
rect 39485 6063 39543 6069
rect 39850 6060 39856 6072
rect 39908 6060 39914 6112
rect 43806 6060 43812 6112
rect 43864 6100 43870 6112
rect 44269 6103 44327 6109
rect 44269 6100 44281 6103
rect 43864 6072 44281 6100
rect 43864 6060 43870 6072
rect 44269 6069 44281 6072
rect 44315 6100 44327 6103
rect 44726 6100 44732 6112
rect 44315 6072 44732 6100
rect 44315 6069 44327 6072
rect 44269 6063 44327 6069
rect 44726 6060 44732 6072
rect 44784 6060 44790 6112
rect 45922 6100 45928 6112
rect 45883 6072 45928 6100
rect 45922 6060 45928 6072
rect 45980 6060 45986 6112
rect 1104 6010 48852 6032
rect 1104 5958 19606 6010
rect 19658 5958 19670 6010
rect 19722 5958 19734 6010
rect 19786 5958 19798 6010
rect 19850 5958 48852 6010
rect 1104 5936 48852 5958
rect 3237 5899 3295 5905
rect 3237 5865 3249 5899
rect 3283 5896 3295 5899
rect 3326 5896 3332 5908
rect 3283 5868 3332 5896
rect 3283 5865 3295 5868
rect 3237 5859 3295 5865
rect 3326 5856 3332 5868
rect 3384 5856 3390 5908
rect 4614 5896 4620 5908
rect 4575 5868 4620 5896
rect 4614 5856 4620 5868
rect 4672 5856 4678 5908
rect 6914 5856 6920 5908
rect 6972 5896 6978 5908
rect 7285 5899 7343 5905
rect 7285 5896 7297 5899
rect 6972 5868 7297 5896
rect 6972 5856 6978 5868
rect 7285 5865 7297 5868
rect 7331 5865 7343 5899
rect 7285 5859 7343 5865
rect 9953 5899 10011 5905
rect 9953 5865 9965 5899
rect 9999 5896 10011 5899
rect 10226 5896 10232 5908
rect 9999 5868 10232 5896
rect 9999 5865 10011 5868
rect 9953 5859 10011 5865
rect 10226 5856 10232 5868
rect 10284 5856 10290 5908
rect 11974 5896 11980 5908
rect 11935 5868 11980 5896
rect 11974 5856 11980 5868
rect 12032 5856 12038 5908
rect 13354 5856 13360 5908
rect 13412 5896 13418 5908
rect 13909 5899 13967 5905
rect 13909 5896 13921 5899
rect 13412 5868 13921 5896
rect 13412 5856 13418 5868
rect 13909 5865 13921 5868
rect 13955 5896 13967 5899
rect 13998 5896 14004 5908
rect 13955 5868 14004 5896
rect 13955 5865 13967 5868
rect 13909 5859 13967 5865
rect 13998 5856 14004 5868
rect 14056 5896 14062 5908
rect 14461 5899 14519 5905
rect 14461 5896 14473 5899
rect 14056 5868 14473 5896
rect 14056 5856 14062 5868
rect 14461 5865 14473 5868
rect 14507 5865 14519 5899
rect 15470 5896 15476 5908
rect 15431 5868 15476 5896
rect 14461 5859 14519 5865
rect 15470 5856 15476 5868
rect 15528 5856 15534 5908
rect 22094 5856 22100 5908
rect 22152 5896 22158 5908
rect 23019 5899 23077 5905
rect 23019 5896 23031 5899
rect 22152 5868 23031 5896
rect 22152 5856 22158 5868
rect 23019 5865 23031 5868
rect 23065 5896 23077 5899
rect 23106 5896 23112 5908
rect 23065 5868 23112 5896
rect 23065 5865 23077 5868
rect 23019 5859 23077 5865
rect 23106 5856 23112 5868
rect 23164 5856 23170 5908
rect 26237 5899 26295 5905
rect 26237 5865 26249 5899
rect 26283 5896 26295 5899
rect 26510 5896 26516 5908
rect 26283 5868 26516 5896
rect 26283 5865 26295 5868
rect 26237 5859 26295 5865
rect 26510 5856 26516 5868
rect 26568 5856 26574 5908
rect 33686 5856 33692 5908
rect 33744 5896 33750 5908
rect 33781 5899 33839 5905
rect 33781 5896 33793 5899
rect 33744 5868 33793 5896
rect 33744 5856 33750 5868
rect 33781 5865 33793 5868
rect 33827 5865 33839 5899
rect 36262 5896 36268 5908
rect 36223 5868 36268 5896
rect 33781 5859 33839 5865
rect 6178 5837 6184 5840
rect 6172 5828 6184 5837
rect 6139 5800 6184 5828
rect 6172 5791 6184 5800
rect 6178 5788 6184 5791
rect 6236 5788 6242 5840
rect 11514 5828 11520 5840
rect 11475 5800 11520 5828
rect 11514 5788 11520 5800
rect 11572 5788 11578 5840
rect 12796 5831 12854 5837
rect 12796 5797 12808 5831
rect 12842 5828 12854 5831
rect 12894 5828 12900 5840
rect 12842 5800 12900 5828
rect 12842 5797 12854 5800
rect 12796 5791 12854 5797
rect 12894 5788 12900 5800
rect 12952 5788 12958 5840
rect 16016 5831 16074 5837
rect 16016 5797 16028 5831
rect 16062 5828 16074 5831
rect 16114 5828 16120 5840
rect 16062 5800 16120 5828
rect 16062 5797 16074 5800
rect 16016 5791 16074 5797
rect 16114 5788 16120 5800
rect 16172 5788 16178 5840
rect 18230 5828 18236 5840
rect 17972 5800 18236 5828
rect 8202 5720 8208 5772
rect 8260 5760 8266 5772
rect 8389 5763 8447 5769
rect 8389 5760 8401 5763
rect 8260 5732 8401 5760
rect 8260 5720 8266 5732
rect 8389 5729 8401 5732
rect 8435 5760 8447 5763
rect 9214 5760 9220 5772
rect 8435 5732 9220 5760
rect 8435 5729 8447 5732
rect 8389 5723 8447 5729
rect 9214 5720 9220 5732
rect 9272 5720 9278 5772
rect 10042 5720 10048 5772
rect 10100 5760 10106 5772
rect 10229 5763 10287 5769
rect 10229 5760 10241 5763
rect 10100 5732 10241 5760
rect 10100 5720 10106 5732
rect 10229 5729 10241 5732
rect 10275 5729 10287 5763
rect 11330 5760 11336 5772
rect 11291 5732 11336 5760
rect 10229 5723 10287 5729
rect 11330 5720 11336 5732
rect 11388 5720 11394 5772
rect 12434 5720 12440 5772
rect 12492 5760 12498 5772
rect 12529 5763 12587 5769
rect 12529 5760 12541 5763
rect 12492 5732 12541 5760
rect 12492 5720 12498 5732
rect 12529 5729 12541 5732
rect 12575 5729 12587 5763
rect 15746 5760 15752 5772
rect 15659 5732 15752 5760
rect 12529 5723 12587 5729
rect 15746 5720 15752 5732
rect 15804 5760 15810 5772
rect 17678 5760 17684 5772
rect 15804 5732 17684 5760
rect 15804 5720 15810 5732
rect 17678 5720 17684 5732
rect 17736 5760 17742 5772
rect 17972 5760 18000 5800
rect 18230 5788 18236 5800
rect 18288 5788 18294 5840
rect 20717 5831 20775 5837
rect 20717 5797 20729 5831
rect 20763 5828 20775 5831
rect 20898 5828 20904 5840
rect 20763 5800 20904 5828
rect 20763 5797 20775 5800
rect 20717 5791 20775 5797
rect 20898 5788 20904 5800
rect 20956 5828 20962 5840
rect 21453 5831 21511 5837
rect 21453 5828 21465 5831
rect 20956 5800 21465 5828
rect 20956 5788 20962 5800
rect 21453 5797 21465 5800
rect 21499 5797 21511 5831
rect 21453 5791 21511 5797
rect 21542 5788 21548 5840
rect 21600 5828 21606 5840
rect 21600 5800 21645 5828
rect 21600 5788 21606 5800
rect 26602 5788 26608 5840
rect 26660 5828 26666 5840
rect 26780 5831 26838 5837
rect 26780 5828 26792 5831
rect 26660 5800 26792 5828
rect 26660 5788 26666 5800
rect 26780 5797 26792 5800
rect 26826 5828 26838 5831
rect 27062 5828 27068 5840
rect 26826 5800 27068 5828
rect 26826 5797 26838 5800
rect 26780 5791 26838 5797
rect 27062 5788 27068 5800
rect 27120 5828 27126 5840
rect 27522 5828 27528 5840
rect 27120 5800 27528 5828
rect 27120 5788 27126 5800
rect 27522 5788 27528 5800
rect 27580 5788 27586 5840
rect 29086 5788 29092 5840
rect 29144 5828 29150 5840
rect 29426 5831 29484 5837
rect 29426 5828 29438 5831
rect 29144 5800 29438 5828
rect 29144 5788 29150 5800
rect 29426 5797 29438 5800
rect 29472 5797 29484 5831
rect 29426 5791 29484 5797
rect 18506 5769 18512 5772
rect 18489 5763 18512 5769
rect 18489 5760 18501 5763
rect 17736 5732 18000 5760
rect 18064 5732 18501 5760
rect 17736 5720 17742 5732
rect 4617 5695 4675 5701
rect 4617 5661 4629 5695
rect 4663 5661 4675 5695
rect 4617 5655 4675 5661
rect 4632 5624 4660 5655
rect 4706 5652 4712 5704
rect 4764 5692 4770 5704
rect 5902 5692 5908 5704
rect 4764 5664 4809 5692
rect 5815 5664 5908 5692
rect 4764 5652 4770 5664
rect 5902 5652 5908 5664
rect 5960 5652 5966 5704
rect 11606 5692 11612 5704
rect 11567 5664 11612 5692
rect 11606 5652 11612 5664
rect 11664 5652 11670 5704
rect 4798 5624 4804 5636
rect 4632 5596 4804 5624
rect 4798 5584 4804 5596
rect 4856 5584 4862 5636
rect 4157 5559 4215 5565
rect 4157 5525 4169 5559
rect 4203 5556 4215 5559
rect 5718 5556 5724 5568
rect 4203 5528 5724 5556
rect 4203 5525 4215 5528
rect 4157 5519 4215 5525
rect 5718 5516 5724 5528
rect 5776 5516 5782 5568
rect 5920 5556 5948 5652
rect 11054 5624 11060 5636
rect 11015 5596 11060 5624
rect 11054 5584 11060 5596
rect 11112 5584 11118 5636
rect 6270 5556 6276 5568
rect 5920 5528 6276 5556
rect 6270 5516 6276 5528
rect 6328 5516 6334 5568
rect 8294 5556 8300 5568
rect 8255 5528 8300 5556
rect 8294 5516 8300 5528
rect 8352 5516 8358 5568
rect 8573 5559 8631 5565
rect 8573 5525 8585 5559
rect 8619 5556 8631 5559
rect 8754 5556 8760 5568
rect 8619 5528 8760 5556
rect 8619 5525 8631 5528
rect 8573 5519 8631 5525
rect 8754 5516 8760 5528
rect 8812 5516 8818 5568
rect 8846 5516 8852 5568
rect 8904 5556 8910 5568
rect 8941 5559 8999 5565
rect 8941 5556 8953 5559
rect 8904 5528 8953 5556
rect 8904 5516 8910 5528
rect 8941 5525 8953 5528
rect 8987 5525 8999 5559
rect 9490 5556 9496 5568
rect 9451 5528 9496 5556
rect 8941 5519 8999 5525
rect 9490 5516 9496 5528
rect 9548 5516 9554 5568
rect 18064 5565 18092 5732
rect 18489 5729 18501 5732
rect 18564 5760 18570 5772
rect 18564 5732 18637 5760
rect 18489 5723 18512 5729
rect 18506 5720 18512 5723
rect 18564 5720 18570 5732
rect 20530 5720 20536 5772
rect 20588 5760 20594 5772
rect 21269 5763 21327 5769
rect 21269 5760 21281 5763
rect 20588 5732 21281 5760
rect 20588 5720 20594 5732
rect 21269 5729 21281 5732
rect 21315 5729 21327 5763
rect 21269 5723 21327 5729
rect 22094 5720 22100 5772
rect 22152 5760 22158 5772
rect 22465 5763 22523 5769
rect 22465 5760 22477 5763
rect 22152 5732 22477 5760
rect 22152 5720 22158 5732
rect 22465 5729 22477 5732
rect 22511 5760 22523 5763
rect 23290 5760 23296 5772
rect 22511 5732 23296 5760
rect 22511 5729 22523 5732
rect 22465 5723 22523 5729
rect 23290 5720 23296 5732
rect 23348 5720 23354 5772
rect 26418 5720 26424 5772
rect 26476 5760 26482 5772
rect 26513 5763 26571 5769
rect 26513 5760 26525 5763
rect 26476 5732 26525 5760
rect 26476 5720 26482 5732
rect 26513 5729 26525 5732
rect 26559 5760 26571 5763
rect 27154 5760 27160 5772
rect 26559 5732 27160 5760
rect 26559 5729 26571 5732
rect 26513 5723 26571 5729
rect 27154 5720 27160 5732
rect 27212 5760 27218 5772
rect 28994 5760 29000 5772
rect 27212 5732 29000 5760
rect 27212 5720 27218 5732
rect 28994 5720 29000 5732
rect 29052 5760 29058 5772
rect 29181 5763 29239 5769
rect 29181 5760 29193 5763
rect 29052 5732 29193 5760
rect 29052 5720 29058 5732
rect 29181 5729 29193 5732
rect 29227 5729 29239 5763
rect 29181 5723 29239 5729
rect 32306 5720 32312 5772
rect 32364 5760 32370 5772
rect 32657 5763 32715 5769
rect 32657 5760 32669 5763
rect 32364 5732 32669 5760
rect 32364 5720 32370 5732
rect 32657 5729 32669 5732
rect 32703 5729 32715 5763
rect 33796 5760 33824 5859
rect 36262 5856 36268 5868
rect 36320 5856 36326 5908
rect 38194 5856 38200 5908
rect 38252 5896 38258 5908
rect 42058 5896 42064 5908
rect 38252 5868 38297 5896
rect 42019 5868 42064 5896
rect 38252 5856 38258 5868
rect 42058 5856 42064 5868
rect 42116 5856 42122 5908
rect 43806 5896 43812 5908
rect 43767 5868 43812 5896
rect 43806 5856 43812 5868
rect 43864 5856 43870 5908
rect 44177 5899 44235 5905
rect 44177 5865 44189 5899
rect 44223 5896 44235 5899
rect 44358 5896 44364 5908
rect 44223 5868 44364 5896
rect 44223 5865 44235 5868
rect 44177 5859 44235 5865
rect 44358 5856 44364 5868
rect 44416 5856 44422 5908
rect 37734 5788 37740 5840
rect 37792 5788 37798 5840
rect 35152 5763 35210 5769
rect 35152 5760 35164 5763
rect 33796 5732 35164 5760
rect 32657 5723 32715 5729
rect 35152 5729 35164 5732
rect 35198 5760 35210 5763
rect 35434 5760 35440 5772
rect 35198 5732 35440 5760
rect 35198 5729 35210 5732
rect 35152 5723 35210 5729
rect 35434 5720 35440 5732
rect 35492 5720 35498 5772
rect 37553 5763 37611 5769
rect 37553 5729 37565 5763
rect 37599 5760 37611 5763
rect 37752 5760 37780 5788
rect 40678 5760 40684 5772
rect 37599 5732 38240 5760
rect 40639 5732 40684 5760
rect 37599 5729 37611 5732
rect 37553 5723 37611 5729
rect 18230 5692 18236 5704
rect 18191 5664 18236 5692
rect 18230 5652 18236 5664
rect 18288 5652 18294 5704
rect 22554 5692 22560 5704
rect 22112 5664 22560 5692
rect 20990 5624 20996 5636
rect 20951 5596 20996 5624
rect 20990 5584 20996 5596
rect 21048 5584 21054 5636
rect 22112 5633 22140 5664
rect 22554 5652 22560 5664
rect 22612 5652 22618 5704
rect 23014 5692 23020 5704
rect 22975 5664 23020 5692
rect 23014 5652 23020 5664
rect 23072 5652 23078 5704
rect 31846 5652 31852 5704
rect 31904 5692 31910 5704
rect 32401 5695 32459 5701
rect 32401 5692 32413 5695
rect 31904 5664 32413 5692
rect 31904 5652 31910 5664
rect 32401 5661 32413 5664
rect 32447 5661 32459 5695
rect 32401 5655 32459 5661
rect 22097 5627 22155 5633
rect 22097 5593 22109 5627
rect 22143 5593 22155 5627
rect 22097 5587 22155 5593
rect 17129 5559 17187 5565
rect 17129 5525 17141 5559
rect 17175 5556 17187 5559
rect 18049 5559 18107 5565
rect 18049 5556 18061 5559
rect 17175 5528 18061 5556
rect 17175 5525 17187 5528
rect 17129 5519 17187 5525
rect 18049 5525 18061 5528
rect 18095 5525 18107 5559
rect 18049 5519 18107 5525
rect 19613 5559 19671 5565
rect 19613 5525 19625 5559
rect 19659 5556 19671 5559
rect 19978 5556 19984 5568
rect 19659 5528 19984 5556
rect 19659 5525 19671 5528
rect 19613 5519 19671 5525
rect 19978 5516 19984 5528
rect 20036 5556 20042 5568
rect 20622 5556 20628 5568
rect 20036 5528 20628 5556
rect 20036 5516 20042 5528
rect 20622 5516 20628 5528
rect 20680 5516 20686 5568
rect 24026 5516 24032 5568
rect 24084 5556 24090 5568
rect 24397 5559 24455 5565
rect 24397 5556 24409 5559
rect 24084 5528 24409 5556
rect 24084 5516 24090 5528
rect 24397 5525 24409 5528
rect 24443 5525 24455 5559
rect 24397 5519 24455 5525
rect 27614 5516 27620 5568
rect 27672 5556 27678 5568
rect 27893 5559 27951 5565
rect 27893 5556 27905 5559
rect 27672 5528 27905 5556
rect 27672 5516 27678 5528
rect 27893 5525 27905 5528
rect 27939 5525 27951 5559
rect 27893 5519 27951 5525
rect 30561 5559 30619 5565
rect 30561 5525 30573 5559
rect 30607 5556 30619 5559
rect 30742 5556 30748 5568
rect 30607 5528 30748 5556
rect 30607 5525 30619 5528
rect 30561 5519 30619 5525
rect 30742 5516 30748 5528
rect 30800 5516 30806 5568
rect 32416 5556 32444 5655
rect 34606 5652 34612 5704
rect 34664 5692 34670 5704
rect 34885 5695 34943 5701
rect 34885 5692 34897 5695
rect 34664 5664 34897 5692
rect 34664 5652 34670 5664
rect 34885 5661 34897 5664
rect 34931 5661 34943 5695
rect 34885 5655 34943 5661
rect 36538 5652 36544 5704
rect 36596 5692 36602 5704
rect 37090 5692 37096 5704
rect 36596 5664 37096 5692
rect 36596 5652 36602 5664
rect 37090 5652 37096 5664
rect 37148 5692 37154 5704
rect 38212 5701 38240 5732
rect 40678 5720 40684 5732
rect 40736 5720 40742 5772
rect 40954 5769 40960 5772
rect 40948 5760 40960 5769
rect 40915 5732 40960 5760
rect 40948 5723 40960 5732
rect 40954 5720 40960 5723
rect 41012 5720 41018 5772
rect 37737 5695 37795 5701
rect 37737 5692 37749 5695
rect 37148 5664 37749 5692
rect 37148 5652 37154 5664
rect 37737 5661 37749 5664
rect 37783 5661 37795 5695
rect 37737 5655 37795 5661
rect 38197 5695 38255 5701
rect 38197 5661 38209 5695
rect 38243 5661 38255 5695
rect 38470 5692 38476 5704
rect 38431 5664 38476 5692
rect 38197 5655 38255 5661
rect 38470 5652 38476 5664
rect 38528 5652 38534 5704
rect 33042 5556 33048 5568
rect 32416 5528 33048 5556
rect 33042 5516 33048 5528
rect 33100 5516 33106 5568
rect 33594 5516 33600 5568
rect 33652 5556 33658 5568
rect 34330 5556 34336 5568
rect 33652 5528 34336 5556
rect 33652 5516 33658 5528
rect 34330 5516 34336 5528
rect 34388 5516 34394 5568
rect 39577 5559 39635 5565
rect 39577 5525 39589 5559
rect 39623 5556 39635 5559
rect 39942 5556 39948 5568
rect 39623 5528 39948 5556
rect 39623 5525 39635 5528
rect 39577 5519 39635 5525
rect 39942 5516 39948 5528
rect 40000 5516 40006 5568
rect 40589 5559 40647 5565
rect 40589 5525 40601 5559
rect 40635 5556 40647 5559
rect 40678 5556 40684 5568
rect 40635 5528 40684 5556
rect 40635 5525 40647 5528
rect 40589 5519 40647 5525
rect 40678 5516 40684 5528
rect 40736 5516 40742 5568
rect 1104 5466 48852 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 34966 5466
rect 35018 5414 35030 5466
rect 35082 5414 35094 5466
rect 35146 5414 35158 5466
rect 35210 5414 48852 5466
rect 1104 5392 48852 5414
rect 3053 5355 3111 5361
rect 3053 5321 3065 5355
rect 3099 5352 3111 5355
rect 3326 5352 3332 5364
rect 3099 5324 3332 5352
rect 3099 5321 3111 5324
rect 3053 5315 3111 5321
rect 3160 5225 3188 5324
rect 3326 5312 3332 5324
rect 3384 5312 3390 5364
rect 4525 5355 4583 5361
rect 4525 5321 4537 5355
rect 4571 5352 4583 5355
rect 4614 5352 4620 5364
rect 4571 5324 4620 5352
rect 4571 5321 4583 5324
rect 4525 5315 4583 5321
rect 4614 5312 4620 5324
rect 4672 5312 4678 5364
rect 6178 5312 6184 5364
rect 6236 5352 6242 5364
rect 6549 5355 6607 5361
rect 6549 5352 6561 5355
rect 6236 5324 6561 5352
rect 6236 5312 6242 5324
rect 6549 5321 6561 5324
rect 6595 5321 6607 5355
rect 6549 5315 6607 5321
rect 7009 5355 7067 5361
rect 7009 5321 7021 5355
rect 7055 5352 7067 5355
rect 8202 5352 8208 5364
rect 7055 5324 8208 5352
rect 7055 5321 7067 5324
rect 7009 5315 7067 5321
rect 8202 5312 8208 5324
rect 8260 5312 8266 5364
rect 9214 5352 9220 5364
rect 9175 5324 9220 5352
rect 9214 5312 9220 5324
rect 9272 5312 9278 5364
rect 11057 5355 11115 5361
rect 11057 5321 11069 5355
rect 11103 5352 11115 5355
rect 11330 5352 11336 5364
rect 11103 5324 11336 5352
rect 11103 5321 11115 5324
rect 11057 5315 11115 5321
rect 11330 5312 11336 5324
rect 11388 5312 11394 5364
rect 11425 5355 11483 5361
rect 11425 5321 11437 5355
rect 11471 5352 11483 5355
rect 11514 5352 11520 5364
rect 11471 5324 11520 5352
rect 11471 5321 11483 5324
rect 11425 5315 11483 5321
rect 11514 5312 11520 5324
rect 11572 5352 11578 5364
rect 11793 5355 11851 5361
rect 11793 5352 11805 5355
rect 11572 5324 11805 5352
rect 11572 5312 11578 5324
rect 11793 5321 11805 5324
rect 11839 5321 11851 5355
rect 11793 5315 11851 5321
rect 12434 5312 12440 5364
rect 12492 5352 12498 5364
rect 12989 5355 13047 5361
rect 12989 5352 13001 5355
rect 12492 5324 13001 5352
rect 12492 5312 12498 5324
rect 12989 5321 13001 5324
rect 13035 5352 13047 5355
rect 13541 5355 13599 5361
rect 13541 5352 13553 5355
rect 13035 5324 13553 5352
rect 13035 5321 13047 5324
rect 12989 5315 13047 5321
rect 13541 5321 13553 5324
rect 13587 5321 13599 5355
rect 15746 5352 15752 5364
rect 15707 5324 15752 5352
rect 13541 5315 13599 5321
rect 3145 5219 3203 5225
rect 3145 5185 3157 5219
rect 3191 5185 3203 5219
rect 8220 5216 8248 5312
rect 8297 5287 8355 5293
rect 8297 5253 8309 5287
rect 8343 5284 8355 5287
rect 9582 5284 9588 5296
rect 8343 5256 9588 5284
rect 8343 5253 8355 5256
rect 8297 5247 8355 5253
rect 9582 5244 9588 5256
rect 9640 5244 9646 5296
rect 11348 5284 11376 5312
rect 12621 5287 12679 5293
rect 12621 5284 12633 5287
rect 11348 5256 12633 5284
rect 12621 5253 12633 5256
rect 12667 5253 12679 5287
rect 12621 5247 12679 5253
rect 13556 5228 13584 5315
rect 15746 5312 15752 5324
rect 15804 5312 15810 5364
rect 17402 5352 17408 5364
rect 17363 5324 17408 5352
rect 17402 5312 17408 5324
rect 17460 5312 17466 5364
rect 17865 5355 17923 5361
rect 17865 5321 17877 5355
rect 17911 5352 17923 5355
rect 18046 5352 18052 5364
rect 17911 5324 18052 5352
rect 17911 5321 17923 5324
rect 17865 5315 17923 5321
rect 18046 5312 18052 5324
rect 18104 5312 18110 5364
rect 18230 5312 18236 5364
rect 18288 5352 18294 5364
rect 19061 5355 19119 5361
rect 19061 5352 19073 5355
rect 18288 5324 19073 5352
rect 18288 5312 18294 5324
rect 19061 5321 19073 5324
rect 19107 5352 19119 5355
rect 20530 5352 20536 5364
rect 19107 5324 20208 5352
rect 20491 5324 20536 5352
rect 19107 5321 19119 5324
rect 19061 5315 19119 5321
rect 8665 5219 8723 5225
rect 8665 5216 8677 5219
rect 8220 5188 8677 5216
rect 3145 5179 3203 5185
rect 8665 5185 8677 5188
rect 8711 5185 8723 5219
rect 13538 5216 13544 5228
rect 13451 5188 13544 5216
rect 8665 5179 8723 5185
rect 13538 5176 13544 5188
rect 13596 5216 13602 5228
rect 13725 5219 13783 5225
rect 13725 5216 13737 5219
rect 13596 5188 13737 5216
rect 13596 5176 13602 5188
rect 13725 5185 13737 5188
rect 13771 5185 13783 5219
rect 18064 5216 18092 5312
rect 18141 5287 18199 5293
rect 18141 5253 18153 5287
rect 18187 5284 18199 5287
rect 19426 5284 19432 5296
rect 18187 5256 19432 5284
rect 18187 5253 18199 5256
rect 18141 5247 18199 5253
rect 19426 5244 19432 5256
rect 19484 5244 19490 5296
rect 20180 5284 20208 5324
rect 20530 5312 20536 5324
rect 20588 5312 20594 5364
rect 23106 5352 23112 5364
rect 23067 5324 23112 5352
rect 23106 5312 23112 5324
rect 23164 5312 23170 5364
rect 23474 5352 23480 5364
rect 23435 5324 23480 5352
rect 23474 5312 23480 5324
rect 23532 5312 23538 5364
rect 23750 5352 23756 5364
rect 23711 5324 23756 5352
rect 23750 5312 23756 5324
rect 23808 5312 23814 5364
rect 26237 5355 26295 5361
rect 26237 5321 26249 5355
rect 26283 5352 26295 5355
rect 26878 5352 26884 5364
rect 26283 5324 26884 5352
rect 26283 5321 26295 5324
rect 26237 5315 26295 5321
rect 26878 5312 26884 5324
rect 26936 5312 26942 5364
rect 27154 5352 27160 5364
rect 27115 5324 27160 5352
rect 27154 5312 27160 5324
rect 27212 5312 27218 5364
rect 27341 5355 27399 5361
rect 27341 5321 27353 5355
rect 27387 5352 27399 5355
rect 27617 5355 27675 5361
rect 27617 5352 27629 5355
rect 27387 5324 27629 5352
rect 27387 5321 27399 5324
rect 27341 5315 27399 5321
rect 27617 5321 27629 5324
rect 27663 5352 27675 5355
rect 28442 5352 28448 5364
rect 27663 5324 28448 5352
rect 27663 5321 27675 5324
rect 27617 5315 27675 5321
rect 28442 5312 28448 5324
rect 28500 5312 28506 5364
rect 28721 5355 28779 5361
rect 28721 5321 28733 5355
rect 28767 5352 28779 5355
rect 29086 5352 29092 5364
rect 28767 5324 29092 5352
rect 28767 5321 28779 5324
rect 28721 5315 28779 5321
rect 29086 5312 29092 5324
rect 29144 5312 29150 5364
rect 33042 5312 33048 5364
rect 33100 5352 33106 5364
rect 33229 5355 33287 5361
rect 33229 5352 33241 5355
rect 33100 5324 33241 5352
rect 33100 5312 33106 5324
rect 33229 5321 33241 5324
rect 33275 5352 33287 5355
rect 34606 5352 34612 5364
rect 33275 5324 34612 5352
rect 33275 5321 33287 5324
rect 33229 5315 33287 5321
rect 34606 5312 34612 5324
rect 34664 5352 34670 5364
rect 35069 5355 35127 5361
rect 35069 5352 35081 5355
rect 34664 5324 35081 5352
rect 34664 5312 34670 5324
rect 35069 5321 35081 5324
rect 35115 5321 35127 5355
rect 35434 5352 35440 5364
rect 35395 5324 35440 5352
rect 35069 5315 35127 5321
rect 35434 5312 35440 5324
rect 35492 5312 35498 5364
rect 35989 5355 36047 5361
rect 35989 5321 36001 5355
rect 36035 5352 36047 5355
rect 37182 5352 37188 5364
rect 36035 5324 37188 5352
rect 36035 5321 36047 5324
rect 35989 5315 36047 5321
rect 20901 5287 20959 5293
rect 20901 5284 20913 5287
rect 20180 5256 20913 5284
rect 20901 5253 20913 5256
rect 20947 5253 20959 5287
rect 20901 5247 20959 5253
rect 18509 5219 18567 5225
rect 18509 5216 18521 5219
rect 18064 5188 18521 5216
rect 13725 5179 13783 5185
rect 18509 5185 18521 5188
rect 18555 5185 18567 5219
rect 18509 5179 18567 5185
rect 5629 5151 5687 5157
rect 5629 5148 5641 5151
rect 5552 5120 5641 5148
rect 3326 5040 3332 5092
rect 3384 5089 3390 5092
rect 3384 5083 3448 5089
rect 3384 5049 3402 5083
rect 3436 5080 3448 5083
rect 4062 5080 4068 5092
rect 3436 5052 4068 5080
rect 3436 5049 3448 5052
rect 3384 5043 3448 5049
rect 3384 5040 3390 5043
rect 4062 5040 4068 5052
rect 4120 5040 4126 5092
rect 5552 5024 5580 5120
rect 5629 5117 5641 5120
rect 5675 5117 5687 5151
rect 6822 5148 6828 5160
rect 6783 5120 6828 5148
rect 5629 5111 5687 5117
rect 6822 5108 6828 5120
rect 6880 5148 6886 5160
rect 7377 5151 7435 5157
rect 7377 5148 7389 5151
rect 6880 5120 7389 5148
rect 6880 5108 6886 5120
rect 7377 5117 7389 5120
rect 7423 5117 7435 5151
rect 7377 5111 7435 5117
rect 10689 5151 10747 5157
rect 10689 5117 10701 5151
rect 10735 5148 10747 5151
rect 11238 5148 11244 5160
rect 10735 5120 11244 5148
rect 10735 5117 10747 5120
rect 10689 5111 10747 5117
rect 11238 5108 11244 5120
rect 11296 5108 11302 5160
rect 13998 5157 14004 5160
rect 12437 5151 12495 5157
rect 12437 5148 12449 5151
rect 12176 5120 12449 5148
rect 8846 5080 8852 5092
rect 8807 5052 8852 5080
rect 8846 5040 8852 5052
rect 8904 5040 8910 5092
rect 4154 4972 4160 5024
rect 4212 5012 4218 5024
rect 4798 5012 4804 5024
rect 4212 4984 4804 5012
rect 4212 4972 4218 4984
rect 4798 4972 4804 4984
rect 4856 5012 4862 5024
rect 5077 5015 5135 5021
rect 5077 5012 5089 5015
rect 4856 4984 5089 5012
rect 4856 4972 4862 4984
rect 5077 4981 5089 4984
rect 5123 4981 5135 5015
rect 5534 5012 5540 5024
rect 5495 4984 5540 5012
rect 5077 4975 5135 4981
rect 5534 4972 5540 4984
rect 5592 4972 5598 5024
rect 5810 5012 5816 5024
rect 5771 4984 5816 5012
rect 5810 4972 5816 4984
rect 5868 4972 5874 5024
rect 6270 5012 6276 5024
rect 6231 4984 6276 5012
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 8113 5015 8171 5021
rect 8113 4981 8125 5015
rect 8159 5012 8171 5015
rect 8754 5012 8760 5024
rect 8159 4984 8760 5012
rect 8159 4981 8171 4984
rect 8113 4975 8171 4981
rect 8754 4972 8760 4984
rect 8812 4972 8818 5024
rect 10321 5015 10379 5021
rect 10321 4981 10333 5015
rect 10367 5012 10379 5015
rect 11606 5012 11612 5024
rect 10367 4984 11612 5012
rect 10367 4981 10379 4984
rect 10321 4975 10379 4981
rect 11606 4972 11612 4984
rect 11664 4972 11670 5024
rect 11698 4972 11704 5024
rect 11756 5012 11762 5024
rect 12176 5021 12204 5120
rect 12437 5117 12449 5120
rect 12483 5117 12495 5151
rect 13992 5148 14004 5157
rect 13959 5120 14004 5148
rect 12437 5111 12495 5117
rect 13992 5111 14004 5120
rect 13998 5108 14004 5111
rect 14056 5108 14062 5160
rect 19797 5151 19855 5157
rect 19797 5148 19809 5151
rect 19628 5120 19809 5148
rect 18506 5040 18512 5092
rect 18564 5080 18570 5092
rect 18693 5083 18751 5089
rect 18693 5080 18705 5083
rect 18564 5052 18705 5080
rect 18564 5040 18570 5052
rect 18693 5049 18705 5052
rect 18739 5049 18751 5083
rect 18693 5043 18751 5049
rect 12161 5015 12219 5021
rect 12161 5012 12173 5015
rect 11756 4984 12173 5012
rect 11756 4972 11762 4984
rect 12161 4981 12173 4984
rect 12207 4981 12219 5015
rect 15102 5012 15108 5024
rect 15063 4984 15108 5012
rect 12161 4975 12219 4981
rect 15102 4972 15108 4984
rect 15160 4972 15166 5024
rect 16114 5012 16120 5024
rect 16075 4984 16120 5012
rect 16114 4972 16120 4984
rect 16172 4972 16178 5024
rect 17402 4972 17408 5024
rect 17460 5012 17466 5024
rect 18601 5015 18659 5021
rect 18601 5012 18613 5015
rect 17460 4984 18613 5012
rect 17460 4972 17466 4984
rect 18601 4981 18613 4984
rect 18647 4981 18659 5015
rect 18601 4975 18659 4981
rect 19334 4972 19340 5024
rect 19392 5012 19398 5024
rect 19628 5021 19656 5120
rect 19797 5117 19809 5120
rect 19843 5117 19855 5151
rect 20916 5148 20944 5247
rect 23492 5216 23520 5312
rect 25958 5244 25964 5296
rect 26016 5284 26022 5296
rect 26602 5284 26608 5296
rect 26016 5256 26608 5284
rect 26016 5244 26022 5256
rect 26602 5244 26608 5256
rect 26660 5244 26666 5296
rect 29365 5287 29423 5293
rect 29365 5284 29377 5287
rect 26712 5256 29377 5284
rect 24121 5219 24179 5225
rect 24121 5216 24133 5219
rect 23492 5188 24133 5216
rect 24121 5185 24133 5188
rect 24167 5185 24179 5219
rect 24121 5179 24179 5185
rect 24210 5176 24216 5228
rect 24268 5216 24274 5228
rect 24305 5219 24363 5225
rect 24305 5216 24317 5219
rect 24268 5188 24317 5216
rect 24268 5176 24274 5188
rect 24305 5185 24317 5188
rect 24351 5216 24363 5219
rect 24762 5216 24768 5228
rect 24351 5188 24768 5216
rect 24351 5185 24363 5188
rect 24305 5179 24363 5185
rect 24762 5176 24768 5188
rect 24820 5176 24826 5228
rect 26712 5225 26740 5256
rect 29365 5253 29377 5256
rect 29411 5253 29423 5287
rect 29365 5247 29423 5253
rect 25317 5219 25375 5225
rect 25317 5185 25329 5219
rect 25363 5216 25375 5219
rect 26697 5219 26755 5225
rect 26697 5216 26709 5219
rect 25363 5188 26709 5216
rect 25363 5185 25375 5188
rect 25317 5179 25375 5185
rect 26697 5185 26709 5188
rect 26743 5185 26755 5219
rect 26697 5179 26755 5185
rect 26789 5219 26847 5225
rect 26789 5185 26801 5219
rect 26835 5216 26847 5219
rect 27341 5219 27399 5225
rect 27341 5216 27353 5219
rect 26835 5188 27353 5216
rect 26835 5185 26847 5188
rect 26789 5179 26847 5185
rect 27341 5185 27353 5188
rect 27387 5185 27399 5219
rect 28994 5216 29000 5228
rect 28955 5188 29000 5216
rect 27341 5179 27399 5185
rect 21082 5148 21088 5160
rect 20916 5120 21088 5148
rect 19797 5111 19855 5117
rect 21082 5108 21088 5120
rect 21140 5108 21146 5160
rect 25685 5151 25743 5157
rect 25685 5117 25697 5151
rect 25731 5148 25743 5151
rect 26602 5148 26608 5160
rect 25731 5120 26608 5148
rect 25731 5117 25743 5120
rect 25685 5111 25743 5117
rect 26602 5108 26608 5120
rect 26660 5148 26666 5160
rect 26660 5120 26740 5148
rect 26660 5108 26666 5120
rect 21352 5083 21410 5089
rect 21352 5049 21364 5083
rect 21398 5080 21410 5083
rect 21542 5080 21548 5092
rect 21398 5052 21548 5080
rect 21398 5049 21410 5052
rect 21352 5043 21410 5049
rect 21542 5040 21548 5052
rect 21600 5040 21606 5092
rect 22738 5080 22744 5092
rect 22480 5052 22744 5080
rect 19613 5015 19671 5021
rect 19613 5012 19625 5015
rect 19392 4984 19625 5012
rect 19392 4972 19398 4984
rect 19613 4981 19625 4984
rect 19659 4981 19671 5015
rect 19978 5012 19984 5024
rect 19939 4984 19984 5012
rect 19613 4975 19671 4981
rect 19978 4972 19984 4984
rect 20036 4972 20042 5024
rect 22480 5021 22508 5052
rect 22738 5040 22744 5052
rect 22796 5080 22802 5092
rect 23658 5080 23664 5092
rect 22796 5052 23664 5080
rect 22796 5040 22802 5052
rect 23658 5040 23664 5052
rect 23716 5040 23722 5092
rect 26712 5089 26740 5120
rect 26697 5083 26755 5089
rect 26697 5049 26709 5083
rect 26743 5049 26755 5083
rect 26697 5043 26755 5049
rect 22465 5015 22523 5021
rect 22465 4981 22477 5015
rect 22511 4981 22523 5015
rect 22465 4975 22523 4981
rect 23566 4972 23572 5024
rect 23624 5012 23630 5024
rect 24213 5015 24271 5021
rect 24213 5012 24225 5015
rect 23624 4984 24225 5012
rect 23624 4972 23630 4984
rect 24213 4981 24225 4984
rect 24259 5012 24271 5015
rect 24673 5015 24731 5021
rect 24673 5012 24685 5015
rect 24259 4984 24685 5012
rect 24259 4981 24271 4984
rect 24213 4975 24271 4981
rect 24673 4981 24685 4984
rect 24719 4981 24731 5015
rect 25958 5012 25964 5024
rect 25919 4984 25964 5012
rect 24673 4975 24731 4981
rect 25958 4972 25964 4984
rect 26016 4972 26022 5024
rect 26050 4972 26056 5024
rect 26108 5012 26114 5024
rect 26804 5012 26832 5179
rect 28994 5176 29000 5188
rect 29052 5176 29058 5228
rect 29914 5216 29920 5228
rect 29875 5188 29920 5216
rect 29914 5176 29920 5188
rect 29972 5176 29978 5228
rect 36096 5225 36124 5324
rect 37182 5312 37188 5324
rect 37240 5312 37246 5364
rect 38654 5352 38660 5364
rect 38615 5324 38660 5352
rect 38654 5312 38660 5324
rect 38712 5312 38718 5364
rect 36081 5219 36139 5225
rect 36081 5185 36093 5219
rect 36127 5185 36139 5219
rect 36081 5179 36139 5185
rect 29012 5148 29040 5176
rect 31113 5151 31171 5157
rect 31113 5148 31125 5151
rect 29012 5120 31125 5148
rect 31113 5117 31125 5120
rect 31159 5148 31171 5151
rect 31297 5151 31355 5157
rect 31297 5148 31309 5151
rect 31159 5120 31309 5148
rect 31159 5117 31171 5120
rect 31113 5111 31171 5117
rect 31297 5117 31309 5120
rect 31343 5148 31355 5151
rect 31846 5148 31852 5160
rect 31343 5120 31852 5148
rect 31343 5117 31355 5120
rect 31297 5111 31355 5117
rect 31846 5108 31852 5120
rect 31904 5108 31910 5160
rect 29641 5083 29699 5089
rect 29641 5049 29653 5083
rect 29687 5080 29699 5083
rect 30742 5080 30748 5092
rect 29687 5052 30748 5080
rect 29687 5049 29699 5052
rect 29641 5043 29699 5049
rect 30742 5040 30748 5052
rect 30800 5080 30806 5092
rect 31386 5080 31392 5092
rect 30800 5052 31392 5080
rect 30800 5040 30806 5052
rect 31386 5040 31392 5052
rect 31444 5080 31450 5092
rect 31542 5083 31600 5089
rect 31542 5080 31554 5083
rect 31444 5052 31554 5080
rect 31444 5040 31450 5052
rect 31542 5049 31554 5052
rect 31588 5049 31600 5083
rect 33597 5083 33655 5089
rect 33597 5080 33609 5083
rect 31542 5043 31600 5049
rect 32692 5052 33609 5080
rect 26108 4984 26832 5012
rect 26108 4972 26114 4984
rect 29086 4972 29092 5024
rect 29144 5012 29150 5024
rect 29825 5015 29883 5021
rect 29825 5012 29837 5015
rect 29144 4984 29837 5012
rect 29144 4972 29150 4984
rect 29825 4981 29837 4984
rect 29871 5012 29883 5015
rect 30285 5015 30343 5021
rect 30285 5012 30297 5015
rect 29871 4984 30297 5012
rect 29871 4981 29883 4984
rect 29825 4975 29883 4981
rect 30285 4981 30297 4984
rect 30331 4981 30343 5015
rect 30285 4975 30343 4981
rect 32306 4972 32312 5024
rect 32364 5012 32370 5024
rect 32692 5021 32720 5052
rect 33597 5049 33609 5052
rect 33643 5049 33655 5083
rect 33597 5043 33655 5049
rect 32677 5015 32735 5021
rect 32677 5012 32689 5015
rect 32364 4984 32689 5012
rect 32364 4972 32370 4984
rect 32677 4981 32689 4984
rect 32723 4981 32735 5015
rect 32677 4975 32735 4981
rect 34606 4972 34612 5024
rect 34664 5012 34670 5024
rect 36096 5012 36124 5179
rect 40313 5151 40371 5157
rect 40313 5117 40325 5151
rect 40359 5148 40371 5151
rect 40497 5151 40555 5157
rect 40497 5148 40509 5151
rect 40359 5120 40509 5148
rect 40359 5117 40371 5120
rect 40313 5111 40371 5117
rect 40497 5117 40509 5120
rect 40543 5148 40555 5151
rect 40586 5148 40592 5160
rect 40543 5120 40592 5148
rect 40543 5117 40555 5120
rect 40497 5111 40555 5117
rect 40586 5108 40592 5120
rect 40644 5108 40650 5160
rect 36262 5040 36268 5092
rect 36320 5089 36326 5092
rect 36320 5083 36384 5089
rect 36320 5049 36338 5083
rect 36372 5049 36384 5083
rect 36320 5043 36384 5049
rect 36320 5040 36326 5043
rect 37366 5040 37372 5092
rect 37424 5080 37430 5092
rect 38381 5083 38439 5089
rect 38381 5080 38393 5083
rect 37424 5052 38393 5080
rect 37424 5040 37430 5052
rect 38381 5049 38393 5052
rect 38427 5080 38439 5083
rect 38470 5080 38476 5092
rect 38427 5052 38476 5080
rect 38427 5049 38439 5052
rect 38381 5043 38439 5049
rect 38470 5040 38476 5052
rect 38528 5080 38534 5092
rect 38933 5083 38991 5089
rect 38933 5080 38945 5083
rect 38528 5052 38945 5080
rect 38528 5040 38534 5052
rect 38933 5049 38945 5052
rect 38979 5049 38991 5083
rect 38933 5043 38991 5049
rect 39209 5083 39267 5089
rect 39209 5049 39221 5083
rect 39255 5049 39267 5083
rect 39209 5043 39267 5049
rect 37458 5012 37464 5024
rect 34664 4984 36124 5012
rect 37419 4984 37464 5012
rect 34664 4972 34670 4984
rect 37458 4972 37464 4984
rect 37516 4972 37522 5024
rect 38105 5015 38163 5021
rect 38105 4981 38117 5015
rect 38151 5012 38163 5015
rect 38194 5012 38200 5024
rect 38151 4984 38200 5012
rect 38151 4981 38163 4984
rect 38105 4975 38163 4981
rect 38194 4972 38200 4984
rect 38252 4972 38258 5024
rect 39114 5012 39120 5024
rect 39075 4984 39120 5012
rect 39114 4972 39120 4984
rect 39172 4972 39178 5024
rect 39224 5012 39252 5043
rect 40678 5040 40684 5092
rect 40736 5089 40742 5092
rect 40736 5083 40800 5089
rect 40736 5049 40754 5083
rect 40788 5049 40800 5083
rect 40736 5043 40800 5049
rect 40736 5040 40742 5043
rect 39669 5015 39727 5021
rect 39669 5012 39681 5015
rect 39224 4984 39681 5012
rect 39669 4981 39681 4984
rect 39715 5012 39727 5015
rect 40954 5012 40960 5024
rect 39715 4984 40960 5012
rect 39715 4981 39727 4984
rect 39669 4975 39727 4981
rect 40954 4972 40960 4984
rect 41012 5012 41018 5024
rect 41877 5015 41935 5021
rect 41877 5012 41889 5015
rect 41012 4984 41889 5012
rect 41012 4972 41018 4984
rect 41877 4981 41889 4984
rect 41923 4981 41935 5015
rect 41877 4975 41935 4981
rect 1104 4922 48852 4944
rect 1104 4870 19606 4922
rect 19658 4870 19670 4922
rect 19722 4870 19734 4922
rect 19786 4870 19798 4922
rect 19850 4870 48852 4922
rect 1104 4848 48852 4870
rect 3237 4811 3295 4817
rect 3237 4777 3249 4811
rect 3283 4808 3295 4811
rect 3326 4808 3332 4820
rect 3283 4780 3332 4808
rect 3283 4777 3295 4780
rect 3237 4771 3295 4777
rect 3326 4768 3332 4780
rect 3384 4768 3390 4820
rect 4341 4811 4399 4817
rect 4341 4777 4353 4811
rect 4387 4808 4399 4811
rect 4614 4808 4620 4820
rect 4387 4780 4620 4808
rect 4387 4777 4399 4780
rect 4341 4771 4399 4777
rect 4614 4768 4620 4780
rect 4672 4768 4678 4820
rect 5626 4768 5632 4820
rect 5684 4808 5690 4820
rect 6089 4811 6147 4817
rect 6089 4808 6101 4811
rect 5684 4780 6101 4808
rect 5684 4768 5690 4780
rect 6089 4777 6101 4780
rect 6135 4808 6147 4811
rect 6178 4808 6184 4820
rect 6135 4780 6184 4808
rect 6135 4777 6147 4780
rect 6089 4771 6147 4777
rect 6178 4768 6184 4780
rect 6236 4768 6242 4820
rect 7834 4808 7840 4820
rect 7795 4780 7840 4808
rect 7834 4768 7840 4780
rect 7892 4768 7898 4820
rect 11698 4808 11704 4820
rect 11659 4780 11704 4808
rect 11698 4768 11704 4780
rect 11756 4768 11762 4820
rect 12437 4811 12495 4817
rect 12437 4777 12449 4811
rect 12483 4808 12495 4811
rect 12894 4808 12900 4820
rect 12483 4780 12900 4808
rect 12483 4777 12495 4780
rect 12437 4771 12495 4777
rect 12894 4768 12900 4780
rect 12952 4768 12958 4820
rect 13814 4768 13820 4820
rect 13872 4808 13878 4820
rect 14185 4811 14243 4817
rect 14185 4808 14197 4811
rect 13872 4780 14197 4808
rect 13872 4768 13878 4780
rect 14185 4777 14197 4780
rect 14231 4777 14243 4811
rect 15838 4808 15844 4820
rect 15799 4780 15844 4808
rect 14185 4771 14243 4777
rect 15838 4768 15844 4780
rect 15896 4768 15902 4820
rect 18325 4811 18383 4817
rect 18325 4777 18337 4811
rect 18371 4808 18383 4811
rect 18506 4808 18512 4820
rect 18371 4780 18512 4808
rect 18371 4777 18383 4780
rect 18325 4771 18383 4777
rect 18506 4768 18512 4780
rect 18564 4768 18570 4820
rect 20717 4811 20775 4817
rect 20717 4777 20729 4811
rect 20763 4808 20775 4811
rect 21542 4808 21548 4820
rect 20763 4780 21548 4808
rect 20763 4777 20775 4780
rect 20717 4771 20775 4777
rect 21542 4768 21548 4780
rect 21600 4808 21606 4820
rect 21913 4811 21971 4817
rect 21913 4808 21925 4811
rect 21600 4780 21925 4808
rect 21600 4768 21606 4780
rect 21913 4777 21925 4780
rect 21959 4777 21971 4811
rect 22554 4808 22560 4820
rect 22515 4780 22560 4808
rect 21913 4771 21971 4777
rect 22554 4768 22560 4780
rect 22612 4808 22618 4820
rect 23014 4808 23020 4820
rect 22612 4780 23020 4808
rect 22612 4768 22618 4780
rect 23014 4768 23020 4780
rect 23072 4808 23078 4820
rect 23569 4811 23627 4817
rect 23072 4780 23428 4808
rect 23072 4768 23078 4780
rect 5718 4700 5724 4752
rect 5776 4740 5782 4752
rect 5905 4743 5963 4749
rect 5905 4740 5917 4743
rect 5776 4712 5917 4740
rect 5776 4700 5782 4712
rect 5905 4709 5917 4712
rect 5951 4709 5963 4743
rect 7852 4740 7880 4768
rect 23400 4752 23428 4780
rect 23569 4777 23581 4811
rect 23615 4808 23627 4811
rect 23750 4808 23756 4820
rect 23615 4780 23756 4808
rect 23615 4777 23627 4780
rect 23569 4771 23627 4777
rect 23750 4768 23756 4780
rect 23808 4808 23814 4820
rect 24026 4808 24032 4820
rect 23808 4780 24032 4808
rect 23808 4768 23814 4780
rect 24026 4768 24032 4780
rect 24084 4768 24090 4820
rect 24121 4811 24179 4817
rect 24121 4777 24133 4811
rect 24167 4808 24179 4811
rect 24210 4808 24216 4820
rect 24167 4780 24216 4808
rect 24167 4777 24179 4780
rect 24121 4771 24179 4777
rect 24210 4768 24216 4780
rect 24268 4768 24274 4820
rect 24946 4808 24952 4820
rect 24907 4780 24952 4808
rect 24946 4768 24952 4780
rect 25004 4808 25010 4820
rect 26050 4808 26056 4820
rect 25004 4780 26056 4808
rect 25004 4768 25010 4780
rect 26050 4768 26056 4780
rect 26108 4768 26114 4820
rect 27522 4808 27528 4820
rect 26896 4780 27528 4808
rect 5905 4703 5963 4709
rect 6196 4712 7880 4740
rect 6086 4632 6092 4684
rect 6144 4672 6150 4684
rect 6196 4681 6224 4712
rect 8294 4700 8300 4752
rect 8352 4740 8358 4752
rect 8573 4743 8631 4749
rect 8573 4740 8585 4743
rect 8352 4712 8585 4740
rect 8352 4700 8358 4712
rect 8573 4709 8585 4712
rect 8619 4709 8631 4743
rect 8573 4703 8631 4709
rect 16666 4700 16672 4752
rect 16724 4740 16730 4752
rect 17129 4743 17187 4749
rect 17129 4740 17141 4743
rect 16724 4712 17141 4740
rect 16724 4700 16730 4712
rect 17129 4709 17141 4712
rect 17175 4709 17187 4743
rect 21450 4740 21456 4752
rect 21411 4712 21456 4740
rect 17129 4703 17187 4709
rect 21450 4700 21456 4712
rect 21508 4740 21514 4752
rect 22002 4740 22008 4752
rect 21508 4712 22008 4740
rect 21508 4700 21514 4712
rect 22002 4700 22008 4712
rect 22060 4700 22066 4752
rect 23382 4740 23388 4752
rect 23295 4712 23388 4740
rect 23382 4700 23388 4712
rect 23440 4700 23446 4752
rect 23658 4700 23664 4752
rect 23716 4740 23722 4752
rect 26896 4749 26924 4780
rect 27522 4768 27528 4780
rect 27580 4768 27586 4820
rect 30558 4808 30564 4820
rect 30519 4780 30564 4808
rect 30558 4768 30564 4780
rect 30616 4768 30622 4820
rect 31386 4808 31392 4820
rect 31347 4780 31392 4808
rect 31386 4768 31392 4780
rect 31444 4768 31450 4820
rect 32490 4808 32496 4820
rect 32451 4780 32496 4808
rect 32490 4768 32496 4780
rect 32548 4768 32554 4820
rect 33594 4808 33600 4820
rect 33555 4780 33600 4808
rect 33594 4768 33600 4780
rect 33652 4768 33658 4820
rect 36173 4811 36231 4817
rect 36173 4777 36185 4811
rect 36219 4808 36231 4811
rect 36262 4808 36268 4820
rect 36219 4780 36268 4808
rect 36219 4777 36231 4780
rect 36173 4771 36231 4777
rect 36262 4768 36268 4780
rect 36320 4768 36326 4820
rect 37090 4808 37096 4820
rect 37051 4780 37096 4808
rect 37090 4768 37096 4780
rect 37148 4768 37154 4820
rect 38749 4811 38807 4817
rect 38749 4808 38761 4811
rect 38120 4780 38761 4808
rect 38120 4752 38148 4780
rect 38749 4777 38761 4780
rect 38795 4808 38807 4811
rect 39114 4808 39120 4820
rect 38795 4780 39120 4808
rect 38795 4777 38807 4780
rect 38749 4771 38807 4777
rect 39114 4768 39120 4780
rect 39172 4768 39178 4820
rect 40586 4808 40592 4820
rect 40547 4780 40592 4808
rect 40586 4768 40592 4780
rect 40644 4768 40650 4820
rect 40954 4808 40960 4820
rect 40915 4780 40960 4808
rect 40954 4768 40960 4780
rect 41012 4768 41018 4820
rect 26329 4743 26387 4749
rect 23716 4712 23761 4740
rect 23716 4700 23722 4712
rect 26329 4709 26341 4743
rect 26375 4740 26387 4743
rect 26881 4743 26939 4749
rect 26881 4740 26893 4743
rect 26375 4712 26893 4740
rect 26375 4709 26387 4712
rect 26329 4703 26387 4709
rect 26881 4709 26893 4712
rect 26927 4709 26939 4743
rect 27062 4740 27068 4752
rect 27023 4712 27068 4740
rect 26881 4703 26939 4709
rect 27062 4700 27068 4712
rect 27120 4700 27126 4752
rect 27157 4743 27215 4749
rect 27157 4709 27169 4743
rect 27203 4740 27215 4743
rect 28997 4743 29055 4749
rect 28997 4740 29009 4743
rect 27203 4712 29009 4740
rect 27203 4709 27215 4712
rect 27157 4703 27215 4709
rect 28997 4709 29009 4712
rect 29043 4709 29055 4743
rect 38102 4740 38108 4752
rect 38063 4712 38108 4740
rect 28997 4703 29055 4709
rect 6181 4675 6239 4681
rect 6181 4672 6193 4675
rect 6144 4644 6193 4672
rect 6144 4632 6150 4644
rect 6181 4641 6193 4644
rect 6227 4641 6239 4675
rect 8665 4675 8723 4681
rect 8665 4672 8677 4675
rect 6181 4635 6239 4641
rect 7484 4644 8677 4672
rect 5629 4539 5687 4545
rect 5629 4505 5641 4539
rect 5675 4536 5687 4539
rect 6822 4536 6828 4548
rect 5675 4508 6828 4536
rect 5675 4505 5687 4508
rect 5629 4499 5687 4505
rect 6822 4496 6828 4508
rect 6880 4496 6886 4548
rect 2682 4468 2688 4480
rect 2643 4440 2688 4468
rect 2682 4428 2688 4440
rect 2740 4428 2746 4480
rect 4706 4468 4712 4480
rect 4667 4440 4712 4468
rect 4706 4428 4712 4440
rect 4764 4428 4770 4480
rect 5261 4471 5319 4477
rect 5261 4437 5273 4471
rect 5307 4468 5319 4471
rect 5350 4468 5356 4480
rect 5307 4440 5356 4468
rect 5307 4437 5319 4440
rect 5261 4431 5319 4437
rect 5350 4428 5356 4440
rect 5408 4428 5414 4480
rect 7098 4428 7104 4480
rect 7156 4468 7162 4480
rect 7484 4477 7512 4644
rect 8665 4641 8677 4644
rect 8711 4672 8723 4675
rect 8846 4672 8852 4684
rect 8711 4644 8852 4672
rect 8711 4641 8723 4644
rect 8665 4635 8723 4641
rect 8846 4632 8852 4644
rect 8904 4632 8910 4684
rect 10045 4675 10103 4681
rect 10045 4641 10057 4675
rect 10091 4672 10103 4675
rect 10318 4672 10324 4684
rect 10091 4644 10324 4672
rect 10091 4641 10103 4644
rect 10045 4635 10103 4641
rect 10318 4632 10324 4644
rect 10376 4632 10382 4684
rect 11514 4672 11520 4684
rect 11475 4644 11520 4672
rect 11514 4632 11520 4644
rect 11572 4632 11578 4684
rect 15289 4675 15347 4681
rect 15289 4641 15301 4675
rect 15335 4641 15347 4675
rect 15289 4635 15347 4641
rect 8570 4604 8576 4616
rect 8531 4576 8576 4604
rect 8570 4564 8576 4576
rect 8628 4564 8634 4616
rect 11790 4604 11796 4616
rect 11751 4576 11796 4604
rect 11790 4564 11796 4576
rect 11848 4564 11854 4616
rect 14093 4607 14151 4613
rect 14093 4604 14105 4607
rect 13464 4576 14105 4604
rect 8113 4539 8171 4545
rect 8113 4505 8125 4539
rect 8159 4536 8171 4539
rect 8202 4536 8208 4548
rect 8159 4508 8208 4536
rect 8159 4505 8171 4508
rect 8113 4499 8171 4505
rect 8202 4496 8208 4508
rect 8260 4496 8266 4548
rect 11238 4536 11244 4548
rect 11199 4508 11244 4536
rect 11238 4496 11244 4508
rect 11296 4496 11302 4548
rect 13464 4480 13492 4576
rect 14093 4573 14105 4576
rect 14139 4573 14151 4607
rect 14093 4567 14151 4573
rect 14277 4607 14335 4613
rect 14277 4573 14289 4607
rect 14323 4604 14335 4607
rect 15010 4604 15016 4616
rect 14323 4576 15016 4604
rect 14323 4573 14335 4576
rect 14277 4567 14335 4573
rect 15010 4564 15016 4576
rect 15068 4564 15074 4616
rect 13725 4539 13783 4545
rect 13725 4505 13737 4539
rect 13771 4536 13783 4539
rect 15304 4536 15332 4635
rect 16942 4632 16948 4684
rect 17000 4672 17006 4684
rect 17218 4672 17224 4684
rect 17000 4644 17224 4672
rect 17000 4632 17006 4644
rect 17218 4632 17224 4644
rect 17276 4672 17282 4684
rect 18601 4675 18659 4681
rect 18601 4672 18613 4675
rect 17276 4644 18613 4672
rect 17276 4632 17282 4644
rect 18601 4641 18613 4644
rect 18647 4672 18659 4675
rect 18690 4672 18696 4684
rect 18647 4644 18696 4672
rect 18647 4641 18659 4644
rect 18601 4635 18659 4641
rect 18690 4632 18696 4644
rect 18748 4632 18754 4684
rect 19702 4672 19708 4684
rect 19663 4644 19708 4672
rect 19702 4632 19708 4644
rect 19760 4632 19766 4684
rect 20714 4632 20720 4684
rect 20772 4672 20778 4684
rect 20772 4644 21588 4672
rect 20772 4632 20778 4644
rect 21560 4616 21588 4644
rect 24578 4632 24584 4684
rect 24636 4672 24642 4684
rect 24765 4675 24823 4681
rect 24765 4672 24777 4675
rect 24636 4644 24777 4672
rect 24636 4632 24642 4644
rect 24765 4641 24777 4644
rect 24811 4641 24823 4675
rect 24765 4635 24823 4641
rect 26970 4632 26976 4684
rect 27028 4672 27034 4684
rect 27172 4672 27200 4703
rect 38102 4700 38108 4712
rect 38160 4700 38166 4752
rect 38286 4740 38292 4752
rect 38247 4712 38292 4740
rect 38286 4700 38292 4712
rect 38344 4700 38350 4752
rect 29454 4681 29460 4684
rect 29448 4672 29460 4681
rect 27028 4644 27200 4672
rect 29415 4644 29460 4672
rect 27028 4632 27034 4644
rect 17126 4604 17132 4616
rect 17087 4576 17132 4604
rect 17126 4564 17132 4576
rect 17184 4564 17190 4616
rect 19613 4607 19671 4613
rect 19613 4573 19625 4607
rect 19659 4604 19671 4607
rect 20622 4604 20628 4616
rect 19659 4576 20628 4604
rect 19659 4573 19671 4576
rect 19613 4567 19671 4573
rect 20622 4564 20628 4576
rect 20680 4564 20686 4616
rect 21358 4604 21364 4616
rect 21319 4576 21364 4604
rect 21358 4564 21364 4576
rect 21416 4564 21422 4616
rect 21542 4604 21548 4616
rect 21503 4576 21548 4604
rect 21542 4564 21548 4576
rect 21600 4564 21606 4616
rect 25590 4604 25596 4616
rect 25551 4576 25596 4604
rect 25590 4564 25596 4576
rect 25648 4564 25654 4616
rect 16206 4536 16212 4548
rect 13771 4508 16212 4536
rect 13771 4505 13783 4508
rect 13725 4499 13783 4505
rect 16206 4496 16212 4508
rect 16264 4496 16270 4548
rect 20349 4539 20407 4545
rect 20349 4505 20361 4539
rect 20395 4536 20407 4539
rect 20714 4536 20720 4548
rect 20395 4508 20720 4536
rect 20395 4505 20407 4508
rect 20349 4499 20407 4505
rect 20714 4496 20720 4508
rect 20772 4496 20778 4548
rect 20898 4496 20904 4548
rect 20956 4536 20962 4548
rect 20993 4539 21051 4545
rect 20993 4536 21005 4539
rect 20956 4508 21005 4536
rect 20956 4496 20962 4508
rect 20993 4505 21005 4508
rect 21039 4505 21051 4539
rect 20993 4499 21051 4505
rect 23109 4539 23167 4545
rect 23109 4505 23121 4539
rect 23155 4536 23167 4539
rect 23566 4536 23572 4548
rect 23155 4508 23572 4536
rect 23155 4505 23167 4508
rect 23109 4499 23167 4505
rect 23566 4496 23572 4508
rect 23624 4496 23630 4548
rect 26602 4536 26608 4548
rect 26563 4508 26608 4536
rect 26602 4496 26608 4508
rect 26660 4496 26666 4548
rect 7469 4471 7527 4477
rect 7469 4468 7481 4471
rect 7156 4440 7481 4468
rect 7156 4428 7162 4440
rect 7469 4437 7481 4440
rect 7515 4437 7527 4471
rect 10226 4468 10232 4480
rect 10187 4440 10232 4468
rect 7469 4431 7527 4437
rect 10226 4428 10232 4440
rect 10284 4428 10290 4480
rect 11054 4468 11060 4480
rect 11015 4440 11060 4468
rect 11054 4428 11060 4440
rect 11112 4428 11118 4480
rect 12802 4468 12808 4480
rect 12763 4440 12808 4468
rect 12802 4428 12808 4440
rect 12860 4428 12866 4480
rect 13170 4468 13176 4480
rect 13131 4440 13176 4468
rect 13170 4428 13176 4440
rect 13228 4428 13234 4480
rect 13446 4468 13452 4480
rect 13407 4440 13452 4468
rect 13446 4428 13452 4440
rect 13504 4428 13510 4480
rect 13814 4428 13820 4480
rect 13872 4468 13878 4480
rect 14090 4468 14096 4480
rect 13872 4440 14096 4468
rect 13872 4428 13878 4440
rect 14090 4428 14096 4440
rect 14148 4468 14154 4480
rect 14645 4471 14703 4477
rect 14645 4468 14657 4471
rect 14148 4440 14657 4468
rect 14148 4428 14154 4440
rect 14645 4437 14657 4440
rect 14691 4437 14703 4471
rect 15010 4468 15016 4480
rect 14971 4440 15016 4468
rect 14645 4431 14703 4437
rect 15010 4428 15016 4440
rect 15068 4428 15074 4480
rect 15470 4468 15476 4480
rect 15431 4440 15476 4468
rect 15470 4428 15476 4440
rect 15528 4428 15534 4480
rect 16669 4471 16727 4477
rect 16669 4437 16681 4471
rect 16715 4468 16727 4471
rect 17954 4468 17960 4480
rect 16715 4440 17960 4468
rect 16715 4437 16727 4440
rect 16669 4431 16727 4437
rect 17954 4428 17960 4440
rect 18012 4428 18018 4480
rect 19889 4471 19947 4477
rect 19889 4437 19901 4471
rect 19935 4468 19947 4471
rect 20530 4468 20536 4480
rect 19935 4440 20536 4468
rect 19935 4437 19947 4440
rect 19889 4431 19947 4437
rect 20530 4428 20536 4440
rect 20588 4428 20594 4480
rect 24394 4468 24400 4480
rect 24355 4440 24400 4468
rect 24394 4428 24400 4440
rect 24452 4428 24458 4480
rect 25866 4468 25872 4480
rect 25827 4440 25872 4468
rect 25866 4428 25872 4440
rect 25924 4468 25930 4480
rect 27172 4468 27200 4644
rect 29448 4635 29460 4644
rect 29454 4632 29460 4635
rect 29512 4632 29518 4684
rect 32122 4672 32128 4684
rect 32083 4644 32128 4672
rect 32122 4632 32128 4644
rect 32180 4632 32186 4684
rect 32306 4672 32312 4684
rect 32267 4644 32312 4672
rect 32306 4632 32312 4644
rect 32364 4632 32370 4684
rect 33134 4632 33140 4684
rect 33192 4672 33198 4684
rect 33413 4675 33471 4681
rect 33413 4672 33425 4675
rect 33192 4644 33425 4672
rect 33192 4632 33198 4644
rect 33413 4641 33425 4644
rect 33459 4641 33471 4675
rect 33413 4635 33471 4641
rect 37458 4632 37464 4684
rect 37516 4672 37522 4684
rect 38381 4675 38439 4681
rect 38381 4672 38393 4675
rect 37516 4644 38393 4672
rect 37516 4632 37522 4644
rect 38381 4641 38393 4644
rect 38427 4641 38439 4675
rect 38381 4635 38439 4641
rect 28994 4564 29000 4616
rect 29052 4604 29058 4616
rect 29181 4607 29239 4613
rect 29181 4604 29193 4607
rect 29052 4576 29193 4604
rect 29052 4564 29058 4576
rect 29181 4573 29193 4576
rect 29227 4573 29239 4607
rect 29181 4567 29239 4573
rect 31846 4536 31852 4548
rect 31807 4508 31852 4536
rect 31846 4496 31852 4508
rect 31904 4496 31910 4548
rect 37366 4496 37372 4548
rect 37424 4536 37430 4548
rect 37461 4539 37519 4545
rect 37461 4536 37473 4539
rect 37424 4508 37473 4536
rect 37424 4496 37430 4508
rect 37461 4505 37473 4508
rect 37507 4505 37519 4539
rect 37461 4499 37519 4505
rect 27706 4468 27712 4480
rect 25924 4440 27200 4468
rect 27667 4440 27712 4468
rect 25924 4428 25930 4440
rect 27706 4428 27712 4440
rect 27764 4428 27770 4480
rect 28169 4471 28227 4477
rect 28169 4437 28181 4471
rect 28215 4468 28227 4471
rect 28350 4468 28356 4480
rect 28215 4440 28356 4468
rect 28215 4437 28227 4440
rect 28169 4431 28227 4437
rect 28350 4428 28356 4440
rect 28408 4428 28414 4480
rect 32861 4471 32919 4477
rect 32861 4437 32873 4471
rect 32907 4468 32919 4471
rect 33042 4468 33048 4480
rect 32907 4440 33048 4468
rect 32907 4437 32919 4440
rect 32861 4431 32919 4437
rect 33042 4428 33048 4440
rect 33100 4428 33106 4480
rect 33226 4468 33232 4480
rect 33187 4440 33232 4468
rect 33226 4428 33232 4440
rect 33284 4428 33290 4480
rect 37826 4468 37832 4480
rect 37787 4440 37832 4468
rect 37826 4428 37832 4440
rect 37884 4428 37890 4480
rect 40494 4428 40500 4480
rect 40552 4468 40558 4480
rect 41233 4471 41291 4477
rect 41233 4468 41245 4471
rect 40552 4440 41245 4468
rect 40552 4428 40558 4440
rect 41233 4437 41245 4440
rect 41279 4437 41291 4471
rect 41233 4431 41291 4437
rect 1104 4378 48852 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 34966 4378
rect 35018 4326 35030 4378
rect 35082 4326 35094 4378
rect 35146 4326 35158 4378
rect 35210 4326 48852 4378
rect 1104 4304 48852 4326
rect 6178 4264 6184 4276
rect 6139 4236 6184 4264
rect 6178 4224 6184 4236
rect 6236 4224 6242 4276
rect 7193 4267 7251 4273
rect 7193 4233 7205 4267
rect 7239 4264 7251 4267
rect 7834 4264 7840 4276
rect 7239 4236 7840 4264
rect 7239 4233 7251 4236
rect 7193 4227 7251 4233
rect 7834 4224 7840 4236
rect 7892 4224 7898 4276
rect 8294 4224 8300 4276
rect 8352 4264 8358 4276
rect 8570 4264 8576 4276
rect 8352 4236 8576 4264
rect 8352 4224 8358 4236
rect 8570 4224 8576 4236
rect 8628 4264 8634 4276
rect 9861 4267 9919 4273
rect 9861 4264 9873 4267
rect 8628 4236 9873 4264
rect 8628 4224 8634 4236
rect 9861 4233 9873 4236
rect 9907 4233 9919 4267
rect 9861 4227 9919 4233
rect 10965 4267 11023 4273
rect 10965 4233 10977 4267
rect 11011 4264 11023 4267
rect 11241 4267 11299 4273
rect 11241 4264 11253 4267
rect 11011 4236 11253 4264
rect 11011 4233 11023 4236
rect 10965 4227 11023 4233
rect 11241 4233 11253 4236
rect 11287 4264 11299 4267
rect 11790 4264 11796 4276
rect 11287 4236 11796 4264
rect 11287 4233 11299 4236
rect 11241 4227 11299 4233
rect 11790 4224 11796 4236
rect 11848 4224 11854 4276
rect 12805 4267 12863 4273
rect 12805 4233 12817 4267
rect 12851 4264 12863 4267
rect 13446 4264 13452 4276
rect 12851 4236 13452 4264
rect 12851 4233 12863 4236
rect 12805 4227 12863 4233
rect 13446 4224 13452 4236
rect 13504 4224 13510 4276
rect 16206 4264 16212 4276
rect 16167 4236 16212 4264
rect 16206 4224 16212 4236
rect 16264 4224 16270 4276
rect 16666 4264 16672 4276
rect 16627 4236 16672 4264
rect 16666 4224 16672 4236
rect 16724 4224 16730 4276
rect 17126 4224 17132 4276
rect 17184 4264 17190 4276
rect 17313 4267 17371 4273
rect 17313 4264 17325 4267
rect 17184 4236 17325 4264
rect 17184 4224 17190 4236
rect 17313 4233 17325 4236
rect 17359 4233 17371 4267
rect 17313 4227 17371 4233
rect 20993 4267 21051 4273
rect 20993 4233 21005 4267
rect 21039 4264 21051 4267
rect 21450 4264 21456 4276
rect 21039 4236 21456 4264
rect 21039 4233 21051 4236
rect 20993 4227 21051 4233
rect 21450 4224 21456 4236
rect 21508 4224 21514 4276
rect 22738 4264 22744 4276
rect 22699 4236 22744 4264
rect 22738 4224 22744 4236
rect 22796 4224 22802 4276
rect 23382 4264 23388 4276
rect 23343 4236 23388 4264
rect 23382 4224 23388 4236
rect 23440 4224 23446 4276
rect 24949 4267 25007 4273
rect 24949 4233 24961 4267
rect 24995 4264 25007 4267
rect 25866 4264 25872 4276
rect 24995 4236 25872 4264
rect 24995 4233 25007 4236
rect 24949 4227 25007 4233
rect 25866 4224 25872 4236
rect 25924 4224 25930 4276
rect 28994 4264 29000 4276
rect 28955 4236 29000 4264
rect 28994 4224 29000 4236
rect 29052 4224 29058 4276
rect 33134 4224 33140 4276
rect 33192 4264 33198 4276
rect 33965 4267 34023 4273
rect 33965 4264 33977 4267
rect 33192 4236 33977 4264
rect 33192 4224 33198 4236
rect 33965 4233 33977 4236
rect 34011 4233 34023 4267
rect 33965 4227 34023 4233
rect 37369 4267 37427 4273
rect 37369 4233 37381 4267
rect 37415 4264 37427 4267
rect 37458 4264 37464 4276
rect 37415 4236 37464 4264
rect 37415 4233 37427 4236
rect 37369 4227 37427 4233
rect 37458 4224 37464 4236
rect 37516 4224 37522 4276
rect 38102 4224 38108 4276
rect 38160 4264 38166 4276
rect 38289 4267 38347 4273
rect 38289 4264 38301 4267
rect 38160 4236 38301 4264
rect 38160 4224 38166 4236
rect 38289 4233 38301 4236
rect 38335 4233 38347 4267
rect 38289 4227 38347 4233
rect 5166 4156 5172 4208
rect 5224 4196 5230 4208
rect 5261 4199 5319 4205
rect 5261 4196 5273 4199
rect 5224 4168 5273 4196
rect 5224 4156 5230 4168
rect 5261 4165 5273 4168
rect 5307 4165 5319 4199
rect 5261 4159 5319 4165
rect 5350 4156 5356 4208
rect 5408 4196 5414 4208
rect 5408 4168 5488 4196
rect 5408 4156 5414 4168
rect 5460 4128 5488 4168
rect 5810 4156 5816 4208
rect 5868 4196 5874 4208
rect 8205 4199 8263 4205
rect 5868 4168 6868 4196
rect 5868 4156 5874 4168
rect 5626 4128 5632 4140
rect 5460 4100 5632 4128
rect 5626 4088 5632 4100
rect 5684 4088 5690 4140
rect 6840 4128 6868 4168
rect 8205 4165 8217 4199
rect 8251 4165 8263 4199
rect 8205 4159 8263 4165
rect 7929 4131 7987 4137
rect 7929 4128 7941 4131
rect 6840 4100 7941 4128
rect 7929 4097 7941 4100
rect 7975 4128 7987 4131
rect 8110 4128 8116 4140
rect 7975 4100 8116 4128
rect 7975 4097 7987 4100
rect 7929 4091 7987 4097
rect 8110 4088 8116 4100
rect 8168 4088 8174 4140
rect 8220 4128 8248 4159
rect 11514 4156 11520 4208
rect 11572 4196 11578 4208
rect 11974 4196 11980 4208
rect 11572 4168 11980 4196
rect 11572 4156 11578 4168
rect 11974 4156 11980 4168
rect 12032 4156 12038 4208
rect 21358 4196 21364 4208
rect 20640 4168 21364 4196
rect 9493 4131 9551 4137
rect 9493 4128 9505 4131
rect 8220 4100 9505 4128
rect 9493 4097 9505 4100
rect 9539 4128 9551 4131
rect 11698 4128 11704 4140
rect 9539 4100 9720 4128
rect 11659 4100 11704 4128
rect 9539 4097 9551 4100
rect 9493 4091 9551 4097
rect 9692 4069 9720 4100
rect 11698 4088 11704 4100
rect 11756 4088 11762 4140
rect 13170 4128 13176 4140
rect 13131 4100 13176 4128
rect 13170 4088 13176 4100
rect 13228 4088 13234 4140
rect 13354 4128 13360 4140
rect 13315 4100 13360 4128
rect 13354 4088 13360 4100
rect 13412 4088 13418 4140
rect 13817 4131 13875 4137
rect 13817 4097 13829 4131
rect 13863 4128 13875 4131
rect 18601 4131 18659 4137
rect 13863 4100 14412 4128
rect 13863 4097 13875 4100
rect 13817 4091 13875 4097
rect 2593 4063 2651 4069
rect 2593 4029 2605 4063
rect 2639 4029 2651 4063
rect 2593 4023 2651 4029
rect 7009 4063 7067 4069
rect 7009 4029 7021 4063
rect 7055 4060 7067 4063
rect 8481 4063 8539 4069
rect 7055 4032 7696 4060
rect 7055 4029 7067 4032
rect 7009 4023 7067 4029
rect 2608 3936 2636 4023
rect 2774 3952 2780 4004
rect 2832 4001 2838 4004
rect 2832 3995 2896 4001
rect 2832 3961 2850 3995
rect 2884 3992 2896 3995
rect 4062 3992 4068 4004
rect 2884 3964 4068 3992
rect 2884 3961 2896 3964
rect 2832 3955 2896 3961
rect 2832 3952 2838 3955
rect 4062 3952 4068 3964
rect 4120 3952 4126 4004
rect 4706 3992 4712 4004
rect 4619 3964 4712 3992
rect 4706 3952 4712 3964
rect 4764 3992 4770 4004
rect 5810 3992 5816 4004
rect 4764 3964 5816 3992
rect 4764 3952 4770 3964
rect 5810 3952 5816 3964
rect 5868 3952 5874 4004
rect 2501 3927 2559 3933
rect 2501 3893 2513 3927
rect 2547 3924 2559 3927
rect 2590 3924 2596 3936
rect 2547 3896 2596 3924
rect 2547 3893 2559 3896
rect 2501 3887 2559 3893
rect 2590 3884 2596 3896
rect 2648 3884 2654 3936
rect 2958 3884 2964 3936
rect 3016 3924 3022 3936
rect 3973 3927 4031 3933
rect 3973 3924 3985 3927
rect 3016 3896 3985 3924
rect 3016 3884 3022 3896
rect 3973 3893 3985 3896
rect 4019 3893 4031 3927
rect 5074 3924 5080 3936
rect 5035 3896 5080 3924
rect 3973 3887 4031 3893
rect 5074 3884 5080 3896
rect 5132 3924 5138 3936
rect 7668 3933 7696 4032
rect 8481 4029 8493 4063
rect 8527 4060 8539 4063
rect 9677 4063 9735 4069
rect 8527 4032 9260 4060
rect 8527 4029 8539 4032
rect 8481 4023 8539 4029
rect 8754 3992 8760 4004
rect 8715 3964 8760 3992
rect 8754 3952 8760 3964
rect 8812 3952 8818 4004
rect 9232 3936 9260 4032
rect 9677 4029 9689 4063
rect 9723 4029 9735 4063
rect 11054 4060 11060 4072
rect 10967 4032 11060 4060
rect 9677 4023 9735 4029
rect 11054 4020 11060 4032
rect 11112 4060 11118 4072
rect 12342 4060 12348 4072
rect 11112 4032 12348 4060
rect 11112 4020 11118 4032
rect 12342 4020 12348 4032
rect 12400 4020 12406 4072
rect 12802 4020 12808 4072
rect 12860 4060 12866 4072
rect 13832 4060 13860 4091
rect 14277 4063 14335 4069
rect 14277 4060 14289 4063
rect 12860 4032 13860 4060
rect 14108 4032 14289 4060
rect 12860 4020 12866 4032
rect 13280 4001 13308 4032
rect 13265 3995 13323 4001
rect 13265 3961 13277 3995
rect 13311 3961 13323 3995
rect 13265 3955 13323 3961
rect 13538 3952 13544 4004
rect 13596 3992 13602 4004
rect 14108 4001 14136 4032
rect 14277 4029 14289 4032
rect 14323 4029 14335 4063
rect 14384 4060 14412 4100
rect 18601 4097 18613 4131
rect 18647 4128 18659 4131
rect 19061 4131 19119 4137
rect 19061 4128 19073 4131
rect 18647 4100 19073 4128
rect 18647 4097 18659 4100
rect 18601 4091 18659 4097
rect 19061 4097 19073 4100
rect 19107 4128 19119 4131
rect 19426 4128 19432 4140
rect 19107 4100 19432 4128
rect 19107 4097 19119 4100
rect 19061 4091 19119 4097
rect 19426 4088 19432 4100
rect 19484 4088 19490 4140
rect 19518 4088 19524 4140
rect 19576 4128 19582 4140
rect 20533 4131 20591 4137
rect 20533 4128 20545 4131
rect 19576 4100 20545 4128
rect 19576 4088 19582 4100
rect 20533 4097 20545 4100
rect 20579 4128 20591 4131
rect 20640 4128 20668 4168
rect 21358 4156 21364 4168
rect 21416 4156 21422 4208
rect 32306 4196 32312 4208
rect 31680 4168 32312 4196
rect 20579 4100 20668 4128
rect 20579 4097 20591 4100
rect 20533 4091 20591 4097
rect 20714 4088 20720 4140
rect 20772 4128 20778 4140
rect 21729 4131 21787 4137
rect 21729 4128 21741 4131
rect 20772 4100 21741 4128
rect 20772 4088 20778 4100
rect 21729 4097 21741 4100
rect 21775 4097 21787 4131
rect 21729 4091 21787 4097
rect 25869 4131 25927 4137
rect 25869 4097 25881 4131
rect 25915 4128 25927 4131
rect 25958 4128 25964 4140
rect 25915 4100 25964 4128
rect 25915 4097 25927 4100
rect 25869 4091 25927 4097
rect 25958 4088 25964 4100
rect 26016 4088 26022 4140
rect 27706 4088 27712 4140
rect 27764 4128 27770 4140
rect 28261 4131 28319 4137
rect 28261 4128 28273 4131
rect 27764 4100 28273 4128
rect 27764 4088 27770 4100
rect 28261 4097 28273 4100
rect 28307 4128 28319 4131
rect 29546 4128 29552 4140
rect 28307 4100 29552 4128
rect 28307 4097 28319 4100
rect 28261 4091 28319 4097
rect 29546 4088 29552 4100
rect 29604 4088 29610 4140
rect 31389 4131 31447 4137
rect 31389 4097 31401 4131
rect 31435 4128 31447 4131
rect 31680 4128 31708 4168
rect 32306 4156 32312 4168
rect 32364 4156 32370 4208
rect 33594 4128 33600 4140
rect 31435 4100 31708 4128
rect 32968 4100 33600 4128
rect 31435 4097 31447 4100
rect 31389 4091 31447 4097
rect 14544 4063 14602 4069
rect 14544 4060 14556 4063
rect 14384 4032 14556 4060
rect 14277 4023 14335 4029
rect 14544 4029 14556 4032
rect 14590 4060 14602 4063
rect 15102 4060 15108 4072
rect 14590 4032 15108 4060
rect 14590 4029 14602 4032
rect 14544 4023 14602 4029
rect 15102 4020 15108 4032
rect 15160 4020 15166 4072
rect 16761 4063 16819 4069
rect 16761 4029 16773 4063
rect 16807 4060 16819 4063
rect 16850 4060 16856 4072
rect 16807 4032 16856 4060
rect 16807 4029 16819 4032
rect 16761 4023 16819 4029
rect 16850 4020 16856 4032
rect 16908 4020 16914 4072
rect 17770 4020 17776 4072
rect 17828 4060 17834 4072
rect 18123 4063 18181 4069
rect 18123 4060 18135 4063
rect 17828 4032 18135 4060
rect 17828 4020 17834 4032
rect 18123 4029 18135 4032
rect 18169 4029 18181 4063
rect 18690 4060 18696 4072
rect 18651 4032 18696 4060
rect 18123 4023 18181 4029
rect 18690 4020 18696 4032
rect 18748 4020 18754 4072
rect 19334 4020 19340 4072
rect 19392 4060 19398 4072
rect 19702 4060 19708 4072
rect 19392 4032 19708 4060
rect 19392 4020 19398 4032
rect 19702 4020 19708 4032
rect 19760 4020 19766 4072
rect 19981 4063 20039 4069
rect 19981 4029 19993 4063
rect 20027 4060 20039 4063
rect 20254 4060 20260 4072
rect 20027 4032 20260 4060
rect 20027 4029 20039 4032
rect 19981 4023 20039 4029
rect 20254 4020 20260 4032
rect 20312 4060 20318 4072
rect 21159 4063 21217 4069
rect 21159 4060 21171 4063
rect 20312 4032 21171 4060
rect 20312 4020 20318 4032
rect 21159 4029 21171 4032
rect 21205 4029 21217 4063
rect 21159 4023 21217 4029
rect 23566 4020 23572 4072
rect 23624 4060 23630 4072
rect 23661 4063 23719 4069
rect 23661 4060 23673 4063
rect 23624 4032 23673 4060
rect 23624 4020 23630 4032
rect 23661 4029 23673 4032
rect 23707 4060 23719 4063
rect 24213 4063 24271 4069
rect 24213 4060 24225 4063
rect 23707 4032 24225 4060
rect 23707 4029 23719 4032
rect 23661 4023 23719 4029
rect 24213 4029 24225 4032
rect 24259 4029 24271 4063
rect 24762 4060 24768 4072
rect 24723 4032 24768 4060
rect 24213 4023 24271 4029
rect 24762 4020 24768 4032
rect 24820 4060 24826 4072
rect 25317 4063 25375 4069
rect 25317 4060 25329 4063
rect 24820 4032 25329 4060
rect 24820 4020 24826 4032
rect 25317 4029 25329 4032
rect 25363 4029 25375 4063
rect 25317 4023 25375 4029
rect 27525 4063 27583 4069
rect 27525 4029 27537 4063
rect 27571 4060 27583 4063
rect 27571 4032 28212 4060
rect 27571 4029 27583 4032
rect 27525 4023 27583 4029
rect 14093 3995 14151 4001
rect 14093 3992 14105 3995
rect 13596 3964 14105 3992
rect 13596 3952 13602 3964
rect 14093 3961 14105 3964
rect 14139 3961 14151 3995
rect 19720 3992 19748 4020
rect 19720 3964 20300 3992
rect 14093 3955 14151 3961
rect 5721 3927 5779 3933
rect 5721 3924 5733 3927
rect 5132 3896 5733 3924
rect 5132 3884 5138 3896
rect 5721 3893 5733 3896
rect 5767 3893 5779 3927
rect 5721 3887 5779 3893
rect 7653 3927 7711 3933
rect 7653 3893 7665 3927
rect 7699 3924 7711 3927
rect 7742 3924 7748 3936
rect 7699 3896 7748 3924
rect 7699 3893 7711 3896
rect 7653 3887 7711 3893
rect 7742 3884 7748 3896
rect 7800 3884 7806 3936
rect 8294 3884 8300 3936
rect 8352 3924 8358 3936
rect 8665 3927 8723 3933
rect 8665 3924 8677 3927
rect 8352 3896 8677 3924
rect 8352 3884 8358 3896
rect 8665 3893 8677 3896
rect 8711 3893 8723 3927
rect 9214 3924 9220 3936
rect 9175 3896 9220 3924
rect 8665 3887 8723 3893
rect 9214 3884 9220 3896
rect 9272 3884 9278 3936
rect 10318 3924 10324 3936
rect 10279 3896 10324 3924
rect 10318 3884 10324 3896
rect 10376 3884 10382 3936
rect 15654 3924 15660 3936
rect 15615 3896 15660 3924
rect 15654 3884 15660 3896
rect 15712 3884 15718 3936
rect 16942 3924 16948 3936
rect 16903 3896 16948 3924
rect 16942 3884 16948 3896
rect 17000 3884 17006 3936
rect 17862 3924 17868 3936
rect 17823 3896 17868 3924
rect 17862 3884 17868 3896
rect 17920 3924 17926 3936
rect 18598 3924 18604 3936
rect 17920 3896 18604 3924
rect 17920 3884 17926 3896
rect 18598 3884 18604 3896
rect 18656 3884 18662 3936
rect 20162 3924 20168 3936
rect 20123 3896 20168 3924
rect 20162 3884 20168 3896
rect 20220 3884 20226 3936
rect 20272 3924 20300 3964
rect 20806 3952 20812 4004
rect 20864 3992 20870 4004
rect 21453 3995 21511 4001
rect 21453 3992 21465 3995
rect 20864 3964 21465 3992
rect 20864 3952 20870 3964
rect 21453 3961 21465 3964
rect 21499 3961 21511 3995
rect 24946 3992 24952 4004
rect 21453 3955 21511 3961
rect 23860 3964 24952 3992
rect 21637 3927 21695 3933
rect 21637 3924 21649 3927
rect 20272 3896 21649 3924
rect 21637 3893 21649 3896
rect 21683 3924 21695 3927
rect 22097 3927 22155 3933
rect 22097 3924 22109 3927
rect 21683 3896 22109 3924
rect 21683 3893 21695 3896
rect 21637 3887 21695 3893
rect 22097 3893 22109 3896
rect 22143 3893 22155 3927
rect 23106 3924 23112 3936
rect 23067 3896 23112 3924
rect 22097 3887 22155 3893
rect 23106 3884 23112 3896
rect 23164 3884 23170 3936
rect 23860 3933 23888 3964
rect 24946 3952 24952 3964
rect 25004 3952 25010 4004
rect 26234 3952 26240 4004
rect 26292 3992 26298 4004
rect 26292 3964 26337 3992
rect 26292 3952 26298 3964
rect 27614 3952 27620 4004
rect 27672 3992 27678 4004
rect 27985 3995 28043 4001
rect 27985 3992 27997 3995
rect 27672 3964 27997 3992
rect 27672 3952 27678 3964
rect 27985 3961 27997 3964
rect 28031 3961 28043 3995
rect 27985 3955 28043 3961
rect 28184 3936 28212 4032
rect 28994 4020 29000 4072
rect 29052 4060 29058 4072
rect 29270 4060 29276 4072
rect 29052 4032 29276 4060
rect 29052 4020 29058 4032
rect 29270 4020 29276 4032
rect 29328 4060 29334 4072
rect 29825 4063 29883 4069
rect 29825 4060 29837 4063
rect 29328 4032 29837 4060
rect 29328 4020 29334 4032
rect 29825 4029 29837 4032
rect 29871 4029 29883 4063
rect 30374 4060 30380 4072
rect 30335 4032 30380 4060
rect 29825 4023 29883 4029
rect 30374 4020 30380 4032
rect 30432 4060 30438 4072
rect 30929 4063 30987 4069
rect 30929 4060 30941 4063
rect 30432 4032 30941 4060
rect 30432 4020 30438 4032
rect 30929 4029 30941 4032
rect 30975 4029 30987 4063
rect 30929 4023 30987 4029
rect 30282 3992 30288 4004
rect 29472 3964 30288 3992
rect 23845 3927 23903 3933
rect 23845 3893 23857 3927
rect 23891 3893 23903 3927
rect 24578 3924 24584 3936
rect 24539 3896 24584 3924
rect 23845 3887 23903 3893
rect 24578 3884 24584 3896
rect 24636 3884 24642 3936
rect 26326 3924 26332 3936
rect 26287 3896 26332 3924
rect 26326 3884 26332 3896
rect 26384 3884 26390 3936
rect 26602 3884 26608 3936
rect 26660 3924 26666 3936
rect 26789 3927 26847 3933
rect 26789 3924 26801 3927
rect 26660 3896 26801 3924
rect 26660 3884 26666 3896
rect 26789 3893 26801 3896
rect 26835 3893 26847 3927
rect 26789 3887 26847 3893
rect 27699 3927 27757 3933
rect 27699 3893 27711 3927
rect 27745 3924 27757 3927
rect 28074 3924 28080 3936
rect 27745 3896 28080 3924
rect 27745 3893 27757 3896
rect 27699 3887 27757 3893
rect 28074 3884 28080 3896
rect 28132 3884 28138 3936
rect 28166 3884 28172 3936
rect 28224 3924 28230 3936
rect 28626 3924 28632 3936
rect 28224 3896 28269 3924
rect 28587 3896 28632 3924
rect 28224 3884 28230 3896
rect 28626 3884 28632 3896
rect 28684 3884 28690 3936
rect 29472 3933 29500 3964
rect 30282 3952 30288 3964
rect 30340 3952 30346 4004
rect 32582 3992 32588 4004
rect 30576 3964 32588 3992
rect 30576 3933 30604 3964
rect 32582 3952 32588 3964
rect 32640 3992 32646 4004
rect 32968 4001 32996 4100
rect 33594 4088 33600 4100
rect 33652 4088 33658 4140
rect 38013 4131 38071 4137
rect 38013 4097 38025 4131
rect 38059 4128 38071 4131
rect 38286 4128 38292 4140
rect 38059 4100 38292 4128
rect 38059 4097 38071 4100
rect 38013 4091 38071 4097
rect 38286 4088 38292 4100
rect 38344 4088 38350 4140
rect 39850 4128 39856 4140
rect 39811 4100 39856 4128
rect 39850 4088 39856 4100
rect 39908 4128 39914 4140
rect 40402 4128 40408 4140
rect 39908 4100 40408 4128
rect 39908 4088 39914 4100
rect 40402 4088 40408 4100
rect 40460 4128 40466 4140
rect 40957 4131 41015 4137
rect 40957 4128 40969 4131
rect 40460 4100 40969 4128
rect 40460 4088 40466 4100
rect 40957 4097 40969 4100
rect 41003 4097 41015 4131
rect 40957 4091 41015 4097
rect 40494 4060 40500 4072
rect 40455 4032 40500 4060
rect 40494 4020 40500 4032
rect 40552 4020 40558 4072
rect 40770 4060 40776 4072
rect 40604 4032 40776 4060
rect 32953 3995 33011 4001
rect 32953 3992 32965 3995
rect 32640 3964 32965 3992
rect 32640 3952 32646 3964
rect 32953 3961 32965 3964
rect 32999 3961 33011 3995
rect 32953 3955 33011 3961
rect 33226 3952 33232 4004
rect 33284 3992 33290 4004
rect 33284 3964 33329 3992
rect 33284 3952 33290 3964
rect 40034 3952 40040 4004
rect 40092 3992 40098 4004
rect 40604 3992 40632 4032
rect 40770 4020 40776 4032
rect 40828 4060 40834 4072
rect 41233 4063 41291 4069
rect 41233 4060 41245 4063
rect 40828 4032 41245 4060
rect 40828 4020 40834 4032
rect 41233 4029 41245 4032
rect 41279 4029 41291 4063
rect 41233 4023 41291 4029
rect 40092 3964 40632 3992
rect 40092 3952 40098 3964
rect 29457 3927 29515 3933
rect 29457 3893 29469 3927
rect 29503 3893 29515 3927
rect 29457 3887 29515 3893
rect 30561 3927 30619 3933
rect 30561 3893 30573 3927
rect 30607 3893 30619 3927
rect 31478 3924 31484 3936
rect 31439 3896 31484 3924
rect 30561 3887 30619 3893
rect 31478 3884 31484 3896
rect 31536 3884 31542 3936
rect 32122 3924 32128 3936
rect 32083 3896 32128 3924
rect 32122 3884 32128 3896
rect 32180 3884 32186 3936
rect 32667 3927 32725 3933
rect 32667 3893 32679 3927
rect 32713 3924 32725 3927
rect 33042 3924 33048 3936
rect 32713 3896 33048 3924
rect 32713 3893 32725 3896
rect 32667 3887 32725 3893
rect 33042 3884 33048 3896
rect 33100 3884 33106 3936
rect 33134 3884 33140 3936
rect 33192 3924 33198 3936
rect 33962 3924 33968 3936
rect 33192 3896 33968 3924
rect 33192 3884 33198 3896
rect 33962 3884 33968 3896
rect 34020 3884 34026 3936
rect 34882 3924 34888 3936
rect 34843 3896 34888 3924
rect 34882 3884 34888 3896
rect 34940 3884 34946 3936
rect 37366 3884 37372 3936
rect 37424 3924 37430 3936
rect 37461 3927 37519 3933
rect 37461 3924 37473 3927
rect 37424 3896 37473 3924
rect 37424 3884 37430 3896
rect 37461 3893 37473 3896
rect 37507 3893 37519 3927
rect 39390 3924 39396 3936
rect 39351 3896 39396 3924
rect 37461 3887 37519 3893
rect 39390 3884 39396 3896
rect 39448 3884 39454 3936
rect 40313 3927 40371 3933
rect 40313 3893 40325 3927
rect 40359 3924 40371 3927
rect 40959 3927 41017 3933
rect 40959 3924 40971 3927
rect 40359 3896 40971 3924
rect 40359 3893 40371 3896
rect 40313 3887 40371 3893
rect 40959 3893 40971 3896
rect 41005 3924 41017 3927
rect 41046 3924 41052 3936
rect 41005 3896 41052 3924
rect 41005 3893 41017 3896
rect 40959 3887 41017 3893
rect 41046 3884 41052 3896
rect 41104 3884 41110 3936
rect 42334 3924 42340 3936
rect 42295 3896 42340 3924
rect 42334 3884 42340 3896
rect 42392 3884 42398 3936
rect 1104 3834 48852 3856
rect 1104 3782 19606 3834
rect 19658 3782 19670 3834
rect 19722 3782 19734 3834
rect 19786 3782 19798 3834
rect 19850 3782 48852 3834
rect 1104 3760 48852 3782
rect 2314 3720 2320 3732
rect 2227 3692 2320 3720
rect 2314 3680 2320 3692
rect 2372 3720 2378 3732
rect 2958 3720 2964 3732
rect 2372 3692 2964 3720
rect 2372 3680 2378 3692
rect 2958 3680 2964 3692
rect 3016 3680 3022 3732
rect 3881 3723 3939 3729
rect 3881 3720 3893 3723
rect 3068 3692 3893 3720
rect 3068 3661 3096 3692
rect 3881 3689 3893 3692
rect 3927 3720 3939 3723
rect 4614 3720 4620 3732
rect 3927 3692 4620 3720
rect 3927 3689 3939 3692
rect 3881 3683 3939 3689
rect 4614 3680 4620 3692
rect 4672 3680 4678 3732
rect 5718 3720 5724 3732
rect 5679 3692 5724 3720
rect 5718 3680 5724 3692
rect 5776 3680 5782 3732
rect 6086 3720 6092 3732
rect 6047 3692 6092 3720
rect 6086 3680 6092 3692
rect 6144 3680 6150 3732
rect 8202 3720 8208 3732
rect 8163 3692 8208 3720
rect 8202 3680 8208 3692
rect 8260 3680 8266 3732
rect 13630 3720 13636 3732
rect 13591 3692 13636 3720
rect 13630 3680 13636 3692
rect 13688 3680 13694 3732
rect 15470 3680 15476 3732
rect 15528 3720 15534 3732
rect 15933 3723 15991 3729
rect 15933 3720 15945 3723
rect 15528 3692 15945 3720
rect 15528 3680 15534 3692
rect 15933 3689 15945 3692
rect 15979 3720 15991 3723
rect 16758 3720 16764 3732
rect 15979 3692 16764 3720
rect 15979 3689 15991 3692
rect 15933 3683 15991 3689
rect 16758 3680 16764 3692
rect 16816 3680 16822 3732
rect 17218 3720 17224 3732
rect 17179 3692 17224 3720
rect 17218 3680 17224 3692
rect 17276 3680 17282 3732
rect 18598 3680 18604 3732
rect 18656 3720 18662 3732
rect 19245 3723 19303 3729
rect 19245 3720 19257 3723
rect 18656 3692 19257 3720
rect 18656 3680 18662 3692
rect 19245 3689 19257 3692
rect 19291 3689 19303 3723
rect 19245 3683 19303 3689
rect 19426 3680 19432 3732
rect 19484 3720 19490 3732
rect 19797 3723 19855 3729
rect 19797 3720 19809 3723
rect 19484 3692 19809 3720
rect 19484 3680 19490 3692
rect 19797 3689 19809 3692
rect 19843 3720 19855 3723
rect 20070 3720 20076 3732
rect 19843 3692 20076 3720
rect 19843 3689 19855 3692
rect 19797 3683 19855 3689
rect 20070 3680 20076 3692
rect 20128 3680 20134 3732
rect 20254 3720 20260 3732
rect 20215 3692 20260 3720
rect 20254 3680 20260 3692
rect 20312 3680 20318 3732
rect 20714 3680 20720 3732
rect 20772 3720 20778 3732
rect 21085 3723 21143 3729
rect 21085 3720 21097 3723
rect 20772 3692 21097 3720
rect 20772 3680 20778 3692
rect 21085 3689 21097 3692
rect 21131 3689 21143 3723
rect 21542 3720 21548 3732
rect 21503 3692 21548 3720
rect 21085 3683 21143 3689
rect 21542 3680 21548 3692
rect 21600 3680 21606 3732
rect 22087 3723 22145 3729
rect 22087 3689 22099 3723
rect 22133 3720 22145 3723
rect 24305 3723 24363 3729
rect 24305 3720 24317 3723
rect 22133 3692 24317 3720
rect 22133 3689 22145 3692
rect 22087 3683 22145 3689
rect 24305 3689 24317 3692
rect 24351 3720 24363 3723
rect 24394 3720 24400 3732
rect 24351 3692 24400 3720
rect 24351 3689 24363 3692
rect 24305 3683 24363 3689
rect 24394 3680 24400 3692
rect 24452 3680 24458 3732
rect 25501 3723 25559 3729
rect 25501 3689 25513 3723
rect 25547 3720 25559 3723
rect 26142 3720 26148 3732
rect 25547 3692 26148 3720
rect 25547 3689 25559 3692
rect 25501 3683 25559 3689
rect 26142 3680 26148 3692
rect 26200 3680 26206 3732
rect 26234 3680 26240 3732
rect 26292 3720 26298 3732
rect 26970 3720 26976 3732
rect 26292 3692 26976 3720
rect 26292 3680 26298 3692
rect 26970 3680 26976 3692
rect 27028 3720 27034 3732
rect 27065 3723 27123 3729
rect 27065 3720 27077 3723
rect 27028 3692 27077 3720
rect 27028 3680 27034 3692
rect 27065 3689 27077 3692
rect 27111 3689 27123 3723
rect 29454 3720 29460 3732
rect 29367 3692 29460 3720
rect 27065 3683 27123 3689
rect 29454 3680 29460 3692
rect 29512 3680 29518 3732
rect 30466 3720 30472 3732
rect 30427 3692 30472 3720
rect 30466 3680 30472 3692
rect 30524 3680 30530 3732
rect 32587 3723 32645 3729
rect 32587 3689 32599 3723
rect 32633 3720 32645 3723
rect 32674 3720 32680 3732
rect 32633 3692 32680 3720
rect 32633 3689 32645 3692
rect 32587 3683 32645 3689
rect 32674 3680 32680 3692
rect 32732 3680 32738 3732
rect 33962 3720 33968 3732
rect 33923 3692 33968 3720
rect 33962 3680 33968 3692
rect 34020 3680 34026 3732
rect 34514 3720 34520 3732
rect 34475 3692 34520 3720
rect 34514 3680 34520 3692
rect 34572 3720 34578 3732
rect 35621 3723 35679 3729
rect 35621 3720 35633 3723
rect 34572 3692 35633 3720
rect 34572 3680 34578 3692
rect 35621 3689 35633 3692
rect 35667 3689 35679 3723
rect 35621 3683 35679 3689
rect 37093 3723 37151 3729
rect 37093 3689 37105 3723
rect 37139 3720 37151 3723
rect 37826 3720 37832 3732
rect 37139 3692 37832 3720
rect 37139 3689 37151 3692
rect 37093 3683 37151 3689
rect 37826 3680 37832 3692
rect 37884 3720 37890 3732
rect 38289 3723 38347 3729
rect 38289 3720 38301 3723
rect 37884 3692 38301 3720
rect 37884 3680 37890 3692
rect 38289 3689 38301 3692
rect 38335 3689 38347 3723
rect 40770 3720 40776 3732
rect 40731 3692 40776 3720
rect 38289 3683 38347 3689
rect 40770 3680 40776 3692
rect 40828 3680 40834 3732
rect 3053 3655 3111 3661
rect 3053 3621 3065 3655
rect 3099 3621 3111 3655
rect 3053 3615 3111 3621
rect 4706 3612 4712 3664
rect 4764 3652 4770 3664
rect 5169 3655 5227 3661
rect 5169 3652 5181 3655
rect 4764 3624 5181 3652
rect 4764 3612 4770 3624
rect 5169 3621 5181 3624
rect 5215 3621 5227 3655
rect 5169 3615 5227 3621
rect 5626 3612 5632 3664
rect 5684 3652 5690 3664
rect 6426 3655 6484 3661
rect 6426 3652 6438 3655
rect 5684 3624 6438 3652
rect 5684 3612 5690 3624
rect 6426 3621 6438 3624
rect 6472 3621 6484 3655
rect 6426 3615 6484 3621
rect 9490 3612 9496 3664
rect 9548 3652 9554 3664
rect 10229 3655 10287 3661
rect 10229 3652 10241 3655
rect 9548 3624 10241 3652
rect 9548 3612 9554 3624
rect 10229 3621 10241 3624
rect 10275 3621 10287 3655
rect 10229 3615 10287 3621
rect 13170 3612 13176 3664
rect 13228 3652 13234 3664
rect 15013 3655 15071 3661
rect 15013 3652 15025 3655
rect 13228 3624 15025 3652
rect 13228 3612 13234 3624
rect 15013 3621 15025 3624
rect 15059 3652 15071 3655
rect 15654 3652 15660 3664
rect 15059 3624 15660 3652
rect 15059 3621 15071 3624
rect 15013 3615 15071 3621
rect 15654 3612 15660 3624
rect 15712 3612 15718 3664
rect 15838 3612 15844 3664
rect 15896 3652 15902 3664
rect 16025 3655 16083 3661
rect 16025 3652 16037 3655
rect 15896 3624 16037 3652
rect 15896 3612 15902 3624
rect 16025 3621 16037 3624
rect 16071 3621 16083 3655
rect 16025 3615 16083 3621
rect 17126 3612 17132 3664
rect 17184 3652 17190 3664
rect 18110 3655 18168 3661
rect 18110 3652 18122 3655
rect 17184 3624 18122 3652
rect 17184 3612 17190 3624
rect 18110 3621 18122 3624
rect 18156 3621 18168 3655
rect 18110 3615 18168 3621
rect 20162 3612 20168 3664
rect 20220 3652 20226 3664
rect 21821 3655 21879 3661
rect 21821 3652 21833 3655
rect 20220 3624 21833 3652
rect 20220 3612 20226 3624
rect 21821 3621 21833 3624
rect 21867 3652 21879 3655
rect 22557 3655 22615 3661
rect 22557 3652 22569 3655
rect 21867 3624 22569 3652
rect 21867 3621 21879 3624
rect 21821 3615 21879 3621
rect 22557 3621 22569 3624
rect 22603 3621 22615 3655
rect 22557 3615 22615 3621
rect 23661 3655 23719 3661
rect 23661 3621 23673 3655
rect 23707 3652 23719 3655
rect 23934 3652 23940 3664
rect 23707 3624 23940 3652
rect 23707 3621 23719 3624
rect 23661 3615 23719 3621
rect 23934 3612 23940 3624
rect 23992 3652 23998 3664
rect 24121 3655 24179 3661
rect 24121 3652 24133 3655
rect 23992 3624 24133 3652
rect 23992 3612 23998 3624
rect 24121 3621 24133 3624
rect 24167 3621 24179 3655
rect 24121 3615 24179 3621
rect 26326 3612 26332 3664
rect 26384 3652 26390 3664
rect 26881 3655 26939 3661
rect 26881 3652 26893 3655
rect 26384 3624 26893 3652
rect 26384 3612 26390 3624
rect 26881 3621 26893 3624
rect 26927 3621 26939 3655
rect 28626 3652 28632 3664
rect 26881 3615 26939 3621
rect 27172 3624 28632 3652
rect 4525 3587 4583 3593
rect 4525 3553 4537 3587
rect 4571 3584 4583 3587
rect 5261 3587 5319 3593
rect 5261 3584 5273 3587
rect 4571 3556 5273 3584
rect 4571 3553 4583 3556
rect 4525 3547 4583 3553
rect 5261 3553 5273 3556
rect 5307 3584 5319 3587
rect 6086 3584 6092 3596
rect 5307 3556 6092 3584
rect 5307 3553 5319 3556
rect 5261 3547 5319 3553
rect 6086 3544 6092 3556
rect 6144 3544 6150 3596
rect 9125 3587 9183 3593
rect 9125 3553 9137 3587
rect 9171 3584 9183 3587
rect 10045 3587 10103 3593
rect 10045 3584 10057 3587
rect 9171 3556 10057 3584
rect 9171 3553 9183 3556
rect 9125 3547 9183 3553
rect 10045 3553 10057 3556
rect 10091 3584 10103 3587
rect 11149 3587 11207 3593
rect 11149 3584 11161 3587
rect 10091 3556 11161 3584
rect 10091 3553 10103 3556
rect 10045 3547 10103 3553
rect 11149 3553 11161 3556
rect 11195 3584 11207 3587
rect 11238 3584 11244 3596
rect 11195 3556 11244 3584
rect 11195 3553 11207 3556
rect 11149 3547 11207 3553
rect 11238 3544 11244 3556
rect 11296 3584 11302 3596
rect 11589 3587 11647 3593
rect 11589 3584 11601 3587
rect 11296 3556 11601 3584
rect 11296 3544 11302 3556
rect 11589 3553 11601 3556
rect 11635 3553 11647 3587
rect 13814 3584 13820 3596
rect 13775 3556 13820 3584
rect 11589 3547 11647 3553
rect 13814 3544 13820 3556
rect 13872 3544 13878 3596
rect 14737 3587 14795 3593
rect 14737 3553 14749 3587
rect 14783 3584 14795 3587
rect 15749 3587 15807 3593
rect 15749 3584 15761 3587
rect 14783 3556 15761 3584
rect 14783 3553 14795 3556
rect 14737 3547 14795 3553
rect 15749 3553 15761 3556
rect 15795 3584 15807 3587
rect 16942 3584 16948 3596
rect 15795 3556 16948 3584
rect 15795 3553 15807 3556
rect 15749 3547 15807 3553
rect 16942 3544 16948 3556
rect 17000 3544 17006 3596
rect 17678 3544 17684 3596
rect 17736 3584 17742 3596
rect 17865 3587 17923 3593
rect 17865 3584 17877 3587
rect 17736 3556 17877 3584
rect 17736 3544 17742 3556
rect 17865 3553 17877 3556
rect 17911 3553 17923 3587
rect 17865 3547 17923 3553
rect 20714 3544 20720 3596
rect 20772 3584 20778 3596
rect 20901 3587 20959 3593
rect 20901 3584 20913 3587
rect 20772 3556 20913 3584
rect 20772 3544 20778 3556
rect 20901 3553 20913 3556
rect 20947 3584 20959 3587
rect 22094 3584 22100 3596
rect 20947 3556 22100 3584
rect 20947 3553 20959 3556
rect 20901 3547 20959 3553
rect 22094 3544 22100 3556
rect 22152 3544 22158 3596
rect 22370 3584 22376 3596
rect 22331 3556 22376 3584
rect 22370 3544 22376 3556
rect 22428 3544 22434 3596
rect 23474 3544 23480 3596
rect 23532 3584 23538 3596
rect 24397 3587 24455 3593
rect 24397 3584 24409 3587
rect 23532 3556 24409 3584
rect 23532 3544 23538 3556
rect 24397 3553 24409 3556
rect 24443 3553 24455 3587
rect 24397 3547 24455 3553
rect 25317 3587 25375 3593
rect 25317 3553 25329 3587
rect 25363 3584 25375 3587
rect 25590 3584 25596 3596
rect 25363 3556 25596 3584
rect 25363 3553 25375 3556
rect 25317 3547 25375 3553
rect 25590 3544 25596 3556
rect 25648 3544 25654 3596
rect 27172 3593 27200 3624
rect 28626 3612 28632 3624
rect 28684 3652 28690 3664
rect 29472 3652 29500 3680
rect 28684 3624 29500 3652
rect 28684 3612 28690 3624
rect 34882 3612 34888 3664
rect 34940 3652 34946 3664
rect 35250 3652 35256 3664
rect 34940 3624 35256 3652
rect 34940 3612 34946 3624
rect 35250 3612 35256 3624
rect 35308 3652 35314 3664
rect 35437 3655 35495 3661
rect 35437 3652 35449 3655
rect 35308 3624 35449 3652
rect 35308 3612 35314 3624
rect 35437 3621 35449 3624
rect 35483 3621 35495 3655
rect 37458 3652 37464 3664
rect 37419 3624 37464 3652
rect 35437 3615 35495 3621
rect 37458 3612 37464 3624
rect 37516 3612 37522 3664
rect 39390 3612 39396 3664
rect 39448 3652 39454 3664
rect 40037 3655 40095 3661
rect 40037 3652 40049 3655
rect 39448 3624 40049 3652
rect 39448 3612 39454 3624
rect 40037 3621 40049 3624
rect 40083 3621 40095 3655
rect 40218 3652 40224 3664
rect 40179 3624 40224 3652
rect 40037 3615 40095 3621
rect 40218 3612 40224 3624
rect 40276 3612 40282 3664
rect 25961 3587 26019 3593
rect 25961 3553 25973 3587
rect 26007 3584 26019 3587
rect 27157 3587 27215 3593
rect 27157 3584 27169 3587
rect 26007 3556 27169 3584
rect 26007 3553 26019 3556
rect 25961 3547 26019 3553
rect 27157 3553 27169 3556
rect 27203 3553 27215 3587
rect 27157 3547 27215 3553
rect 27706 3544 27712 3596
rect 27764 3584 27770 3596
rect 28350 3593 28356 3596
rect 28344 3584 28356 3593
rect 27764 3556 28356 3584
rect 27764 3544 27770 3556
rect 28344 3547 28356 3556
rect 28408 3584 28414 3596
rect 29086 3584 29092 3596
rect 28408 3556 29092 3584
rect 28350 3544 28356 3547
rect 28408 3544 28414 3556
rect 29086 3544 29092 3556
rect 29144 3544 29150 3596
rect 30926 3584 30932 3596
rect 30887 3556 30932 3584
rect 30926 3544 30932 3556
rect 30984 3544 30990 3596
rect 31938 3584 31944 3596
rect 31851 3556 31944 3584
rect 31938 3544 31944 3556
rect 31996 3584 32002 3596
rect 32861 3587 32919 3593
rect 32861 3584 32873 3587
rect 31996 3556 32873 3584
rect 31996 3544 32002 3556
rect 32861 3553 32873 3556
rect 32907 3553 32919 3587
rect 32861 3547 32919 3553
rect 37366 3544 37372 3596
rect 37424 3584 37430 3596
rect 38105 3587 38163 3593
rect 38105 3584 38117 3587
rect 37424 3556 38117 3584
rect 37424 3544 37430 3556
rect 38105 3553 38117 3556
rect 38151 3553 38163 3587
rect 38105 3547 38163 3553
rect 39209 3587 39267 3593
rect 39209 3553 39221 3587
rect 39255 3584 39267 3587
rect 40236 3584 40264 3612
rect 39255 3556 40264 3584
rect 41233 3587 41291 3593
rect 39255 3553 39267 3556
rect 39209 3547 39267 3553
rect 41233 3553 41245 3587
rect 41279 3553 41291 3587
rect 41233 3547 41291 3553
rect 2961 3519 3019 3525
rect 2961 3516 2973 3519
rect 1688 3488 2973 3516
rect 1688 3392 1716 3488
rect 2961 3485 2973 3488
rect 3007 3485 3019 3519
rect 5166 3516 5172 3528
rect 5127 3488 5172 3516
rect 2961 3479 3019 3485
rect 2498 3448 2504 3460
rect 2459 3420 2504 3448
rect 2498 3408 2504 3420
rect 2556 3408 2562 3460
rect 2976 3448 3004 3479
rect 5166 3476 5172 3488
rect 5224 3476 5230 3528
rect 6178 3516 6184 3528
rect 6139 3488 6184 3516
rect 6178 3476 6184 3488
rect 6236 3476 6242 3528
rect 9582 3476 9588 3528
rect 9640 3516 9646 3528
rect 10321 3519 10379 3525
rect 10321 3516 10333 3519
rect 9640 3488 10333 3516
rect 9640 3476 9646 3488
rect 10321 3485 10333 3488
rect 10367 3516 10379 3519
rect 10689 3519 10747 3525
rect 10689 3516 10701 3519
rect 10367 3488 10701 3516
rect 10367 3485 10379 3488
rect 10321 3479 10379 3485
rect 10689 3485 10701 3488
rect 10735 3485 10747 3519
rect 11330 3516 11336 3528
rect 11291 3488 11336 3516
rect 10689 3479 10747 3485
rect 11330 3476 11336 3488
rect 11388 3476 11394 3528
rect 15102 3476 15108 3528
rect 15160 3516 15166 3528
rect 15838 3516 15844 3528
rect 15160 3488 15844 3516
rect 15160 3476 15166 3488
rect 15838 3476 15844 3488
rect 15896 3476 15902 3528
rect 22649 3519 22707 3525
rect 22649 3485 22661 3519
rect 22695 3516 22707 3519
rect 22830 3516 22836 3528
rect 22695 3488 22836 3516
rect 22695 3485 22707 3488
rect 22649 3479 22707 3485
rect 22830 3476 22836 3488
rect 22888 3516 22894 3528
rect 23750 3516 23756 3528
rect 22888 3488 23756 3516
rect 22888 3476 22894 3488
rect 23750 3476 23756 3488
rect 23808 3476 23814 3528
rect 26329 3519 26387 3525
rect 26329 3485 26341 3519
rect 26375 3516 26387 3519
rect 26418 3516 26424 3528
rect 26375 3488 26424 3516
rect 26375 3485 26387 3488
rect 26329 3479 26387 3485
rect 26418 3476 26424 3488
rect 26476 3476 26482 3528
rect 28077 3519 28135 3525
rect 28077 3485 28089 3519
rect 28123 3485 28135 3519
rect 28077 3479 28135 3485
rect 4709 3451 4767 3457
rect 2976 3420 3556 3448
rect 3528 3392 3556 3420
rect 4709 3417 4721 3451
rect 4755 3448 4767 3451
rect 5442 3448 5448 3460
rect 4755 3420 5448 3448
rect 4755 3417 4767 3420
rect 4709 3411 4767 3417
rect 5442 3408 5448 3420
rect 5500 3408 5506 3460
rect 9214 3408 9220 3460
rect 9272 3448 9278 3460
rect 9769 3451 9827 3457
rect 9769 3448 9781 3451
rect 9272 3420 9781 3448
rect 9272 3408 9278 3420
rect 9769 3417 9781 3420
rect 9815 3417 9827 3451
rect 15470 3448 15476 3460
rect 15431 3420 15476 3448
rect 9769 3411 9827 3417
rect 15470 3408 15476 3420
rect 15528 3408 15534 3460
rect 20714 3448 20720 3460
rect 20675 3420 20720 3448
rect 20714 3408 20720 3420
rect 20772 3408 20778 3460
rect 23842 3448 23848 3460
rect 23803 3420 23848 3448
rect 23842 3408 23848 3420
rect 23900 3408 23906 3460
rect 26602 3448 26608 3460
rect 26563 3420 26608 3448
rect 26602 3408 26608 3420
rect 26660 3408 26666 3460
rect 27614 3448 27620 3460
rect 27575 3420 27620 3448
rect 27614 3408 27620 3420
rect 27672 3408 27678 3460
rect 1670 3380 1676 3392
rect 1631 3352 1676 3380
rect 1670 3340 1676 3352
rect 1728 3340 1734 3392
rect 3510 3380 3516 3392
rect 3471 3352 3516 3380
rect 3510 3340 3516 3352
rect 3568 3340 3574 3392
rect 7561 3383 7619 3389
rect 7561 3349 7573 3383
rect 7607 3380 7619 3383
rect 7650 3380 7656 3392
rect 7607 3352 7656 3380
rect 7607 3349 7619 3352
rect 7561 3343 7619 3349
rect 7650 3340 7656 3352
rect 7708 3340 7714 3392
rect 8294 3340 8300 3392
rect 8352 3380 8358 3392
rect 8481 3383 8539 3389
rect 8481 3380 8493 3383
rect 8352 3352 8493 3380
rect 8352 3340 8358 3352
rect 8481 3349 8493 3352
rect 8527 3349 8539 3383
rect 9490 3380 9496 3392
rect 9451 3352 9496 3380
rect 8481 3343 8539 3349
rect 9490 3340 9496 3352
rect 9548 3340 9554 3392
rect 12710 3380 12716 3392
rect 12623 3352 12716 3380
rect 12710 3340 12716 3352
rect 12768 3380 12774 3392
rect 13265 3383 13323 3389
rect 13265 3380 13277 3383
rect 12768 3352 13277 3380
rect 12768 3340 12774 3352
rect 13265 3349 13277 3352
rect 13311 3349 13323 3383
rect 13265 3343 13323 3349
rect 14001 3383 14059 3389
rect 14001 3349 14013 3383
rect 14047 3380 14059 3383
rect 15010 3380 15016 3392
rect 14047 3352 15016 3380
rect 14047 3349 14059 3352
rect 14001 3343 14059 3349
rect 15010 3340 15016 3352
rect 15068 3380 15074 3392
rect 16482 3380 16488 3392
rect 15068 3352 16488 3380
rect 15068 3340 15074 3352
rect 16482 3340 16488 3352
rect 16540 3340 16546 3392
rect 16850 3380 16856 3392
rect 16811 3352 16856 3380
rect 16850 3340 16856 3352
rect 16908 3340 16914 3392
rect 17770 3380 17776 3392
rect 17731 3352 17776 3380
rect 17770 3340 17776 3352
rect 17828 3340 17834 3392
rect 23293 3383 23351 3389
rect 23293 3349 23305 3383
rect 23339 3380 23351 3383
rect 23474 3380 23480 3392
rect 23339 3352 23480 3380
rect 23339 3349 23351 3352
rect 23293 3343 23351 3349
rect 23474 3340 23480 3352
rect 23532 3340 23538 3392
rect 24854 3380 24860 3392
rect 24767 3352 24860 3380
rect 24854 3340 24860 3352
rect 24912 3380 24918 3392
rect 25133 3383 25191 3389
rect 25133 3380 25145 3383
rect 24912 3352 25145 3380
rect 24912 3340 24918 3352
rect 25133 3349 25145 3352
rect 25179 3349 25191 3383
rect 28092 3380 28120 3479
rect 31846 3476 31852 3528
rect 31904 3516 31910 3528
rect 32125 3519 32183 3525
rect 32125 3516 32137 3519
rect 31904 3488 32137 3516
rect 31904 3476 31910 3488
rect 32125 3485 32137 3488
rect 32171 3485 32183 3519
rect 32582 3516 32588 3528
rect 32543 3488 32588 3516
rect 32125 3479 32183 3485
rect 32582 3476 32588 3488
rect 32640 3476 32646 3528
rect 34977 3519 35035 3525
rect 34977 3485 34989 3519
rect 35023 3516 35035 3519
rect 35342 3516 35348 3528
rect 35023 3488 35348 3516
rect 35023 3485 35035 3488
rect 34977 3479 35035 3485
rect 35342 3476 35348 3488
rect 35400 3516 35406 3528
rect 35713 3519 35771 3525
rect 35713 3516 35725 3519
rect 35400 3488 35725 3516
rect 35400 3476 35406 3488
rect 35713 3485 35725 3488
rect 35759 3485 35771 3519
rect 35713 3479 35771 3485
rect 38381 3519 38439 3525
rect 38381 3485 38393 3519
rect 38427 3516 38439 3519
rect 38562 3516 38568 3528
rect 38427 3488 38568 3516
rect 38427 3485 38439 3488
rect 38381 3479 38439 3485
rect 38562 3476 38568 3488
rect 38620 3476 38626 3528
rect 39577 3519 39635 3525
rect 39577 3485 39589 3519
rect 39623 3516 39635 3519
rect 40313 3519 40371 3525
rect 40313 3516 40325 3519
rect 39623 3488 40325 3516
rect 39623 3485 39635 3488
rect 39577 3479 39635 3485
rect 40313 3485 40325 3488
rect 40359 3516 40371 3519
rect 40678 3516 40684 3528
rect 40359 3488 40684 3516
rect 40359 3485 40371 3488
rect 40313 3479 40371 3485
rect 40678 3476 40684 3488
rect 40736 3476 40742 3528
rect 31481 3451 31539 3457
rect 31481 3448 31493 3451
rect 30392 3420 31493 3448
rect 30392 3392 30420 3420
rect 31481 3417 31493 3420
rect 31527 3417 31539 3451
rect 41248 3448 41276 3547
rect 41785 3451 41843 3457
rect 41785 3448 41797 3451
rect 31481 3411 31539 3417
rect 39776 3420 41797 3448
rect 39776 3392 39804 3420
rect 41785 3417 41797 3420
rect 41831 3417 41843 3451
rect 41785 3411 41843 3417
rect 28810 3380 28816 3392
rect 28092 3352 28816 3380
rect 25133 3343 25191 3349
rect 28810 3340 28816 3352
rect 28868 3340 28874 3392
rect 30193 3383 30251 3389
rect 30193 3349 30205 3383
rect 30239 3380 30251 3383
rect 30374 3380 30380 3392
rect 30239 3352 30380 3380
rect 30239 3349 30251 3352
rect 30193 3343 30251 3349
rect 30374 3340 30380 3352
rect 30432 3340 30438 3392
rect 31110 3380 31116 3392
rect 31071 3352 31116 3380
rect 31110 3340 31116 3352
rect 31168 3340 31174 3392
rect 34514 3340 34520 3392
rect 34572 3380 34578 3392
rect 35161 3383 35219 3389
rect 35161 3380 35173 3383
rect 34572 3352 35173 3380
rect 34572 3340 34578 3352
rect 35161 3349 35173 3352
rect 35207 3349 35219 3383
rect 37826 3380 37832 3392
rect 37787 3352 37832 3380
rect 35161 3343 35219 3349
rect 37826 3340 37832 3352
rect 37884 3340 37890 3392
rect 39758 3380 39764 3392
rect 39719 3352 39764 3380
rect 39758 3340 39764 3352
rect 39816 3340 39822 3392
rect 41046 3380 41052 3392
rect 41007 3352 41052 3380
rect 41046 3340 41052 3352
rect 41104 3340 41110 3392
rect 41138 3340 41144 3392
rect 41196 3380 41202 3392
rect 41417 3383 41475 3389
rect 41417 3380 41429 3383
rect 41196 3352 41429 3380
rect 41196 3340 41202 3352
rect 41417 3349 41429 3352
rect 41463 3349 41475 3383
rect 41417 3343 41475 3349
rect 1104 3290 48852 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 34966 3290
rect 35018 3238 35030 3290
rect 35082 3238 35094 3290
rect 35146 3238 35158 3290
rect 35210 3238 48852 3290
rect 1104 3216 48852 3238
rect 2314 3176 2320 3188
rect 2275 3148 2320 3176
rect 2314 3136 2320 3148
rect 2372 3136 2378 3188
rect 3510 3136 3516 3188
rect 3568 3176 3574 3188
rect 4157 3179 4215 3185
rect 4157 3176 4169 3179
rect 3568 3148 4169 3176
rect 3568 3136 3574 3148
rect 4157 3145 4169 3148
rect 4203 3145 4215 3179
rect 4706 3176 4712 3188
rect 4667 3148 4712 3176
rect 4157 3139 4215 3145
rect 4706 3136 4712 3148
rect 4764 3136 4770 3188
rect 5166 3176 5172 3188
rect 5127 3148 5172 3176
rect 5166 3136 5172 3148
rect 5224 3136 5230 3188
rect 5537 3179 5595 3185
rect 5537 3145 5549 3179
rect 5583 3176 5595 3179
rect 5810 3176 5816 3188
rect 5583 3148 5816 3176
rect 5583 3145 5595 3148
rect 5537 3139 5595 3145
rect 5810 3136 5816 3148
rect 5868 3176 5874 3188
rect 8478 3176 8484 3188
rect 5868 3148 8484 3176
rect 5868 3136 5874 3148
rect 8478 3136 8484 3148
rect 8536 3136 8542 3188
rect 11238 3176 11244 3188
rect 11199 3148 11244 3176
rect 11238 3136 11244 3148
rect 11296 3136 11302 3188
rect 13814 3136 13820 3188
rect 13872 3176 13878 3188
rect 14090 3176 14096 3188
rect 13872 3148 14096 3176
rect 13872 3136 13878 3148
rect 14090 3136 14096 3148
rect 14148 3176 14154 3188
rect 14369 3179 14427 3185
rect 14369 3176 14381 3179
rect 14148 3148 14381 3176
rect 14148 3136 14154 3148
rect 14369 3145 14381 3148
rect 14415 3145 14427 3179
rect 16390 3176 16396 3188
rect 16303 3148 16396 3176
rect 14369 3139 14427 3145
rect 16390 3136 16396 3148
rect 16448 3176 16454 3188
rect 16666 3176 16672 3188
rect 16448 3148 16672 3176
rect 16448 3136 16454 3148
rect 16666 3136 16672 3148
rect 16724 3136 16730 3188
rect 16850 3136 16856 3188
rect 16908 3176 16914 3188
rect 18141 3179 18199 3185
rect 18141 3176 18153 3179
rect 16908 3148 18153 3176
rect 16908 3136 16914 3148
rect 18141 3145 18153 3148
rect 18187 3145 18199 3179
rect 18141 3139 18199 3145
rect 20714 3136 20720 3188
rect 20772 3176 20778 3188
rect 21729 3179 21787 3185
rect 21729 3176 21741 3179
rect 20772 3148 21741 3176
rect 20772 3136 20778 3148
rect 21729 3145 21741 3148
rect 21775 3176 21787 3179
rect 22370 3176 22376 3188
rect 21775 3148 22376 3176
rect 21775 3145 21787 3148
rect 21729 3139 21787 3145
rect 22370 3136 22376 3148
rect 22428 3136 22434 3188
rect 23477 3179 23535 3185
rect 23477 3145 23489 3179
rect 23523 3176 23535 3179
rect 23658 3176 23664 3188
rect 23523 3148 23664 3176
rect 23523 3145 23535 3148
rect 23477 3139 23535 3145
rect 23658 3136 23664 3148
rect 23716 3136 23722 3188
rect 26050 3176 26056 3188
rect 26011 3148 26056 3176
rect 26050 3136 26056 3148
rect 26108 3136 26114 3188
rect 26510 3176 26516 3188
rect 26252 3148 26516 3176
rect 16758 3068 16764 3120
rect 16816 3108 16822 3120
rect 16945 3111 17003 3117
rect 16945 3108 16957 3111
rect 16816 3080 16957 3108
rect 16816 3068 16822 3080
rect 16945 3077 16957 3080
rect 16991 3077 17003 3111
rect 16945 3071 17003 3077
rect 17126 3068 17132 3120
rect 17184 3108 17190 3120
rect 17310 3108 17316 3120
rect 17184 3080 17316 3108
rect 17184 3068 17190 3080
rect 17310 3068 17316 3080
rect 17368 3108 17374 3120
rect 17405 3111 17463 3117
rect 17405 3108 17417 3111
rect 17368 3080 17417 3108
rect 17368 3068 17374 3080
rect 17405 3077 17417 3080
rect 17451 3077 17463 3111
rect 17405 3071 17463 3077
rect 17678 3068 17684 3120
rect 17736 3108 17742 3120
rect 17773 3111 17831 3117
rect 17773 3108 17785 3111
rect 17736 3080 17785 3108
rect 17736 3068 17742 3080
rect 17773 3077 17785 3080
rect 17819 3108 17831 3111
rect 18046 3108 18052 3120
rect 17819 3080 18052 3108
rect 17819 3077 17831 3080
rect 17773 3071 17831 3077
rect 18046 3068 18052 3080
rect 18104 3108 18110 3120
rect 19613 3111 19671 3117
rect 19613 3108 19625 3111
rect 18104 3080 19625 3108
rect 18104 3068 18110 3080
rect 19613 3077 19625 3080
rect 19659 3108 19671 3111
rect 19659 3080 19840 3108
rect 19659 3077 19671 3080
rect 19613 3071 19671 3077
rect 16482 3000 16488 3052
rect 16540 3040 16546 3052
rect 17696 3040 17724 3068
rect 18690 3040 18696 3052
rect 16540 3012 17724 3040
rect 18651 3012 18696 3040
rect 16540 3000 16546 3012
rect 18690 3000 18696 3012
rect 18748 3000 18754 3052
rect 19812 3049 19840 3080
rect 22094 3068 22100 3120
rect 22152 3108 22158 3120
rect 22649 3111 22707 3117
rect 22649 3108 22661 3111
rect 22152 3080 22661 3108
rect 22152 3068 22158 3080
rect 22649 3077 22661 3080
rect 22695 3077 22707 3111
rect 22649 3071 22707 3077
rect 23676 3049 23704 3136
rect 26252 3049 26280 3148
rect 26510 3136 26516 3148
rect 26568 3136 26574 3188
rect 28077 3179 28135 3185
rect 28077 3145 28089 3179
rect 28123 3176 28135 3179
rect 28166 3176 28172 3188
rect 28123 3148 28172 3176
rect 28123 3145 28135 3148
rect 28077 3139 28135 3145
rect 28166 3136 28172 3148
rect 28224 3136 28230 3188
rect 28721 3179 28779 3185
rect 28721 3145 28733 3179
rect 28767 3176 28779 3179
rect 28902 3176 28908 3188
rect 28767 3148 28908 3176
rect 28767 3145 28779 3148
rect 28721 3139 28779 3145
rect 28902 3136 28908 3148
rect 28960 3176 28966 3188
rect 29362 3176 29368 3188
rect 28960 3148 29368 3176
rect 28960 3136 28966 3148
rect 29362 3136 29368 3148
rect 29420 3136 29426 3188
rect 29546 3176 29552 3188
rect 29507 3148 29552 3176
rect 29546 3136 29552 3148
rect 29604 3136 29610 3188
rect 30926 3136 30932 3188
rect 30984 3176 30990 3188
rect 31113 3179 31171 3185
rect 31113 3176 31125 3179
rect 30984 3148 31125 3176
rect 30984 3136 30990 3148
rect 31113 3145 31125 3148
rect 31159 3176 31171 3179
rect 31662 3176 31668 3188
rect 31159 3148 31668 3176
rect 31159 3145 31171 3148
rect 31113 3139 31171 3145
rect 31662 3136 31668 3148
rect 31720 3136 31726 3188
rect 33594 3176 33600 3188
rect 33555 3148 33600 3176
rect 33594 3136 33600 3148
rect 33652 3136 33658 3188
rect 34606 3176 34612 3188
rect 34567 3148 34612 3176
rect 34606 3136 34612 3148
rect 34664 3136 34670 3188
rect 36909 3179 36967 3185
rect 36909 3145 36921 3179
rect 36955 3176 36967 3179
rect 37366 3176 37372 3188
rect 36955 3148 37372 3176
rect 36955 3145 36967 3148
rect 36909 3139 36967 3145
rect 37366 3136 37372 3148
rect 37424 3136 37430 3188
rect 39390 3136 39396 3188
rect 39448 3176 39454 3188
rect 39669 3179 39727 3185
rect 39669 3176 39681 3179
rect 39448 3148 39681 3176
rect 39448 3136 39454 3148
rect 39669 3145 39681 3148
rect 39715 3145 39727 3179
rect 39669 3139 39727 3145
rect 40313 3179 40371 3185
rect 40313 3145 40325 3179
rect 40359 3176 40371 3179
rect 40494 3176 40500 3188
rect 40359 3148 40500 3176
rect 40359 3145 40371 3148
rect 40313 3139 40371 3145
rect 40494 3136 40500 3148
rect 40552 3136 40558 3188
rect 40678 3136 40684 3188
rect 40736 3176 40742 3188
rect 41877 3179 41935 3185
rect 41877 3176 41889 3179
rect 40736 3148 41889 3176
rect 40736 3136 40742 3148
rect 41877 3145 41889 3148
rect 41923 3145 41935 3179
rect 41877 3139 41935 3145
rect 29086 3108 29092 3120
rect 29047 3080 29092 3108
rect 29086 3068 29092 3080
rect 29144 3068 29150 3120
rect 30190 3108 30196 3120
rect 30151 3080 30196 3108
rect 30190 3068 30196 3080
rect 30248 3068 30254 3120
rect 19797 3043 19855 3049
rect 19797 3009 19809 3043
rect 19843 3009 19855 3043
rect 19797 3003 19855 3009
rect 23661 3043 23719 3049
rect 23661 3009 23673 3043
rect 23707 3009 23719 3043
rect 23661 3003 23719 3009
rect 26237 3043 26295 3049
rect 26237 3009 26249 3043
rect 26283 3009 26295 3043
rect 26237 3003 26295 3009
rect 2590 2972 2596 2984
rect 2503 2944 2596 2972
rect 2590 2932 2596 2944
rect 2648 2972 2654 2984
rect 2777 2975 2835 2981
rect 2777 2972 2789 2975
rect 2648 2944 2789 2972
rect 2648 2932 2654 2944
rect 2777 2941 2789 2944
rect 2823 2941 2835 2975
rect 2777 2935 2835 2941
rect 5629 2975 5687 2981
rect 5629 2941 5641 2975
rect 5675 2972 5687 2975
rect 6273 2975 6331 2981
rect 6273 2972 6285 2975
rect 5675 2944 6285 2972
rect 5675 2941 5687 2944
rect 5629 2935 5687 2941
rect 6273 2941 6285 2944
rect 6319 2972 6331 2975
rect 7190 2972 7196 2984
rect 6319 2944 7196 2972
rect 6319 2941 6331 2944
rect 6273 2935 6331 2941
rect 7190 2932 7196 2944
rect 7248 2932 7254 2984
rect 7650 2981 7656 2984
rect 7377 2975 7435 2981
rect 7377 2941 7389 2975
rect 7423 2941 7435 2975
rect 7644 2972 7656 2981
rect 7611 2944 7656 2972
rect 7377 2935 7435 2941
rect 7644 2935 7656 2944
rect 1486 2796 1492 2848
rect 1544 2836 1550 2848
rect 2608 2845 2636 2932
rect 2958 2864 2964 2916
rect 3016 2913 3022 2916
rect 3016 2907 3080 2913
rect 3016 2873 3034 2907
rect 3068 2873 3080 2907
rect 3016 2867 3080 2873
rect 3016 2864 3022 2867
rect 1581 2839 1639 2845
rect 1581 2836 1593 2839
rect 1544 2808 1593 2836
rect 1544 2796 1550 2808
rect 1581 2805 1593 2808
rect 1627 2836 1639 2839
rect 2593 2839 2651 2845
rect 2593 2836 2605 2839
rect 1627 2808 2605 2836
rect 1627 2805 1639 2808
rect 1581 2799 1639 2805
rect 2593 2805 2605 2808
rect 2639 2805 2651 2839
rect 2593 2799 2651 2805
rect 5350 2796 5356 2848
rect 5408 2836 5414 2848
rect 6178 2836 6184 2848
rect 5408 2808 6184 2836
rect 5408 2796 5414 2808
rect 6178 2796 6184 2808
rect 6236 2836 6242 2848
rect 6549 2839 6607 2845
rect 6549 2836 6561 2839
rect 6236 2808 6561 2836
rect 6236 2796 6242 2808
rect 6549 2805 6561 2808
rect 6595 2836 6607 2839
rect 7193 2839 7251 2845
rect 7193 2836 7205 2839
rect 6595 2808 7205 2836
rect 6595 2805 6607 2808
rect 6549 2799 6607 2805
rect 7193 2805 7205 2808
rect 7239 2836 7251 2839
rect 7392 2836 7420 2935
rect 7650 2932 7656 2935
rect 7708 2932 7714 2984
rect 9766 2932 9772 2984
rect 9824 2972 9830 2984
rect 9861 2975 9919 2981
rect 9861 2972 9873 2975
rect 9824 2944 9873 2972
rect 9824 2932 9830 2944
rect 9861 2941 9873 2944
rect 9907 2972 9919 2975
rect 11330 2972 11336 2984
rect 9907 2944 11336 2972
rect 9907 2941 9919 2944
rect 9861 2935 9919 2941
rect 11330 2932 11336 2944
rect 11388 2972 11394 2984
rect 12710 2981 12716 2984
rect 11793 2975 11851 2981
rect 11793 2972 11805 2975
rect 11388 2944 11805 2972
rect 11388 2932 11394 2944
rect 11793 2941 11805 2944
rect 11839 2972 11851 2975
rect 12161 2975 12219 2981
rect 12161 2972 12173 2975
rect 11839 2944 12173 2972
rect 11839 2941 11851 2944
rect 11793 2935 11851 2941
rect 12161 2941 12173 2944
rect 12207 2972 12219 2975
rect 12437 2975 12495 2981
rect 12437 2972 12449 2975
rect 12207 2944 12449 2972
rect 12207 2941 12219 2944
rect 12161 2935 12219 2941
rect 12437 2941 12449 2944
rect 12483 2941 12495 2975
rect 12704 2972 12716 2981
rect 12671 2944 12716 2972
rect 12437 2935 12495 2941
rect 12704 2935 12716 2944
rect 9401 2907 9459 2913
rect 9401 2873 9413 2907
rect 9447 2904 9459 2907
rect 9490 2904 9496 2916
rect 9447 2876 9496 2904
rect 9447 2873 9459 2876
rect 9401 2867 9459 2873
rect 9490 2864 9496 2876
rect 9548 2904 9554 2916
rect 10128 2907 10186 2913
rect 10128 2904 10140 2907
rect 9548 2876 10140 2904
rect 9548 2864 9554 2876
rect 10128 2873 10140 2876
rect 10174 2904 10186 2907
rect 11146 2904 11152 2916
rect 10174 2876 11152 2904
rect 10174 2873 10186 2876
rect 10128 2867 10186 2873
rect 11146 2864 11152 2876
rect 11204 2864 11210 2916
rect 12452 2904 12480 2935
rect 12710 2932 12716 2935
rect 12768 2932 12774 2984
rect 15013 2975 15071 2981
rect 15013 2941 15025 2975
rect 15059 2941 15071 2975
rect 15013 2935 15071 2941
rect 15280 2975 15338 2981
rect 15280 2941 15292 2975
rect 15326 2972 15338 2975
rect 15654 2972 15660 2984
rect 15326 2944 15660 2972
rect 15326 2941 15338 2944
rect 15280 2935 15338 2941
rect 13538 2904 13544 2916
rect 12452 2876 13544 2904
rect 13538 2864 13544 2876
rect 13596 2904 13602 2916
rect 14829 2907 14887 2913
rect 14829 2904 14841 2907
rect 13596 2876 14841 2904
rect 13596 2864 13602 2876
rect 14829 2873 14841 2876
rect 14875 2904 14887 2907
rect 15028 2904 15056 2935
rect 15654 2932 15660 2944
rect 15712 2932 15718 2984
rect 17770 2932 17776 2984
rect 17828 2972 17834 2984
rect 18417 2975 18475 2981
rect 18417 2972 18429 2975
rect 17828 2944 18429 2972
rect 17828 2932 17834 2944
rect 18417 2941 18429 2944
rect 18463 2941 18475 2975
rect 19061 2975 19119 2981
rect 19061 2972 19073 2975
rect 18417 2935 18475 2941
rect 18616 2944 19073 2972
rect 14875 2876 15056 2904
rect 14875 2873 14887 2876
rect 14829 2867 14887 2873
rect 17954 2864 17960 2916
rect 18012 2904 18018 2916
rect 18616 2913 18644 2944
rect 19061 2941 19073 2944
rect 19107 2941 19119 2975
rect 19061 2935 19119 2941
rect 18601 2907 18659 2913
rect 18601 2904 18613 2907
rect 18012 2876 18613 2904
rect 18012 2864 18018 2876
rect 18601 2873 18613 2876
rect 18647 2873 18659 2907
rect 19812 2904 19840 3003
rect 26418 3000 26424 3052
rect 26476 3000 26482 3052
rect 26602 3000 26608 3052
rect 26660 3040 26666 3052
rect 26697 3043 26755 3049
rect 26697 3040 26709 3043
rect 26660 3012 26709 3040
rect 26660 3000 26666 3012
rect 26697 3009 26709 3012
rect 26743 3009 26755 3043
rect 26697 3003 26755 3009
rect 30374 3000 30380 3052
rect 30432 3040 30438 3052
rect 30745 3043 30803 3049
rect 30745 3040 30757 3043
rect 30432 3012 30757 3040
rect 30432 3000 30438 3012
rect 30745 3009 30757 3012
rect 30791 3040 30803 3043
rect 34624 3040 34652 3136
rect 36262 3108 36268 3120
rect 36223 3080 36268 3108
rect 36262 3068 36268 3080
rect 36320 3068 36326 3120
rect 40512 3049 40540 3136
rect 34885 3043 34943 3049
rect 34885 3040 34897 3043
rect 30791 3012 31800 3040
rect 34624 3012 34897 3040
rect 30791 3009 30803 3012
rect 30745 3003 30803 3009
rect 20070 2981 20076 2984
rect 20064 2972 20076 2981
rect 20031 2944 20076 2972
rect 20064 2935 20076 2944
rect 20070 2932 20076 2935
rect 20128 2932 20134 2984
rect 22465 2975 22523 2981
rect 22465 2972 22477 2975
rect 22112 2944 22477 2972
rect 20714 2904 20720 2916
rect 19812 2876 20720 2904
rect 18601 2867 18659 2873
rect 20714 2864 20720 2876
rect 20772 2864 20778 2916
rect 22112 2913 22140 2944
rect 22465 2941 22477 2944
rect 22511 2941 22523 2975
rect 22465 2935 22523 2941
rect 23750 2932 23756 2984
rect 23808 2972 23814 2984
rect 23928 2975 23986 2981
rect 23928 2972 23940 2975
rect 23808 2944 23940 2972
rect 23808 2932 23814 2944
rect 23928 2941 23940 2944
rect 23974 2972 23986 2975
rect 24854 2972 24860 2984
rect 23974 2944 24860 2972
rect 23974 2941 23986 2944
rect 23928 2935 23986 2941
rect 24854 2932 24860 2944
rect 24912 2932 24918 2984
rect 26436 2972 26464 3000
rect 26973 2975 27031 2981
rect 26973 2972 26985 2975
rect 26436 2944 26985 2972
rect 26973 2941 26985 2944
rect 27019 2972 27031 2975
rect 27246 2972 27252 2984
rect 27019 2944 27252 2972
rect 27019 2941 27031 2944
rect 26973 2935 27031 2941
rect 27246 2932 27252 2944
rect 27304 2932 27310 2984
rect 30009 2975 30067 2981
rect 30009 2941 30021 2975
rect 30055 2972 30067 2975
rect 30469 2975 30527 2981
rect 30469 2972 30481 2975
rect 30055 2944 30481 2972
rect 30055 2941 30067 2944
rect 30009 2935 30067 2941
rect 30469 2941 30481 2944
rect 30515 2972 30527 2975
rect 31478 2972 31484 2984
rect 30515 2944 31484 2972
rect 30515 2941 30527 2944
rect 30469 2935 30527 2941
rect 31478 2932 31484 2944
rect 31536 2932 31542 2984
rect 31665 2975 31723 2981
rect 31665 2941 31677 2975
rect 31711 2941 31723 2975
rect 31772 2972 31800 3012
rect 34885 3009 34897 3012
rect 34931 3040 34943 3043
rect 37369 3043 37427 3049
rect 37369 3040 37381 3043
rect 34931 3012 35020 3040
rect 34931 3009 34943 3012
rect 34885 3003 34943 3009
rect 31921 2975 31979 2981
rect 31921 2972 31933 2975
rect 31772 2944 31933 2972
rect 31665 2935 31723 2941
rect 31921 2941 31933 2944
rect 31967 2941 31979 2975
rect 34992 2972 35020 3012
rect 37292 3012 37381 3040
rect 34992 2944 35480 2972
rect 31921 2935 31979 2941
rect 22097 2907 22155 2913
rect 22097 2904 22109 2907
rect 21192 2876 22109 2904
rect 21192 2848 21220 2876
rect 22097 2873 22109 2876
rect 22143 2873 22155 2907
rect 22278 2904 22284 2916
rect 22239 2876 22284 2904
rect 22097 2867 22155 2873
rect 22278 2864 22284 2876
rect 22336 2904 22342 2916
rect 22925 2907 22983 2913
rect 22925 2904 22937 2907
rect 22336 2876 22937 2904
rect 22336 2864 22342 2876
rect 22925 2873 22937 2876
rect 22971 2873 22983 2907
rect 22925 2867 22983 2873
rect 29362 2864 29368 2916
rect 29420 2904 29426 2916
rect 31573 2907 31631 2913
rect 31573 2904 31585 2907
rect 29420 2876 31585 2904
rect 29420 2864 29426 2876
rect 31573 2873 31585 2876
rect 31619 2904 31631 2907
rect 31680 2904 31708 2935
rect 31754 2904 31760 2916
rect 31619 2876 31760 2904
rect 31619 2873 31631 2876
rect 31573 2867 31631 2873
rect 31754 2864 31760 2876
rect 31812 2864 31818 2916
rect 34238 2864 34244 2916
rect 34296 2904 34302 2916
rect 34333 2907 34391 2913
rect 34333 2904 34345 2907
rect 34296 2876 34345 2904
rect 34296 2864 34302 2876
rect 34333 2873 34345 2876
rect 34379 2904 34391 2907
rect 35152 2907 35210 2913
rect 35152 2904 35164 2907
rect 34379 2876 35164 2904
rect 34379 2873 34391 2876
rect 34333 2867 34391 2873
rect 35152 2873 35164 2876
rect 35198 2904 35210 2907
rect 35342 2904 35348 2916
rect 35198 2876 35348 2904
rect 35198 2873 35210 2876
rect 35152 2867 35210 2873
rect 35342 2864 35348 2876
rect 35400 2864 35406 2916
rect 35452 2904 35480 2944
rect 37292 2916 37320 3012
rect 37369 3009 37381 3012
rect 37415 3009 37427 3043
rect 37369 3003 37427 3009
rect 40497 3043 40555 3049
rect 40497 3009 40509 3043
rect 40543 3009 40555 3043
rect 40497 3003 40555 3009
rect 37458 2932 37464 2984
rect 37516 2972 37522 2984
rect 37625 2975 37683 2981
rect 37625 2972 37637 2975
rect 37516 2944 37637 2972
rect 37516 2932 37522 2944
rect 37625 2941 37637 2944
rect 37671 2941 37683 2975
rect 37625 2935 37683 2941
rect 37274 2904 37280 2916
rect 35452 2876 37280 2904
rect 37274 2864 37280 2876
rect 37332 2864 37338 2916
rect 40034 2864 40040 2916
rect 40092 2904 40098 2916
rect 40742 2907 40800 2913
rect 40742 2904 40754 2907
rect 40092 2876 40754 2904
rect 40092 2864 40098 2876
rect 40742 2873 40754 2876
rect 40788 2904 40800 2907
rect 41046 2904 41052 2916
rect 40788 2876 41052 2904
rect 40788 2873 40800 2876
rect 40742 2867 40800 2873
rect 41046 2864 41052 2876
rect 41104 2904 41110 2916
rect 41322 2904 41328 2916
rect 41104 2876 41328 2904
rect 41104 2864 41110 2876
rect 41322 2864 41328 2876
rect 41380 2864 41386 2916
rect 8754 2836 8760 2848
rect 7239 2808 7420 2836
rect 8715 2808 8760 2836
rect 7239 2805 7251 2808
rect 7193 2799 7251 2805
rect 8754 2796 8760 2808
rect 8812 2796 8818 2848
rect 9766 2836 9772 2848
rect 9727 2808 9772 2836
rect 9766 2796 9772 2808
rect 9824 2796 9830 2848
rect 13817 2839 13875 2845
rect 13817 2805 13829 2839
rect 13863 2836 13875 2839
rect 13906 2836 13912 2848
rect 13863 2808 13912 2836
rect 13863 2805 13875 2808
rect 13817 2799 13875 2805
rect 13906 2796 13912 2808
rect 13964 2796 13970 2848
rect 21174 2836 21180 2848
rect 21135 2808 21180 2836
rect 21174 2796 21180 2808
rect 21232 2796 21238 2848
rect 24762 2796 24768 2848
rect 24820 2836 24826 2848
rect 25041 2839 25099 2845
rect 25041 2836 25053 2839
rect 24820 2808 25053 2836
rect 24820 2796 24826 2808
rect 25041 2805 25053 2808
rect 25087 2805 25099 2839
rect 25590 2836 25596 2848
rect 25551 2808 25596 2836
rect 25041 2799 25099 2805
rect 25590 2796 25596 2808
rect 25648 2796 25654 2848
rect 26050 2796 26056 2848
rect 26108 2836 26114 2848
rect 26699 2839 26757 2845
rect 26699 2836 26711 2839
rect 26108 2808 26711 2836
rect 26108 2796 26114 2808
rect 26699 2805 26711 2808
rect 26745 2836 26757 2839
rect 26786 2836 26792 2848
rect 26745 2808 26792 2836
rect 26745 2805 26757 2808
rect 26699 2799 26757 2805
rect 26786 2796 26792 2808
rect 26844 2796 26850 2848
rect 30466 2796 30472 2848
rect 30524 2836 30530 2848
rect 30653 2839 30711 2845
rect 30653 2836 30665 2839
rect 30524 2808 30665 2836
rect 30524 2796 30530 2808
rect 30653 2805 30665 2808
rect 30699 2805 30711 2839
rect 30653 2799 30711 2805
rect 33045 2839 33103 2845
rect 33045 2805 33057 2839
rect 33091 2836 33103 2839
rect 33134 2836 33140 2848
rect 33091 2808 33140 2836
rect 33091 2805 33103 2808
rect 33045 2799 33103 2805
rect 33134 2796 33140 2808
rect 33192 2796 33198 2848
rect 38562 2796 38568 2848
rect 38620 2836 38626 2848
rect 38749 2839 38807 2845
rect 38749 2836 38761 2839
rect 38620 2808 38761 2836
rect 38620 2796 38626 2808
rect 38749 2805 38761 2808
rect 38795 2836 38807 2839
rect 39301 2839 39359 2845
rect 39301 2836 39313 2839
rect 38795 2808 39313 2836
rect 38795 2805 38807 2808
rect 38749 2799 38807 2805
rect 39301 2805 39313 2808
rect 39347 2805 39359 2839
rect 39301 2799 39359 2805
rect 1104 2746 48852 2768
rect 1104 2694 19606 2746
rect 19658 2694 19670 2746
rect 19722 2694 19734 2746
rect 19786 2694 19798 2746
rect 19850 2694 48852 2746
rect 1104 2672 48852 2694
rect 2869 2635 2927 2641
rect 2869 2601 2881 2635
rect 2915 2632 2927 2635
rect 2915 2604 3556 2632
rect 2915 2601 2927 2604
rect 2869 2595 2927 2601
rect 1670 2524 1676 2576
rect 1728 2573 1734 2576
rect 3528 2573 3556 2604
rect 5626 2592 5632 2644
rect 5684 2632 5690 2644
rect 5721 2635 5779 2641
rect 5721 2632 5733 2635
rect 5684 2604 5733 2632
rect 5684 2592 5690 2604
rect 5721 2601 5733 2604
rect 5767 2632 5779 2635
rect 6273 2635 6331 2641
rect 6273 2632 6285 2635
rect 5767 2604 6285 2632
rect 5767 2601 5779 2604
rect 5721 2595 5779 2601
rect 6273 2601 6285 2604
rect 6319 2601 6331 2635
rect 7098 2632 7104 2644
rect 7059 2604 7104 2632
rect 6273 2595 6331 2601
rect 7098 2592 7104 2604
rect 7156 2592 7162 2644
rect 7558 2632 7564 2644
rect 7519 2604 7564 2632
rect 7558 2592 7564 2604
rect 7616 2592 7622 2644
rect 7650 2592 7656 2644
rect 7708 2632 7714 2644
rect 7837 2635 7895 2641
rect 7837 2632 7849 2635
rect 7708 2604 7849 2632
rect 7708 2592 7714 2604
rect 7837 2601 7849 2604
rect 7883 2632 7895 2635
rect 8573 2635 8631 2641
rect 8573 2632 8585 2635
rect 7883 2604 8585 2632
rect 7883 2601 7895 2604
rect 7837 2595 7895 2601
rect 8573 2601 8585 2604
rect 8619 2632 8631 2635
rect 9033 2635 9091 2641
rect 9033 2632 9045 2635
rect 8619 2604 9045 2632
rect 8619 2601 8631 2604
rect 8573 2595 8631 2601
rect 9033 2601 9045 2604
rect 9079 2601 9091 2635
rect 11146 2632 11152 2644
rect 11107 2604 11152 2632
rect 9033 2595 9091 2601
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 12526 2592 12532 2644
rect 12584 2632 12590 2644
rect 12989 2635 13047 2641
rect 12989 2632 13001 2635
rect 12584 2604 13001 2632
rect 12584 2592 12590 2604
rect 12989 2601 13001 2604
rect 13035 2601 13047 2635
rect 12989 2595 13047 2601
rect 14461 2635 14519 2641
rect 14461 2601 14473 2635
rect 14507 2632 14519 2635
rect 15102 2632 15108 2644
rect 14507 2604 15108 2632
rect 14507 2601 14519 2604
rect 14461 2595 14519 2601
rect 15102 2592 15108 2604
rect 15160 2592 15166 2644
rect 17129 2635 17187 2641
rect 17129 2601 17141 2635
rect 17175 2632 17187 2635
rect 17310 2632 17316 2644
rect 17175 2604 17316 2632
rect 17175 2601 17187 2604
rect 17129 2595 17187 2601
rect 17310 2592 17316 2604
rect 17368 2592 17374 2644
rect 17773 2635 17831 2641
rect 17773 2601 17785 2635
rect 17819 2632 17831 2635
rect 17862 2632 17868 2644
rect 17819 2604 17868 2632
rect 17819 2601 17831 2604
rect 17773 2595 17831 2601
rect 17862 2592 17868 2604
rect 17920 2592 17926 2644
rect 18046 2632 18052 2644
rect 18007 2604 18052 2632
rect 18046 2592 18052 2604
rect 18104 2592 18110 2644
rect 19981 2635 20039 2641
rect 19981 2601 19993 2635
rect 20027 2632 20039 2635
rect 20070 2632 20076 2644
rect 20027 2604 20076 2632
rect 20027 2601 20039 2604
rect 19981 2595 20039 2601
rect 20070 2592 20076 2604
rect 20128 2592 20134 2644
rect 20625 2635 20683 2641
rect 20625 2601 20637 2635
rect 20671 2632 20683 2635
rect 21174 2632 21180 2644
rect 20671 2604 21180 2632
rect 20671 2601 20683 2604
rect 20625 2595 20683 2601
rect 21174 2592 21180 2604
rect 21232 2592 21238 2644
rect 22830 2632 22836 2644
rect 22791 2604 22836 2632
rect 22830 2592 22836 2604
rect 22888 2592 22894 2644
rect 23474 2632 23480 2644
rect 23435 2604 23480 2632
rect 23474 2592 23480 2604
rect 23532 2592 23538 2644
rect 23658 2592 23664 2644
rect 23716 2632 23722 2644
rect 23753 2635 23811 2641
rect 23753 2632 23765 2635
rect 23716 2604 23765 2632
rect 23716 2592 23722 2604
rect 23753 2601 23765 2604
rect 23799 2601 23811 2635
rect 25682 2632 25688 2644
rect 25643 2604 25688 2632
rect 23753 2595 23811 2601
rect 25682 2592 25688 2604
rect 25740 2592 25746 2644
rect 26326 2592 26332 2644
rect 26384 2632 26390 2644
rect 26513 2635 26571 2641
rect 26513 2632 26525 2635
rect 26384 2604 26525 2632
rect 26384 2592 26390 2604
rect 26513 2601 26525 2604
rect 26559 2601 26571 2635
rect 27893 2635 27951 2641
rect 27893 2632 27905 2635
rect 26513 2595 26571 2601
rect 27264 2604 27905 2632
rect 1728 2567 1792 2573
rect 1728 2533 1746 2567
rect 1780 2533 1792 2567
rect 1728 2527 1792 2533
rect 3513 2567 3571 2573
rect 3513 2533 3525 2567
rect 3559 2564 3571 2567
rect 4608 2567 4666 2573
rect 4608 2564 4620 2567
rect 3559 2536 4620 2564
rect 3559 2533 3571 2536
rect 3513 2527 3571 2533
rect 4608 2533 4620 2536
rect 4654 2564 4666 2567
rect 5074 2564 5080 2576
rect 4654 2536 5080 2564
rect 4654 2533 4666 2536
rect 4608 2527 4666 2533
rect 1728 2524 1734 2527
rect 5074 2524 5080 2536
rect 5132 2524 5138 2576
rect 1486 2496 1492 2508
rect 1447 2468 1492 2496
rect 1486 2456 1492 2468
rect 1544 2456 1550 2508
rect 2590 2456 2596 2508
rect 2648 2496 2654 2508
rect 3789 2499 3847 2505
rect 3789 2496 3801 2499
rect 2648 2468 3801 2496
rect 2648 2456 2654 2468
rect 3789 2465 3801 2468
rect 3835 2496 3847 2499
rect 4341 2499 4399 2505
rect 4341 2496 4353 2499
rect 3835 2468 4353 2496
rect 3835 2465 3847 2468
rect 3789 2459 3847 2465
rect 4341 2465 4353 2468
rect 4387 2496 4399 2499
rect 5350 2496 5356 2508
rect 4387 2468 5356 2496
rect 4387 2465 4399 2468
rect 4341 2459 4399 2465
rect 5350 2456 5356 2468
rect 5408 2456 5414 2508
rect 6917 2499 6975 2505
rect 6917 2465 6929 2499
rect 6963 2496 6975 2499
rect 7576 2496 7604 2592
rect 8389 2567 8447 2573
rect 8389 2533 8401 2567
rect 8435 2564 8447 2567
rect 8754 2564 8760 2576
rect 8435 2536 8760 2564
rect 8435 2533 8447 2536
rect 8389 2527 8447 2533
rect 6963 2468 7604 2496
rect 6963 2465 6975 2468
rect 6917 2459 6975 2465
rect 6733 2431 6791 2437
rect 6733 2397 6745 2431
rect 6779 2428 6791 2431
rect 8404 2428 8432 2527
rect 8754 2524 8760 2536
rect 8812 2564 8818 2576
rect 10036 2567 10094 2573
rect 10036 2564 10048 2567
rect 8812 2536 10048 2564
rect 8812 2524 8818 2536
rect 10036 2533 10048 2536
rect 10082 2564 10094 2567
rect 11701 2567 11759 2573
rect 11701 2564 11713 2567
rect 10082 2536 11713 2564
rect 10082 2533 10094 2536
rect 10036 2527 10094 2533
rect 11701 2533 11713 2536
rect 11747 2533 11759 2567
rect 11701 2527 11759 2533
rect 12437 2567 12495 2573
rect 12437 2533 12449 2567
rect 12483 2564 12495 2567
rect 12710 2564 12716 2576
rect 12483 2536 12716 2564
rect 12483 2533 12495 2536
rect 12437 2527 12495 2533
rect 12710 2524 12716 2536
rect 12768 2564 12774 2576
rect 12805 2567 12863 2573
rect 12805 2564 12817 2567
rect 12768 2536 12817 2564
rect 12768 2524 12774 2536
rect 12805 2533 12817 2536
rect 12851 2533 12863 2567
rect 12805 2527 12863 2533
rect 14185 2567 14243 2573
rect 14185 2533 14197 2567
rect 14231 2564 14243 2567
rect 16482 2564 16488 2576
rect 14231 2536 15240 2564
rect 14231 2533 14243 2536
rect 14185 2527 14243 2533
rect 8478 2456 8484 2508
rect 8536 2496 8542 2508
rect 8665 2499 8723 2505
rect 8665 2496 8677 2499
rect 8536 2468 8677 2496
rect 8536 2456 8542 2468
rect 8665 2465 8677 2468
rect 8711 2496 8723 2499
rect 9582 2496 9588 2508
rect 8711 2468 9588 2496
rect 8711 2465 8723 2468
rect 8665 2459 8723 2465
rect 9582 2456 9588 2468
rect 9640 2456 9646 2508
rect 11422 2456 11428 2508
rect 11480 2496 11486 2508
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 11480 2468 12633 2496
rect 11480 2456 11486 2468
rect 12621 2465 12633 2468
rect 12667 2465 12679 2499
rect 12621 2459 12679 2465
rect 14277 2499 14335 2505
rect 14277 2465 14289 2499
rect 14323 2496 14335 2499
rect 14323 2468 14964 2496
rect 14323 2465 14335 2468
rect 14277 2459 14335 2465
rect 6779 2400 8432 2428
rect 9493 2431 9551 2437
rect 6779 2397 6791 2400
rect 6733 2391 6791 2397
rect 9493 2397 9505 2431
rect 9539 2428 9551 2431
rect 9766 2428 9772 2440
rect 9539 2400 9772 2428
rect 9539 2397 9551 2400
rect 9493 2391 9551 2397
rect 9766 2388 9772 2400
rect 9824 2388 9830 2440
rect 12636 2428 12664 2459
rect 13265 2431 13323 2437
rect 13265 2428 13277 2431
rect 12636 2400 13277 2428
rect 13265 2397 13277 2400
rect 13311 2397 13323 2431
rect 13265 2391 13323 2397
rect 8113 2363 8171 2369
rect 8113 2329 8125 2363
rect 8159 2360 8171 2363
rect 8202 2360 8208 2372
rect 8159 2332 8208 2360
rect 8159 2329 8171 2332
rect 8113 2323 8171 2329
rect 8202 2320 8208 2332
rect 8260 2320 8266 2372
rect 7742 2252 7748 2304
rect 7800 2292 7806 2304
rect 8754 2292 8760 2304
rect 7800 2264 8760 2292
rect 7800 2252 7806 2264
rect 8754 2252 8760 2264
rect 8812 2252 8818 2304
rect 14936 2301 14964 2468
rect 15212 2428 15240 2536
rect 15764 2536 16488 2564
rect 15764 2505 15792 2536
rect 16482 2524 16488 2536
rect 16540 2524 16546 2576
rect 17880 2564 17908 2592
rect 18846 2567 18904 2573
rect 18846 2564 18858 2567
rect 17880 2536 18858 2564
rect 18846 2533 18858 2536
rect 18892 2533 18904 2567
rect 18846 2527 18904 2533
rect 20714 2524 20720 2576
rect 20772 2564 20778 2576
rect 20901 2567 20959 2573
rect 20901 2564 20913 2567
rect 20772 2536 20913 2564
rect 20772 2524 20778 2536
rect 20901 2533 20913 2536
rect 20947 2533 20959 2567
rect 21192 2564 21220 2592
rect 21698 2567 21756 2573
rect 21698 2564 21710 2567
rect 21192 2536 21710 2564
rect 20901 2527 20959 2533
rect 21698 2533 21710 2536
rect 21744 2533 21756 2567
rect 23492 2564 23520 2592
rect 27264 2576 27292 2604
rect 27893 2601 27905 2604
rect 27939 2601 27951 2635
rect 27893 2595 27951 2601
rect 29362 2592 29368 2644
rect 29420 2632 29426 2644
rect 29457 2635 29515 2641
rect 29457 2632 29469 2635
rect 29420 2604 29469 2632
rect 29420 2592 29426 2604
rect 29457 2601 29469 2604
rect 29503 2601 29515 2635
rect 29457 2595 29515 2601
rect 24550 2567 24608 2573
rect 24550 2564 24562 2567
rect 23492 2536 24562 2564
rect 21698 2527 21756 2533
rect 24550 2533 24562 2536
rect 24596 2564 24608 2567
rect 24762 2564 24768 2576
rect 24596 2536 24768 2564
rect 24596 2533 24608 2536
rect 24550 2527 24608 2533
rect 15289 2499 15347 2505
rect 15289 2465 15301 2499
rect 15335 2496 15347 2499
rect 15749 2499 15807 2505
rect 15749 2496 15761 2499
rect 15335 2468 15761 2496
rect 15335 2465 15347 2468
rect 15289 2459 15347 2465
rect 15749 2465 15761 2468
rect 15795 2465 15807 2499
rect 16005 2499 16063 2505
rect 16005 2496 16017 2499
rect 15749 2459 15807 2465
rect 15856 2468 16017 2496
rect 15856 2428 15884 2468
rect 16005 2465 16017 2468
rect 16051 2496 16063 2499
rect 16390 2496 16396 2508
rect 16051 2468 16396 2496
rect 16051 2465 16063 2468
rect 16005 2459 16063 2465
rect 16390 2456 16396 2468
rect 16448 2456 16454 2508
rect 18046 2456 18052 2508
rect 18104 2496 18110 2508
rect 18601 2499 18659 2505
rect 18601 2496 18613 2499
rect 18104 2468 18613 2496
rect 18104 2456 18110 2468
rect 18601 2465 18613 2468
rect 18647 2465 18659 2499
rect 20916 2496 20944 2527
rect 24762 2524 24768 2536
rect 24820 2524 24826 2576
rect 27246 2564 27252 2576
rect 27207 2536 27252 2564
rect 27246 2524 27252 2536
rect 27304 2524 27310 2576
rect 27433 2567 27491 2573
rect 27433 2533 27445 2567
rect 27479 2564 27491 2567
rect 27614 2564 27620 2576
rect 27479 2536 27620 2564
rect 27479 2533 27491 2536
rect 27433 2527 27491 2533
rect 27614 2524 27620 2536
rect 27672 2564 27678 2576
rect 28261 2567 28319 2573
rect 28261 2564 28273 2567
rect 27672 2536 28273 2564
rect 27672 2524 27678 2536
rect 28261 2533 28273 2536
rect 28307 2533 28319 2567
rect 28261 2527 28319 2533
rect 21453 2499 21511 2505
rect 21453 2496 21465 2499
rect 20916 2468 21465 2496
rect 18601 2459 18659 2465
rect 21453 2465 21465 2468
rect 21499 2465 21511 2499
rect 21453 2459 21511 2465
rect 23658 2456 23664 2508
rect 23716 2496 23722 2508
rect 24305 2499 24363 2505
rect 24305 2496 24317 2499
rect 23716 2468 24317 2496
rect 23716 2456 23722 2468
rect 24305 2465 24317 2468
rect 24351 2465 24363 2499
rect 24305 2459 24363 2465
rect 27525 2499 27583 2505
rect 27525 2465 27537 2499
rect 27571 2496 27583 2499
rect 27706 2496 27712 2508
rect 27571 2468 27712 2496
rect 27571 2465 27583 2468
rect 27525 2459 27583 2465
rect 27706 2456 27712 2468
rect 27764 2456 27770 2508
rect 28442 2496 28448 2508
rect 28403 2468 28448 2496
rect 28442 2456 28448 2468
rect 28500 2496 28506 2508
rect 28997 2499 29055 2505
rect 28997 2496 29009 2499
rect 28500 2468 29009 2496
rect 28500 2456 28506 2468
rect 28997 2465 29009 2468
rect 29043 2465 29055 2499
rect 29472 2496 29500 2595
rect 30374 2592 30380 2644
rect 30432 2632 30438 2644
rect 31113 2635 31171 2641
rect 31113 2632 31125 2635
rect 30432 2604 31125 2632
rect 30432 2592 30438 2604
rect 31113 2601 31125 2604
rect 31159 2601 31171 2635
rect 31754 2632 31760 2644
rect 31715 2604 31760 2632
rect 31113 2595 31171 2601
rect 31754 2592 31760 2604
rect 31812 2592 31818 2644
rect 32217 2635 32275 2641
rect 32217 2601 32229 2635
rect 32263 2632 32275 2635
rect 32674 2632 32680 2644
rect 32263 2604 32680 2632
rect 32263 2601 32275 2604
rect 32217 2595 32275 2601
rect 32674 2592 32680 2604
rect 32732 2592 32738 2644
rect 34238 2632 34244 2644
rect 34199 2604 34244 2632
rect 34238 2592 34244 2604
rect 34296 2592 34302 2644
rect 35161 2635 35219 2641
rect 35161 2601 35173 2635
rect 35207 2632 35219 2635
rect 35250 2632 35256 2644
rect 35207 2604 35256 2632
rect 35207 2601 35219 2604
rect 35161 2595 35219 2601
rect 35250 2592 35256 2604
rect 35308 2592 35314 2644
rect 37274 2592 37280 2644
rect 37332 2632 37338 2644
rect 37921 2635 37979 2641
rect 37921 2632 37933 2635
rect 37332 2604 37933 2632
rect 37332 2592 37338 2604
rect 37921 2601 37933 2604
rect 37967 2632 37979 2635
rect 38013 2635 38071 2641
rect 38013 2632 38025 2635
rect 37967 2604 38025 2632
rect 37967 2601 37979 2604
rect 37921 2595 37979 2601
rect 38013 2601 38025 2604
rect 38059 2601 38071 2635
rect 38013 2595 38071 2601
rect 39669 2635 39727 2641
rect 39669 2601 39681 2635
rect 39715 2632 39727 2635
rect 40034 2632 40040 2644
rect 39715 2604 40040 2632
rect 39715 2601 39727 2604
rect 39669 2595 39727 2601
rect 40034 2592 40040 2604
rect 40092 2592 40098 2644
rect 40402 2592 40408 2644
rect 40460 2632 40466 2644
rect 40497 2635 40555 2641
rect 40497 2632 40509 2635
rect 40460 2604 40509 2632
rect 40460 2592 40466 2604
rect 40497 2601 40509 2604
rect 40543 2601 40555 2635
rect 40497 2595 40555 2601
rect 29546 2524 29552 2576
rect 29604 2564 29610 2576
rect 29978 2567 30036 2573
rect 29978 2564 29990 2567
rect 29604 2536 29990 2564
rect 29604 2524 29610 2536
rect 29978 2533 29990 2536
rect 30024 2533 30036 2567
rect 29978 2527 30036 2533
rect 29733 2499 29791 2505
rect 29733 2496 29745 2499
rect 29472 2468 29745 2496
rect 28997 2459 29055 2465
rect 29733 2465 29745 2468
rect 29779 2465 29791 2499
rect 31772 2496 31800 2592
rect 33134 2573 33140 2576
rect 33128 2564 33140 2573
rect 33047 2536 33140 2564
rect 33128 2527 33140 2536
rect 33192 2564 33198 2576
rect 38562 2573 38568 2576
rect 36357 2567 36415 2573
rect 36357 2564 36369 2567
rect 33192 2536 36369 2564
rect 33134 2524 33140 2527
rect 33192 2524 33198 2536
rect 36357 2533 36369 2536
rect 36403 2533 36415 2567
rect 36357 2527 36415 2533
rect 37737 2567 37795 2573
rect 37737 2533 37749 2567
rect 37783 2564 37795 2567
rect 38534 2567 38568 2573
rect 38534 2564 38546 2567
rect 37783 2536 38546 2564
rect 37783 2533 37795 2536
rect 37737 2527 37795 2533
rect 38534 2533 38546 2536
rect 38620 2564 38626 2576
rect 38620 2536 38682 2564
rect 38534 2527 38568 2533
rect 38562 2524 38568 2527
rect 38620 2524 38626 2536
rect 32861 2499 32919 2505
rect 32861 2496 32873 2499
rect 31772 2468 32873 2496
rect 29733 2459 29791 2465
rect 32861 2465 32873 2468
rect 32907 2465 32919 2499
rect 32861 2459 32919 2465
rect 34514 2456 34520 2508
rect 34572 2496 34578 2508
rect 35437 2499 35495 2505
rect 35437 2496 35449 2499
rect 34572 2468 35449 2496
rect 34572 2456 34578 2468
rect 35437 2465 35449 2468
rect 35483 2496 35495 2499
rect 35989 2499 36047 2505
rect 35989 2496 36001 2499
rect 35483 2468 36001 2496
rect 35483 2465 35495 2468
rect 35437 2459 35495 2465
rect 35989 2465 36001 2468
rect 36035 2465 36047 2499
rect 36630 2496 36636 2508
rect 36591 2468 36636 2496
rect 35989 2459 36047 2465
rect 36630 2456 36636 2468
rect 36688 2496 36694 2508
rect 37090 2496 37096 2508
rect 36688 2468 37096 2496
rect 36688 2456 36694 2468
rect 37090 2456 37096 2468
rect 37148 2496 37154 2508
rect 37185 2499 37243 2505
rect 37185 2496 37197 2499
rect 37148 2468 37197 2496
rect 37148 2456 37154 2468
rect 37185 2465 37197 2468
rect 37231 2465 37243 2499
rect 37185 2459 37243 2465
rect 37921 2499 37979 2505
rect 37921 2465 37933 2499
rect 37967 2496 37979 2499
rect 38289 2499 38347 2505
rect 38289 2496 38301 2499
rect 37967 2468 38301 2496
rect 37967 2465 37979 2468
rect 37921 2459 37979 2465
rect 38289 2465 38301 2468
rect 38335 2465 38347 2499
rect 38289 2459 38347 2465
rect 15212 2400 15884 2428
rect 40512 2428 40540 2595
rect 40957 2567 41015 2573
rect 40957 2533 40969 2567
rect 41003 2564 41015 2567
rect 41693 2567 41751 2573
rect 41693 2564 41705 2567
rect 41003 2536 41705 2564
rect 41003 2533 41015 2536
rect 40957 2527 41015 2533
rect 41693 2533 41705 2536
rect 41739 2564 41751 2567
rect 42334 2564 42340 2576
rect 41739 2536 42340 2564
rect 41739 2533 41751 2536
rect 41693 2527 41751 2533
rect 42334 2524 42340 2536
rect 42392 2564 42398 2576
rect 42392 2536 44864 2564
rect 42392 2524 42398 2536
rect 41414 2456 41420 2508
rect 41472 2496 41478 2508
rect 41785 2499 41843 2505
rect 41785 2496 41797 2499
rect 41472 2468 41797 2496
rect 41472 2456 41478 2468
rect 41785 2465 41797 2468
rect 41831 2496 41843 2499
rect 42153 2499 42211 2505
rect 42153 2496 42165 2499
rect 41831 2468 42165 2496
rect 41831 2465 41843 2468
rect 41785 2459 41843 2465
rect 42153 2465 42165 2468
rect 42199 2465 42211 2499
rect 42153 2459 42211 2465
rect 42426 2456 42432 2508
rect 42484 2496 42490 2508
rect 42702 2496 42708 2508
rect 42484 2468 42708 2496
rect 42484 2456 42490 2468
rect 42702 2456 42708 2468
rect 42760 2496 42766 2508
rect 44836 2505 44864 2536
rect 43257 2499 43315 2505
rect 43257 2496 43269 2499
rect 42760 2468 43269 2496
rect 42760 2456 42766 2468
rect 43257 2465 43269 2468
rect 43303 2465 43315 2499
rect 43257 2459 43315 2465
rect 44821 2499 44879 2505
rect 44821 2465 44833 2499
rect 44867 2496 44879 2499
rect 45186 2496 45192 2508
rect 44867 2468 45192 2496
rect 44867 2465 44879 2468
rect 44821 2459 44879 2465
rect 45186 2456 45192 2468
rect 45244 2456 45250 2508
rect 41601 2431 41659 2437
rect 41601 2428 41613 2431
rect 40512 2400 41613 2428
rect 41601 2397 41613 2400
rect 41647 2397 41659 2431
rect 41601 2391 41659 2397
rect 26970 2360 26976 2372
rect 26931 2332 26976 2360
rect 26970 2320 26976 2332
rect 27028 2320 27034 2372
rect 27614 2320 27620 2372
rect 27672 2360 27678 2372
rect 28629 2363 28687 2369
rect 28629 2360 28641 2363
rect 27672 2332 28641 2360
rect 27672 2320 27678 2332
rect 28629 2329 28641 2332
rect 28675 2329 28687 2363
rect 28629 2323 28687 2329
rect 36817 2363 36875 2369
rect 36817 2329 36829 2363
rect 36863 2360 36875 2363
rect 38194 2360 38200 2372
rect 36863 2332 38200 2360
rect 36863 2329 36875 2332
rect 36817 2323 36875 2329
rect 38194 2320 38200 2332
rect 38252 2320 38258 2372
rect 40218 2320 40224 2372
rect 40276 2360 40282 2372
rect 41233 2363 41291 2369
rect 41233 2360 41245 2363
rect 40276 2332 41245 2360
rect 40276 2320 40282 2332
rect 41233 2329 41245 2332
rect 41279 2329 41291 2363
rect 41233 2323 41291 2329
rect 42889 2363 42947 2369
rect 42889 2329 42901 2363
rect 42935 2360 42947 2363
rect 43806 2360 43812 2372
rect 42935 2332 43812 2360
rect 42935 2329 42947 2332
rect 42889 2323 42947 2329
rect 43806 2320 43812 2332
rect 43864 2320 43870 2372
rect 45005 2363 45063 2369
rect 45005 2329 45017 2363
rect 45051 2360 45063 2363
rect 46474 2360 46480 2372
rect 45051 2332 46480 2360
rect 45051 2329 45063 2332
rect 45005 2323 45063 2329
rect 46474 2320 46480 2332
rect 46532 2320 46538 2372
rect 14921 2295 14979 2301
rect 14921 2261 14933 2295
rect 14967 2292 14979 2295
rect 15470 2292 15476 2304
rect 14967 2264 15476 2292
rect 14967 2261 14979 2264
rect 14921 2255 14979 2261
rect 15470 2252 15476 2264
rect 15528 2252 15534 2304
rect 35621 2295 35679 2301
rect 35621 2261 35633 2295
rect 35667 2292 35679 2295
rect 35710 2292 35716 2304
rect 35667 2264 35716 2292
rect 35667 2261 35679 2264
rect 35621 2255 35679 2261
rect 35710 2252 35716 2264
rect 35768 2252 35774 2304
rect 45186 2252 45192 2304
rect 45244 2292 45250 2304
rect 45373 2295 45431 2301
rect 45373 2292 45385 2295
rect 45244 2264 45385 2292
rect 45244 2252 45250 2264
rect 45373 2261 45385 2264
rect 45419 2261 45431 2295
rect 45373 2255 45431 2261
rect 1104 2202 48852 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 34966 2202
rect 35018 2150 35030 2202
rect 35082 2150 35094 2202
rect 35146 2150 35158 2202
rect 35210 2150 48852 2202
rect 1104 2128 48852 2150
rect 4706 552 4712 604
rect 4764 592 4770 604
rect 4982 592 4988 604
rect 4764 564 4988 592
rect 4764 552 4770 564
rect 4982 552 4988 564
rect 5040 552 5046 604
<< via1 >>
rect 19606 47302 19658 47354
rect 19670 47302 19722 47354
rect 19734 47302 19786 47354
rect 19798 47302 19850 47354
rect 4246 46758 4298 46810
rect 4310 46758 4362 46810
rect 4374 46758 4426 46810
rect 4438 46758 4490 46810
rect 34966 46758 35018 46810
rect 35030 46758 35082 46810
rect 35094 46758 35146 46810
rect 35158 46758 35210 46810
rect 19606 46214 19658 46266
rect 19670 46214 19722 46266
rect 19734 46214 19786 46266
rect 19798 46214 19850 46266
rect 4246 45670 4298 45722
rect 4310 45670 4362 45722
rect 4374 45670 4426 45722
rect 4438 45670 4490 45722
rect 34966 45670 35018 45722
rect 35030 45670 35082 45722
rect 35094 45670 35146 45722
rect 35158 45670 35210 45722
rect 46940 45543 46992 45552
rect 46940 45509 46949 45543
rect 46949 45509 46983 45543
rect 46983 45509 46992 45543
rect 46940 45500 46992 45509
rect 46756 45407 46808 45416
rect 46756 45373 46765 45407
rect 46765 45373 46799 45407
rect 46799 45373 46808 45407
rect 46756 45364 46808 45373
rect 19606 45126 19658 45178
rect 19670 45126 19722 45178
rect 19734 45126 19786 45178
rect 19798 45126 19850 45178
rect 4246 44582 4298 44634
rect 4310 44582 4362 44634
rect 4374 44582 4426 44634
rect 4438 44582 4490 44634
rect 34966 44582 35018 44634
rect 35030 44582 35082 44634
rect 35094 44582 35146 44634
rect 35158 44582 35210 44634
rect 46940 44523 46992 44532
rect 46940 44489 46949 44523
rect 46949 44489 46983 44523
rect 46983 44489 46992 44523
rect 46940 44480 46992 44489
rect 47400 44523 47452 44532
rect 47400 44489 47409 44523
rect 47409 44489 47443 44523
rect 47443 44489 47452 44523
rect 47400 44480 47452 44489
rect 46112 44276 46164 44328
rect 47400 44276 47452 44328
rect 19606 44038 19658 44090
rect 19670 44038 19722 44090
rect 19734 44038 19786 44090
rect 19798 44038 19850 44090
rect 4246 43494 4298 43546
rect 4310 43494 4362 43546
rect 4374 43494 4426 43546
rect 4438 43494 4490 43546
rect 34966 43494 35018 43546
rect 35030 43494 35082 43546
rect 35094 43494 35146 43546
rect 35158 43494 35210 43546
rect 19606 42950 19658 43002
rect 19670 42950 19722 43002
rect 19734 42950 19786 43002
rect 19798 42950 19850 43002
rect 4246 42406 4298 42458
rect 4310 42406 4362 42458
rect 4374 42406 4426 42458
rect 4438 42406 4490 42458
rect 34966 42406 35018 42458
rect 35030 42406 35082 42458
rect 35094 42406 35146 42458
rect 35158 42406 35210 42458
rect 19606 41862 19658 41914
rect 19670 41862 19722 41914
rect 19734 41862 19786 41914
rect 19798 41862 19850 41914
rect 46940 41803 46992 41812
rect 46940 41769 46949 41803
rect 46949 41769 46983 41803
rect 46983 41769 46992 41803
rect 46940 41760 46992 41769
rect 46756 41667 46808 41676
rect 46756 41633 46765 41667
rect 46765 41633 46799 41667
rect 46799 41633 46808 41667
rect 46756 41624 46808 41633
rect 4246 41318 4298 41370
rect 4310 41318 4362 41370
rect 4374 41318 4426 41370
rect 4438 41318 4490 41370
rect 34966 41318 35018 41370
rect 35030 41318 35082 41370
rect 35094 41318 35146 41370
rect 35158 41318 35210 41370
rect 46756 40919 46808 40928
rect 46756 40885 46765 40919
rect 46765 40885 46799 40919
rect 46799 40885 46808 40919
rect 46756 40876 46808 40885
rect 19606 40774 19658 40826
rect 19670 40774 19722 40826
rect 19734 40774 19786 40826
rect 19798 40774 19850 40826
rect 4246 40230 4298 40282
rect 4310 40230 4362 40282
rect 4374 40230 4426 40282
rect 4438 40230 4490 40282
rect 34966 40230 35018 40282
rect 35030 40230 35082 40282
rect 35094 40230 35146 40282
rect 35158 40230 35210 40282
rect 46296 40060 46348 40112
rect 46756 40060 46808 40112
rect 19606 39686 19658 39738
rect 19670 39686 19722 39738
rect 19734 39686 19786 39738
rect 19798 39686 19850 39738
rect 4246 39142 4298 39194
rect 4310 39142 4362 39194
rect 4374 39142 4426 39194
rect 4438 39142 4490 39194
rect 34966 39142 35018 39194
rect 35030 39142 35082 39194
rect 35094 39142 35146 39194
rect 35158 39142 35210 39194
rect 19606 38598 19658 38650
rect 19670 38598 19722 38650
rect 19734 38598 19786 38650
rect 19798 38598 19850 38650
rect 46940 38539 46992 38548
rect 46940 38505 46949 38539
rect 46949 38505 46983 38539
rect 46983 38505 46992 38539
rect 46940 38496 46992 38505
rect 46756 38403 46808 38412
rect 46756 38369 46765 38403
rect 46765 38369 46799 38403
rect 46799 38369 46808 38403
rect 46756 38360 46808 38369
rect 4246 38054 4298 38106
rect 4310 38054 4362 38106
rect 4374 38054 4426 38106
rect 4438 38054 4490 38106
rect 34966 38054 35018 38106
rect 35030 38054 35082 38106
rect 35094 38054 35146 38106
rect 35158 38054 35210 38106
rect 45652 37612 45704 37664
rect 46756 37655 46808 37664
rect 46756 37621 46765 37655
rect 46765 37621 46799 37655
rect 46799 37621 46808 37655
rect 46756 37612 46808 37621
rect 19606 37510 19658 37562
rect 19670 37510 19722 37562
rect 19734 37510 19786 37562
rect 19798 37510 19850 37562
rect 4246 36966 4298 37018
rect 4310 36966 4362 37018
rect 4374 36966 4426 37018
rect 4438 36966 4490 37018
rect 34966 36966 35018 37018
rect 35030 36966 35082 37018
rect 35094 36966 35146 37018
rect 35158 36966 35210 37018
rect 19606 36422 19658 36474
rect 19670 36422 19722 36474
rect 19734 36422 19786 36474
rect 19798 36422 19850 36474
rect 4246 35878 4298 35930
rect 4310 35878 4362 35930
rect 4374 35878 4426 35930
rect 4438 35878 4490 35930
rect 34966 35878 35018 35930
rect 35030 35878 35082 35930
rect 35094 35878 35146 35930
rect 35158 35878 35210 35930
rect 19606 35334 19658 35386
rect 19670 35334 19722 35386
rect 19734 35334 19786 35386
rect 19798 35334 19850 35386
rect 46940 35275 46992 35284
rect 46940 35241 46949 35275
rect 46949 35241 46983 35275
rect 46983 35241 46992 35275
rect 46940 35232 46992 35241
rect 46756 35139 46808 35148
rect 46756 35105 46765 35139
rect 46765 35105 46799 35139
rect 46799 35105 46808 35139
rect 46756 35096 46808 35105
rect 4246 34790 4298 34842
rect 4310 34790 4362 34842
rect 4374 34790 4426 34842
rect 4438 34790 4490 34842
rect 34966 34790 35018 34842
rect 35030 34790 35082 34842
rect 35094 34790 35146 34842
rect 35158 34790 35210 34842
rect 46756 34731 46808 34740
rect 46756 34697 46765 34731
rect 46765 34697 46799 34731
rect 46799 34697 46808 34731
rect 46756 34688 46808 34697
rect 19606 34246 19658 34298
rect 19670 34246 19722 34298
rect 19734 34246 19786 34298
rect 19798 34246 19850 34298
rect 4246 33702 4298 33754
rect 4310 33702 4362 33754
rect 4374 33702 4426 33754
rect 4438 33702 4490 33754
rect 34966 33702 35018 33754
rect 35030 33702 35082 33754
rect 35094 33702 35146 33754
rect 35158 33702 35210 33754
rect 19606 33158 19658 33210
rect 19670 33158 19722 33210
rect 19734 33158 19786 33210
rect 19798 33158 19850 33210
rect 4246 32614 4298 32666
rect 4310 32614 4362 32666
rect 4374 32614 4426 32666
rect 4438 32614 4490 32666
rect 34966 32614 35018 32666
rect 35030 32614 35082 32666
rect 35094 32614 35146 32666
rect 35158 32614 35210 32666
rect 19606 32070 19658 32122
rect 19670 32070 19722 32122
rect 19734 32070 19786 32122
rect 19798 32070 19850 32122
rect 46940 32011 46992 32020
rect 46940 31977 46949 32011
rect 46949 31977 46983 32011
rect 46983 31977 46992 32011
rect 46940 31968 46992 31977
rect 46756 31875 46808 31884
rect 46756 31841 46765 31875
rect 46765 31841 46799 31875
rect 46799 31841 46808 31875
rect 46756 31832 46808 31841
rect 42340 31628 42392 31680
rect 4246 31526 4298 31578
rect 4310 31526 4362 31578
rect 4374 31526 4426 31578
rect 4438 31526 4490 31578
rect 34966 31526 35018 31578
rect 35030 31526 35082 31578
rect 35094 31526 35146 31578
rect 35158 31526 35210 31578
rect 42616 31220 42668 31272
rect 42340 31195 42392 31204
rect 42340 31161 42374 31195
rect 42374 31161 42392 31195
rect 42340 31152 42392 31161
rect 43444 31127 43496 31136
rect 43444 31093 43453 31127
rect 43453 31093 43487 31127
rect 43487 31093 43496 31127
rect 43444 31084 43496 31093
rect 46756 31127 46808 31136
rect 46756 31093 46765 31127
rect 46765 31093 46799 31127
rect 46799 31093 46808 31127
rect 46756 31084 46808 31093
rect 19606 30982 19658 31034
rect 19670 30982 19722 31034
rect 19734 30982 19786 31034
rect 19798 30982 19850 31034
rect 42340 30880 42392 30932
rect 42064 30855 42116 30864
rect 42064 30821 42073 30855
rect 42073 30821 42107 30855
rect 42107 30821 42116 30855
rect 42064 30812 42116 30821
rect 41880 30744 41932 30796
rect 43628 30787 43680 30796
rect 43628 30753 43662 30787
rect 43662 30753 43680 30787
rect 43628 30744 43680 30753
rect 45560 30744 45612 30796
rect 42340 30719 42392 30728
rect 42340 30685 42349 30719
rect 42349 30685 42383 30719
rect 42383 30685 42392 30719
rect 42340 30676 42392 30685
rect 42616 30676 42668 30728
rect 43352 30719 43404 30728
rect 43352 30685 43361 30719
rect 43361 30685 43395 30719
rect 43395 30685 43404 30719
rect 43352 30676 43404 30685
rect 45836 30719 45888 30728
rect 45836 30685 45845 30719
rect 45845 30685 45879 30719
rect 45879 30685 45888 30719
rect 45836 30676 45888 30685
rect 47216 30651 47268 30660
rect 47216 30617 47225 30651
rect 47225 30617 47259 30651
rect 47259 30617 47268 30651
rect 47216 30608 47268 30617
rect 41788 30583 41840 30592
rect 41788 30549 41797 30583
rect 41797 30549 41831 30583
rect 41831 30549 41840 30583
rect 41788 30540 41840 30549
rect 46204 30540 46256 30592
rect 4246 30438 4298 30490
rect 4310 30438 4362 30490
rect 4374 30438 4426 30490
rect 4438 30438 4490 30490
rect 34966 30438 35018 30490
rect 35030 30438 35082 30490
rect 35094 30438 35146 30490
rect 35158 30438 35210 30490
rect 41880 30336 41932 30388
rect 42064 30379 42116 30388
rect 42064 30345 42073 30379
rect 42073 30345 42107 30379
rect 42107 30345 42116 30379
rect 42064 30336 42116 30345
rect 42616 30379 42668 30388
rect 42616 30345 42625 30379
rect 42625 30345 42659 30379
rect 42659 30345 42668 30379
rect 42616 30336 42668 30345
rect 45928 30336 45980 30388
rect 46756 30336 46808 30388
rect 41696 30200 41748 30252
rect 45560 30268 45612 30320
rect 42800 30132 42852 30184
rect 43444 30132 43496 30184
rect 45836 30132 45888 30184
rect 46204 30132 46256 30184
rect 41420 30039 41472 30048
rect 41420 30005 41429 30039
rect 41429 30005 41463 30039
rect 41463 30005 41472 30039
rect 44088 30039 44140 30048
rect 41420 29996 41472 30005
rect 44088 30005 44097 30039
rect 44097 30005 44131 30039
rect 44131 30005 44140 30039
rect 44088 29996 44140 30005
rect 45192 29996 45244 30048
rect 45836 30039 45888 30048
rect 45836 30005 45845 30039
rect 45845 30005 45879 30039
rect 45879 30005 45888 30039
rect 45836 29996 45888 30005
rect 47492 30039 47544 30048
rect 47492 30005 47501 30039
rect 47501 30005 47535 30039
rect 47535 30005 47544 30039
rect 47492 29996 47544 30005
rect 19606 29894 19658 29946
rect 19670 29894 19722 29946
rect 19734 29894 19786 29946
rect 19798 29894 19850 29946
rect 41880 29792 41932 29844
rect 42800 29835 42852 29844
rect 42800 29801 42809 29835
rect 42809 29801 42843 29835
rect 42843 29801 42852 29835
rect 42800 29792 42852 29801
rect 43352 29792 43404 29844
rect 43628 29792 43680 29844
rect 45008 29792 45060 29844
rect 45560 29792 45612 29844
rect 39580 29724 39632 29776
rect 42432 29724 42484 29776
rect 44088 29724 44140 29776
rect 45836 29724 45888 29776
rect 47492 29724 47544 29776
rect 43352 29656 43404 29708
rect 45192 29699 45244 29708
rect 45192 29665 45201 29699
rect 45201 29665 45235 29699
rect 45235 29665 45244 29699
rect 45192 29656 45244 29665
rect 39028 29588 39080 29640
rect 41420 29588 41472 29640
rect 42064 29588 42116 29640
rect 42340 29631 42392 29640
rect 42340 29597 42349 29631
rect 42349 29597 42383 29631
rect 42383 29597 42392 29631
rect 42340 29588 42392 29597
rect 40224 29452 40276 29504
rect 42340 29452 42392 29504
rect 4246 29350 4298 29402
rect 4310 29350 4362 29402
rect 4374 29350 4426 29402
rect 4438 29350 4490 29402
rect 34966 29350 35018 29402
rect 35030 29350 35082 29402
rect 35094 29350 35146 29402
rect 35158 29350 35210 29402
rect 39580 29291 39632 29300
rect 39580 29257 39589 29291
rect 39589 29257 39623 29291
rect 39623 29257 39632 29291
rect 39580 29248 39632 29257
rect 41880 29248 41932 29300
rect 42064 29248 42116 29300
rect 45100 29248 45152 29300
rect 45192 29248 45244 29300
rect 45560 29248 45612 29300
rect 45836 29291 45888 29300
rect 45836 29257 45845 29291
rect 45845 29257 45879 29291
rect 45879 29257 45888 29291
rect 45836 29248 45888 29257
rect 46940 29291 46992 29300
rect 46940 29257 46949 29291
rect 46949 29257 46983 29291
rect 46983 29257 46992 29291
rect 46940 29248 46992 29257
rect 41328 29180 41380 29232
rect 42892 29180 42944 29232
rect 44916 29180 44968 29232
rect 41236 29112 41288 29164
rect 40224 29044 40276 29096
rect 39396 28976 39448 29028
rect 40316 28976 40368 29028
rect 41236 28976 41288 29028
rect 42340 29044 42392 29096
rect 42800 29112 42852 29164
rect 45008 29155 45060 29164
rect 45008 29121 45017 29155
rect 45017 29121 45051 29155
rect 45051 29121 45060 29155
rect 45008 29112 45060 29121
rect 41696 28976 41748 29028
rect 41788 28976 41840 29028
rect 45836 29044 45888 29096
rect 39028 28908 39080 28960
rect 39212 28908 39264 28960
rect 40224 28951 40276 28960
rect 40224 28917 40233 28951
rect 40233 28917 40267 28951
rect 40267 28917 40276 28951
rect 40224 28908 40276 28917
rect 45100 29019 45152 29028
rect 45100 28985 45109 29019
rect 45109 28985 45143 29019
rect 45143 28985 45152 29019
rect 45100 28976 45152 28985
rect 45468 28976 45520 29028
rect 45744 28976 45796 29028
rect 47308 29019 47360 29028
rect 47308 28985 47317 29019
rect 47317 28985 47351 29019
rect 47351 28985 47360 29019
rect 47308 28976 47360 28985
rect 45192 28908 45244 28960
rect 19606 28806 19658 28858
rect 19670 28806 19722 28858
rect 19734 28806 19786 28858
rect 19798 28806 19850 28858
rect 40316 28747 40368 28756
rect 40316 28713 40325 28747
rect 40325 28713 40359 28747
rect 40359 28713 40368 28747
rect 40316 28704 40368 28713
rect 41236 28747 41288 28756
rect 41236 28713 41245 28747
rect 41245 28713 41279 28747
rect 41279 28713 41288 28747
rect 41236 28704 41288 28713
rect 42432 28747 42484 28756
rect 42432 28713 42441 28747
rect 42441 28713 42475 28747
rect 42475 28713 42484 28747
rect 42432 28704 42484 28713
rect 42800 28747 42852 28756
rect 42800 28713 42809 28747
rect 42809 28713 42843 28747
rect 42843 28713 42852 28747
rect 42800 28704 42852 28713
rect 41972 28679 42024 28688
rect 41972 28645 41981 28679
rect 41981 28645 42015 28679
rect 42015 28645 42024 28679
rect 41972 28636 42024 28645
rect 45100 28679 45152 28688
rect 45100 28645 45109 28679
rect 45109 28645 45143 28679
rect 45143 28645 45152 28679
rect 45100 28636 45152 28645
rect 39028 28568 39080 28620
rect 39212 28611 39264 28620
rect 39212 28577 39246 28611
rect 39246 28577 39264 28611
rect 39212 28568 39264 28577
rect 42064 28611 42116 28620
rect 42064 28577 42073 28611
rect 42073 28577 42107 28611
rect 42107 28577 42116 28611
rect 42064 28568 42116 28577
rect 42892 28568 42944 28620
rect 43996 28568 44048 28620
rect 44916 28611 44968 28620
rect 44916 28577 44925 28611
rect 44925 28577 44959 28611
rect 44959 28577 44968 28611
rect 44916 28568 44968 28577
rect 45560 28568 45612 28620
rect 46388 28611 46440 28620
rect 46388 28577 46422 28611
rect 46422 28577 46440 28611
rect 46388 28568 46440 28577
rect 41880 28543 41932 28552
rect 41880 28509 41889 28543
rect 41889 28509 41923 28543
rect 41923 28509 41932 28543
rect 41880 28500 41932 28509
rect 45192 28543 45244 28552
rect 45192 28509 45201 28543
rect 45201 28509 45235 28543
rect 45235 28509 45244 28543
rect 45192 28500 45244 28509
rect 40316 28432 40368 28484
rect 45744 28432 45796 28484
rect 41512 28407 41564 28416
rect 41512 28373 41521 28407
rect 41521 28373 41555 28407
rect 41555 28373 41564 28407
rect 41512 28364 41564 28373
rect 43536 28407 43588 28416
rect 43536 28373 43545 28407
rect 43545 28373 43579 28407
rect 43579 28373 43588 28407
rect 43536 28364 43588 28373
rect 44640 28407 44692 28416
rect 44640 28373 44649 28407
rect 44649 28373 44683 28407
rect 44683 28373 44692 28407
rect 44640 28364 44692 28373
rect 47492 28407 47544 28416
rect 47492 28373 47501 28407
rect 47501 28373 47535 28407
rect 47535 28373 47544 28407
rect 47492 28364 47544 28373
rect 4246 28262 4298 28314
rect 4310 28262 4362 28314
rect 4374 28262 4426 28314
rect 4438 28262 4490 28314
rect 34966 28262 35018 28314
rect 35030 28262 35082 28314
rect 35094 28262 35146 28314
rect 35158 28262 35210 28314
rect 39212 28160 39264 28212
rect 43996 28203 44048 28212
rect 43996 28169 44005 28203
rect 44005 28169 44039 28203
rect 44039 28169 44048 28203
rect 43996 28160 44048 28169
rect 45100 28160 45152 28212
rect 42892 28092 42944 28144
rect 43168 28024 43220 28076
rect 45560 28092 45612 28144
rect 46204 28024 46256 28076
rect 47492 28067 47544 28076
rect 47492 28033 47501 28067
rect 47501 28033 47535 28067
rect 47535 28033 47544 28067
rect 47492 28024 47544 28033
rect 39120 27956 39172 28008
rect 41144 27956 41196 28008
rect 44548 27999 44600 28008
rect 44548 27965 44557 27999
rect 44557 27965 44591 27999
rect 44591 27965 44600 27999
rect 44548 27956 44600 27965
rect 46388 27956 46440 28008
rect 43536 27931 43588 27940
rect 43536 27897 43545 27931
rect 43545 27897 43579 27931
rect 43579 27897 43588 27931
rect 43536 27888 43588 27897
rect 39120 27820 39172 27872
rect 39948 27863 40000 27872
rect 39948 27829 39957 27863
rect 39957 27829 39991 27863
rect 39991 27829 40000 27863
rect 39948 27820 40000 27829
rect 41880 27863 41932 27872
rect 41880 27829 41889 27863
rect 41889 27829 41923 27863
rect 41923 27829 41932 27863
rect 41880 27820 41932 27829
rect 42800 27820 42852 27872
rect 44088 27888 44140 27940
rect 46940 27956 46992 28008
rect 45468 27820 45520 27872
rect 47400 27888 47452 27940
rect 19606 27718 19658 27770
rect 19670 27718 19722 27770
rect 19734 27718 19786 27770
rect 19798 27718 19850 27770
rect 39948 27616 40000 27668
rect 41972 27616 42024 27668
rect 42800 27616 42852 27668
rect 43168 27616 43220 27668
rect 44916 27616 44968 27668
rect 46940 27659 46992 27668
rect 46940 27625 46949 27659
rect 46949 27625 46983 27659
rect 46983 27625 46992 27659
rect 46940 27616 46992 27625
rect 39396 27591 39448 27600
rect 39396 27557 39430 27591
rect 39430 27557 39448 27591
rect 39396 27548 39448 27557
rect 41420 27548 41472 27600
rect 43260 27548 43312 27600
rect 41512 27480 41564 27532
rect 44640 27480 44692 27532
rect 45560 27523 45612 27532
rect 45560 27489 45569 27523
rect 45569 27489 45603 27523
rect 45603 27489 45612 27523
rect 45560 27480 45612 27489
rect 46204 27480 46256 27532
rect 38108 27412 38160 27464
rect 39120 27455 39172 27464
rect 39120 27421 39129 27455
rect 39129 27421 39163 27455
rect 39163 27421 39172 27455
rect 39120 27412 39172 27421
rect 42248 27455 42300 27464
rect 42248 27421 42257 27455
rect 42257 27421 42291 27455
rect 42291 27421 42300 27455
rect 42248 27412 42300 27421
rect 41696 27387 41748 27396
rect 41696 27353 41705 27387
rect 41705 27353 41739 27387
rect 41739 27353 41748 27387
rect 41696 27344 41748 27353
rect 38292 27319 38344 27328
rect 38292 27285 38301 27319
rect 38301 27285 38335 27319
rect 38335 27285 38344 27319
rect 38292 27276 38344 27285
rect 44272 27319 44324 27328
rect 44272 27285 44281 27319
rect 44281 27285 44315 27319
rect 44315 27285 44324 27319
rect 44272 27276 44324 27285
rect 45192 27276 45244 27328
rect 4246 27174 4298 27226
rect 4310 27174 4362 27226
rect 4374 27174 4426 27226
rect 4438 27174 4490 27226
rect 34966 27174 35018 27226
rect 35030 27174 35082 27226
rect 35094 27174 35146 27226
rect 35158 27174 35210 27226
rect 38108 27115 38160 27124
rect 38108 27081 38117 27115
rect 38117 27081 38151 27115
rect 38151 27081 38160 27115
rect 38108 27072 38160 27081
rect 38384 27115 38436 27124
rect 38384 27081 38393 27115
rect 38393 27081 38427 27115
rect 38427 27081 38436 27115
rect 38384 27072 38436 27081
rect 39396 27072 39448 27124
rect 43260 27115 43312 27124
rect 43260 27081 43269 27115
rect 43269 27081 43303 27115
rect 43303 27081 43312 27115
rect 43260 27072 43312 27081
rect 44640 27072 44692 27124
rect 45560 27115 45612 27124
rect 45560 27081 45569 27115
rect 45569 27081 45603 27115
rect 45603 27081 45612 27115
rect 45560 27072 45612 27081
rect 46204 27072 46256 27124
rect 43904 27047 43956 27056
rect 43904 27013 43913 27047
rect 43913 27013 43947 27047
rect 43947 27013 43956 27047
rect 43904 27004 43956 27013
rect 44272 26979 44324 26988
rect 44272 26945 44281 26979
rect 44281 26945 44315 26979
rect 44315 26945 44324 26979
rect 44272 26936 44324 26945
rect 38660 26868 38712 26920
rect 39120 26868 39172 26920
rect 41420 26868 41472 26920
rect 35900 26800 35952 26852
rect 38384 26800 38436 26852
rect 41880 26800 41932 26852
rect 44088 26800 44140 26852
rect 35992 26732 36044 26784
rect 37188 26775 37240 26784
rect 37188 26741 37197 26775
rect 37197 26741 37231 26775
rect 37231 26741 37240 26775
rect 37188 26732 37240 26741
rect 38292 26732 38344 26784
rect 42432 26732 42484 26784
rect 45008 26732 45060 26784
rect 45284 26775 45336 26784
rect 45284 26741 45293 26775
rect 45293 26741 45327 26775
rect 45327 26741 45336 26775
rect 45284 26732 45336 26741
rect 19606 26630 19658 26682
rect 19670 26630 19722 26682
rect 19734 26630 19786 26682
rect 19798 26630 19850 26682
rect 35900 26571 35952 26580
rect 35900 26537 35909 26571
rect 35909 26537 35943 26571
rect 35943 26537 35952 26571
rect 35900 26528 35952 26537
rect 38384 26571 38436 26580
rect 38384 26537 38393 26571
rect 38393 26537 38427 26571
rect 38427 26537 38436 26571
rect 38384 26528 38436 26537
rect 38568 26528 38620 26580
rect 41512 26528 41564 26580
rect 41880 26503 41932 26512
rect 41880 26469 41889 26503
rect 41889 26469 41923 26503
rect 41923 26469 41932 26503
rect 41880 26460 41932 26469
rect 44732 26460 44784 26512
rect 38752 26435 38804 26444
rect 38752 26401 38786 26435
rect 38786 26401 38804 26435
rect 38752 26392 38804 26401
rect 40684 26392 40736 26444
rect 43352 26435 43404 26444
rect 43352 26401 43361 26435
rect 43361 26401 43395 26435
rect 43395 26401 43404 26435
rect 43904 26435 43956 26444
rect 43352 26392 43404 26401
rect 43904 26401 43913 26435
rect 43913 26401 43947 26435
rect 43947 26401 43956 26435
rect 43904 26392 43956 26401
rect 44548 26392 44600 26444
rect 45560 26392 45612 26444
rect 46848 26392 46900 26444
rect 36728 26231 36780 26240
rect 36728 26197 36737 26231
rect 36737 26197 36771 26231
rect 36771 26197 36780 26231
rect 36728 26188 36780 26197
rect 37096 26188 37148 26240
rect 41328 26256 41380 26308
rect 41604 26256 41656 26308
rect 41972 26367 42024 26376
rect 41972 26333 41981 26367
rect 41981 26333 42015 26367
rect 42015 26333 42024 26367
rect 41972 26324 42024 26333
rect 45192 26367 45244 26376
rect 45192 26333 45201 26367
rect 45201 26333 45235 26367
rect 45235 26333 45244 26367
rect 45192 26324 45244 26333
rect 38660 26188 38712 26240
rect 42432 26231 42484 26240
rect 42432 26197 42441 26231
rect 42441 26197 42475 26231
rect 42475 26197 42484 26231
rect 42432 26188 42484 26197
rect 44640 26231 44692 26240
rect 44640 26197 44649 26231
rect 44649 26197 44683 26231
rect 44683 26197 44692 26231
rect 44640 26188 44692 26197
rect 47492 26231 47544 26240
rect 47492 26197 47501 26231
rect 47501 26197 47535 26231
rect 47535 26197 47544 26231
rect 47492 26188 47544 26197
rect 4246 26086 4298 26138
rect 4310 26086 4362 26138
rect 4374 26086 4426 26138
rect 4438 26086 4490 26138
rect 34966 26086 35018 26138
rect 35030 26086 35082 26138
rect 35094 26086 35146 26138
rect 35158 26086 35210 26138
rect 38384 25984 38436 26036
rect 38660 26027 38712 26036
rect 38660 25993 38669 26027
rect 38669 25993 38703 26027
rect 38703 25993 38712 26027
rect 38660 25984 38712 25993
rect 38752 25984 38804 26036
rect 41604 26027 41656 26036
rect 41604 25993 41613 26027
rect 41613 25993 41647 26027
rect 41647 25993 41656 26027
rect 41604 25984 41656 25993
rect 41972 25984 42024 26036
rect 45008 26027 45060 26036
rect 45008 25993 45017 26027
rect 45017 25993 45051 26027
rect 45051 25993 45060 26027
rect 45008 25984 45060 25993
rect 45560 25984 45612 26036
rect 40592 25959 40644 25968
rect 40592 25925 40601 25959
rect 40601 25925 40635 25959
rect 40635 25925 40644 25959
rect 40592 25916 40644 25925
rect 41420 25916 41472 25968
rect 42248 25916 42300 25968
rect 40684 25848 40736 25900
rect 44548 25916 44600 25968
rect 35992 25780 36044 25832
rect 36728 25780 36780 25832
rect 38568 25780 38620 25832
rect 35992 25687 36044 25696
rect 35992 25653 36001 25687
rect 36001 25653 36035 25687
rect 36035 25653 36044 25687
rect 35992 25644 36044 25653
rect 36360 25644 36412 25696
rect 37096 25712 37148 25764
rect 44640 25780 44692 25832
rect 46204 25780 46256 25832
rect 47492 25780 47544 25832
rect 41328 25712 41380 25764
rect 42432 25712 42484 25764
rect 43536 25712 43588 25764
rect 44732 25644 44784 25696
rect 46848 25644 46900 25696
rect 47400 25644 47452 25696
rect 19606 25542 19658 25594
rect 19670 25542 19722 25594
rect 19734 25542 19786 25594
rect 19798 25542 19850 25594
rect 35992 25440 36044 25492
rect 36176 25440 36228 25492
rect 40684 25483 40736 25492
rect 40684 25449 40693 25483
rect 40693 25449 40727 25483
rect 40727 25449 40736 25483
rect 40684 25440 40736 25449
rect 41880 25440 41932 25492
rect 44548 25483 44600 25492
rect 44548 25449 44557 25483
rect 44557 25449 44591 25483
rect 44591 25449 44600 25483
rect 44548 25440 44600 25449
rect 44640 25440 44692 25492
rect 46940 25483 46992 25492
rect 46940 25449 46949 25483
rect 46949 25449 46983 25483
rect 46983 25449 46992 25483
rect 46940 25440 46992 25449
rect 37832 25372 37884 25424
rect 38568 25372 38620 25424
rect 39580 25415 39632 25424
rect 39580 25381 39614 25415
rect 39614 25381 39632 25415
rect 39580 25372 39632 25381
rect 41972 25372 42024 25424
rect 43444 25372 43496 25424
rect 46020 25372 46072 25424
rect 36268 25347 36320 25356
rect 36268 25313 36277 25347
rect 36277 25313 36311 25347
rect 36311 25313 36320 25347
rect 36268 25304 36320 25313
rect 38660 25304 38712 25356
rect 43536 25347 43588 25356
rect 36912 25236 36964 25288
rect 38200 25279 38252 25288
rect 38200 25245 38209 25279
rect 38209 25245 38243 25279
rect 38243 25245 38252 25279
rect 38200 25236 38252 25245
rect 43536 25313 43545 25347
rect 43545 25313 43579 25347
rect 43579 25313 43588 25347
rect 43536 25304 43588 25313
rect 46756 25347 46808 25356
rect 46756 25313 46765 25347
rect 46765 25313 46799 25347
rect 46799 25313 46808 25347
rect 47308 25347 47360 25356
rect 46756 25304 46808 25313
rect 47308 25313 47317 25347
rect 47317 25313 47351 25347
rect 47351 25313 47360 25347
rect 47308 25304 47360 25313
rect 42616 25236 42668 25288
rect 35992 25211 36044 25220
rect 35992 25177 36001 25211
rect 36001 25177 36035 25211
rect 36035 25177 36044 25211
rect 35992 25168 36044 25177
rect 38292 25168 38344 25220
rect 44732 25168 44784 25220
rect 45836 25279 45888 25288
rect 45836 25245 45845 25279
rect 45845 25245 45879 25279
rect 45879 25245 45888 25279
rect 45836 25236 45888 25245
rect 47400 25236 47452 25288
rect 42340 25143 42392 25152
rect 42340 25109 42349 25143
rect 42349 25109 42383 25143
rect 42383 25109 42392 25143
rect 42340 25100 42392 25109
rect 46388 25100 46440 25152
rect 46848 25100 46900 25152
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 34966 24998 35018 25050
rect 35030 24998 35082 25050
rect 35094 24998 35146 25050
rect 35158 24998 35210 25050
rect 36912 24939 36964 24948
rect 36912 24905 36921 24939
rect 36921 24905 36955 24939
rect 36955 24905 36964 24939
rect 36912 24896 36964 24905
rect 37832 24939 37884 24948
rect 37832 24905 37841 24939
rect 37841 24905 37875 24939
rect 37875 24905 37884 24939
rect 37832 24896 37884 24905
rect 38200 24939 38252 24948
rect 38200 24905 38209 24939
rect 38209 24905 38243 24939
rect 38243 24905 38252 24939
rect 38200 24896 38252 24905
rect 38660 24896 38712 24948
rect 39580 24896 39632 24948
rect 42340 24896 42392 24948
rect 43536 24896 43588 24948
rect 45560 24896 45612 24948
rect 38752 24760 38804 24812
rect 36360 24692 36412 24744
rect 38660 24735 38712 24744
rect 38660 24701 38669 24735
rect 38669 24701 38703 24735
rect 38703 24701 38712 24735
rect 38660 24692 38712 24701
rect 35808 24667 35860 24676
rect 35808 24633 35842 24667
rect 35842 24633 35860 24667
rect 35808 24624 35860 24633
rect 43352 24692 43404 24744
rect 35440 24599 35492 24608
rect 35440 24565 35449 24599
rect 35449 24565 35483 24599
rect 35483 24565 35492 24599
rect 35440 24556 35492 24565
rect 39120 24556 39172 24608
rect 42064 24556 42116 24608
rect 42340 24556 42392 24608
rect 46020 24624 46072 24676
rect 46388 24667 46440 24676
rect 46388 24633 46422 24667
rect 46422 24633 46440 24667
rect 46388 24624 46440 24633
rect 46848 24624 46900 24676
rect 42892 24556 42944 24608
rect 43444 24599 43496 24608
rect 43444 24565 43453 24599
rect 43453 24565 43487 24599
rect 43487 24565 43496 24599
rect 43444 24556 43496 24565
rect 46940 24556 46992 24608
rect 19606 24454 19658 24506
rect 19670 24454 19722 24506
rect 19734 24454 19786 24506
rect 19798 24454 19850 24506
rect 36268 24352 36320 24404
rect 38568 24352 38620 24404
rect 41880 24352 41932 24404
rect 42340 24352 42392 24404
rect 42616 24395 42668 24404
rect 42616 24361 42625 24395
rect 42625 24361 42659 24395
rect 42659 24361 42668 24395
rect 42616 24352 42668 24361
rect 45836 24352 45888 24404
rect 46848 24395 46900 24404
rect 46848 24361 46857 24395
rect 46857 24361 46891 24395
rect 46891 24361 46900 24395
rect 46848 24352 46900 24361
rect 36636 24327 36688 24336
rect 36636 24293 36645 24327
rect 36645 24293 36679 24327
rect 36679 24293 36688 24327
rect 36636 24284 36688 24293
rect 35808 24216 35860 24268
rect 37188 24284 37240 24336
rect 42064 24216 42116 24268
rect 46020 24216 46072 24268
rect 35716 24148 35768 24200
rect 37188 24148 37240 24200
rect 45468 24191 45520 24200
rect 45468 24157 45477 24191
rect 45477 24157 45511 24191
rect 45511 24157 45520 24191
rect 45468 24148 45520 24157
rect 36176 24123 36228 24132
rect 36176 24089 36185 24123
rect 36185 24089 36219 24123
rect 36219 24089 36228 24123
rect 36176 24080 36228 24089
rect 30472 24012 30524 24064
rect 41604 24012 41656 24064
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 34966 23910 35018 23962
rect 35030 23910 35082 23962
rect 35094 23910 35146 23962
rect 35158 23910 35210 23962
rect 31300 23851 31352 23860
rect 31300 23817 31309 23851
rect 31309 23817 31343 23851
rect 31343 23817 31352 23851
rect 31300 23808 31352 23817
rect 35808 23808 35860 23860
rect 41052 23851 41104 23860
rect 41052 23817 41061 23851
rect 41061 23817 41095 23851
rect 41095 23817 41104 23851
rect 41052 23808 41104 23817
rect 42064 23851 42116 23860
rect 42064 23817 42073 23851
rect 42073 23817 42107 23851
rect 42107 23817 42116 23851
rect 42064 23808 42116 23817
rect 42248 23808 42300 23860
rect 35716 23740 35768 23792
rect 41604 23715 41656 23724
rect 41604 23681 41613 23715
rect 41613 23681 41647 23715
rect 41647 23681 41656 23715
rect 41604 23672 41656 23681
rect 35440 23604 35492 23656
rect 31668 23536 31720 23588
rect 31852 23579 31904 23588
rect 31852 23545 31861 23579
rect 31861 23545 31895 23579
rect 31895 23545 31904 23579
rect 31852 23536 31904 23545
rect 30472 23468 30524 23520
rect 35808 23468 35860 23520
rect 36912 23604 36964 23656
rect 42248 23604 42300 23656
rect 42616 23604 42668 23656
rect 41420 23536 41472 23588
rect 37280 23468 37332 23520
rect 38476 23468 38528 23520
rect 38660 23511 38712 23520
rect 38660 23477 38669 23511
rect 38669 23477 38703 23511
rect 38703 23477 38712 23511
rect 38660 23468 38712 23477
rect 41052 23468 41104 23520
rect 44088 23468 44140 23520
rect 44640 23468 44692 23520
rect 45468 23511 45520 23520
rect 45468 23477 45477 23511
rect 45477 23477 45511 23511
rect 45511 23477 45520 23511
rect 45468 23468 45520 23477
rect 46020 23468 46072 23520
rect 19606 23366 19658 23418
rect 19670 23366 19722 23418
rect 19734 23366 19786 23418
rect 19798 23366 19850 23418
rect 31760 23264 31812 23316
rect 36912 23264 36964 23316
rect 38200 23264 38252 23316
rect 38936 23264 38988 23316
rect 41420 23264 41472 23316
rect 42616 23307 42668 23316
rect 42616 23273 42625 23307
rect 42625 23273 42659 23307
rect 42659 23273 42668 23307
rect 42616 23264 42668 23273
rect 46020 23307 46072 23316
rect 46020 23273 46029 23307
rect 46029 23273 46063 23307
rect 46063 23273 46072 23307
rect 46020 23264 46072 23273
rect 47032 23264 47084 23316
rect 31852 23196 31904 23248
rect 33232 23196 33284 23248
rect 38660 23171 38712 23180
rect 38660 23137 38669 23171
rect 38669 23137 38703 23171
rect 38703 23137 38712 23171
rect 38660 23128 38712 23137
rect 38752 23128 38804 23180
rect 39856 23128 39908 23180
rect 44916 23171 44968 23180
rect 44916 23137 44950 23171
rect 44950 23137 44968 23171
rect 44916 23128 44968 23137
rect 47308 23128 47360 23180
rect 34060 23103 34112 23112
rect 34060 23069 34069 23103
rect 34069 23069 34103 23103
rect 34103 23069 34112 23103
rect 34060 23060 34112 23069
rect 34612 23060 34664 23112
rect 39028 23060 39080 23112
rect 39120 23103 39172 23112
rect 39120 23069 39129 23103
rect 39129 23069 39163 23103
rect 39163 23069 39172 23103
rect 44640 23103 44692 23112
rect 39120 23060 39172 23069
rect 44640 23069 44649 23103
rect 44649 23069 44683 23103
rect 44683 23069 44692 23103
rect 44640 23060 44692 23069
rect 33600 23035 33652 23044
rect 33600 23001 33609 23035
rect 33609 23001 33643 23035
rect 33643 23001 33652 23035
rect 33600 22992 33652 23001
rect 36176 22967 36228 22976
rect 36176 22933 36185 22967
rect 36185 22933 36219 22967
rect 36219 22933 36228 22967
rect 36176 22924 36228 22933
rect 40500 22967 40552 22976
rect 40500 22933 40509 22967
rect 40509 22933 40543 22967
rect 40543 22933 40552 22967
rect 40500 22924 40552 22933
rect 41328 22924 41380 22976
rect 44088 22924 44140 22976
rect 46664 22967 46716 22976
rect 46664 22933 46673 22967
rect 46673 22933 46707 22967
rect 46707 22933 46716 22967
rect 46664 22924 46716 22933
rect 46940 22967 46992 22976
rect 46940 22933 46949 22967
rect 46949 22933 46983 22967
rect 46983 22933 46992 22967
rect 46940 22924 46992 22933
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 34966 22822 35018 22874
rect 35030 22822 35082 22874
rect 35094 22822 35146 22874
rect 35158 22822 35210 22874
rect 34060 22720 34112 22772
rect 34612 22695 34664 22704
rect 34612 22661 34621 22695
rect 34621 22661 34655 22695
rect 34655 22661 34664 22695
rect 34612 22652 34664 22661
rect 31852 22584 31904 22636
rect 37372 22720 37424 22772
rect 39120 22720 39172 22772
rect 39856 22763 39908 22772
rect 39856 22729 39865 22763
rect 39865 22729 39899 22763
rect 39899 22729 39908 22763
rect 39856 22720 39908 22729
rect 42616 22720 42668 22772
rect 44916 22763 44968 22772
rect 44916 22729 44925 22763
rect 44925 22729 44959 22763
rect 44959 22729 44968 22763
rect 44916 22720 44968 22729
rect 46296 22763 46348 22772
rect 46296 22729 46305 22763
rect 46305 22729 46339 22763
rect 46339 22729 46348 22763
rect 46296 22720 46348 22729
rect 38568 22695 38620 22704
rect 38568 22661 38577 22695
rect 38577 22661 38611 22695
rect 38611 22661 38620 22695
rect 38568 22652 38620 22661
rect 47308 22695 47360 22704
rect 47308 22661 47317 22695
rect 47317 22661 47351 22695
rect 47351 22661 47360 22695
rect 47308 22652 47360 22661
rect 32404 22516 32456 22568
rect 29552 22423 29604 22432
rect 29552 22389 29561 22423
rect 29561 22389 29595 22423
rect 29595 22389 29604 22423
rect 29552 22380 29604 22389
rect 32220 22423 32272 22432
rect 32220 22389 32229 22423
rect 32229 22389 32263 22423
rect 32263 22389 32272 22423
rect 32220 22380 32272 22389
rect 33600 22380 33652 22432
rect 35808 22380 35860 22432
rect 38476 22584 38528 22636
rect 46664 22584 46716 22636
rect 46848 22627 46900 22636
rect 46848 22593 46857 22627
rect 46857 22593 46891 22627
rect 46891 22593 46900 22627
rect 46848 22584 46900 22593
rect 37188 22516 37240 22568
rect 38200 22516 38252 22568
rect 39028 22516 39080 22568
rect 38660 22448 38712 22500
rect 37280 22380 37332 22432
rect 38936 22380 38988 22432
rect 40408 22380 40460 22432
rect 44640 22516 44692 22568
rect 46112 22516 46164 22568
rect 41328 22448 41380 22500
rect 41604 22448 41656 22500
rect 44088 22448 44140 22500
rect 45100 22448 45152 22500
rect 45560 22380 45612 22432
rect 46940 22380 46992 22432
rect 19606 22278 19658 22330
rect 19670 22278 19722 22330
rect 19734 22278 19786 22330
rect 19798 22278 19850 22330
rect 29552 22176 29604 22228
rect 29920 22176 29972 22228
rect 31760 22176 31812 22228
rect 32220 22176 32272 22228
rect 33048 22176 33100 22228
rect 34612 22176 34664 22228
rect 37372 22176 37424 22228
rect 38568 22176 38620 22228
rect 38752 22176 38804 22228
rect 32404 22151 32456 22160
rect 32404 22117 32413 22151
rect 32413 22117 32447 22151
rect 32447 22117 32456 22151
rect 32404 22108 32456 22117
rect 33600 22108 33652 22160
rect 39856 22176 39908 22228
rect 45100 22219 45152 22228
rect 45100 22185 45109 22219
rect 45109 22185 45143 22219
rect 45143 22185 45152 22219
rect 45100 22176 45152 22185
rect 41512 22151 41564 22160
rect 30288 22040 30340 22092
rect 36452 22083 36504 22092
rect 36452 22049 36461 22083
rect 36461 22049 36495 22083
rect 36495 22049 36504 22083
rect 36452 22040 36504 22049
rect 36544 22040 36596 22092
rect 37188 22040 37240 22092
rect 37556 22040 37608 22092
rect 41512 22117 41521 22151
rect 41521 22117 41555 22151
rect 41555 22117 41564 22151
rect 41512 22108 41564 22117
rect 43904 22151 43956 22160
rect 43904 22117 43913 22151
rect 43913 22117 43947 22151
rect 43947 22117 43956 22151
rect 43904 22108 43956 22117
rect 27988 21972 28040 22024
rect 28908 22015 28960 22024
rect 28908 21981 28917 22015
rect 28917 21981 28951 22015
rect 28951 21981 28960 22015
rect 28908 21972 28960 21981
rect 33048 21972 33100 22024
rect 33508 21972 33560 22024
rect 28264 21836 28316 21888
rect 31208 21879 31260 21888
rect 31208 21845 31217 21879
rect 31217 21845 31251 21879
rect 31251 21845 31260 21879
rect 31208 21836 31260 21845
rect 33232 21836 33284 21888
rect 37556 21836 37608 21888
rect 38200 21972 38252 22024
rect 40776 22040 40828 22092
rect 41328 22083 41380 22092
rect 41328 22049 41337 22083
rect 41337 22049 41371 22083
rect 41371 22049 41380 22083
rect 41328 22040 41380 22049
rect 43444 22040 43496 22092
rect 44916 22108 44968 22160
rect 45560 22040 45612 22092
rect 46848 22040 46900 22092
rect 38660 22015 38712 22024
rect 38660 21981 38669 22015
rect 38669 21981 38703 22015
rect 38703 21981 38712 22015
rect 38660 21972 38712 21981
rect 41604 22015 41656 22024
rect 41604 21981 41613 22015
rect 41613 21981 41647 22015
rect 41647 21981 41656 22015
rect 41604 21972 41656 21981
rect 46112 22015 46164 22024
rect 46112 21981 46121 22015
rect 46121 21981 46155 22015
rect 46155 21981 46164 22015
rect 46112 21972 46164 21981
rect 41052 21947 41104 21956
rect 41052 21913 41061 21947
rect 41061 21913 41095 21947
rect 41095 21913 41104 21947
rect 41052 21904 41104 21913
rect 47492 21947 47544 21956
rect 47492 21913 47501 21947
rect 47501 21913 47535 21947
rect 47535 21913 47544 21947
rect 47492 21904 47544 21913
rect 38292 21836 38344 21888
rect 38752 21836 38804 21888
rect 42340 21836 42392 21888
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 34966 21734 35018 21786
rect 35030 21734 35082 21786
rect 35094 21734 35146 21786
rect 35158 21734 35210 21786
rect 28908 21632 28960 21684
rect 29736 21632 29788 21684
rect 32404 21632 32456 21684
rect 37372 21632 37424 21684
rect 37556 21675 37608 21684
rect 37556 21641 37565 21675
rect 37565 21641 37599 21675
rect 37599 21641 37608 21675
rect 37556 21632 37608 21641
rect 38660 21675 38712 21684
rect 38660 21641 38669 21675
rect 38669 21641 38703 21675
rect 38703 21641 38712 21675
rect 38660 21632 38712 21641
rect 41420 21632 41472 21684
rect 43444 21675 43496 21684
rect 43444 21641 43453 21675
rect 43453 21641 43487 21675
rect 43487 21641 43496 21675
rect 43444 21632 43496 21641
rect 44916 21632 44968 21684
rect 45560 21675 45612 21684
rect 45560 21641 45569 21675
rect 45569 21641 45603 21675
rect 45603 21641 45612 21675
rect 45560 21632 45612 21641
rect 46848 21632 46900 21684
rect 27896 21564 27948 21616
rect 28264 21539 28316 21548
rect 28264 21505 28273 21539
rect 28273 21505 28307 21539
rect 28307 21505 28316 21539
rect 28264 21496 28316 21505
rect 27988 21471 28040 21480
rect 27988 21437 27997 21471
rect 27997 21437 28031 21471
rect 28031 21437 28040 21471
rect 27988 21428 28040 21437
rect 43168 21564 43220 21616
rect 43904 21564 43956 21616
rect 29920 21539 29972 21548
rect 29920 21505 29929 21539
rect 29929 21505 29963 21539
rect 29963 21505 29972 21539
rect 29920 21496 29972 21505
rect 41328 21496 41380 21548
rect 41972 21496 42024 21548
rect 44180 21496 44232 21548
rect 46112 21539 46164 21548
rect 46112 21505 46121 21539
rect 46121 21505 46155 21539
rect 46155 21505 46164 21539
rect 46112 21496 46164 21505
rect 29644 21403 29696 21412
rect 29644 21369 29653 21403
rect 29653 21369 29687 21403
rect 29687 21369 29696 21403
rect 29644 21360 29696 21369
rect 29736 21360 29788 21412
rect 31208 21428 31260 21480
rect 33600 21428 33652 21480
rect 31668 21360 31720 21412
rect 33508 21360 33560 21412
rect 35808 21428 35860 21480
rect 40776 21471 40828 21480
rect 40776 21437 40785 21471
rect 40785 21437 40819 21471
rect 40819 21437 40828 21471
rect 40776 21428 40828 21437
rect 35532 21403 35584 21412
rect 35532 21369 35566 21403
rect 35566 21369 35584 21403
rect 35532 21360 35584 21369
rect 36452 21360 36504 21412
rect 42800 21428 42852 21480
rect 44088 21403 44140 21412
rect 44088 21369 44097 21403
rect 44097 21369 44131 21403
rect 44131 21369 44140 21403
rect 44088 21360 44140 21369
rect 46388 21403 46440 21412
rect 46388 21369 46422 21403
rect 46422 21369 46440 21403
rect 46388 21360 46440 21369
rect 29828 21335 29880 21344
rect 29828 21301 29837 21335
rect 29837 21301 29871 21335
rect 29871 21301 29880 21335
rect 29828 21292 29880 21301
rect 36636 21335 36688 21344
rect 36636 21301 36645 21335
rect 36645 21301 36679 21335
rect 36679 21301 36688 21335
rect 36636 21292 36688 21301
rect 38200 21335 38252 21344
rect 38200 21301 38209 21335
rect 38209 21301 38243 21335
rect 38243 21301 38252 21335
rect 38200 21292 38252 21301
rect 40776 21292 40828 21344
rect 44180 21292 44232 21344
rect 19606 21190 19658 21242
rect 19670 21190 19722 21242
rect 19734 21190 19786 21242
rect 19798 21190 19850 21242
rect 36452 21088 36504 21140
rect 36544 21131 36596 21140
rect 36544 21097 36553 21131
rect 36553 21097 36587 21131
rect 36587 21097 36596 21131
rect 36544 21088 36596 21097
rect 41420 21088 41472 21140
rect 41604 21131 41656 21140
rect 41604 21097 41613 21131
rect 41613 21097 41647 21131
rect 41647 21097 41656 21131
rect 41604 21088 41656 21097
rect 42340 21131 42392 21140
rect 42340 21097 42349 21131
rect 42349 21097 42383 21131
rect 42383 21097 42392 21131
rect 42340 21088 42392 21097
rect 43168 21131 43220 21140
rect 43168 21097 43177 21131
rect 43177 21097 43211 21131
rect 43211 21097 43220 21131
rect 43168 21088 43220 21097
rect 43444 21131 43496 21140
rect 43444 21097 43453 21131
rect 43453 21097 43487 21131
rect 43487 21097 43496 21131
rect 43444 21088 43496 21097
rect 44088 21088 44140 21140
rect 46112 21131 46164 21140
rect 46112 21097 46121 21131
rect 46121 21097 46155 21131
rect 46155 21097 46164 21131
rect 46112 21088 46164 21097
rect 47216 21088 47268 21140
rect 30932 21063 30984 21072
rect 30932 21029 30941 21063
rect 30941 21029 30975 21063
rect 30975 21029 30984 21063
rect 30932 21020 30984 21029
rect 31208 21020 31260 21072
rect 35532 21020 35584 21072
rect 44640 21020 44692 21072
rect 28080 20952 28132 21004
rect 32496 20952 32548 21004
rect 44180 20952 44232 21004
rect 46756 20995 46808 21004
rect 46756 20961 46765 20995
rect 46765 20961 46799 20995
rect 46799 20961 46808 20995
rect 46756 20952 46808 20961
rect 27252 20884 27304 20936
rect 27620 20884 27672 20936
rect 27896 20927 27948 20936
rect 27896 20893 27905 20927
rect 27905 20893 27939 20927
rect 27939 20893 27948 20927
rect 27896 20884 27948 20893
rect 30472 20859 30524 20868
rect 30472 20825 30481 20859
rect 30481 20825 30515 20859
rect 30515 20825 30524 20859
rect 30472 20816 30524 20825
rect 29828 20748 29880 20800
rect 30380 20748 30432 20800
rect 32864 20927 32916 20936
rect 32864 20893 32873 20927
rect 32873 20893 32907 20927
rect 32907 20893 32916 20927
rect 32864 20884 32916 20893
rect 33048 20884 33100 20936
rect 40316 20927 40368 20936
rect 40316 20893 40325 20927
rect 40325 20893 40359 20927
rect 40359 20893 40368 20927
rect 40316 20884 40368 20893
rect 45100 20927 45152 20936
rect 45100 20893 45109 20927
rect 45109 20893 45143 20927
rect 45143 20893 45152 20927
rect 45100 20884 45152 20893
rect 46388 20884 46440 20936
rect 45468 20816 45520 20868
rect 32772 20748 32824 20800
rect 34244 20791 34296 20800
rect 34244 20757 34253 20791
rect 34253 20757 34287 20791
rect 34287 20757 34296 20791
rect 34244 20748 34296 20757
rect 38016 20791 38068 20800
rect 38016 20757 38025 20791
rect 38025 20757 38059 20791
rect 38059 20757 38068 20791
rect 38016 20748 38068 20757
rect 38292 20791 38344 20800
rect 38292 20757 38301 20791
rect 38301 20757 38335 20791
rect 38335 20757 38344 20791
rect 38292 20748 38344 20757
rect 40776 20791 40828 20800
rect 40776 20757 40785 20791
rect 40785 20757 40819 20791
rect 40819 20757 40828 20791
rect 40776 20748 40828 20757
rect 41328 20748 41380 20800
rect 44180 20748 44232 20800
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 34966 20646 35018 20698
rect 35030 20646 35082 20698
rect 35094 20646 35146 20698
rect 35158 20646 35210 20698
rect 27896 20544 27948 20596
rect 30932 20544 30984 20596
rect 33048 20544 33100 20596
rect 33232 20587 33284 20596
rect 33232 20553 33241 20587
rect 33241 20553 33275 20587
rect 33275 20553 33284 20587
rect 33232 20544 33284 20553
rect 34704 20544 34756 20596
rect 35808 20544 35860 20596
rect 40316 20587 40368 20596
rect 31024 20519 31076 20528
rect 31024 20485 31033 20519
rect 31033 20485 31067 20519
rect 31067 20485 31076 20519
rect 31024 20476 31076 20485
rect 32404 20519 32456 20528
rect 32404 20485 32413 20519
rect 32413 20485 32447 20519
rect 32447 20485 32456 20519
rect 32404 20476 32456 20485
rect 40316 20553 40325 20587
rect 40325 20553 40359 20587
rect 40359 20553 40368 20587
rect 40316 20544 40368 20553
rect 40592 20587 40644 20596
rect 40592 20553 40601 20587
rect 40601 20553 40635 20587
rect 40635 20553 40644 20587
rect 40592 20544 40644 20553
rect 41420 20544 41472 20596
rect 28080 20408 28132 20460
rect 37740 20408 37792 20460
rect 42800 20544 42852 20596
rect 44180 20544 44232 20596
rect 46756 20587 46808 20596
rect 46756 20553 46765 20587
rect 46765 20553 46799 20587
rect 46799 20553 46808 20587
rect 46756 20544 46808 20553
rect 44640 20519 44692 20528
rect 44640 20485 44649 20519
rect 44649 20485 44683 20519
rect 44683 20485 44692 20519
rect 44640 20476 44692 20485
rect 29736 20340 29788 20392
rect 29920 20383 29972 20392
rect 29920 20349 29954 20383
rect 29954 20349 29972 20383
rect 29920 20340 29972 20349
rect 38016 20340 38068 20392
rect 40684 20340 40736 20392
rect 42248 20383 42300 20392
rect 42248 20349 42257 20383
rect 42257 20349 42291 20383
rect 42291 20349 42300 20383
rect 42248 20340 42300 20349
rect 42432 20408 42484 20460
rect 42984 20451 43036 20460
rect 42984 20417 42993 20451
rect 42993 20417 43027 20451
rect 43027 20417 43036 20451
rect 42984 20408 43036 20417
rect 43996 20408 44048 20460
rect 32864 20272 32916 20324
rect 33232 20272 33284 20324
rect 33600 20272 33652 20324
rect 41604 20272 41656 20324
rect 27252 20204 27304 20256
rect 27436 20247 27488 20256
rect 27436 20213 27445 20247
rect 27445 20213 27479 20247
rect 27479 20213 27488 20247
rect 27436 20204 27488 20213
rect 34244 20204 34296 20256
rect 34520 20204 34572 20256
rect 35440 20204 35492 20256
rect 37188 20204 37240 20256
rect 39304 20247 39356 20256
rect 39304 20213 39313 20247
rect 39313 20213 39347 20247
rect 39347 20213 39356 20247
rect 39304 20204 39356 20213
rect 39856 20247 39908 20256
rect 39856 20213 39865 20247
rect 39865 20213 39899 20247
rect 39899 20213 39908 20247
rect 39856 20204 39908 20213
rect 40592 20204 40644 20256
rect 19606 20102 19658 20154
rect 19670 20102 19722 20154
rect 19734 20102 19786 20154
rect 19798 20102 19850 20154
rect 29920 20000 29972 20052
rect 30932 20000 30984 20052
rect 31208 20043 31260 20052
rect 31208 20009 31217 20043
rect 31217 20009 31251 20043
rect 31251 20009 31260 20043
rect 31208 20000 31260 20009
rect 33232 20043 33284 20052
rect 33232 20009 33241 20043
rect 33241 20009 33275 20043
rect 33275 20009 33284 20043
rect 33232 20000 33284 20009
rect 33600 20043 33652 20052
rect 33600 20009 33609 20043
rect 33609 20009 33643 20043
rect 33643 20009 33652 20043
rect 33600 20000 33652 20009
rect 38016 20000 38068 20052
rect 38660 20000 38712 20052
rect 41604 20043 41656 20052
rect 41604 20009 41613 20043
rect 41613 20009 41647 20043
rect 41647 20009 41656 20043
rect 41604 20000 41656 20009
rect 42248 20000 42300 20052
rect 45100 20000 45152 20052
rect 47400 20043 47452 20052
rect 47400 20009 47409 20043
rect 47409 20009 47443 20043
rect 47443 20009 47452 20043
rect 47400 20000 47452 20009
rect 32772 19975 32824 19984
rect 32772 19941 32781 19975
rect 32781 19941 32815 19975
rect 32815 19941 32824 19975
rect 32772 19932 32824 19941
rect 39304 19932 39356 19984
rect 40224 19932 40276 19984
rect 42156 19932 42208 19984
rect 42984 19932 43036 19984
rect 32128 19907 32180 19916
rect 32128 19873 32137 19907
rect 32137 19873 32171 19907
rect 32171 19873 32180 19907
rect 32128 19864 32180 19873
rect 34612 19864 34664 19916
rect 34980 19907 35032 19916
rect 34980 19873 35014 19907
rect 35014 19873 35032 19907
rect 34980 19864 35032 19873
rect 37740 19907 37792 19916
rect 37740 19873 37749 19907
rect 37749 19873 37783 19907
rect 37783 19873 37792 19907
rect 37740 19864 37792 19873
rect 38384 19864 38436 19916
rect 45008 19907 45060 19916
rect 45008 19873 45042 19907
rect 45042 19873 45060 19907
rect 45008 19864 45060 19873
rect 47308 19864 47360 19916
rect 29920 19796 29972 19848
rect 30380 19796 30432 19848
rect 34428 19796 34480 19848
rect 34704 19839 34756 19848
rect 34704 19805 34713 19839
rect 34713 19805 34747 19839
rect 34747 19805 34756 19839
rect 34704 19796 34756 19805
rect 43720 19839 43772 19848
rect 34704 19660 34756 19712
rect 36084 19703 36136 19712
rect 36084 19669 36093 19703
rect 36093 19669 36127 19703
rect 36127 19669 36136 19703
rect 36084 19660 36136 19669
rect 43720 19805 43729 19839
rect 43729 19805 43763 19839
rect 43763 19805 43772 19839
rect 43720 19796 43772 19805
rect 44732 19839 44784 19848
rect 44732 19805 44741 19839
rect 44741 19805 44775 19839
rect 44775 19805 44784 19839
rect 44732 19796 44784 19805
rect 40408 19660 40460 19712
rect 44180 19660 44232 19712
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 34966 19558 35018 19610
rect 35030 19558 35082 19610
rect 35094 19558 35146 19610
rect 35158 19558 35210 19610
rect 31208 19456 31260 19508
rect 37740 19499 37792 19508
rect 37740 19465 37749 19499
rect 37749 19465 37783 19499
rect 37783 19465 37792 19499
rect 37740 19456 37792 19465
rect 40592 19499 40644 19508
rect 40592 19465 40601 19499
rect 40601 19465 40635 19499
rect 40635 19465 40644 19499
rect 40592 19456 40644 19465
rect 43720 19456 43772 19508
rect 47308 19499 47360 19508
rect 47308 19465 47317 19499
rect 47317 19465 47351 19499
rect 47351 19465 47360 19499
rect 47308 19456 47360 19465
rect 31024 19388 31076 19440
rect 29736 19363 29788 19372
rect 29736 19329 29745 19363
rect 29745 19329 29779 19363
rect 29779 19329 29788 19363
rect 29736 19320 29788 19329
rect 35440 19320 35492 19372
rect 38660 19363 38712 19372
rect 38660 19329 38669 19363
rect 38669 19329 38703 19363
rect 38703 19329 38712 19363
rect 38660 19320 38712 19329
rect 40224 19320 40276 19372
rect 30196 19184 30248 19236
rect 32220 19295 32272 19304
rect 32220 19261 32229 19295
rect 32229 19261 32263 19295
rect 32263 19261 32272 19295
rect 32220 19252 32272 19261
rect 34428 19252 34480 19304
rect 34704 19295 34756 19304
rect 34704 19261 34713 19295
rect 34713 19261 34747 19295
rect 34747 19261 34756 19295
rect 34704 19252 34756 19261
rect 34796 19252 34848 19304
rect 35348 19252 35400 19304
rect 38568 19252 38620 19304
rect 33600 19159 33652 19168
rect 33600 19125 33609 19159
rect 33609 19125 33643 19159
rect 33643 19125 33652 19159
rect 33600 19116 33652 19125
rect 44180 19363 44232 19372
rect 44180 19329 44189 19363
rect 44189 19329 44223 19363
rect 44223 19329 44232 19363
rect 44180 19320 44232 19329
rect 45008 19320 45060 19372
rect 44088 19252 44140 19304
rect 37188 19184 37240 19236
rect 35624 19116 35676 19168
rect 36912 19159 36964 19168
rect 36912 19125 36921 19159
rect 36921 19125 36955 19159
rect 36955 19125 36964 19159
rect 36912 19116 36964 19125
rect 37832 19116 37884 19168
rect 39120 19116 39172 19168
rect 40408 19116 40460 19168
rect 40960 19184 41012 19236
rect 42156 19184 42208 19236
rect 43444 19116 43496 19168
rect 44732 19116 44784 19168
rect 46112 19116 46164 19168
rect 19606 19014 19658 19066
rect 19670 19014 19722 19066
rect 19734 19014 19786 19066
rect 19798 19014 19850 19066
rect 34612 18955 34664 18964
rect 34612 18921 34621 18955
rect 34621 18921 34655 18955
rect 34655 18921 34664 18955
rect 34612 18912 34664 18921
rect 38660 18912 38712 18964
rect 40224 18955 40276 18964
rect 40224 18921 40233 18955
rect 40233 18921 40267 18955
rect 40267 18921 40276 18955
rect 40224 18912 40276 18921
rect 40776 18955 40828 18964
rect 40776 18921 40787 18955
rect 40787 18921 40821 18955
rect 40821 18921 40828 18955
rect 42156 18955 42208 18964
rect 40776 18912 40828 18921
rect 42156 18921 42165 18955
rect 42165 18921 42199 18955
rect 42199 18921 42208 18955
rect 42156 18912 42208 18921
rect 45008 18955 45060 18964
rect 45008 18921 45017 18955
rect 45017 18921 45051 18955
rect 45051 18921 45060 18955
rect 45008 18912 45060 18921
rect 29368 18844 29420 18896
rect 30196 18887 30248 18896
rect 30196 18853 30205 18887
rect 30205 18853 30239 18887
rect 30239 18853 30248 18887
rect 30196 18844 30248 18853
rect 34520 18844 34572 18896
rect 35348 18844 35400 18896
rect 35624 18887 35676 18896
rect 35624 18853 35633 18887
rect 35633 18853 35667 18887
rect 35667 18853 35676 18887
rect 35624 18844 35676 18853
rect 36084 18844 36136 18896
rect 36912 18844 36964 18896
rect 29920 18819 29972 18828
rect 29920 18785 29929 18819
rect 29929 18785 29963 18819
rect 29963 18785 29972 18819
rect 29920 18776 29972 18785
rect 38108 18819 38160 18828
rect 38108 18785 38117 18819
rect 38117 18785 38151 18819
rect 38151 18785 38160 18819
rect 38108 18776 38160 18785
rect 40224 18776 40276 18828
rect 44364 18776 44416 18828
rect 45560 18776 45612 18828
rect 46940 18776 46992 18828
rect 34520 18708 34572 18760
rect 38384 18751 38436 18760
rect 38384 18717 38393 18751
rect 38393 18717 38427 18751
rect 38427 18717 38436 18751
rect 38384 18708 38436 18717
rect 39948 18708 40000 18760
rect 40684 18708 40736 18760
rect 40960 18708 41012 18760
rect 43628 18751 43680 18760
rect 30288 18640 30340 18692
rect 37832 18683 37884 18692
rect 37832 18649 37841 18683
rect 37841 18649 37875 18683
rect 37875 18649 37884 18683
rect 37832 18640 37884 18649
rect 43628 18717 43637 18751
rect 43637 18717 43671 18751
rect 43671 18717 43680 18751
rect 43628 18708 43680 18717
rect 46112 18751 46164 18760
rect 46112 18717 46121 18751
rect 46121 18717 46155 18751
rect 46155 18717 46164 18751
rect 46112 18708 46164 18717
rect 30104 18572 30156 18624
rect 31760 18572 31812 18624
rect 32128 18572 32180 18624
rect 35256 18572 35308 18624
rect 40500 18572 40552 18624
rect 42892 18615 42944 18624
rect 42892 18581 42901 18615
rect 42901 18581 42935 18615
rect 42935 18581 42944 18615
rect 42892 18572 42944 18581
rect 47492 18615 47544 18624
rect 47492 18581 47501 18615
rect 47501 18581 47535 18615
rect 47535 18581 47544 18615
rect 47492 18572 47544 18581
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 34966 18470 35018 18522
rect 35030 18470 35082 18522
rect 35094 18470 35146 18522
rect 35158 18470 35210 18522
rect 29920 18368 29972 18420
rect 35624 18368 35676 18420
rect 36912 18368 36964 18420
rect 35348 18300 35400 18352
rect 37832 18368 37884 18420
rect 38108 18411 38160 18420
rect 38108 18377 38117 18411
rect 38117 18377 38151 18411
rect 38151 18377 38160 18411
rect 38108 18368 38160 18377
rect 39948 18411 40000 18420
rect 39948 18377 39957 18411
rect 39957 18377 39991 18411
rect 39991 18377 40000 18411
rect 39948 18368 40000 18377
rect 40776 18411 40828 18420
rect 40776 18377 40785 18411
rect 40785 18377 40819 18411
rect 40819 18377 40828 18411
rect 40776 18368 40828 18377
rect 41972 18411 42024 18420
rect 41972 18377 41981 18411
rect 41981 18377 42015 18411
rect 42015 18377 42024 18411
rect 41972 18368 42024 18377
rect 43628 18368 43680 18420
rect 43996 18368 44048 18420
rect 44364 18411 44416 18420
rect 44364 18377 44373 18411
rect 44373 18377 44407 18411
rect 44407 18377 44416 18411
rect 44364 18368 44416 18377
rect 45560 18411 45612 18420
rect 45560 18377 45569 18411
rect 45569 18377 45603 18411
rect 45603 18377 45612 18411
rect 45560 18368 45612 18377
rect 46112 18368 46164 18420
rect 40224 18343 40276 18352
rect 40224 18309 40233 18343
rect 40233 18309 40267 18343
rect 40267 18309 40276 18343
rect 40224 18300 40276 18309
rect 34428 18232 34480 18284
rect 42892 18232 42944 18284
rect 29736 18164 29788 18216
rect 34796 18164 34848 18216
rect 35348 18164 35400 18216
rect 35808 18164 35860 18216
rect 35992 18207 36044 18216
rect 35992 18173 36015 18207
rect 36015 18173 36044 18207
rect 35992 18164 36044 18173
rect 44088 18300 44140 18352
rect 30104 18096 30156 18148
rect 43260 18139 43312 18148
rect 43260 18105 43269 18139
rect 43269 18105 43303 18139
rect 43303 18105 43312 18139
rect 43260 18096 43312 18105
rect 46388 18139 46440 18148
rect 46388 18105 46422 18139
rect 46422 18105 46440 18139
rect 46388 18096 46440 18105
rect 29368 18028 29420 18080
rect 30196 18028 30248 18080
rect 35808 18028 35860 18080
rect 37188 18028 37240 18080
rect 38384 18028 38436 18080
rect 39120 18028 39172 18080
rect 41052 18071 41104 18080
rect 41052 18037 41061 18071
rect 41061 18037 41095 18071
rect 41095 18037 41104 18071
rect 41052 18028 41104 18037
rect 42984 18028 43036 18080
rect 46940 18028 46992 18080
rect 19606 17926 19658 17978
rect 19670 17926 19722 17978
rect 19734 17926 19786 17978
rect 19798 17926 19850 17978
rect 30196 17756 30248 17808
rect 30564 17799 30616 17808
rect 30564 17765 30573 17799
rect 30573 17765 30607 17799
rect 30607 17765 30616 17799
rect 30564 17756 30616 17765
rect 30748 17799 30800 17808
rect 30748 17765 30757 17799
rect 30757 17765 30791 17799
rect 30791 17765 30800 17799
rect 30748 17756 30800 17765
rect 35992 17867 36044 17876
rect 35992 17833 36001 17867
rect 36001 17833 36035 17867
rect 36035 17833 36044 17867
rect 35992 17824 36044 17833
rect 41144 17867 41196 17876
rect 41144 17833 41153 17867
rect 41153 17833 41187 17867
rect 41187 17833 41196 17867
rect 41144 17824 41196 17833
rect 44088 17824 44140 17876
rect 46112 17824 46164 17876
rect 29092 17731 29144 17740
rect 29092 17697 29101 17731
rect 29101 17697 29135 17731
rect 29135 17697 29144 17731
rect 29092 17688 29144 17697
rect 30104 17731 30156 17740
rect 30104 17697 30113 17731
rect 30113 17697 30147 17731
rect 30147 17697 30156 17731
rect 34704 17756 34756 17808
rect 35256 17756 35308 17808
rect 43168 17756 43220 17808
rect 43996 17799 44048 17808
rect 43996 17765 44005 17799
rect 44005 17765 44039 17799
rect 44039 17765 44048 17799
rect 43996 17756 44048 17765
rect 45744 17799 45796 17808
rect 45744 17765 45753 17799
rect 45753 17765 45787 17799
rect 45787 17765 45796 17799
rect 45744 17756 45796 17765
rect 46756 17799 46808 17808
rect 46756 17765 46765 17799
rect 46765 17765 46799 17799
rect 46799 17765 46808 17799
rect 46756 17756 46808 17765
rect 46940 17799 46992 17808
rect 46940 17765 46949 17799
rect 46949 17765 46983 17799
rect 46983 17765 46992 17799
rect 46940 17756 46992 17765
rect 32220 17731 32272 17740
rect 30104 17688 30156 17697
rect 32220 17697 32229 17731
rect 32229 17697 32263 17731
rect 32263 17697 32272 17731
rect 32220 17688 32272 17697
rect 32312 17688 32364 17740
rect 42064 17731 42116 17740
rect 34520 17620 34572 17672
rect 35256 17620 35308 17672
rect 35532 17663 35584 17672
rect 35532 17629 35541 17663
rect 35541 17629 35575 17663
rect 35575 17629 35584 17663
rect 35532 17620 35584 17629
rect 42064 17697 42073 17731
rect 42073 17697 42107 17731
rect 42107 17697 42116 17731
rect 42064 17688 42116 17697
rect 43720 17731 43772 17740
rect 43720 17697 43729 17731
rect 43729 17697 43763 17731
rect 43763 17697 43772 17731
rect 43720 17688 43772 17697
rect 45560 17731 45612 17740
rect 45560 17697 45569 17731
rect 45569 17697 45603 17731
rect 45603 17697 45612 17731
rect 45560 17688 45612 17697
rect 46388 17688 46440 17740
rect 42616 17620 42668 17672
rect 29368 17552 29420 17604
rect 35440 17552 35492 17604
rect 43444 17595 43496 17604
rect 43444 17561 43453 17595
rect 43453 17561 43487 17595
rect 43487 17561 43496 17595
rect 43444 17552 43496 17561
rect 46480 17552 46532 17604
rect 31944 17527 31996 17536
rect 31944 17493 31953 17527
rect 31953 17493 31987 17527
rect 31987 17493 31996 17527
rect 31944 17484 31996 17493
rect 41604 17527 41656 17536
rect 41604 17493 41613 17527
rect 41613 17493 41647 17527
rect 41647 17493 41656 17527
rect 41604 17484 41656 17493
rect 42248 17527 42300 17536
rect 42248 17493 42257 17527
rect 42257 17493 42291 17527
rect 42291 17493 42300 17527
rect 42248 17484 42300 17493
rect 43260 17484 43312 17536
rect 45284 17527 45336 17536
rect 45284 17493 45293 17527
rect 45293 17493 45327 17527
rect 45327 17493 45336 17527
rect 45284 17484 45336 17493
rect 47124 17527 47176 17536
rect 47124 17493 47133 17527
rect 47133 17493 47167 17527
rect 47167 17493 47176 17527
rect 47124 17484 47176 17493
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 34966 17382 35018 17434
rect 35030 17382 35082 17434
rect 35094 17382 35146 17434
rect 35158 17382 35210 17434
rect 30748 17280 30800 17332
rect 26516 17255 26568 17264
rect 26516 17221 26525 17255
rect 26525 17221 26559 17255
rect 26559 17221 26568 17255
rect 26516 17212 26568 17221
rect 30564 17212 30616 17264
rect 32220 17280 32272 17332
rect 34704 17323 34756 17332
rect 34704 17289 34713 17323
rect 34713 17289 34747 17323
rect 34747 17289 34756 17323
rect 34704 17280 34756 17289
rect 35256 17280 35308 17332
rect 42064 17280 42116 17332
rect 42616 17323 42668 17332
rect 42616 17289 42625 17323
rect 42625 17289 42659 17323
rect 42659 17289 42668 17323
rect 42616 17280 42668 17289
rect 42984 17323 43036 17332
rect 42984 17289 42993 17323
rect 42993 17289 43027 17323
rect 43027 17289 43036 17323
rect 42984 17280 43036 17289
rect 43720 17323 43772 17332
rect 43720 17289 43729 17323
rect 43729 17289 43763 17323
rect 43763 17289 43772 17323
rect 43720 17280 43772 17289
rect 44088 17323 44140 17332
rect 44088 17289 44097 17323
rect 44097 17289 44131 17323
rect 44131 17289 44140 17323
rect 44088 17280 44140 17289
rect 45560 17280 45612 17332
rect 46112 17280 46164 17332
rect 46388 17280 46440 17332
rect 35532 17255 35584 17264
rect 35532 17221 35541 17255
rect 35541 17221 35575 17255
rect 35575 17221 35584 17255
rect 35532 17212 35584 17221
rect 31852 17187 31904 17196
rect 31852 17153 31861 17187
rect 31861 17153 31895 17187
rect 31895 17153 31904 17187
rect 31852 17144 31904 17153
rect 41328 17144 41380 17196
rect 41604 17187 41656 17196
rect 41604 17153 41613 17187
rect 41613 17153 41647 17187
rect 41647 17153 41656 17187
rect 41604 17144 41656 17153
rect 23756 17119 23808 17128
rect 23756 17085 23765 17119
rect 23765 17085 23799 17119
rect 23799 17085 23808 17119
rect 23756 17076 23808 17085
rect 26792 17119 26844 17128
rect 26792 17085 26801 17119
rect 26801 17085 26835 17119
rect 26835 17085 26844 17119
rect 26792 17076 26844 17085
rect 27160 17076 27212 17128
rect 30472 17076 30524 17128
rect 31944 17076 31996 17128
rect 23480 17051 23532 17060
rect 23480 17017 23489 17051
rect 23489 17017 23523 17051
rect 23523 17017 23532 17051
rect 23480 17008 23532 17017
rect 26884 17008 26936 17060
rect 25780 16940 25832 16992
rect 29092 16940 29144 16992
rect 30564 16940 30616 16992
rect 37280 17076 37332 17128
rect 42708 17076 42760 17128
rect 42984 17076 43036 17128
rect 44548 17076 44600 17128
rect 37740 17008 37792 17060
rect 40040 17008 40092 17060
rect 45744 17008 45796 17060
rect 46572 17008 46624 17060
rect 32312 16940 32364 16992
rect 38660 16940 38712 16992
rect 44180 16940 44232 16992
rect 19606 16838 19658 16890
rect 19670 16838 19722 16890
rect 19734 16838 19786 16890
rect 19798 16838 19850 16890
rect 31852 16779 31904 16788
rect 26884 16668 26936 16720
rect 27160 16711 27212 16720
rect 27160 16677 27194 16711
rect 27194 16677 27212 16711
rect 29920 16711 29972 16720
rect 27160 16668 27212 16677
rect 29920 16677 29929 16711
rect 29929 16677 29963 16711
rect 29963 16677 29972 16711
rect 29920 16668 29972 16677
rect 23756 16600 23808 16652
rect 28816 16643 28868 16652
rect 28816 16609 28825 16643
rect 28825 16609 28859 16643
rect 28859 16609 28868 16643
rect 28816 16600 28868 16609
rect 30012 16643 30064 16652
rect 30012 16609 30021 16643
rect 30021 16609 30055 16643
rect 30055 16609 30064 16643
rect 30012 16600 30064 16609
rect 25320 16532 25372 16584
rect 26884 16575 26936 16584
rect 26884 16541 26893 16575
rect 26893 16541 26927 16575
rect 26927 16541 26936 16575
rect 26884 16532 26936 16541
rect 29368 16532 29420 16584
rect 31852 16745 31861 16779
rect 31861 16745 31895 16779
rect 31895 16745 31904 16779
rect 31852 16736 31904 16745
rect 31944 16736 31996 16788
rect 33692 16736 33744 16788
rect 37280 16779 37332 16788
rect 37280 16745 37289 16779
rect 37289 16745 37323 16779
rect 37323 16745 37332 16779
rect 37280 16736 37332 16745
rect 39396 16736 39448 16788
rect 34428 16668 34480 16720
rect 38568 16711 38620 16720
rect 38568 16677 38602 16711
rect 38602 16677 38620 16711
rect 38568 16668 38620 16677
rect 41420 16736 41472 16788
rect 42984 16736 43036 16788
rect 45284 16736 45336 16788
rect 46572 16779 46624 16788
rect 46572 16745 46581 16779
rect 46581 16745 46615 16779
rect 46615 16745 46624 16779
rect 46572 16736 46624 16745
rect 46756 16736 46808 16788
rect 42248 16668 42300 16720
rect 43812 16668 43864 16720
rect 32128 16643 32180 16652
rect 32128 16609 32137 16643
rect 32137 16609 32171 16643
rect 32171 16609 32180 16643
rect 32128 16600 32180 16609
rect 32312 16643 32364 16652
rect 32312 16609 32321 16643
rect 32321 16609 32355 16643
rect 32355 16609 32364 16643
rect 32312 16600 32364 16609
rect 33784 16643 33836 16652
rect 33784 16609 33793 16643
rect 33793 16609 33827 16643
rect 33827 16609 33836 16643
rect 33784 16600 33836 16609
rect 34060 16643 34112 16652
rect 34060 16609 34094 16643
rect 34094 16609 34112 16643
rect 43168 16643 43220 16652
rect 34060 16600 34112 16609
rect 43168 16609 43177 16643
rect 43177 16609 43211 16643
rect 43211 16609 43220 16643
rect 43168 16600 43220 16609
rect 43720 16643 43772 16652
rect 43720 16609 43729 16643
rect 43729 16609 43763 16643
rect 43763 16609 43772 16643
rect 43720 16600 43772 16609
rect 45560 16668 45612 16720
rect 46112 16668 46164 16720
rect 45468 16643 45520 16652
rect 45468 16609 45502 16643
rect 45502 16609 45520 16643
rect 45468 16600 45520 16609
rect 30656 16532 30708 16584
rect 38292 16575 38344 16584
rect 38292 16541 38301 16575
rect 38301 16541 38335 16575
rect 38335 16541 38344 16575
rect 38292 16532 38344 16541
rect 40408 16532 40460 16584
rect 40776 16575 40828 16584
rect 40776 16541 40785 16575
rect 40785 16541 40819 16575
rect 40819 16541 40828 16575
rect 40776 16532 40828 16541
rect 43996 16575 44048 16584
rect 43996 16541 44005 16575
rect 44005 16541 44039 16575
rect 44039 16541 44048 16575
rect 43996 16532 44048 16541
rect 29000 16396 29052 16448
rect 30472 16439 30524 16448
rect 30472 16405 30481 16439
rect 30481 16405 30515 16439
rect 30515 16405 30524 16439
rect 30472 16396 30524 16405
rect 31484 16439 31536 16448
rect 31484 16405 31493 16439
rect 31493 16405 31527 16439
rect 31527 16405 31536 16439
rect 31484 16396 31536 16405
rect 33968 16396 34020 16448
rect 44548 16396 44600 16448
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 34966 16294 35018 16346
rect 35030 16294 35082 16346
rect 35094 16294 35146 16346
rect 35158 16294 35210 16346
rect 25320 16235 25372 16244
rect 25320 16201 25329 16235
rect 25329 16201 25363 16235
rect 25363 16201 25372 16235
rect 25320 16192 25372 16201
rect 26792 16192 26844 16244
rect 29000 16235 29052 16244
rect 29000 16201 29009 16235
rect 29009 16201 29043 16235
rect 29043 16201 29052 16235
rect 29000 16192 29052 16201
rect 29368 16235 29420 16244
rect 29368 16201 29377 16235
rect 29377 16201 29411 16235
rect 29411 16201 29420 16235
rect 29368 16192 29420 16201
rect 30380 16235 30432 16244
rect 30380 16201 30389 16235
rect 30389 16201 30423 16235
rect 30423 16201 30432 16235
rect 30380 16192 30432 16201
rect 30472 16192 30524 16244
rect 32312 16192 32364 16244
rect 33784 16192 33836 16244
rect 38660 16235 38712 16244
rect 31760 16124 31812 16176
rect 33508 16124 33560 16176
rect 31300 16099 31352 16108
rect 31300 16065 31309 16099
rect 31309 16065 31343 16099
rect 31343 16065 31352 16099
rect 31300 16056 31352 16065
rect 31484 16099 31536 16108
rect 31484 16065 31493 16099
rect 31493 16065 31527 16099
rect 31527 16065 31536 16099
rect 31484 16056 31536 16065
rect 33692 16099 33744 16108
rect 33692 16065 33701 16099
rect 33701 16065 33735 16099
rect 33735 16065 33744 16099
rect 33692 16056 33744 16065
rect 25780 16031 25832 16040
rect 25780 15997 25814 16031
rect 25814 15997 25832 16031
rect 25780 15988 25832 15997
rect 28816 15988 28868 16040
rect 27620 15920 27672 15972
rect 29552 15920 29604 15972
rect 34060 16124 34112 16176
rect 38660 16201 38669 16235
rect 38669 16201 38703 16235
rect 38703 16201 38712 16235
rect 38660 16192 38712 16201
rect 39948 16192 40000 16244
rect 43812 16235 43864 16244
rect 43812 16201 43821 16235
rect 43821 16201 43855 16235
rect 43855 16201 43864 16235
rect 43812 16192 43864 16201
rect 44548 16235 44600 16244
rect 44548 16201 44557 16235
rect 44557 16201 44591 16235
rect 44591 16201 44600 16235
rect 44548 16192 44600 16201
rect 45560 16235 45612 16244
rect 45560 16201 45569 16235
rect 45569 16201 45603 16235
rect 45603 16201 45612 16235
rect 45560 16192 45612 16201
rect 39396 16099 39448 16108
rect 39396 16065 39405 16099
rect 39405 16065 39439 16099
rect 39439 16065 39448 16099
rect 39396 16056 39448 16065
rect 43996 16056 44048 16108
rect 45284 16056 45336 16108
rect 30288 15920 30340 15972
rect 33968 15920 34020 15972
rect 34336 15920 34388 15972
rect 35716 15920 35768 15972
rect 38660 15920 38712 15972
rect 40776 15988 40828 16040
rect 41236 15988 41288 16040
rect 41420 15988 41472 16040
rect 40868 15920 40920 15972
rect 44548 15920 44600 15972
rect 26608 15852 26660 15904
rect 26884 15852 26936 15904
rect 28172 15852 28224 15904
rect 28356 15895 28408 15904
rect 28356 15861 28365 15895
rect 28365 15861 28399 15895
rect 28399 15861 28408 15895
rect 28356 15852 28408 15861
rect 29000 15852 29052 15904
rect 30380 15852 30432 15904
rect 30564 15852 30616 15904
rect 32128 15852 32180 15904
rect 32956 15852 33008 15904
rect 37924 15852 37976 15904
rect 38292 15895 38344 15904
rect 38292 15861 38301 15895
rect 38301 15861 38335 15895
rect 38335 15861 38344 15895
rect 38292 15852 38344 15861
rect 42064 15895 42116 15904
rect 42064 15861 42073 15895
rect 42073 15861 42107 15895
rect 42107 15861 42116 15895
rect 42064 15852 42116 15861
rect 43168 15895 43220 15904
rect 43168 15861 43177 15895
rect 43177 15861 43211 15895
rect 43211 15861 43220 15895
rect 43168 15852 43220 15861
rect 43444 15895 43496 15904
rect 43444 15861 43453 15895
rect 43453 15861 43487 15895
rect 43487 15861 43496 15895
rect 43444 15852 43496 15861
rect 44272 15895 44324 15904
rect 44272 15861 44281 15895
rect 44281 15861 44315 15895
rect 44315 15861 44324 15895
rect 44272 15852 44324 15861
rect 44824 15852 44876 15904
rect 45560 15920 45612 15972
rect 47492 15988 47544 16040
rect 46572 15920 46624 15972
rect 46388 15852 46440 15904
rect 19606 15750 19658 15802
rect 19670 15750 19722 15802
rect 19734 15750 19786 15802
rect 19798 15750 19850 15802
rect 25780 15648 25832 15700
rect 26792 15648 26844 15700
rect 29552 15691 29604 15700
rect 29552 15657 29561 15691
rect 29561 15657 29595 15691
rect 29595 15657 29604 15691
rect 29552 15648 29604 15657
rect 31300 15691 31352 15700
rect 31300 15657 31309 15691
rect 31309 15657 31343 15691
rect 31343 15657 31352 15691
rect 31300 15648 31352 15657
rect 38660 15648 38712 15700
rect 39396 15648 39448 15700
rect 40776 15648 40828 15700
rect 41236 15691 41288 15700
rect 41236 15657 41245 15691
rect 41245 15657 41279 15691
rect 41279 15657 41288 15691
rect 41236 15648 41288 15657
rect 43444 15648 43496 15700
rect 44180 15648 44232 15700
rect 44548 15691 44600 15700
rect 44548 15657 44557 15691
rect 44557 15657 44591 15691
rect 44591 15657 44600 15691
rect 44548 15648 44600 15657
rect 45468 15648 45520 15700
rect 47492 15691 47544 15700
rect 47492 15657 47501 15691
rect 47501 15657 47535 15691
rect 47535 15657 47544 15691
rect 47492 15648 47544 15657
rect 28632 15580 28684 15632
rect 29000 15580 29052 15632
rect 33048 15580 33100 15632
rect 35256 15580 35308 15632
rect 38200 15580 38252 15632
rect 41144 15580 41196 15632
rect 42064 15580 42116 15632
rect 43076 15580 43128 15632
rect 44088 15580 44140 15632
rect 28172 15555 28224 15564
rect 28172 15521 28181 15555
rect 28181 15521 28215 15555
rect 28215 15521 28224 15555
rect 28172 15512 28224 15521
rect 30656 15555 30708 15564
rect 30656 15521 30665 15555
rect 30665 15521 30699 15555
rect 30699 15521 30708 15555
rect 30656 15512 30708 15521
rect 31300 15512 31352 15564
rect 34796 15512 34848 15564
rect 35716 15512 35768 15564
rect 46112 15555 46164 15564
rect 46112 15521 46121 15555
rect 46121 15521 46155 15555
rect 46155 15521 46164 15555
rect 46112 15512 46164 15521
rect 46388 15555 46440 15564
rect 46388 15521 46422 15555
rect 46422 15521 46440 15555
rect 46388 15512 46440 15521
rect 33508 15487 33560 15496
rect 33508 15453 33517 15487
rect 33517 15453 33551 15487
rect 33551 15453 33560 15487
rect 33508 15444 33560 15453
rect 34428 15444 34480 15496
rect 40868 15444 40920 15496
rect 43996 15487 44048 15496
rect 30656 15308 30708 15360
rect 30840 15351 30892 15360
rect 30840 15317 30849 15351
rect 30849 15317 30883 15351
rect 30883 15317 30892 15351
rect 30840 15308 30892 15317
rect 32312 15351 32364 15360
rect 32312 15317 32321 15351
rect 32321 15317 32355 15351
rect 32355 15317 32364 15351
rect 32312 15308 32364 15317
rect 33140 15308 33192 15360
rect 34428 15351 34480 15360
rect 34428 15317 34437 15351
rect 34437 15317 34471 15351
rect 34471 15317 34480 15351
rect 34428 15308 34480 15317
rect 41328 15308 41380 15360
rect 43996 15453 44005 15487
rect 44005 15453 44039 15487
rect 44039 15453 44048 15487
rect 43996 15444 44048 15453
rect 43260 15376 43312 15428
rect 42340 15308 42392 15360
rect 44824 15351 44876 15360
rect 44824 15317 44833 15351
rect 44833 15317 44867 15351
rect 44867 15317 44876 15351
rect 44824 15308 44876 15317
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 34966 15206 35018 15258
rect 35030 15206 35082 15258
rect 35094 15206 35146 15258
rect 35158 15206 35210 15258
rect 28172 15147 28224 15156
rect 28172 15113 28181 15147
rect 28181 15113 28215 15147
rect 28215 15113 28224 15147
rect 28172 15104 28224 15113
rect 28632 15147 28684 15156
rect 28632 15113 28641 15147
rect 28641 15113 28675 15147
rect 28675 15113 28684 15147
rect 28632 15104 28684 15113
rect 30380 15147 30432 15156
rect 30380 15113 30389 15147
rect 30389 15113 30423 15147
rect 30423 15113 30432 15147
rect 30380 15104 30432 15113
rect 31300 15147 31352 15156
rect 31300 15113 31309 15147
rect 31309 15113 31343 15147
rect 31343 15113 31352 15147
rect 31300 15104 31352 15113
rect 31760 15104 31812 15156
rect 33048 15104 33100 15156
rect 33140 15104 33192 15156
rect 32312 14968 32364 15020
rect 30656 14943 30708 14952
rect 30656 14909 30665 14943
rect 30665 14909 30699 14943
rect 30699 14909 30708 14943
rect 30656 14900 30708 14909
rect 31944 14900 31996 14952
rect 34796 15104 34848 15156
rect 40776 15147 40828 15156
rect 40776 15113 40785 15147
rect 40785 15113 40819 15147
rect 40819 15113 40828 15147
rect 40776 15104 40828 15113
rect 41144 15147 41196 15156
rect 41144 15113 41153 15147
rect 41153 15113 41187 15147
rect 41187 15113 41196 15147
rect 41144 15104 41196 15113
rect 43076 15147 43128 15156
rect 43076 15113 43085 15147
rect 43085 15113 43119 15147
rect 43119 15113 43128 15147
rect 43076 15104 43128 15113
rect 44180 15147 44232 15156
rect 44180 15113 44189 15147
rect 44189 15113 44223 15147
rect 44223 15113 44232 15147
rect 44180 15104 44232 15113
rect 46112 15104 46164 15156
rect 46848 15104 46900 15156
rect 40868 15036 40920 15088
rect 42524 15036 42576 15088
rect 46940 15079 46992 15088
rect 46940 15045 46949 15079
rect 46949 15045 46983 15079
rect 46983 15045 46992 15079
rect 46940 15036 46992 15045
rect 30840 14875 30892 14884
rect 30840 14841 30849 14875
rect 30849 14841 30883 14875
rect 30883 14841 30892 14875
rect 30840 14832 30892 14841
rect 35164 14943 35216 14952
rect 35164 14909 35173 14943
rect 35173 14909 35207 14943
rect 35207 14909 35216 14943
rect 35164 14900 35216 14909
rect 37924 14943 37976 14952
rect 27620 14807 27672 14816
rect 27620 14773 27629 14807
rect 27629 14773 27663 14807
rect 27663 14773 27672 14807
rect 27620 14764 27672 14773
rect 30288 14764 30340 14816
rect 31668 14807 31720 14816
rect 31668 14773 31677 14807
rect 31677 14773 31711 14807
rect 31711 14773 31720 14807
rect 35256 14832 35308 14884
rect 36268 14832 36320 14884
rect 31668 14764 31720 14773
rect 37648 14764 37700 14816
rect 37924 14909 37933 14943
rect 37933 14909 37967 14943
rect 37967 14909 37976 14943
rect 37924 14900 37976 14909
rect 38200 14943 38252 14952
rect 38200 14909 38234 14943
rect 38234 14909 38252 14943
rect 38200 14900 38252 14909
rect 41420 14900 41472 14952
rect 41788 14900 41840 14952
rect 42340 14900 42392 14952
rect 42800 14900 42852 14952
rect 43260 14900 43312 14952
rect 44456 14900 44508 14952
rect 44824 14900 44876 14952
rect 46848 14900 46900 14952
rect 41972 14875 42024 14884
rect 41972 14841 41981 14875
rect 41981 14841 42015 14875
rect 42015 14841 42024 14875
rect 41972 14832 42024 14841
rect 39304 14807 39356 14816
rect 39304 14773 39313 14807
rect 39313 14773 39347 14807
rect 39347 14773 39356 14807
rect 39304 14764 39356 14773
rect 41788 14764 41840 14816
rect 42616 14807 42668 14816
rect 42616 14773 42625 14807
rect 42625 14773 42659 14807
rect 42659 14773 42668 14807
rect 42616 14764 42668 14773
rect 46388 14832 46440 14884
rect 46848 14764 46900 14816
rect 19606 14662 19658 14714
rect 19670 14662 19722 14714
rect 19734 14662 19786 14714
rect 19798 14662 19850 14714
rect 28356 14560 28408 14612
rect 27528 14492 27580 14544
rect 29368 14492 29420 14544
rect 30656 14560 30708 14612
rect 31668 14560 31720 14612
rect 31944 14603 31996 14612
rect 31944 14569 31953 14603
rect 31953 14569 31987 14603
rect 31987 14569 31996 14603
rect 31944 14560 31996 14569
rect 32312 14560 32364 14612
rect 33508 14560 33560 14612
rect 34796 14560 34848 14612
rect 39120 14603 39172 14612
rect 39120 14569 39129 14603
rect 39129 14569 39163 14603
rect 39163 14569 39172 14603
rect 39120 14560 39172 14569
rect 41972 14560 42024 14612
rect 42248 14603 42300 14612
rect 42248 14569 42257 14603
rect 42257 14569 42291 14603
rect 42291 14569 42300 14603
rect 42248 14560 42300 14569
rect 43996 14560 44048 14612
rect 30012 14492 30064 14544
rect 26608 14467 26660 14476
rect 26608 14433 26617 14467
rect 26617 14433 26651 14467
rect 26651 14433 26660 14467
rect 26608 14424 26660 14433
rect 26884 14467 26936 14476
rect 26884 14433 26918 14467
rect 26918 14433 26936 14467
rect 26884 14424 26936 14433
rect 29736 14424 29788 14476
rect 30932 14467 30984 14476
rect 8392 14331 8444 14340
rect 8392 14297 8401 14331
rect 8401 14297 8435 14331
rect 8435 14297 8444 14331
rect 8392 14288 8444 14297
rect 30932 14433 30941 14467
rect 30941 14433 30975 14467
rect 30975 14433 30984 14467
rect 30932 14424 30984 14433
rect 32128 14424 32180 14476
rect 39304 14492 39356 14544
rect 40868 14535 40920 14544
rect 40868 14501 40877 14535
rect 40877 14501 40911 14535
rect 40911 14501 40920 14535
rect 40868 14492 40920 14501
rect 42800 14492 42852 14544
rect 43076 14492 43128 14544
rect 44088 14492 44140 14544
rect 44456 14535 44508 14544
rect 44456 14501 44465 14535
rect 44465 14501 44499 14535
rect 44499 14501 44508 14535
rect 44456 14492 44508 14501
rect 38292 14424 38344 14476
rect 42524 14424 42576 14476
rect 47216 14424 47268 14476
rect 37648 14356 37700 14408
rect 40684 14399 40736 14408
rect 40684 14365 40693 14399
rect 40693 14365 40727 14399
rect 40727 14365 40736 14399
rect 40684 14356 40736 14365
rect 44272 14399 44324 14408
rect 44272 14365 44281 14399
rect 44281 14365 44315 14399
rect 44315 14365 44324 14399
rect 44272 14356 44324 14365
rect 32312 14288 32364 14340
rect 34520 14288 34572 14340
rect 42616 14288 42668 14340
rect 43168 14288 43220 14340
rect 46756 14288 46808 14340
rect 19800 14263 19852 14272
rect 19800 14229 19809 14263
rect 19809 14229 19843 14263
rect 19843 14229 19852 14263
rect 19800 14220 19852 14229
rect 27988 14263 28040 14272
rect 27988 14229 27997 14263
rect 27997 14229 28031 14263
rect 28031 14229 28040 14263
rect 27988 14220 28040 14229
rect 31576 14263 31628 14272
rect 31576 14229 31585 14263
rect 31585 14229 31619 14263
rect 31619 14229 31628 14263
rect 31576 14220 31628 14229
rect 33600 14220 33652 14272
rect 33968 14263 34020 14272
rect 33968 14229 33977 14263
rect 33977 14229 34011 14263
rect 34011 14229 34020 14263
rect 33968 14220 34020 14229
rect 35256 14263 35308 14272
rect 35256 14229 35265 14263
rect 35265 14229 35299 14263
rect 35299 14229 35308 14263
rect 35256 14220 35308 14229
rect 43628 14263 43680 14272
rect 43628 14229 43637 14263
rect 43637 14229 43671 14263
rect 43671 14229 43680 14263
rect 43628 14220 43680 14229
rect 46572 14263 46624 14272
rect 46572 14229 46581 14263
rect 46581 14229 46615 14263
rect 46615 14229 46624 14263
rect 46572 14220 46624 14229
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 34966 14118 35018 14170
rect 35030 14118 35082 14170
rect 35094 14118 35146 14170
rect 35158 14118 35210 14170
rect 26608 14059 26660 14068
rect 26608 14025 26617 14059
rect 26617 14025 26651 14059
rect 26651 14025 26660 14059
rect 26608 14016 26660 14025
rect 26884 14016 26936 14068
rect 29736 14059 29788 14068
rect 29736 14025 29745 14059
rect 29745 14025 29779 14059
rect 29779 14025 29788 14059
rect 29736 14016 29788 14025
rect 30932 14016 30984 14068
rect 36268 14059 36320 14068
rect 36268 14025 36277 14059
rect 36277 14025 36311 14059
rect 36311 14025 36320 14059
rect 36268 14016 36320 14025
rect 39304 14016 39356 14068
rect 41788 14016 41840 14068
rect 42524 14059 42576 14068
rect 42524 14025 42533 14059
rect 42533 14025 42567 14059
rect 42567 14025 42576 14059
rect 42524 14016 42576 14025
rect 43076 14059 43128 14068
rect 43076 14025 43085 14059
rect 43085 14025 43119 14059
rect 43119 14025 43128 14059
rect 43076 14016 43128 14025
rect 44272 14016 44324 14068
rect 47216 14059 47268 14068
rect 47216 14025 47225 14059
rect 47225 14025 47259 14059
rect 47259 14025 47268 14059
rect 47216 14016 47268 14025
rect 19340 13948 19392 14000
rect 29368 13948 29420 14000
rect 20260 13923 20312 13932
rect 20260 13889 20269 13923
rect 20269 13889 20303 13923
rect 20303 13889 20312 13923
rect 20260 13880 20312 13889
rect 28632 13880 28684 13932
rect 30288 13923 30340 13932
rect 8300 13855 8352 13864
rect 8300 13821 8309 13855
rect 8309 13821 8343 13855
rect 8343 13821 8352 13855
rect 8300 13812 8352 13821
rect 8392 13812 8444 13864
rect 20628 13812 20680 13864
rect 27620 13812 27672 13864
rect 30288 13889 30297 13923
rect 30297 13889 30331 13923
rect 30331 13889 30340 13923
rect 30288 13880 30340 13889
rect 19800 13744 19852 13796
rect 27988 13744 28040 13796
rect 31576 13812 31628 13864
rect 32312 13923 32364 13932
rect 32312 13889 32321 13923
rect 32321 13889 32355 13923
rect 32355 13889 32364 13923
rect 32312 13880 32364 13889
rect 32864 13880 32916 13932
rect 33968 13948 34020 14000
rect 34428 13948 34480 14000
rect 40040 13880 40092 13932
rect 32128 13812 32180 13864
rect 33600 13855 33652 13864
rect 33600 13821 33609 13855
rect 33609 13821 33643 13855
rect 33643 13821 33652 13855
rect 33600 13812 33652 13821
rect 34796 13812 34848 13864
rect 35164 13855 35216 13864
rect 35164 13821 35198 13855
rect 35198 13821 35216 13855
rect 31024 13744 31076 13796
rect 33876 13744 33928 13796
rect 35164 13812 35216 13821
rect 35716 13812 35768 13864
rect 37648 13812 37700 13864
rect 46756 13880 46808 13932
rect 35256 13744 35308 13796
rect 36268 13744 36320 13796
rect 39212 13744 39264 13796
rect 41328 13812 41380 13864
rect 40684 13744 40736 13796
rect 4712 13676 4764 13728
rect 8760 13676 8812 13728
rect 27436 13719 27488 13728
rect 27436 13685 27445 13719
rect 27445 13685 27479 13719
rect 27479 13685 27488 13719
rect 43628 13812 43680 13864
rect 45468 13812 45520 13864
rect 46572 13812 46624 13864
rect 44732 13744 44784 13796
rect 47032 13744 47084 13796
rect 28632 13719 28684 13728
rect 27436 13676 27488 13685
rect 28632 13685 28641 13719
rect 28641 13685 28675 13719
rect 28675 13685 28684 13719
rect 28632 13676 28684 13685
rect 29920 13676 29972 13728
rect 32220 13719 32272 13728
rect 32220 13685 32229 13719
rect 32229 13685 32263 13719
rect 32263 13685 32272 13719
rect 32220 13676 32272 13685
rect 33784 13719 33836 13728
rect 33784 13685 33793 13719
rect 33793 13685 33827 13719
rect 33827 13685 33836 13719
rect 33784 13676 33836 13685
rect 37372 13719 37424 13728
rect 37372 13685 37381 13719
rect 37381 13685 37415 13719
rect 37415 13685 37424 13719
rect 37372 13676 37424 13685
rect 38292 13719 38344 13728
rect 38292 13685 38301 13719
rect 38301 13685 38335 13719
rect 38335 13685 38344 13719
rect 38292 13676 38344 13685
rect 43352 13719 43404 13728
rect 43352 13685 43361 13719
rect 43361 13685 43395 13719
rect 43395 13685 43404 13719
rect 43352 13676 43404 13685
rect 44916 13719 44968 13728
rect 44916 13685 44925 13719
rect 44925 13685 44959 13719
rect 44959 13685 44968 13719
rect 44916 13676 44968 13685
rect 46388 13676 46440 13728
rect 19606 13574 19658 13626
rect 19670 13574 19722 13626
rect 19734 13574 19786 13626
rect 19798 13574 19850 13626
rect 4804 13472 4856 13524
rect 5632 13472 5684 13524
rect 29368 13515 29420 13524
rect 29368 13481 29377 13515
rect 29377 13481 29411 13515
rect 29411 13481 29420 13515
rect 29368 13472 29420 13481
rect 31024 13515 31076 13524
rect 31024 13481 31033 13515
rect 31033 13481 31067 13515
rect 31067 13481 31076 13515
rect 31024 13472 31076 13481
rect 33232 13472 33284 13524
rect 34520 13472 34572 13524
rect 40684 13515 40736 13524
rect 40684 13481 40693 13515
rect 40693 13481 40727 13515
rect 40727 13481 40736 13515
rect 40684 13472 40736 13481
rect 43260 13472 43312 13524
rect 44732 13515 44784 13524
rect 44732 13481 44741 13515
rect 44741 13481 44775 13515
rect 44775 13481 44784 13515
rect 44732 13472 44784 13481
rect 46940 13472 46992 13524
rect 4712 13447 4764 13456
rect 4712 13413 4721 13447
rect 4721 13413 4755 13447
rect 4755 13413 4764 13447
rect 4712 13404 4764 13413
rect 2044 13311 2096 13320
rect 2044 13277 2053 13311
rect 2053 13277 2087 13311
rect 2087 13277 2096 13311
rect 2044 13268 2096 13277
rect 4620 13311 4672 13320
rect 4620 13277 4629 13311
rect 4629 13277 4663 13311
rect 4663 13277 4672 13311
rect 4620 13268 4672 13277
rect 1492 13132 1544 13184
rect 4068 13132 4120 13184
rect 19340 13404 19392 13456
rect 27436 13447 27488 13456
rect 27436 13413 27470 13447
rect 27470 13413 27488 13447
rect 27436 13404 27488 13413
rect 29920 13447 29972 13456
rect 29920 13413 29954 13447
rect 29954 13413 29972 13447
rect 29920 13404 29972 13413
rect 32680 13447 32732 13456
rect 32680 13413 32689 13447
rect 32689 13413 32723 13447
rect 32723 13413 32732 13447
rect 32680 13404 32732 13413
rect 32864 13404 32916 13456
rect 35348 13447 35400 13456
rect 35348 13413 35357 13447
rect 35357 13413 35391 13447
rect 35391 13413 35400 13447
rect 35348 13404 35400 13413
rect 38108 13404 38160 13456
rect 39304 13404 39356 13456
rect 42800 13404 42852 13456
rect 6736 13379 6788 13388
rect 6736 13345 6770 13379
rect 6770 13345 6788 13379
rect 19616 13379 19668 13388
rect 6736 13336 6788 13345
rect 19616 13345 19625 13379
rect 19625 13345 19659 13379
rect 19659 13345 19668 13379
rect 19616 13336 19668 13345
rect 26608 13336 26660 13388
rect 27160 13379 27212 13388
rect 27160 13345 27169 13379
rect 27169 13345 27203 13379
rect 27203 13345 27212 13379
rect 27160 13336 27212 13345
rect 33048 13336 33100 13388
rect 33324 13336 33376 13388
rect 6460 13311 6512 13320
rect 6460 13277 6469 13311
rect 6469 13277 6503 13311
rect 6503 13277 6512 13311
rect 6460 13268 6512 13277
rect 18880 13268 18932 13320
rect 29644 13311 29696 13320
rect 29644 13277 29653 13311
rect 29653 13277 29687 13311
rect 29687 13277 29696 13311
rect 29644 13268 29696 13277
rect 36176 13336 36228 13388
rect 46756 13336 46808 13388
rect 36636 13268 36688 13320
rect 37372 13268 37424 13320
rect 38200 13311 38252 13320
rect 38200 13277 38209 13311
rect 38209 13277 38243 13311
rect 38243 13277 38252 13311
rect 38200 13268 38252 13277
rect 38292 13268 38344 13320
rect 39212 13268 39264 13320
rect 43352 13311 43404 13320
rect 43352 13277 43361 13311
rect 43361 13277 43395 13311
rect 43395 13277 43404 13311
rect 43352 13268 43404 13277
rect 46112 13311 46164 13320
rect 46112 13277 46121 13311
rect 46121 13277 46155 13311
rect 46155 13277 46164 13311
rect 46112 13268 46164 13277
rect 32220 13243 32272 13252
rect 32220 13209 32229 13243
rect 32229 13209 32263 13243
rect 32263 13209 32272 13243
rect 32220 13200 32272 13209
rect 37832 13243 37884 13252
rect 37832 13209 37841 13243
rect 37841 13209 37875 13243
rect 37875 13209 37884 13243
rect 37832 13200 37884 13209
rect 7196 13132 7248 13184
rect 7380 13132 7432 13184
rect 20352 13132 20404 13184
rect 28632 13132 28684 13184
rect 32772 13132 32824 13184
rect 33876 13132 33928 13184
rect 36176 13175 36228 13184
rect 36176 13141 36185 13175
rect 36185 13141 36219 13175
rect 36219 13141 36228 13175
rect 36176 13132 36228 13141
rect 36912 13175 36964 13184
rect 36912 13141 36921 13175
rect 36921 13141 36955 13175
rect 36955 13141 36964 13175
rect 36912 13132 36964 13141
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 34966 13030 35018 13082
rect 35030 13030 35082 13082
rect 35094 13030 35146 13082
rect 35158 13030 35210 13082
rect 5632 12971 5684 12980
rect 5632 12937 5641 12971
rect 5641 12937 5675 12971
rect 5675 12937 5684 12971
rect 5632 12928 5684 12937
rect 6460 12971 6512 12980
rect 6460 12937 6469 12971
rect 6469 12937 6503 12971
rect 6503 12937 6512 12971
rect 6460 12928 6512 12937
rect 7656 12928 7708 12980
rect 19432 12928 19484 12980
rect 19616 12928 19668 12980
rect 27160 12971 27212 12980
rect 27160 12937 27169 12971
rect 27169 12937 27203 12971
rect 27203 12937 27212 12971
rect 27160 12928 27212 12937
rect 27436 12928 27488 12980
rect 29920 12928 29972 12980
rect 32680 12928 32732 12980
rect 36268 12971 36320 12980
rect 36268 12937 36277 12971
rect 36277 12937 36311 12971
rect 36311 12937 36320 12971
rect 36268 12928 36320 12937
rect 38200 12928 38252 12980
rect 39304 12928 39356 12980
rect 6920 12903 6972 12912
rect 6920 12869 6929 12903
rect 6929 12869 6963 12903
rect 6963 12869 6972 12903
rect 6920 12860 6972 12869
rect 31760 12860 31812 12912
rect 32864 12860 32916 12912
rect 39212 12860 39264 12912
rect 39948 12860 40000 12912
rect 43352 12928 43404 12980
rect 44088 12971 44140 12980
rect 44088 12937 44097 12971
rect 44097 12937 44131 12971
rect 44131 12937 44140 12971
rect 44088 12928 44140 12937
rect 42800 12860 42852 12912
rect 6828 12792 6880 12844
rect 7380 12835 7432 12844
rect 7380 12801 7389 12835
rect 7389 12801 7423 12835
rect 7423 12801 7432 12835
rect 7380 12792 7432 12801
rect 20352 12835 20404 12844
rect 20352 12801 20361 12835
rect 20361 12801 20395 12835
rect 20395 12801 20404 12835
rect 20352 12792 20404 12801
rect 41512 12835 41564 12844
rect 41512 12801 41521 12835
rect 41521 12801 41555 12835
rect 41555 12801 41564 12835
rect 41512 12792 41564 12801
rect 44548 12835 44600 12844
rect 44548 12801 44557 12835
rect 44557 12801 44591 12835
rect 44591 12801 44600 12835
rect 44548 12792 44600 12801
rect 44916 12792 44968 12844
rect 1492 12767 1544 12776
rect 1492 12733 1501 12767
rect 1501 12733 1535 12767
rect 1535 12733 1544 12767
rect 1492 12724 1544 12733
rect 2044 12724 2096 12776
rect 4160 12767 4212 12776
rect 4160 12733 4169 12767
rect 4169 12733 4203 12767
rect 4203 12733 4212 12767
rect 4160 12724 4212 12733
rect 6460 12724 6512 12776
rect 7012 12724 7064 12776
rect 7196 12724 7248 12776
rect 8300 12724 8352 12776
rect 8760 12767 8812 12776
rect 5540 12656 5592 12708
rect 2688 12588 2740 12640
rect 6736 12588 6788 12640
rect 7656 12588 7708 12640
rect 8760 12733 8794 12767
rect 8794 12733 8812 12767
rect 8760 12724 8812 12733
rect 19984 12724 20036 12776
rect 20260 12724 20312 12776
rect 32128 12724 32180 12776
rect 32772 12724 32824 12776
rect 33232 12767 33284 12776
rect 33232 12733 33266 12767
rect 33266 12733 33284 12767
rect 33232 12724 33284 12733
rect 34612 12724 34664 12776
rect 36820 12767 36872 12776
rect 36820 12733 36829 12767
rect 36829 12733 36863 12767
rect 36863 12733 36872 12767
rect 36820 12724 36872 12733
rect 36912 12724 36964 12776
rect 41788 12767 41840 12776
rect 9588 12588 9640 12640
rect 18880 12631 18932 12640
rect 18880 12597 18889 12631
rect 18889 12597 18923 12631
rect 18923 12597 18932 12631
rect 18880 12588 18932 12597
rect 20444 12588 20496 12640
rect 20720 12588 20772 12640
rect 29644 12631 29696 12640
rect 29644 12597 29653 12631
rect 29653 12597 29687 12631
rect 29687 12597 29696 12631
rect 29644 12588 29696 12597
rect 31024 12631 31076 12640
rect 31024 12597 31033 12631
rect 31033 12597 31067 12631
rect 31067 12597 31076 12631
rect 33784 12656 33836 12708
rect 35256 12656 35308 12708
rect 37188 12656 37240 12708
rect 41788 12733 41822 12767
rect 41822 12733 41840 12767
rect 41788 12724 41840 12733
rect 43352 12724 43404 12776
rect 44088 12724 44140 12776
rect 45468 12928 45520 12980
rect 46756 12928 46808 12980
rect 46112 12767 46164 12776
rect 31024 12588 31076 12597
rect 33232 12588 33284 12640
rect 38200 12631 38252 12640
rect 38200 12597 38209 12631
rect 38209 12597 38243 12631
rect 38243 12597 38252 12631
rect 38200 12588 38252 12597
rect 41328 12588 41380 12640
rect 41512 12588 41564 12640
rect 44088 12588 44140 12640
rect 44732 12588 44784 12640
rect 45560 12631 45612 12640
rect 45560 12597 45569 12631
rect 45569 12597 45603 12631
rect 45603 12597 45612 12631
rect 46112 12733 46121 12767
rect 46121 12733 46155 12767
rect 46155 12733 46164 12767
rect 46112 12724 46164 12733
rect 46388 12767 46440 12776
rect 46388 12733 46422 12767
rect 46422 12733 46440 12767
rect 46388 12724 46440 12733
rect 45560 12588 45612 12597
rect 19606 12486 19658 12538
rect 19670 12486 19722 12538
rect 19734 12486 19786 12538
rect 19798 12486 19850 12538
rect 4620 12384 4672 12436
rect 5540 12384 5592 12436
rect 6828 12384 6880 12436
rect 7656 12427 7708 12436
rect 7656 12393 7665 12427
rect 7665 12393 7699 12427
rect 7699 12393 7708 12427
rect 7656 12384 7708 12393
rect 8760 12384 8812 12436
rect 19340 12427 19392 12436
rect 19340 12393 19349 12427
rect 19349 12393 19383 12427
rect 19383 12393 19392 12427
rect 19340 12384 19392 12393
rect 19432 12384 19484 12436
rect 20260 12384 20312 12436
rect 22284 12427 22336 12436
rect 22284 12393 22293 12427
rect 22293 12393 22327 12427
rect 22327 12393 22336 12427
rect 22284 12384 22336 12393
rect 29920 12384 29972 12436
rect 31668 12384 31720 12436
rect 33140 12384 33192 12436
rect 34244 12384 34296 12436
rect 35256 12384 35308 12436
rect 38200 12384 38252 12436
rect 41052 12384 41104 12436
rect 44088 12427 44140 12436
rect 44088 12393 44097 12427
rect 44097 12393 44131 12427
rect 44131 12393 44140 12427
rect 44088 12384 44140 12393
rect 47032 12384 47084 12436
rect 2320 12316 2372 12368
rect 2688 12316 2740 12368
rect 4804 12316 4856 12368
rect 7104 12359 7156 12368
rect 7104 12325 7113 12359
rect 7113 12325 7147 12359
rect 7147 12325 7156 12359
rect 7104 12316 7156 12325
rect 18236 12316 18288 12368
rect 20628 12316 20680 12368
rect 20812 12316 20864 12368
rect 21364 12316 21416 12368
rect 29644 12316 29696 12368
rect 32680 12316 32732 12368
rect 36820 12316 36872 12368
rect 37648 12316 37700 12368
rect 38568 12359 38620 12368
rect 38568 12325 38577 12359
rect 38577 12325 38611 12359
rect 38611 12325 38620 12359
rect 38568 12316 38620 12325
rect 39764 12316 39816 12368
rect 45008 12316 45060 12368
rect 45468 12316 45520 12368
rect 1492 12291 1544 12300
rect 1492 12257 1501 12291
rect 1501 12257 1535 12291
rect 1535 12257 1544 12291
rect 1492 12248 1544 12257
rect 4160 12248 4212 12300
rect 6920 12291 6972 12300
rect 6920 12257 6929 12291
rect 6929 12257 6963 12291
rect 6963 12257 6972 12291
rect 6920 12248 6972 12257
rect 9956 12291 10008 12300
rect 9956 12257 9990 12291
rect 9990 12257 10008 12291
rect 9956 12248 10008 12257
rect 17868 12248 17920 12300
rect 19892 12248 19944 12300
rect 27160 12248 27212 12300
rect 28356 12291 28408 12300
rect 28356 12257 28365 12291
rect 28365 12257 28399 12291
rect 28399 12257 28408 12291
rect 28356 12248 28408 12257
rect 28632 12291 28684 12300
rect 28632 12257 28666 12291
rect 28666 12257 28684 12291
rect 28632 12248 28684 12257
rect 38384 12291 38436 12300
rect 3976 12180 4028 12232
rect 38384 12257 38393 12291
rect 38393 12257 38427 12291
rect 38427 12257 38436 12291
rect 38384 12248 38436 12257
rect 41512 12248 41564 12300
rect 44548 12248 44600 12300
rect 45284 12291 45336 12300
rect 45284 12257 45318 12291
rect 45318 12257 45336 12291
rect 45284 12248 45336 12257
rect 47492 12291 47544 12300
rect 47492 12257 47501 12291
rect 47501 12257 47535 12291
rect 47535 12257 47544 12291
rect 47492 12248 47544 12257
rect 6460 12180 6512 12232
rect 9680 12223 9732 12232
rect 9680 12189 9689 12223
rect 9689 12189 9723 12223
rect 9723 12189 9732 12223
rect 9680 12180 9732 12189
rect 18512 12180 18564 12232
rect 20904 12223 20956 12232
rect 20904 12189 20913 12223
rect 20913 12189 20947 12223
rect 20947 12189 20956 12223
rect 20904 12180 20956 12189
rect 32128 12223 32180 12232
rect 32128 12189 32137 12223
rect 32137 12189 32171 12223
rect 32171 12189 32180 12223
rect 32128 12180 32180 12189
rect 33876 12180 33928 12232
rect 34612 12223 34664 12232
rect 34612 12189 34621 12223
rect 34621 12189 34655 12223
rect 34655 12189 34664 12223
rect 34612 12180 34664 12189
rect 37280 12180 37332 12232
rect 39028 12180 39080 12232
rect 40040 12223 40092 12232
rect 40040 12189 40049 12223
rect 40049 12189 40083 12223
rect 40083 12189 40092 12223
rect 40040 12180 40092 12189
rect 40224 12223 40276 12232
rect 40224 12189 40233 12223
rect 40233 12189 40267 12223
rect 40267 12189 40276 12223
rect 40224 12180 40276 12189
rect 45008 12223 45060 12232
rect 45008 12189 45017 12223
rect 45017 12189 45051 12223
rect 45051 12189 45060 12223
rect 45008 12180 45060 12189
rect 38108 12155 38160 12164
rect 38108 12121 38117 12155
rect 38117 12121 38151 12155
rect 38151 12121 38160 12155
rect 38108 12112 38160 12121
rect 46388 12155 46440 12164
rect 46388 12121 46397 12155
rect 46397 12121 46431 12155
rect 46431 12121 46440 12155
rect 46388 12112 46440 12121
rect 2872 12087 2924 12096
rect 2872 12053 2881 12087
rect 2881 12053 2915 12087
rect 2915 12053 2924 12087
rect 2872 12044 2924 12053
rect 3884 12044 3936 12096
rect 5540 12044 5592 12096
rect 11244 12044 11296 12096
rect 13636 12087 13688 12096
rect 13636 12053 13645 12087
rect 13645 12053 13679 12087
rect 13679 12053 13688 12087
rect 13636 12044 13688 12053
rect 16028 12087 16080 12096
rect 16028 12053 16037 12087
rect 16037 12053 16071 12087
rect 16071 12053 16080 12087
rect 16028 12044 16080 12053
rect 18604 12044 18656 12096
rect 19248 12044 19300 12096
rect 19984 12044 20036 12096
rect 20444 12087 20496 12096
rect 20444 12053 20453 12087
rect 20453 12053 20487 12087
rect 20487 12053 20496 12087
rect 20444 12044 20496 12053
rect 23572 12044 23624 12096
rect 33232 12044 33284 12096
rect 39672 12087 39724 12096
rect 39672 12053 39681 12087
rect 39681 12053 39715 12087
rect 39715 12053 39724 12087
rect 39672 12044 39724 12053
rect 40868 12087 40920 12096
rect 40868 12053 40877 12087
rect 40877 12053 40911 12087
rect 40911 12053 40920 12087
rect 40868 12044 40920 12053
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 34966 11942 35018 11994
rect 35030 11942 35082 11994
rect 35094 11942 35146 11994
rect 35158 11942 35210 11994
rect 1492 11840 1544 11892
rect 2872 11883 2924 11892
rect 2872 11849 2881 11883
rect 2881 11849 2915 11883
rect 2915 11849 2924 11883
rect 2872 11840 2924 11849
rect 3976 11840 4028 11892
rect 4804 11883 4856 11892
rect 4804 11849 4813 11883
rect 4813 11849 4847 11883
rect 4847 11849 4856 11883
rect 4804 11840 4856 11849
rect 5540 11883 5592 11892
rect 5540 11849 5549 11883
rect 5549 11849 5583 11883
rect 5583 11849 5592 11883
rect 5540 11840 5592 11849
rect 6920 11840 6972 11892
rect 9956 11840 10008 11892
rect 17868 11883 17920 11892
rect 17868 11849 17877 11883
rect 17877 11849 17911 11883
rect 17911 11849 17920 11883
rect 17868 11840 17920 11849
rect 18236 11883 18288 11892
rect 18236 11849 18245 11883
rect 18245 11849 18279 11883
rect 18279 11849 18288 11883
rect 18236 11840 18288 11849
rect 21364 11883 21416 11892
rect 21364 11849 21373 11883
rect 21373 11849 21407 11883
rect 21407 11849 21416 11883
rect 21364 11840 21416 11849
rect 25044 11883 25096 11892
rect 25044 11849 25053 11883
rect 25053 11849 25087 11883
rect 25087 11849 25096 11883
rect 25044 11840 25096 11849
rect 28356 11883 28408 11892
rect 28356 11849 28365 11883
rect 28365 11849 28399 11883
rect 28399 11849 28408 11883
rect 28356 11840 28408 11849
rect 28632 11840 28684 11892
rect 32128 11883 32180 11892
rect 32128 11849 32137 11883
rect 32137 11849 32171 11883
rect 32171 11849 32180 11883
rect 32128 11840 32180 11849
rect 32680 11840 32732 11892
rect 34244 11883 34296 11892
rect 34244 11849 34253 11883
rect 34253 11849 34287 11883
rect 34287 11849 34296 11883
rect 34244 11840 34296 11849
rect 34612 11883 34664 11892
rect 34612 11849 34621 11883
rect 34621 11849 34655 11883
rect 34655 11849 34664 11883
rect 34612 11840 34664 11849
rect 35256 11840 35308 11892
rect 39028 11883 39080 11892
rect 39028 11849 39037 11883
rect 39037 11849 39071 11883
rect 39071 11849 39080 11883
rect 39028 11840 39080 11849
rect 39764 11840 39816 11892
rect 40040 11883 40092 11892
rect 40040 11849 40049 11883
rect 40049 11849 40083 11883
rect 40083 11849 40092 11883
rect 40040 11840 40092 11849
rect 45284 11840 45336 11892
rect 47492 11883 47544 11892
rect 47492 11849 47501 11883
rect 47501 11849 47535 11883
rect 47535 11849 47544 11883
rect 47492 11840 47544 11849
rect 2780 11772 2832 11824
rect 2412 11704 2464 11756
rect 3424 11815 3476 11824
rect 3424 11781 3433 11815
rect 3433 11781 3467 11815
rect 3467 11781 3476 11815
rect 3424 11772 3476 11781
rect 7104 11772 7156 11824
rect 12440 11772 12492 11824
rect 20904 11772 20956 11824
rect 22192 11772 22244 11824
rect 34520 11772 34572 11824
rect 7656 11704 7708 11756
rect 8760 11704 8812 11756
rect 9680 11704 9732 11756
rect 11888 11704 11940 11756
rect 13544 11747 13596 11756
rect 13544 11713 13553 11747
rect 13553 11713 13587 11747
rect 13587 11713 13596 11747
rect 13544 11704 13596 11713
rect 16028 11704 16080 11756
rect 23664 11747 23716 11756
rect 23664 11713 23673 11747
rect 23673 11713 23707 11747
rect 23707 11713 23716 11747
rect 23664 11704 23716 11713
rect 37648 11747 37700 11756
rect 37648 11713 37657 11747
rect 37657 11713 37691 11747
rect 37691 11713 37700 11747
rect 37648 11704 37700 11713
rect 11152 11636 11204 11688
rect 12348 11636 12400 11688
rect 13636 11636 13688 11688
rect 2320 11611 2372 11620
rect 2320 11577 2329 11611
rect 2329 11577 2363 11611
rect 2363 11577 2372 11611
rect 2320 11568 2372 11577
rect 2688 11568 2740 11620
rect 2780 11568 2832 11620
rect 3976 11611 4028 11620
rect 3976 11577 3985 11611
rect 3985 11577 4019 11611
rect 4019 11577 4028 11611
rect 3976 11568 4028 11577
rect 7196 11568 7248 11620
rect 7840 11568 7892 11620
rect 4068 11500 4120 11552
rect 5816 11543 5868 11552
rect 5816 11509 5825 11543
rect 5825 11509 5859 11543
rect 5859 11509 5868 11543
rect 5816 11500 5868 11509
rect 8392 11500 8444 11552
rect 14924 11543 14976 11552
rect 14924 11509 14933 11543
rect 14933 11509 14967 11543
rect 14967 11509 14976 11543
rect 14924 11500 14976 11509
rect 15476 11543 15528 11552
rect 15476 11509 15485 11543
rect 15485 11509 15519 11543
rect 15519 11509 15528 11543
rect 15476 11500 15528 11509
rect 15844 11543 15896 11552
rect 15844 11509 15853 11543
rect 15853 11509 15887 11543
rect 15887 11509 15896 11543
rect 15844 11500 15896 11509
rect 18144 11500 18196 11552
rect 19248 11611 19300 11620
rect 19248 11577 19282 11611
rect 19282 11577 19300 11611
rect 19248 11568 19300 11577
rect 23572 11568 23624 11620
rect 20628 11500 20680 11552
rect 42708 11636 42760 11688
rect 40868 11568 40920 11620
rect 36084 11500 36136 11552
rect 41144 11543 41196 11552
rect 41144 11509 41153 11543
rect 41153 11509 41187 11543
rect 41187 11509 41196 11543
rect 41144 11500 41196 11509
rect 41512 11500 41564 11552
rect 44180 11500 44232 11552
rect 45008 11543 45060 11552
rect 45008 11509 45017 11543
rect 45017 11509 45051 11543
rect 45051 11509 45060 11543
rect 45008 11500 45060 11509
rect 19606 11398 19658 11450
rect 19670 11398 19722 11450
rect 19734 11398 19786 11450
rect 19798 11398 19850 11450
rect 2412 11339 2464 11348
rect 2412 11305 2421 11339
rect 2421 11305 2455 11339
rect 2455 11305 2464 11339
rect 2412 11296 2464 11305
rect 2688 11339 2740 11348
rect 2688 11305 2697 11339
rect 2697 11305 2731 11339
rect 2731 11305 2740 11339
rect 2688 11296 2740 11305
rect 2780 11296 2832 11348
rect 5448 11339 5500 11348
rect 5448 11305 5481 11339
rect 5481 11305 5500 11339
rect 5448 11296 5500 11305
rect 5816 11296 5868 11348
rect 7656 11296 7708 11348
rect 13084 11296 13136 11348
rect 13636 11296 13688 11348
rect 15844 11296 15896 11348
rect 37280 11296 37332 11348
rect 38384 11339 38436 11348
rect 38384 11305 38393 11339
rect 38393 11305 38427 11339
rect 38427 11305 38436 11339
rect 38384 11296 38436 11305
rect 38568 11296 38620 11348
rect 40868 11296 40920 11348
rect 2320 11228 2372 11280
rect 3424 11160 3476 11212
rect 4620 11160 4672 11212
rect 10692 11160 10744 11212
rect 11888 11228 11940 11280
rect 14924 11228 14976 11280
rect 16028 11228 16080 11280
rect 26240 11228 26292 11280
rect 27528 11228 27580 11280
rect 33692 11228 33744 11280
rect 34244 11228 34296 11280
rect 11612 11203 11664 11212
rect 11612 11169 11646 11203
rect 11646 11169 11664 11203
rect 11612 11160 11664 11169
rect 13544 11160 13596 11212
rect 15660 11203 15712 11212
rect 15660 11169 15669 11203
rect 15669 11169 15703 11203
rect 15703 11169 15712 11203
rect 15660 11160 15712 11169
rect 18420 11203 18472 11212
rect 18420 11169 18454 11203
rect 18454 11169 18472 11203
rect 5908 11092 5960 11144
rect 5540 11024 5592 11076
rect 6460 11067 6512 11076
rect 4988 10956 5040 11008
rect 5448 10956 5500 11008
rect 6460 11033 6469 11067
rect 6469 11033 6503 11067
rect 6503 11033 6512 11067
rect 6460 11024 6512 11033
rect 7472 11024 7524 11076
rect 10416 11067 10468 11076
rect 10416 11033 10425 11067
rect 10425 11033 10459 11067
rect 10459 11033 10468 11067
rect 10416 11024 10468 11033
rect 18420 11160 18472 11169
rect 18144 11135 18196 11144
rect 18144 11101 18153 11135
rect 18153 11101 18187 11135
rect 18187 11101 18196 11135
rect 18144 11092 18196 11101
rect 7196 10956 7248 11008
rect 7840 10999 7892 11008
rect 7840 10965 7849 10999
rect 7849 10965 7883 10999
rect 7883 10965 7892 10999
rect 7840 10956 7892 10965
rect 8484 10999 8536 11008
rect 8484 10965 8493 10999
rect 8493 10965 8527 10999
rect 8527 10965 8536 10999
rect 8484 10956 8536 10965
rect 17776 10956 17828 11008
rect 18512 10956 18564 11008
rect 19248 11024 19300 11076
rect 20904 11024 20956 11076
rect 20720 10956 20772 11008
rect 26608 11203 26660 11212
rect 26608 11169 26617 11203
rect 26617 11169 26651 11203
rect 26651 11169 26660 11203
rect 26608 11160 26660 11169
rect 27160 11160 27212 11212
rect 28356 11160 28408 11212
rect 29644 11160 29696 11212
rect 33968 11160 34020 11212
rect 37740 11203 37792 11212
rect 37740 11169 37749 11203
rect 37749 11169 37783 11203
rect 37783 11169 37792 11203
rect 37740 11160 37792 11169
rect 39672 11160 39724 11212
rect 41328 11228 41380 11280
rect 43628 11228 43680 11280
rect 40960 11203 41012 11212
rect 40960 11169 40994 11203
rect 40994 11169 41012 11203
rect 40960 11160 41012 11169
rect 43076 11160 43128 11212
rect 22192 11135 22244 11144
rect 22192 11101 22201 11135
rect 22201 11101 22235 11135
rect 22235 11101 22244 11135
rect 22192 11092 22244 11101
rect 23572 11067 23624 11076
rect 22192 10956 22244 11008
rect 23112 10956 23164 11008
rect 23572 11033 23581 11067
rect 23581 11033 23615 11067
rect 23615 11033 23624 11067
rect 23572 11024 23624 11033
rect 27988 11067 28040 11076
rect 27988 11033 27997 11067
rect 27997 11033 28031 11067
rect 28031 11033 28040 11067
rect 27988 11024 28040 11033
rect 30472 11067 30524 11076
rect 30472 11033 30481 11067
rect 30481 11033 30515 11067
rect 30515 11033 30524 11067
rect 30472 11024 30524 11033
rect 40224 11024 40276 11076
rect 40592 11024 40644 11076
rect 43168 11067 43220 11076
rect 43168 11033 43177 11067
rect 43177 11033 43211 11067
rect 43211 11033 43220 11067
rect 43168 11024 43220 11033
rect 35348 10956 35400 11008
rect 39580 10956 39632 11008
rect 43444 10999 43496 11008
rect 43444 10965 43453 10999
rect 43453 10965 43487 10999
rect 43487 10965 43496 10999
rect 43444 10956 43496 10965
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 34966 10854 35018 10906
rect 35030 10854 35082 10906
rect 35094 10854 35146 10906
rect 35158 10854 35210 10906
rect 4620 10752 4672 10804
rect 4988 10795 5040 10804
rect 4988 10761 4997 10795
rect 4997 10761 5031 10795
rect 5031 10761 5040 10795
rect 4988 10752 5040 10761
rect 5264 10795 5316 10804
rect 5264 10761 5273 10795
rect 5273 10761 5307 10795
rect 5307 10761 5316 10795
rect 5264 10752 5316 10761
rect 5816 10752 5868 10804
rect 11060 10795 11112 10804
rect 11060 10761 11069 10795
rect 11069 10761 11103 10795
rect 11103 10761 11112 10795
rect 11060 10752 11112 10761
rect 11888 10795 11940 10804
rect 11888 10761 11897 10795
rect 11897 10761 11931 10795
rect 11931 10761 11940 10795
rect 11888 10752 11940 10761
rect 12532 10795 12584 10804
rect 12532 10761 12541 10795
rect 12541 10761 12575 10795
rect 12575 10761 12584 10795
rect 12532 10752 12584 10761
rect 15660 10795 15712 10804
rect 15660 10761 15669 10795
rect 15669 10761 15703 10795
rect 15703 10761 15712 10795
rect 15660 10752 15712 10761
rect 16028 10795 16080 10804
rect 16028 10761 16037 10795
rect 16037 10761 16071 10795
rect 16071 10761 16080 10795
rect 16028 10752 16080 10761
rect 18420 10752 18472 10804
rect 22284 10752 22336 10804
rect 26148 10752 26200 10804
rect 27252 10795 27304 10804
rect 27252 10761 27261 10795
rect 27261 10761 27295 10795
rect 27295 10761 27304 10795
rect 27252 10752 27304 10761
rect 29644 10752 29696 10804
rect 33876 10795 33928 10804
rect 33876 10761 33885 10795
rect 33885 10761 33919 10795
rect 33919 10761 33928 10795
rect 33876 10752 33928 10761
rect 34244 10795 34296 10804
rect 34244 10761 34253 10795
rect 34253 10761 34287 10795
rect 34287 10761 34296 10795
rect 34244 10752 34296 10761
rect 37740 10752 37792 10804
rect 6920 10727 6972 10736
rect 6920 10693 6929 10727
rect 6929 10693 6963 10727
rect 6963 10693 6972 10727
rect 6920 10684 6972 10693
rect 11428 10727 11480 10736
rect 11428 10693 11437 10727
rect 11437 10693 11471 10727
rect 11471 10693 11480 10727
rect 11428 10684 11480 10693
rect 19248 10684 19300 10736
rect 34796 10684 34848 10736
rect 39672 10752 39724 10804
rect 40960 10752 41012 10804
rect 41512 10795 41564 10804
rect 41512 10761 41521 10795
rect 41521 10761 41555 10795
rect 41555 10761 41564 10795
rect 41512 10752 41564 10761
rect 43076 10752 43128 10804
rect 1492 10616 1544 10668
rect 7472 10659 7524 10668
rect 7472 10625 7481 10659
rect 7481 10625 7515 10659
rect 7515 10625 7524 10659
rect 7472 10616 7524 10625
rect 11060 10616 11112 10668
rect 11612 10616 11664 10668
rect 13084 10659 13136 10668
rect 13084 10625 13093 10659
rect 13093 10625 13127 10659
rect 13127 10625 13136 10659
rect 13084 10616 13136 10625
rect 20260 10616 20312 10668
rect 20904 10616 20956 10668
rect 28356 10616 28408 10668
rect 29276 10659 29328 10668
rect 29276 10625 29285 10659
rect 29285 10625 29319 10659
rect 29319 10625 29328 10659
rect 29276 10616 29328 10625
rect 39764 10684 39816 10736
rect 41328 10684 41380 10736
rect 2412 10548 2464 10600
rect 5540 10591 5592 10600
rect 5540 10557 5549 10591
rect 5549 10557 5583 10591
rect 5583 10557 5592 10591
rect 5540 10548 5592 10557
rect 7196 10591 7248 10600
rect 7196 10557 7205 10591
rect 7205 10557 7239 10591
rect 7239 10557 7248 10591
rect 7196 10548 7248 10557
rect 5908 10480 5960 10532
rect 8484 10548 8536 10600
rect 11152 10548 11204 10600
rect 12440 10548 12492 10600
rect 18512 10548 18564 10600
rect 20444 10548 20496 10600
rect 37832 10548 37884 10600
rect 9680 10480 9732 10532
rect 12992 10523 13044 10532
rect 12992 10489 13001 10523
rect 13001 10489 13035 10523
rect 13035 10489 13044 10523
rect 12992 10480 13044 10489
rect 17868 10480 17920 10532
rect 18604 10523 18656 10532
rect 18604 10489 18613 10523
rect 18613 10489 18647 10523
rect 18647 10489 18656 10523
rect 18604 10480 18656 10489
rect 26056 10480 26108 10532
rect 29552 10523 29604 10532
rect 29552 10489 29586 10523
rect 29586 10489 29604 10523
rect 29552 10480 29604 10489
rect 35348 10480 35400 10532
rect 39212 10523 39264 10532
rect 39212 10489 39221 10523
rect 39221 10489 39255 10523
rect 39255 10489 39264 10523
rect 39212 10480 39264 10489
rect 39580 10480 39632 10532
rect 41788 10523 41840 10532
rect 41788 10489 41797 10523
rect 41797 10489 41831 10523
rect 41831 10489 41840 10523
rect 41788 10480 41840 10489
rect 42064 10523 42116 10532
rect 42064 10489 42073 10523
rect 42073 10489 42107 10523
rect 42107 10489 42116 10523
rect 42064 10480 42116 10489
rect 43628 10523 43680 10532
rect 43628 10489 43662 10523
rect 43662 10489 43680 10523
rect 43628 10480 43680 10489
rect 2504 10412 2556 10464
rect 5264 10412 5316 10464
rect 6552 10412 6604 10464
rect 9772 10455 9824 10464
rect 9772 10421 9781 10455
rect 9781 10421 9815 10455
rect 9815 10421 9824 10455
rect 9772 10412 9824 10421
rect 10692 10412 10744 10464
rect 17776 10455 17828 10464
rect 17776 10421 17785 10455
rect 17785 10421 17819 10455
rect 17819 10421 17828 10455
rect 17776 10412 17828 10421
rect 20996 10412 21048 10464
rect 21456 10412 21508 10464
rect 23020 10412 23072 10464
rect 36360 10455 36412 10464
rect 36360 10421 36369 10455
rect 36369 10421 36403 10455
rect 36403 10421 36412 10455
rect 36360 10412 36412 10421
rect 41972 10455 42024 10464
rect 41972 10421 41981 10455
rect 41981 10421 42015 10455
rect 42015 10421 42024 10455
rect 41972 10412 42024 10421
rect 44088 10412 44140 10464
rect 19606 10310 19658 10362
rect 19670 10310 19722 10362
rect 19734 10310 19786 10362
rect 19798 10310 19850 10362
rect 1492 10208 1544 10260
rect 2504 10251 2556 10260
rect 2504 10217 2513 10251
rect 2513 10217 2547 10251
rect 2547 10217 2556 10251
rect 2504 10208 2556 10217
rect 5264 10251 5316 10260
rect 5264 10217 5273 10251
rect 5273 10217 5307 10251
rect 5307 10217 5316 10251
rect 5264 10208 5316 10217
rect 5540 10251 5592 10260
rect 5540 10217 5549 10251
rect 5549 10217 5583 10251
rect 5583 10217 5592 10251
rect 5540 10208 5592 10217
rect 5908 10251 5960 10260
rect 5908 10217 5917 10251
rect 5917 10217 5951 10251
rect 5951 10217 5960 10251
rect 5908 10208 5960 10217
rect 8484 10208 8536 10260
rect 12348 10208 12400 10260
rect 12992 10208 13044 10260
rect 17868 10251 17920 10260
rect 17868 10217 17877 10251
rect 17877 10217 17911 10251
rect 17911 10217 17920 10251
rect 17868 10208 17920 10217
rect 18512 10208 18564 10260
rect 18604 10208 18656 10260
rect 20260 10208 20312 10260
rect 2044 10140 2096 10192
rect 2688 10140 2740 10192
rect 7104 10140 7156 10192
rect 11152 10140 11204 10192
rect 12532 10183 12584 10192
rect 12532 10149 12541 10183
rect 12541 10149 12575 10183
rect 12575 10149 12584 10183
rect 12532 10140 12584 10149
rect 15936 10140 15988 10192
rect 23204 10208 23256 10260
rect 25412 10251 25464 10260
rect 25412 10217 25421 10251
rect 25421 10217 25455 10251
rect 25455 10217 25464 10251
rect 25412 10208 25464 10217
rect 26608 10208 26660 10260
rect 28724 10208 28776 10260
rect 29644 10208 29696 10260
rect 34244 10208 34296 10260
rect 39212 10208 39264 10260
rect 40592 10251 40644 10260
rect 40592 10217 40601 10251
rect 40601 10217 40635 10251
rect 40635 10217 40644 10251
rect 40592 10208 40644 10217
rect 41788 10251 41840 10260
rect 41788 10217 41797 10251
rect 41797 10217 41831 10251
rect 41831 10217 41840 10251
rect 41788 10208 41840 10217
rect 43076 10251 43128 10260
rect 43076 10217 43085 10251
rect 43085 10217 43119 10251
rect 43119 10217 43128 10251
rect 43076 10208 43128 10217
rect 46940 10251 46992 10260
rect 46940 10217 46949 10251
rect 46949 10217 46983 10251
rect 46983 10217 46992 10251
rect 46940 10208 46992 10217
rect 21272 10183 21324 10192
rect 21272 10149 21281 10183
rect 21281 10149 21315 10183
rect 21315 10149 21324 10183
rect 21272 10140 21324 10149
rect 21456 10183 21508 10192
rect 21456 10149 21465 10183
rect 21465 10149 21499 10183
rect 21499 10149 21508 10183
rect 21456 10140 21508 10149
rect 21732 10140 21784 10192
rect 22192 10183 22244 10192
rect 22192 10149 22201 10183
rect 22201 10149 22235 10183
rect 22235 10149 22244 10183
rect 22192 10140 22244 10149
rect 26056 10183 26108 10192
rect 26056 10149 26065 10183
rect 26065 10149 26099 10183
rect 26099 10149 26108 10183
rect 26056 10140 26108 10149
rect 27528 10140 27580 10192
rect 28816 10183 28868 10192
rect 28816 10149 28825 10183
rect 28825 10149 28859 10183
rect 28859 10149 28868 10183
rect 28816 10140 28868 10149
rect 37740 10140 37792 10192
rect 39580 10140 39632 10192
rect 42064 10140 42116 10192
rect 43444 10140 43496 10192
rect 43904 10183 43956 10192
rect 43904 10149 43913 10183
rect 43913 10149 43947 10183
rect 43947 10149 43956 10183
rect 43904 10140 43956 10149
rect 4620 10072 4672 10124
rect 5356 10115 5408 10124
rect 5356 10081 5365 10115
rect 5365 10081 5399 10115
rect 5399 10081 5408 10115
rect 5356 10072 5408 10081
rect 9772 10072 9824 10124
rect 10416 10072 10468 10124
rect 15660 10115 15712 10124
rect 15660 10081 15669 10115
rect 15669 10081 15703 10115
rect 15703 10081 15712 10115
rect 15660 10072 15712 10081
rect 34520 10072 34572 10124
rect 35808 10072 35860 10124
rect 38108 10115 38160 10124
rect 38108 10081 38117 10115
rect 38117 10081 38151 10115
rect 38151 10081 38160 10115
rect 38108 10072 38160 10081
rect 39304 10115 39356 10124
rect 39304 10081 39313 10115
rect 39313 10081 39347 10115
rect 39347 10081 39356 10115
rect 39304 10072 39356 10081
rect 40776 10072 40828 10124
rect 41144 10072 41196 10124
rect 42432 10072 42484 10124
rect 45836 10115 45888 10124
rect 2504 10047 2556 10056
rect 2504 10013 2513 10047
rect 2513 10013 2547 10047
rect 2547 10013 2556 10047
rect 2504 10004 2556 10013
rect 7012 10047 7064 10056
rect 7012 10013 7021 10047
rect 7021 10013 7055 10047
rect 7055 10013 7064 10047
rect 7012 10004 7064 10013
rect 7288 10004 7340 10056
rect 7840 10004 7892 10056
rect 9680 10047 9732 10056
rect 9680 10013 9689 10047
rect 9689 10013 9723 10047
rect 9723 10013 9732 10047
rect 9680 10004 9732 10013
rect 12808 10047 12860 10056
rect 12808 10013 12817 10047
rect 12817 10013 12851 10047
rect 12851 10013 12860 10047
rect 12808 10004 12860 10013
rect 15200 10004 15252 10056
rect 23020 10047 23072 10056
rect 23020 10013 23029 10047
rect 23029 10013 23063 10047
rect 23063 10013 23072 10047
rect 23020 10004 23072 10013
rect 23112 10047 23164 10056
rect 23112 10013 23121 10047
rect 23121 10013 23155 10047
rect 23155 10013 23164 10047
rect 25320 10047 25372 10056
rect 23112 10004 23164 10013
rect 25320 10013 25329 10047
rect 25329 10013 25363 10047
rect 25363 10013 25372 10047
rect 25320 10004 25372 10013
rect 25504 10047 25556 10056
rect 25504 10013 25513 10047
rect 25513 10013 25547 10047
rect 25547 10013 25556 10047
rect 25504 10004 25556 10013
rect 29000 10004 29052 10056
rect 35348 10047 35400 10056
rect 35348 10013 35357 10047
rect 35357 10013 35391 10047
rect 35391 10013 35400 10047
rect 35348 10004 35400 10013
rect 38568 10004 38620 10056
rect 6552 9979 6604 9988
rect 6552 9945 6561 9979
rect 6561 9945 6595 9979
rect 6595 9945 6604 9979
rect 6552 9936 6604 9945
rect 10692 9936 10744 9988
rect 37832 9979 37884 9988
rect 37832 9945 37841 9979
rect 37841 9945 37875 9979
rect 37875 9945 37884 9979
rect 37832 9936 37884 9945
rect 45836 10081 45870 10115
rect 45870 10081 45888 10115
rect 45836 10072 45888 10081
rect 43628 10004 43680 10056
rect 45560 10047 45612 10056
rect 45560 10013 45569 10047
rect 45569 10013 45603 10047
rect 45603 10013 45612 10047
rect 45560 10004 45612 10013
rect 2688 9868 2740 9920
rect 4712 9911 4764 9920
rect 4712 9877 4721 9911
rect 4721 9877 4755 9911
rect 4755 9877 4764 9911
rect 4712 9868 4764 9877
rect 5448 9868 5500 9920
rect 7196 9868 7248 9920
rect 11060 9911 11112 9920
rect 11060 9877 11069 9911
rect 11069 9877 11103 9911
rect 11103 9877 11112 9911
rect 11060 9868 11112 9877
rect 15384 9911 15436 9920
rect 15384 9877 15393 9911
rect 15393 9877 15427 9911
rect 15427 9877 15436 9911
rect 15384 9868 15436 9877
rect 23572 9868 23624 9920
rect 24952 9911 25004 9920
rect 24952 9877 24961 9911
rect 24961 9877 24995 9911
rect 24995 9877 25004 9911
rect 24952 9868 25004 9877
rect 28540 9911 28592 9920
rect 28540 9877 28549 9911
rect 28549 9877 28583 9911
rect 28583 9877 28592 9911
rect 28540 9868 28592 9877
rect 29552 9911 29604 9920
rect 29552 9877 29561 9911
rect 29561 9877 29595 9911
rect 29595 9877 29604 9911
rect 29552 9868 29604 9877
rect 30012 9868 30064 9920
rect 35440 9868 35492 9920
rect 41972 9868 42024 9920
rect 44272 9868 44324 9920
rect 45100 9868 45152 9920
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 34966 9766 35018 9818
rect 35030 9766 35082 9818
rect 35094 9766 35146 9818
rect 35158 9766 35210 9818
rect 2504 9664 2556 9716
rect 5356 9707 5408 9716
rect 5356 9673 5365 9707
rect 5365 9673 5399 9707
rect 5399 9673 5408 9707
rect 5356 9664 5408 9673
rect 5908 9664 5960 9716
rect 7012 9707 7064 9716
rect 7012 9673 7021 9707
rect 7021 9673 7055 9707
rect 7055 9673 7064 9707
rect 7012 9664 7064 9673
rect 8484 9664 8536 9716
rect 12532 9664 12584 9716
rect 12808 9664 12860 9716
rect 15660 9664 15712 9716
rect 2780 9639 2832 9648
rect 2780 9605 2789 9639
rect 2789 9605 2823 9639
rect 2823 9605 2832 9639
rect 2780 9596 2832 9605
rect 4620 9596 4672 9648
rect 2688 9528 2740 9580
rect 21456 9664 21508 9716
rect 21732 9707 21784 9716
rect 21732 9673 21741 9707
rect 21741 9673 21775 9707
rect 21775 9673 21784 9707
rect 21732 9664 21784 9673
rect 23020 9664 23072 9716
rect 23204 9707 23256 9716
rect 23204 9673 23213 9707
rect 23213 9673 23247 9707
rect 23247 9673 23256 9707
rect 23204 9664 23256 9673
rect 16672 9596 16724 9648
rect 21272 9639 21324 9648
rect 21272 9605 21281 9639
rect 21281 9605 21315 9639
rect 21315 9605 21324 9639
rect 21272 9596 21324 9605
rect 21916 9596 21968 9648
rect 23112 9596 23164 9648
rect 24584 9596 24636 9648
rect 25412 9664 25464 9716
rect 27804 9664 27856 9716
rect 28540 9664 28592 9716
rect 28724 9707 28776 9716
rect 28724 9673 28733 9707
rect 28733 9673 28767 9707
rect 28767 9673 28776 9707
rect 28724 9664 28776 9673
rect 28816 9664 28868 9716
rect 27160 9639 27212 9648
rect 27160 9605 27169 9639
rect 27169 9605 27203 9639
rect 27203 9605 27212 9639
rect 27160 9596 27212 9605
rect 29276 9664 29328 9716
rect 1492 9460 1544 9512
rect 2412 9460 2464 9512
rect 4160 9392 4212 9444
rect 4988 9460 5040 9512
rect 12348 9528 12400 9580
rect 34244 9664 34296 9716
rect 34796 9664 34848 9716
rect 37740 9707 37792 9716
rect 34520 9596 34572 9648
rect 30104 9571 30156 9580
rect 30104 9537 30113 9571
rect 30113 9537 30147 9571
rect 30147 9537 30156 9571
rect 30104 9528 30156 9537
rect 37740 9673 37749 9707
rect 37749 9673 37783 9707
rect 37783 9673 37792 9707
rect 37740 9664 37792 9673
rect 40776 9707 40828 9716
rect 40776 9673 40785 9707
rect 40785 9673 40819 9707
rect 40819 9673 40828 9707
rect 40776 9664 40828 9673
rect 41420 9664 41472 9716
rect 41696 9664 41748 9716
rect 43444 9664 43496 9716
rect 42800 9596 42852 9648
rect 43904 9596 43956 9648
rect 46940 9639 46992 9648
rect 46940 9605 46949 9639
rect 46949 9605 46983 9639
rect 46983 9605 46992 9639
rect 46940 9596 46992 9605
rect 47400 9639 47452 9648
rect 47400 9605 47409 9639
rect 47409 9605 47443 9639
rect 47443 9605 47452 9639
rect 47400 9596 47452 9605
rect 35532 9571 35584 9580
rect 35532 9537 35541 9571
rect 35541 9537 35575 9571
rect 35575 9537 35584 9571
rect 35532 9528 35584 9537
rect 41696 9528 41748 9580
rect 42064 9528 42116 9580
rect 7840 9503 7892 9512
rect 7840 9469 7863 9503
rect 7863 9469 7892 9503
rect 3976 9324 4028 9376
rect 4712 9392 4764 9444
rect 6460 9392 6512 9444
rect 7840 9460 7892 9469
rect 15292 9460 15344 9512
rect 15568 9460 15620 9512
rect 9956 9392 10008 9444
rect 6552 9367 6604 9376
rect 6552 9333 6561 9367
rect 6561 9333 6595 9367
rect 6595 9333 6604 9367
rect 6552 9324 6604 9333
rect 7104 9324 7156 9376
rect 9680 9367 9732 9376
rect 9680 9333 9689 9367
rect 9689 9333 9723 9367
rect 9723 9333 9732 9367
rect 9680 9324 9732 9333
rect 10140 9392 10192 9444
rect 10968 9392 11020 9444
rect 14648 9392 14700 9444
rect 25320 9392 25372 9444
rect 26056 9392 26108 9444
rect 40776 9460 40828 9512
rect 43168 9460 43220 9512
rect 44272 9460 44324 9512
rect 45836 9460 45888 9512
rect 46480 9460 46532 9512
rect 30380 9435 30432 9444
rect 30380 9401 30414 9435
rect 30414 9401 30432 9435
rect 30380 9392 30432 9401
rect 36360 9392 36412 9444
rect 42616 9435 42668 9444
rect 42616 9401 42625 9435
rect 42625 9401 42659 9435
rect 42659 9401 42668 9435
rect 42616 9392 42668 9401
rect 44824 9435 44876 9444
rect 44824 9401 44833 9435
rect 44833 9401 44867 9435
rect 44867 9401 44876 9435
rect 44824 9392 44876 9401
rect 45100 9435 45152 9444
rect 45100 9401 45109 9435
rect 45109 9401 45143 9435
rect 45143 9401 45152 9435
rect 45100 9392 45152 9401
rect 15936 9367 15988 9376
rect 15936 9333 15945 9367
rect 15945 9333 15979 9367
rect 15979 9333 15988 9367
rect 15936 9324 15988 9333
rect 24676 9324 24728 9376
rect 26608 9367 26660 9376
rect 26608 9333 26617 9367
rect 26617 9333 26651 9367
rect 26651 9333 26660 9367
rect 26608 9324 26660 9333
rect 27896 9367 27948 9376
rect 27896 9333 27905 9367
rect 27905 9333 27939 9367
rect 27939 9333 27948 9367
rect 27896 9324 27948 9333
rect 28264 9367 28316 9376
rect 28264 9333 28273 9367
rect 28273 9333 28307 9367
rect 28307 9333 28316 9367
rect 28264 9324 28316 9333
rect 30012 9324 30064 9376
rect 36452 9324 36504 9376
rect 38108 9367 38160 9376
rect 38108 9333 38117 9367
rect 38117 9333 38151 9367
rect 38151 9333 38160 9367
rect 38108 9324 38160 9333
rect 38568 9367 38620 9376
rect 38568 9333 38577 9367
rect 38577 9333 38611 9367
rect 38611 9333 38620 9367
rect 38568 9324 38620 9333
rect 38660 9324 38712 9376
rect 39304 9367 39356 9376
rect 39304 9333 39313 9367
rect 39313 9333 39347 9367
rect 39347 9333 39356 9367
rect 39304 9324 39356 9333
rect 42524 9324 42576 9376
rect 45008 9367 45060 9376
rect 45008 9333 45017 9367
rect 45017 9333 45051 9367
rect 45051 9333 45060 9367
rect 45008 9324 45060 9333
rect 45192 9324 45244 9376
rect 45560 9367 45612 9376
rect 45560 9333 45569 9367
rect 45569 9333 45603 9367
rect 45603 9333 45612 9367
rect 45560 9324 45612 9333
rect 19606 9222 19658 9274
rect 19670 9222 19722 9274
rect 19734 9222 19786 9274
rect 19798 9222 19850 9274
rect 1492 9120 1544 9172
rect 2412 9163 2464 9172
rect 2412 9129 2421 9163
rect 2421 9129 2455 9163
rect 2455 9129 2464 9163
rect 2412 9120 2464 9129
rect 2780 9163 2832 9172
rect 2780 9129 2789 9163
rect 2789 9129 2823 9163
rect 2823 9129 2832 9163
rect 7840 9163 7892 9172
rect 2780 9120 2832 9129
rect 7840 9129 7849 9163
rect 7849 9129 7883 9163
rect 7883 9129 7892 9163
rect 7840 9120 7892 9129
rect 8484 9163 8536 9172
rect 8484 9129 8493 9163
rect 8493 9129 8527 9163
rect 8527 9129 8536 9163
rect 8484 9120 8536 9129
rect 10416 9163 10468 9172
rect 10416 9129 10425 9163
rect 10425 9129 10459 9163
rect 10459 9129 10468 9163
rect 10416 9120 10468 9129
rect 16672 9163 16724 9172
rect 16672 9129 16681 9163
rect 16681 9129 16715 9163
rect 16715 9129 16724 9163
rect 16672 9120 16724 9129
rect 26056 9163 26108 9172
rect 26056 9129 26065 9163
rect 26065 9129 26099 9163
rect 26099 9129 26108 9163
rect 26056 9120 26108 9129
rect 26608 9120 26660 9172
rect 29552 9120 29604 9172
rect 30380 9120 30432 9172
rect 35348 9120 35400 9172
rect 35992 9120 36044 9172
rect 36360 9120 36412 9172
rect 40040 9163 40092 9172
rect 4620 9095 4672 9104
rect 4620 9061 4629 9095
rect 4629 9061 4663 9095
rect 4663 9061 4672 9095
rect 4620 9052 4672 9061
rect 2044 8984 2096 9036
rect 5172 8984 5224 9036
rect 7288 9052 7340 9104
rect 10140 9095 10192 9104
rect 10140 9061 10149 9095
rect 10149 9061 10183 9095
rect 10183 9061 10192 9095
rect 10140 9052 10192 9061
rect 12256 9095 12308 9104
rect 12256 9061 12290 9095
rect 12290 9061 12308 9095
rect 12256 9052 12308 9061
rect 24584 9095 24636 9104
rect 24584 9061 24593 9095
rect 24593 9061 24627 9095
rect 24627 9061 24636 9095
rect 24584 9052 24636 9061
rect 27160 9095 27212 9104
rect 27160 9061 27169 9095
rect 27169 9061 27203 9095
rect 27203 9061 27212 9095
rect 27160 9052 27212 9061
rect 27804 9052 27856 9104
rect 28080 9095 28132 9104
rect 28080 9061 28089 9095
rect 28089 9061 28123 9095
rect 28123 9061 28132 9095
rect 28080 9052 28132 9061
rect 29092 9052 29144 9104
rect 30012 9052 30064 9104
rect 35808 9052 35860 9104
rect 38936 9095 38988 9104
rect 6552 8984 6604 9036
rect 15016 8984 15068 9036
rect 15936 8984 15988 9036
rect 18052 9027 18104 9036
rect 18052 8993 18086 9027
rect 18086 8993 18104 9027
rect 18052 8984 18104 8993
rect 22284 9027 22336 9036
rect 22284 8993 22293 9027
rect 22293 8993 22327 9027
rect 22327 8993 22336 9027
rect 22284 8984 22336 8993
rect 22928 8984 22980 9036
rect 29000 8984 29052 9036
rect 30196 8984 30248 9036
rect 30840 8984 30892 9036
rect 31852 8984 31904 9036
rect 6460 8959 6512 8968
rect 4160 8891 4212 8900
rect 4160 8857 4169 8891
rect 4169 8857 4203 8891
rect 4203 8857 4212 8891
rect 4160 8848 4212 8857
rect 6460 8925 6469 8959
rect 6469 8925 6503 8959
rect 6503 8925 6512 8959
rect 6460 8916 6512 8925
rect 11980 8959 12032 8968
rect 11980 8925 11989 8959
rect 11989 8925 12023 8959
rect 12023 8925 12032 8959
rect 11980 8916 12032 8925
rect 15292 8959 15344 8968
rect 15292 8925 15301 8959
rect 15301 8925 15335 8959
rect 15335 8925 15344 8959
rect 15292 8916 15344 8925
rect 17776 8959 17828 8968
rect 17776 8925 17785 8959
rect 17785 8925 17819 8959
rect 17819 8925 17828 8959
rect 17776 8916 17828 8925
rect 20904 8959 20956 8968
rect 20904 8925 20913 8959
rect 20913 8925 20947 8959
rect 20947 8925 20956 8959
rect 20904 8916 20956 8925
rect 24676 8959 24728 8968
rect 24676 8925 24685 8959
rect 24685 8925 24719 8959
rect 24719 8925 24728 8959
rect 24676 8916 24728 8925
rect 27068 8959 27120 8968
rect 27068 8925 27077 8959
rect 27077 8925 27111 8959
rect 27111 8925 27120 8959
rect 27068 8916 27120 8925
rect 28172 8959 28224 8968
rect 28172 8925 28181 8959
rect 28181 8925 28215 8959
rect 28215 8925 28224 8959
rect 28172 8916 28224 8925
rect 30104 8916 30156 8968
rect 31576 8916 31628 8968
rect 36452 8959 36504 8968
rect 36452 8925 36461 8959
rect 36461 8925 36495 8959
rect 36495 8925 36504 8959
rect 36452 8916 36504 8925
rect 38936 9061 38945 9095
rect 38945 9061 38979 9095
rect 38979 9061 38988 9095
rect 38936 9052 38988 9061
rect 39120 9095 39172 9104
rect 39120 9061 39129 9095
rect 39129 9061 39163 9095
rect 39163 9061 39172 9095
rect 39120 9052 39172 9061
rect 40040 9129 40049 9163
rect 40049 9129 40083 9163
rect 40083 9129 40092 9163
rect 41972 9163 42024 9172
rect 40040 9120 40092 9129
rect 41972 9129 41981 9163
rect 41981 9129 42015 9163
rect 42015 9129 42024 9163
rect 41972 9120 42024 9129
rect 42432 9163 42484 9172
rect 42432 9129 42441 9163
rect 42441 9129 42475 9163
rect 42475 9129 42484 9163
rect 42432 9120 42484 9129
rect 44824 9120 44876 9172
rect 46480 9163 46532 9172
rect 46480 9129 46489 9163
rect 46489 9129 46523 9163
rect 46523 9129 46532 9163
rect 46480 9120 46532 9129
rect 40684 9095 40736 9104
rect 40684 9061 40693 9095
rect 40693 9061 40727 9095
rect 40727 9061 40736 9095
rect 40684 9052 40736 9061
rect 40776 9095 40828 9104
rect 40776 9061 40785 9095
rect 40785 9061 40819 9095
rect 40819 9061 40828 9095
rect 40776 9052 40828 9061
rect 45008 9052 45060 9104
rect 45560 9052 45612 9104
rect 38568 8984 38620 9036
rect 40500 9027 40552 9036
rect 40500 8993 40509 9027
rect 40509 8993 40543 9027
rect 40543 8993 40552 9027
rect 40500 8984 40552 8993
rect 42432 8984 42484 9036
rect 36728 8916 36780 8968
rect 39212 8959 39264 8968
rect 39212 8925 39221 8959
rect 39221 8925 39255 8959
rect 39255 8925 39264 8959
rect 39212 8916 39264 8925
rect 44180 8916 44232 8968
rect 44824 8916 44876 8968
rect 45192 8984 45244 9036
rect 4804 8848 4856 8900
rect 13820 8848 13872 8900
rect 15108 8848 15160 8900
rect 27896 8848 27948 8900
rect 38108 8848 38160 8900
rect 38660 8891 38712 8900
rect 38660 8857 38669 8891
rect 38669 8857 38703 8891
rect 38703 8857 38712 8891
rect 38660 8848 38712 8857
rect 12624 8780 12676 8832
rect 14648 8823 14700 8832
rect 14648 8789 14657 8823
rect 14657 8789 14691 8823
rect 14691 8789 14700 8823
rect 14648 8780 14700 8789
rect 17592 8823 17644 8832
rect 17592 8789 17601 8823
rect 17601 8789 17635 8823
rect 17635 8789 17644 8823
rect 17592 8780 17644 8789
rect 17684 8780 17736 8832
rect 20812 8780 20864 8832
rect 26240 8780 26292 8832
rect 29184 8823 29236 8832
rect 29184 8789 29193 8823
rect 29193 8789 29227 8823
rect 29227 8789 29236 8823
rect 29184 8780 29236 8789
rect 30748 8780 30800 8832
rect 32496 8780 32548 8832
rect 43628 8823 43680 8832
rect 43628 8789 43637 8823
rect 43637 8789 43671 8823
rect 43671 8789 43680 8823
rect 43628 8780 43680 8789
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 34966 8678 35018 8730
rect 35030 8678 35082 8730
rect 35094 8678 35146 8730
rect 35158 8678 35210 8730
rect 2044 8619 2096 8628
rect 2044 8585 2053 8619
rect 2053 8585 2087 8619
rect 2087 8585 2096 8619
rect 2044 8576 2096 8585
rect 4620 8576 4672 8628
rect 4804 8619 4856 8628
rect 4804 8585 4813 8619
rect 4813 8585 4847 8619
rect 4847 8585 4856 8619
rect 4804 8576 4856 8585
rect 1492 8508 1544 8560
rect 5172 8551 5224 8560
rect 5172 8517 5181 8551
rect 5181 8517 5215 8551
rect 5215 8517 5224 8551
rect 5172 8508 5224 8517
rect 6552 8576 6604 8628
rect 15016 8619 15068 8628
rect 15016 8585 15025 8619
rect 15025 8585 15059 8619
rect 15059 8585 15068 8619
rect 15016 8576 15068 8585
rect 15292 8619 15344 8628
rect 15292 8585 15301 8619
rect 15301 8585 15335 8619
rect 15335 8585 15344 8619
rect 15292 8576 15344 8585
rect 17776 8619 17828 8628
rect 17776 8585 17785 8619
rect 17785 8585 17819 8619
rect 17819 8585 17828 8619
rect 17776 8576 17828 8585
rect 22284 8576 22336 8628
rect 22928 8619 22980 8628
rect 16396 8551 16448 8560
rect 16396 8517 16405 8551
rect 16405 8517 16439 8551
rect 16439 8517 16448 8551
rect 16396 8508 16448 8517
rect 2780 8415 2832 8424
rect 2780 8381 2814 8415
rect 2814 8381 2832 8415
rect 2780 8372 2832 8381
rect 14648 8440 14700 8492
rect 17684 8440 17736 8492
rect 22928 8585 22937 8619
rect 22937 8585 22971 8619
rect 22971 8585 22980 8619
rect 22928 8576 22980 8585
rect 27068 8576 27120 8628
rect 28080 8576 28132 8628
rect 29184 8576 29236 8628
rect 29552 8619 29604 8628
rect 29552 8585 29561 8619
rect 29561 8585 29595 8619
rect 29595 8585 29604 8619
rect 29552 8576 29604 8585
rect 31576 8619 31628 8628
rect 31576 8585 31585 8619
rect 31585 8585 31619 8619
rect 31619 8585 31628 8619
rect 31576 8576 31628 8585
rect 31944 8576 31996 8628
rect 35992 8619 36044 8628
rect 35992 8585 36001 8619
rect 36001 8585 36035 8619
rect 36035 8585 36044 8619
rect 35992 8576 36044 8585
rect 38936 8619 38988 8628
rect 38936 8585 38945 8619
rect 38945 8585 38979 8619
rect 38979 8585 38988 8619
rect 38936 8576 38988 8585
rect 40500 8576 40552 8628
rect 42432 8619 42484 8628
rect 42432 8585 42441 8619
rect 42441 8585 42475 8619
rect 42475 8585 42484 8619
rect 42432 8576 42484 8585
rect 29092 8551 29144 8560
rect 6460 8304 6512 8356
rect 11980 8372 12032 8424
rect 20812 8415 20864 8424
rect 20812 8381 20846 8415
rect 20846 8381 20864 8415
rect 20812 8372 20864 8381
rect 29092 8517 29101 8551
rect 29101 8517 29135 8551
rect 29135 8517 29144 8551
rect 29092 8508 29144 8517
rect 29368 8508 29420 8560
rect 6920 8304 6972 8356
rect 12532 8304 12584 8356
rect 16948 8347 17000 8356
rect 4068 8236 4120 8288
rect 9680 8236 9732 8288
rect 11980 8236 12032 8288
rect 12900 8236 12952 8288
rect 16948 8313 16957 8347
rect 16957 8313 16991 8347
rect 16991 8313 17000 8347
rect 16948 8304 17000 8313
rect 17592 8304 17644 8356
rect 18512 8304 18564 8356
rect 16856 8279 16908 8288
rect 16856 8245 16865 8279
rect 16865 8245 16899 8279
rect 16899 8245 16908 8279
rect 16856 8236 16908 8245
rect 18604 8236 18656 8288
rect 24676 8372 24728 8424
rect 23940 8347 23992 8356
rect 23940 8313 23974 8347
rect 23974 8313 23992 8347
rect 23940 8304 23992 8313
rect 23848 8236 23900 8288
rect 30748 8440 30800 8492
rect 30840 8483 30892 8492
rect 30840 8449 30849 8483
rect 30849 8449 30883 8483
rect 30883 8449 30892 8483
rect 42800 8551 42852 8560
rect 42800 8517 42809 8551
rect 42809 8517 42843 8551
rect 42843 8517 42852 8551
rect 42800 8508 42852 8517
rect 46940 8551 46992 8560
rect 46940 8517 46949 8551
rect 46949 8517 46983 8551
rect 46983 8517 46992 8551
rect 46940 8508 46992 8517
rect 30840 8440 30892 8449
rect 26516 8304 26568 8356
rect 30748 8347 30800 8356
rect 30748 8313 30757 8347
rect 30757 8313 30791 8347
rect 30791 8313 30800 8347
rect 30748 8304 30800 8313
rect 35532 8372 35584 8424
rect 36544 8372 36596 8424
rect 40316 8372 40368 8424
rect 43628 8483 43680 8492
rect 43628 8449 43637 8483
rect 43637 8449 43671 8483
rect 43671 8449 43680 8483
rect 43628 8440 43680 8449
rect 47400 8483 47452 8492
rect 47400 8449 47409 8483
rect 47409 8449 47443 8483
rect 47443 8449 47452 8483
rect 47400 8440 47452 8449
rect 31852 8304 31904 8356
rect 32496 8304 32548 8356
rect 26608 8236 26660 8288
rect 30288 8236 30340 8288
rect 37832 8279 37884 8288
rect 37832 8245 37841 8279
rect 37841 8245 37875 8279
rect 37875 8245 37884 8279
rect 37832 8236 37884 8245
rect 37924 8236 37976 8288
rect 39120 8304 39172 8356
rect 40316 8279 40368 8288
rect 40316 8245 40325 8279
rect 40325 8245 40359 8279
rect 40359 8245 40368 8279
rect 40316 8236 40368 8245
rect 40684 8236 40736 8288
rect 41604 8304 41656 8356
rect 43076 8304 43128 8356
rect 44824 8236 44876 8288
rect 45560 8279 45612 8288
rect 45560 8245 45569 8279
rect 45569 8245 45603 8279
rect 45603 8245 45612 8279
rect 45560 8236 45612 8245
rect 19606 8134 19658 8186
rect 19670 8134 19722 8186
rect 19734 8134 19786 8186
rect 19798 8134 19850 8186
rect 2044 8032 2096 8084
rect 2688 8032 2740 8084
rect 4804 8032 4856 8084
rect 6552 8075 6604 8084
rect 6552 8041 6561 8075
rect 6561 8041 6595 8075
rect 6595 8041 6604 8075
rect 6552 8032 6604 8041
rect 12256 8032 12308 8084
rect 16856 8032 16908 8084
rect 18052 8032 18104 8084
rect 20260 8032 20312 8084
rect 20812 8032 20864 8084
rect 21180 8032 21232 8084
rect 4620 7964 4672 8016
rect 11244 7964 11296 8016
rect 12532 7964 12584 8016
rect 16396 7964 16448 8016
rect 16488 8007 16540 8016
rect 16488 7973 16497 8007
rect 16497 7973 16531 8007
rect 16531 7973 16540 8007
rect 16948 8007 17000 8016
rect 16488 7964 16540 7973
rect 16948 7973 16957 8007
rect 16957 7973 16991 8007
rect 16991 7973 17000 8007
rect 16948 7964 17000 7973
rect 18604 7964 18656 8016
rect 22008 8032 22060 8084
rect 24676 8075 24728 8084
rect 24676 8041 24685 8075
rect 24685 8041 24719 8075
rect 24719 8041 24728 8075
rect 24676 8032 24728 8041
rect 24952 8032 25004 8084
rect 26516 8032 26568 8084
rect 28172 8032 28224 8084
rect 28448 8075 28500 8084
rect 28448 8041 28457 8075
rect 28457 8041 28491 8075
rect 28491 8041 28500 8075
rect 30288 8075 30340 8084
rect 28448 8032 28500 8041
rect 1952 7896 2004 7948
rect 13820 7896 13872 7948
rect 17776 7896 17828 7948
rect 27068 7964 27120 8016
rect 29368 8007 29420 8016
rect 29368 7973 29377 8007
rect 29377 7973 29411 8007
rect 29411 7973 29420 8007
rect 29368 7964 29420 7973
rect 29552 8007 29604 8016
rect 29552 7973 29561 8007
rect 29561 7973 29595 8007
rect 29595 7973 29604 8007
rect 29552 7964 29604 7973
rect 30288 8041 30297 8075
rect 30297 8041 30331 8075
rect 30331 8041 30340 8075
rect 30288 8032 30340 8041
rect 31576 8032 31628 8084
rect 31852 8032 31904 8084
rect 36452 8075 36504 8084
rect 36452 8041 36461 8075
rect 36461 8041 36495 8075
rect 36495 8041 36504 8075
rect 36452 8032 36504 8041
rect 40500 8032 40552 8084
rect 41604 8075 41656 8084
rect 41604 8041 41613 8075
rect 41613 8041 41647 8075
rect 41647 8041 41656 8075
rect 41604 8032 41656 8041
rect 42524 8032 42576 8084
rect 43628 8032 43680 8084
rect 45560 8032 45612 8084
rect 36728 7964 36780 8016
rect 37832 7964 37884 8016
rect 24952 7896 25004 7948
rect 26608 7896 26660 7948
rect 4068 7871 4120 7880
rect 4068 7837 4077 7871
rect 4077 7837 4111 7871
rect 4111 7837 4120 7871
rect 4068 7828 4120 7837
rect 9312 7828 9364 7880
rect 9680 7871 9732 7880
rect 9680 7837 9689 7871
rect 9689 7837 9723 7871
rect 9723 7837 9732 7871
rect 9680 7828 9732 7837
rect 12900 7871 12952 7880
rect 12900 7837 12909 7871
rect 12909 7837 12943 7871
rect 12943 7837 12952 7871
rect 12900 7828 12952 7837
rect 13084 7871 13136 7880
rect 13084 7837 13093 7871
rect 13093 7837 13127 7871
rect 13127 7837 13136 7871
rect 13084 7828 13136 7837
rect 16580 7871 16632 7880
rect 16580 7837 16589 7871
rect 16589 7837 16623 7871
rect 16623 7837 16632 7871
rect 16580 7828 16632 7837
rect 20996 7828 21048 7880
rect 21456 7828 21508 7880
rect 21640 7871 21692 7880
rect 21640 7837 21649 7871
rect 21649 7837 21683 7871
rect 21683 7837 21692 7871
rect 21640 7828 21692 7837
rect 21916 7871 21968 7880
rect 21916 7837 21925 7871
rect 21925 7837 21959 7871
rect 21959 7837 21968 7871
rect 21916 7828 21968 7837
rect 22008 7828 22060 7880
rect 22100 7828 22152 7880
rect 24584 7828 24636 7880
rect 26148 7828 26200 7880
rect 23940 7760 23992 7812
rect 24768 7760 24820 7812
rect 39948 7896 40000 7948
rect 45376 7896 45428 7948
rect 37740 7871 37792 7880
rect 37740 7837 37749 7871
rect 37749 7837 37783 7871
rect 37783 7837 37792 7871
rect 37740 7828 37792 7837
rect 40224 7871 40276 7880
rect 40224 7837 40233 7871
rect 40233 7837 40267 7871
rect 40267 7837 40276 7871
rect 40224 7828 40276 7837
rect 44824 7871 44876 7880
rect 44824 7837 44833 7871
rect 44833 7837 44867 7871
rect 44867 7837 44876 7871
rect 44824 7828 44876 7837
rect 30656 7760 30708 7812
rect 6920 7735 6972 7744
rect 6920 7701 6929 7735
rect 6929 7701 6963 7735
rect 6963 7701 6972 7735
rect 6920 7692 6972 7701
rect 11796 7692 11848 7744
rect 13820 7692 13872 7744
rect 15016 7735 15068 7744
rect 15016 7701 15025 7735
rect 15025 7701 15059 7735
rect 15059 7701 15068 7735
rect 15016 7692 15068 7701
rect 16028 7735 16080 7744
rect 16028 7701 16037 7735
rect 16037 7701 16071 7735
rect 16071 7701 16080 7735
rect 16028 7692 16080 7701
rect 20812 7692 20864 7744
rect 21640 7692 21692 7744
rect 23296 7692 23348 7744
rect 25320 7692 25372 7744
rect 27620 7692 27672 7744
rect 30748 7735 30800 7744
rect 30748 7701 30757 7735
rect 30757 7701 30791 7735
rect 30791 7701 30800 7735
rect 30748 7692 30800 7701
rect 38384 7692 38436 7744
rect 39948 7692 40000 7744
rect 43076 7735 43128 7744
rect 43076 7701 43085 7735
rect 43085 7701 43119 7735
rect 43119 7701 43128 7735
rect 43076 7692 43128 7701
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 34966 7590 35018 7642
rect 35030 7590 35082 7642
rect 35094 7590 35146 7642
rect 35158 7590 35210 7642
rect 4620 7488 4672 7540
rect 11244 7531 11296 7540
rect 11244 7497 11253 7531
rect 11253 7497 11287 7531
rect 11287 7497 11296 7531
rect 11244 7488 11296 7497
rect 11980 7488 12032 7540
rect 5448 7420 5500 7472
rect 12808 7488 12860 7540
rect 16396 7531 16448 7540
rect 16396 7497 16405 7531
rect 16405 7497 16439 7531
rect 16439 7497 16448 7531
rect 16396 7488 16448 7497
rect 17776 7531 17828 7540
rect 17776 7497 17785 7531
rect 17785 7497 17819 7531
rect 17819 7497 17828 7531
rect 17776 7488 17828 7497
rect 20260 7531 20312 7540
rect 20260 7497 20269 7531
rect 20269 7497 20303 7531
rect 20303 7497 20312 7531
rect 20260 7488 20312 7497
rect 20904 7488 20956 7540
rect 21640 7488 21692 7540
rect 24584 7531 24636 7540
rect 24584 7497 24593 7531
rect 24593 7497 24627 7531
rect 24627 7497 24636 7531
rect 24584 7488 24636 7497
rect 24860 7531 24912 7540
rect 24860 7497 24869 7531
rect 24869 7497 24903 7531
rect 24903 7497 24912 7531
rect 24860 7488 24912 7497
rect 27068 7488 27120 7540
rect 29552 7488 29604 7540
rect 15108 7420 15160 7472
rect 16488 7420 16540 7472
rect 20812 7463 20864 7472
rect 20812 7429 20821 7463
rect 20821 7429 20855 7463
rect 20855 7429 20864 7463
rect 20812 7420 20864 7429
rect 18604 7395 18656 7404
rect 18604 7361 18613 7395
rect 18613 7361 18647 7395
rect 18647 7361 18656 7395
rect 18604 7352 18656 7361
rect 21180 7420 21232 7472
rect 21456 7420 21508 7472
rect 21916 7420 21968 7472
rect 27712 7463 27764 7472
rect 27712 7429 27721 7463
rect 27721 7429 27755 7463
rect 27755 7429 27764 7463
rect 27712 7420 27764 7429
rect 22008 7352 22060 7404
rect 28264 7352 28316 7404
rect 29644 7352 29696 7404
rect 30196 7395 30248 7404
rect 30196 7361 30205 7395
rect 30205 7361 30239 7395
rect 30239 7361 30248 7395
rect 30196 7352 30248 7361
rect 31484 7488 31536 7540
rect 32496 7531 32548 7540
rect 32496 7497 32505 7531
rect 32505 7497 32539 7531
rect 32539 7497 32548 7531
rect 32496 7488 32548 7497
rect 37832 7488 37884 7540
rect 37924 7531 37976 7540
rect 37924 7497 37933 7531
rect 37933 7497 37967 7531
rect 37967 7497 37976 7531
rect 39948 7531 40000 7540
rect 37924 7488 37976 7497
rect 39948 7497 39957 7531
rect 39957 7497 39991 7531
rect 39991 7497 40000 7531
rect 39948 7488 40000 7497
rect 42524 7488 42576 7540
rect 36728 7420 36780 7472
rect 38384 7395 38436 7404
rect 38384 7361 38393 7395
rect 38393 7361 38427 7395
rect 38427 7361 38436 7395
rect 38384 7352 38436 7361
rect 39948 7352 40000 7404
rect 9312 7327 9364 7336
rect 5540 7259 5592 7268
rect 5540 7225 5549 7259
rect 5549 7225 5583 7259
rect 5583 7225 5592 7259
rect 5540 7216 5592 7225
rect 5632 7216 5684 7268
rect 1952 7148 2004 7200
rect 4160 7191 4212 7200
rect 4160 7157 4169 7191
rect 4169 7157 4203 7191
rect 4203 7157 4212 7191
rect 4160 7148 4212 7157
rect 5724 7191 5776 7200
rect 5724 7157 5733 7191
rect 5733 7157 5767 7191
rect 5767 7157 5776 7191
rect 5724 7148 5776 7157
rect 6920 7148 6972 7200
rect 9312 7293 9321 7327
rect 9321 7293 9355 7327
rect 9355 7293 9364 7327
rect 9312 7284 9364 7293
rect 11980 7284 12032 7336
rect 12348 7284 12400 7336
rect 16948 7284 17000 7336
rect 21180 7284 21232 7336
rect 9588 7259 9640 7268
rect 9588 7225 9622 7259
rect 9622 7225 9640 7259
rect 9588 7216 9640 7225
rect 12900 7216 12952 7268
rect 15292 7259 15344 7268
rect 15292 7225 15301 7259
rect 15301 7225 15335 7259
rect 15335 7225 15344 7259
rect 15292 7216 15344 7225
rect 15384 7216 15436 7268
rect 10232 7148 10284 7200
rect 12348 7148 12400 7200
rect 12440 7148 12492 7200
rect 13912 7148 13964 7200
rect 15016 7148 15068 7200
rect 18512 7216 18564 7268
rect 22100 7284 22152 7336
rect 22560 7284 22612 7336
rect 25320 7327 25372 7336
rect 25320 7293 25329 7327
rect 25329 7293 25363 7327
rect 25363 7293 25372 7327
rect 25320 7284 25372 7293
rect 29736 7284 29788 7336
rect 33600 7327 33652 7336
rect 28264 7259 28316 7268
rect 28264 7225 28273 7259
rect 28273 7225 28307 7259
rect 28307 7225 28316 7259
rect 28264 7216 28316 7225
rect 33600 7293 33609 7327
rect 33609 7293 33643 7327
rect 33643 7293 33652 7327
rect 33600 7284 33652 7293
rect 40316 7327 40368 7336
rect 40316 7293 40325 7327
rect 40325 7293 40359 7327
rect 40359 7293 40368 7327
rect 40316 7284 40368 7293
rect 40684 7284 40736 7336
rect 31208 7216 31260 7268
rect 40500 7216 40552 7268
rect 41144 7216 41196 7268
rect 43444 7259 43496 7268
rect 43444 7225 43453 7259
rect 43453 7225 43487 7259
rect 43487 7225 43496 7259
rect 43628 7284 43680 7336
rect 43444 7216 43496 7225
rect 44824 7216 44876 7268
rect 16580 7148 16632 7200
rect 23480 7148 23532 7200
rect 25504 7191 25556 7200
rect 25504 7157 25513 7191
rect 25513 7157 25547 7191
rect 25547 7157 25556 7191
rect 25504 7148 25556 7157
rect 26608 7191 26660 7200
rect 26608 7157 26617 7191
rect 26617 7157 26651 7191
rect 26651 7157 26660 7191
rect 26608 7148 26660 7157
rect 28172 7191 28224 7200
rect 28172 7157 28181 7191
rect 28181 7157 28215 7191
rect 28215 7157 28224 7191
rect 28172 7148 28224 7157
rect 30472 7148 30524 7200
rect 33784 7191 33836 7200
rect 33784 7157 33793 7191
rect 33793 7157 33827 7191
rect 33827 7157 33836 7191
rect 33784 7148 33836 7157
rect 37280 7148 37332 7200
rect 37740 7148 37792 7200
rect 37832 7148 37884 7200
rect 44180 7148 44232 7200
rect 45836 7148 45888 7200
rect 46940 7191 46992 7200
rect 46940 7157 46949 7191
rect 46949 7157 46983 7191
rect 46983 7157 46992 7191
rect 46940 7148 46992 7157
rect 47400 7191 47452 7200
rect 47400 7157 47409 7191
rect 47409 7157 47443 7191
rect 47443 7157 47452 7191
rect 47400 7148 47452 7157
rect 19606 7046 19658 7098
rect 19670 7046 19722 7098
rect 19734 7046 19786 7098
rect 19798 7046 19850 7098
rect 9588 6944 9640 6996
rect 10232 6987 10284 6996
rect 10232 6953 10241 6987
rect 10241 6953 10275 6987
rect 10275 6953 10284 6987
rect 10232 6944 10284 6953
rect 11244 6944 11296 6996
rect 11612 6944 11664 6996
rect 12532 6987 12584 6996
rect 12532 6953 12541 6987
rect 12541 6953 12575 6987
rect 12575 6953 12584 6987
rect 12532 6944 12584 6953
rect 12900 6987 12952 6996
rect 12900 6953 12909 6987
rect 12909 6953 12943 6987
rect 12943 6953 12952 6987
rect 12900 6944 12952 6953
rect 15292 6944 15344 6996
rect 18604 6944 18656 6996
rect 29736 6987 29788 6996
rect 29736 6953 29745 6987
rect 29745 6953 29779 6987
rect 29779 6953 29788 6987
rect 29736 6944 29788 6953
rect 30656 6987 30708 6996
rect 30656 6953 30665 6987
rect 30665 6953 30699 6987
rect 30699 6953 30708 6987
rect 30656 6944 30708 6953
rect 38384 6987 38436 6996
rect 38384 6953 38393 6987
rect 38393 6953 38427 6987
rect 38427 6953 38436 6987
rect 38384 6944 38436 6953
rect 41144 6987 41196 6996
rect 41144 6953 41153 6987
rect 41153 6953 41187 6987
rect 41187 6953 41196 6987
rect 41144 6944 41196 6953
rect 3332 6876 3384 6928
rect 4160 6876 4212 6928
rect 3240 6808 3292 6860
rect 5540 6876 5592 6928
rect 6828 6876 6880 6928
rect 6184 6851 6236 6860
rect 6184 6817 6218 6851
rect 6218 6817 6236 6851
rect 10048 6851 10100 6860
rect 6184 6808 6236 6817
rect 10048 6817 10057 6851
rect 10057 6817 10091 6851
rect 10091 6817 10100 6851
rect 10048 6808 10100 6817
rect 3976 6672 4028 6724
rect 4160 6672 4212 6724
rect 5540 6740 5592 6792
rect 5908 6783 5960 6792
rect 5908 6749 5917 6783
rect 5917 6749 5951 6783
rect 5951 6749 5960 6783
rect 5908 6740 5960 6749
rect 9496 6740 9548 6792
rect 11980 6808 12032 6860
rect 13820 6808 13872 6860
rect 15200 6808 15252 6860
rect 15476 6808 15528 6860
rect 16028 6808 16080 6860
rect 16396 6851 16448 6860
rect 16396 6817 16405 6851
rect 16405 6817 16439 6851
rect 16439 6817 16448 6851
rect 16396 6808 16448 6817
rect 18512 6808 18564 6860
rect 21364 6808 21416 6860
rect 21916 6808 21968 6860
rect 24952 6851 25004 6860
rect 24952 6817 24961 6851
rect 24961 6817 24995 6851
rect 24995 6817 25004 6851
rect 24952 6808 25004 6817
rect 26884 6808 26936 6860
rect 11796 6783 11848 6792
rect 11796 6749 11805 6783
rect 11805 6749 11839 6783
rect 11839 6749 11848 6783
rect 11796 6740 11848 6749
rect 20536 6740 20588 6792
rect 22928 6740 22980 6792
rect 23940 6783 23992 6792
rect 23940 6749 23949 6783
rect 23949 6749 23983 6783
rect 23983 6749 23992 6783
rect 23940 6740 23992 6749
rect 21180 6715 21232 6724
rect 21180 6681 21189 6715
rect 21189 6681 21223 6715
rect 21223 6681 21232 6715
rect 21180 6672 21232 6681
rect 28264 6876 28316 6928
rect 28448 6876 28500 6928
rect 29184 6876 29236 6928
rect 33784 6876 33836 6928
rect 34336 6919 34388 6928
rect 34336 6885 34345 6919
rect 34345 6885 34379 6919
rect 34379 6885 34388 6919
rect 34336 6876 34388 6885
rect 27620 6808 27672 6860
rect 32496 6808 32548 6860
rect 42616 6808 42668 6860
rect 44180 6808 44232 6860
rect 44732 6808 44784 6860
rect 46112 6851 46164 6860
rect 46112 6817 46135 6851
rect 46135 6817 46164 6851
rect 46112 6808 46164 6817
rect 27712 6783 27764 6792
rect 27712 6749 27721 6783
rect 27721 6749 27755 6783
rect 27755 6749 27764 6783
rect 27712 6740 27764 6749
rect 37832 6783 37884 6792
rect 37832 6749 37841 6783
rect 37841 6749 37875 6783
rect 37875 6749 37884 6783
rect 37832 6740 37884 6749
rect 43352 6783 43404 6792
rect 43352 6749 43361 6783
rect 43361 6749 43395 6783
rect 43395 6749 43404 6783
rect 43352 6740 43404 6749
rect 45836 6783 45888 6792
rect 45836 6749 45845 6783
rect 45845 6749 45879 6783
rect 45879 6749 45888 6783
rect 45836 6740 45888 6749
rect 4712 6604 4764 6656
rect 5632 6604 5684 6656
rect 5724 6604 5776 6656
rect 6184 6604 6236 6656
rect 9404 6604 9456 6656
rect 11336 6647 11388 6656
rect 11336 6613 11345 6647
rect 11345 6613 11379 6647
rect 11379 6613 11388 6647
rect 11336 6604 11388 6613
rect 13360 6604 13412 6656
rect 15752 6604 15804 6656
rect 15936 6604 15988 6656
rect 23756 6647 23808 6656
rect 23756 6613 23765 6647
rect 23765 6613 23799 6647
rect 23799 6613 23808 6647
rect 23756 6604 23808 6613
rect 26240 6647 26292 6656
rect 26240 6613 26249 6647
rect 26249 6613 26283 6647
rect 26283 6613 26292 6647
rect 26240 6604 26292 6613
rect 26516 6604 26568 6656
rect 29092 6647 29144 6656
rect 29092 6613 29101 6647
rect 29101 6613 29135 6647
rect 29135 6613 29144 6647
rect 29092 6604 29144 6613
rect 30564 6604 30616 6656
rect 31208 6647 31260 6656
rect 31208 6613 31217 6647
rect 31217 6613 31251 6647
rect 31251 6613 31260 6647
rect 31208 6604 31260 6613
rect 32496 6647 32548 6656
rect 32496 6613 32505 6647
rect 32505 6613 32539 6647
rect 32539 6613 32548 6647
rect 32496 6604 32548 6613
rect 33324 6647 33376 6656
rect 33324 6613 33333 6647
rect 33333 6613 33367 6647
rect 33367 6613 33376 6647
rect 33324 6604 33376 6613
rect 33692 6647 33744 6656
rect 33692 6613 33701 6647
rect 33701 6613 33735 6647
rect 33735 6613 33744 6647
rect 33692 6604 33744 6613
rect 33876 6647 33928 6656
rect 33876 6613 33885 6647
rect 33885 6613 33919 6647
rect 33919 6613 33928 6647
rect 33876 6604 33928 6613
rect 35256 6647 35308 6656
rect 35256 6613 35265 6647
rect 35265 6613 35299 6647
rect 35299 6613 35308 6647
rect 35256 6604 35308 6613
rect 44732 6647 44784 6656
rect 44732 6613 44741 6647
rect 44741 6613 44775 6647
rect 44775 6613 44784 6647
rect 44732 6604 44784 6613
rect 45376 6647 45428 6656
rect 45376 6613 45385 6647
rect 45385 6613 45419 6647
rect 45419 6613 45428 6647
rect 45376 6604 45428 6613
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 34966 6502 35018 6554
rect 35030 6502 35082 6554
rect 35094 6502 35146 6554
rect 35158 6502 35210 6554
rect 3332 6400 3384 6452
rect 6276 6443 6328 6452
rect 6276 6409 6285 6443
rect 6285 6409 6319 6443
rect 6319 6409 6328 6443
rect 6276 6400 6328 6409
rect 9312 6400 9364 6452
rect 8208 6375 8260 6384
rect 8208 6341 8217 6375
rect 8217 6341 8251 6375
rect 8251 6341 8260 6375
rect 8208 6332 8260 6341
rect 9404 6264 9456 6316
rect 10048 6400 10100 6452
rect 11612 6443 11664 6452
rect 11612 6409 11621 6443
rect 11621 6409 11655 6443
rect 11655 6409 11664 6443
rect 11612 6400 11664 6409
rect 11796 6400 11848 6452
rect 16396 6443 16448 6452
rect 16396 6409 16405 6443
rect 16405 6409 16439 6443
rect 16439 6409 16448 6443
rect 16396 6400 16448 6409
rect 17960 6400 18012 6452
rect 18236 6400 18288 6452
rect 13636 6332 13688 6384
rect 16488 6332 16540 6384
rect 15844 6264 15896 6316
rect 21916 6400 21968 6452
rect 22928 6400 22980 6452
rect 23848 6400 23900 6452
rect 24860 6400 24912 6452
rect 25504 6400 25556 6452
rect 7840 6196 7892 6248
rect 4620 6128 4672 6180
rect 8668 6171 8720 6180
rect 8668 6137 8677 6171
rect 8677 6137 8711 6171
rect 8711 6137 8720 6171
rect 8668 6128 8720 6137
rect 10232 6196 10284 6248
rect 13360 6239 13412 6248
rect 13360 6205 13369 6239
rect 13369 6205 13403 6239
rect 13403 6205 13412 6239
rect 13360 6196 13412 6205
rect 15752 6239 15804 6248
rect 15752 6205 15761 6239
rect 15761 6205 15795 6239
rect 15795 6205 15804 6239
rect 15752 6196 15804 6205
rect 23756 6196 23808 6248
rect 13084 6128 13136 6180
rect 15936 6171 15988 6180
rect 15936 6137 15945 6171
rect 15945 6137 15979 6171
rect 15979 6137 15988 6171
rect 15936 6128 15988 6137
rect 19984 6171 20036 6180
rect 19984 6137 20018 6171
rect 20018 6137 20036 6171
rect 19984 6128 20036 6137
rect 21364 6128 21416 6180
rect 26424 6400 26476 6452
rect 26608 6400 26660 6452
rect 27712 6443 27764 6452
rect 27712 6409 27721 6443
rect 27721 6409 27755 6443
rect 27755 6409 27764 6443
rect 27712 6400 27764 6409
rect 29184 6400 29236 6452
rect 31208 6400 31260 6452
rect 33784 6400 33836 6452
rect 42616 6443 42668 6452
rect 42616 6409 42625 6443
rect 42625 6409 42659 6443
rect 42659 6409 42668 6443
rect 42616 6400 42668 6409
rect 43076 6400 43128 6452
rect 46112 6400 46164 6452
rect 26240 6375 26292 6384
rect 26240 6341 26249 6375
rect 26249 6341 26283 6375
rect 26283 6341 26292 6375
rect 26240 6332 26292 6341
rect 33140 6332 33192 6384
rect 35532 6332 35584 6384
rect 37740 6375 37792 6384
rect 37740 6341 37749 6375
rect 37749 6341 37783 6375
rect 37783 6341 37792 6375
rect 37740 6332 37792 6341
rect 43444 6375 43496 6384
rect 43444 6341 43453 6375
rect 43453 6341 43487 6375
rect 43487 6341 43496 6375
rect 43444 6332 43496 6341
rect 32404 6307 32456 6316
rect 32404 6273 32413 6307
rect 32413 6273 32447 6307
rect 32447 6273 32456 6307
rect 32404 6264 32456 6273
rect 33324 6264 33376 6316
rect 36268 6264 36320 6316
rect 26240 6196 26292 6248
rect 26516 6171 26568 6180
rect 3240 6060 3292 6112
rect 4804 6060 4856 6112
rect 5908 6103 5960 6112
rect 5908 6069 5917 6103
rect 5917 6069 5951 6103
rect 5951 6069 5960 6103
rect 5908 6060 5960 6069
rect 6736 6060 6788 6112
rect 12900 6103 12952 6112
rect 12900 6069 12909 6103
rect 12909 6069 12943 6103
rect 12943 6069 12952 6103
rect 12900 6060 12952 6069
rect 13728 6060 13780 6112
rect 14096 6103 14148 6112
rect 14096 6069 14105 6103
rect 14105 6069 14139 6103
rect 14139 6069 14148 6103
rect 14096 6060 14148 6069
rect 18052 6103 18104 6112
rect 18052 6069 18061 6103
rect 18061 6069 18095 6103
rect 18095 6069 18104 6103
rect 18052 6060 18104 6069
rect 21548 6060 21600 6112
rect 26516 6137 26525 6171
rect 26525 6137 26559 6171
rect 26559 6137 26568 6171
rect 26516 6128 26568 6137
rect 27620 6128 27672 6180
rect 29000 6128 29052 6180
rect 30564 6171 30616 6180
rect 30564 6137 30598 6171
rect 30598 6137 30616 6171
rect 30564 6128 30616 6137
rect 33324 6171 33376 6180
rect 33324 6137 33333 6171
rect 33333 6137 33367 6171
rect 33367 6137 33376 6171
rect 33324 6128 33376 6137
rect 35256 6196 35308 6248
rect 33600 6128 33652 6180
rect 26884 6060 26936 6112
rect 29644 6103 29696 6112
rect 29644 6069 29653 6103
rect 29653 6069 29687 6103
rect 29687 6069 29696 6103
rect 29644 6060 29696 6069
rect 29920 6060 29972 6112
rect 33876 6060 33928 6112
rect 37832 6196 37884 6248
rect 45376 6264 45428 6316
rect 39304 6239 39356 6248
rect 39304 6205 39313 6239
rect 39313 6205 39347 6239
rect 39347 6205 39356 6239
rect 39304 6196 39356 6205
rect 44364 6239 44416 6248
rect 44364 6205 44373 6239
rect 44373 6205 44407 6239
rect 44407 6205 44416 6239
rect 44364 6196 44416 6205
rect 38292 6171 38344 6180
rect 38292 6137 38301 6171
rect 38301 6137 38335 6171
rect 38335 6137 38344 6171
rect 38292 6128 38344 6137
rect 38660 6060 38712 6112
rect 39856 6060 39908 6112
rect 43812 6060 43864 6112
rect 44732 6060 44784 6112
rect 45928 6103 45980 6112
rect 45928 6069 45937 6103
rect 45937 6069 45971 6103
rect 45971 6069 45980 6103
rect 45928 6060 45980 6069
rect 19606 5958 19658 6010
rect 19670 5958 19722 6010
rect 19734 5958 19786 6010
rect 19798 5958 19850 6010
rect 3332 5856 3384 5908
rect 4620 5899 4672 5908
rect 4620 5865 4629 5899
rect 4629 5865 4663 5899
rect 4663 5865 4672 5899
rect 4620 5856 4672 5865
rect 6920 5856 6972 5908
rect 10232 5856 10284 5908
rect 11980 5899 12032 5908
rect 11980 5865 11989 5899
rect 11989 5865 12023 5899
rect 12023 5865 12032 5899
rect 11980 5856 12032 5865
rect 13360 5856 13412 5908
rect 14004 5856 14056 5908
rect 15476 5899 15528 5908
rect 15476 5865 15485 5899
rect 15485 5865 15519 5899
rect 15519 5865 15528 5899
rect 15476 5856 15528 5865
rect 22100 5856 22152 5908
rect 23112 5856 23164 5908
rect 26516 5856 26568 5908
rect 33692 5856 33744 5908
rect 36268 5899 36320 5908
rect 6184 5831 6236 5840
rect 6184 5797 6218 5831
rect 6218 5797 6236 5831
rect 6184 5788 6236 5797
rect 11520 5831 11572 5840
rect 11520 5797 11529 5831
rect 11529 5797 11563 5831
rect 11563 5797 11572 5831
rect 11520 5788 11572 5797
rect 12900 5788 12952 5840
rect 16120 5788 16172 5840
rect 8208 5720 8260 5772
rect 9220 5720 9272 5772
rect 10048 5720 10100 5772
rect 11336 5763 11388 5772
rect 11336 5729 11345 5763
rect 11345 5729 11379 5763
rect 11379 5729 11388 5763
rect 11336 5720 11388 5729
rect 12440 5720 12492 5772
rect 15752 5763 15804 5772
rect 15752 5729 15761 5763
rect 15761 5729 15795 5763
rect 15795 5729 15804 5763
rect 15752 5720 15804 5729
rect 17684 5720 17736 5772
rect 18236 5788 18288 5840
rect 20904 5788 20956 5840
rect 21548 5831 21600 5840
rect 21548 5797 21557 5831
rect 21557 5797 21591 5831
rect 21591 5797 21600 5831
rect 21548 5788 21600 5797
rect 26608 5788 26660 5840
rect 27068 5788 27120 5840
rect 27528 5788 27580 5840
rect 29092 5788 29144 5840
rect 18512 5763 18564 5772
rect 4712 5695 4764 5704
rect 4712 5661 4721 5695
rect 4721 5661 4755 5695
rect 4755 5661 4764 5695
rect 5908 5695 5960 5704
rect 4712 5652 4764 5661
rect 5908 5661 5917 5695
rect 5917 5661 5951 5695
rect 5951 5661 5960 5695
rect 5908 5652 5960 5661
rect 11612 5695 11664 5704
rect 11612 5661 11621 5695
rect 11621 5661 11655 5695
rect 11655 5661 11664 5695
rect 11612 5652 11664 5661
rect 4804 5584 4856 5636
rect 5724 5516 5776 5568
rect 11060 5627 11112 5636
rect 11060 5593 11069 5627
rect 11069 5593 11103 5627
rect 11103 5593 11112 5627
rect 11060 5584 11112 5593
rect 6276 5516 6328 5568
rect 8300 5559 8352 5568
rect 8300 5525 8309 5559
rect 8309 5525 8343 5559
rect 8343 5525 8352 5559
rect 8300 5516 8352 5525
rect 8760 5516 8812 5568
rect 8852 5516 8904 5568
rect 9496 5559 9548 5568
rect 9496 5525 9505 5559
rect 9505 5525 9539 5559
rect 9539 5525 9548 5559
rect 9496 5516 9548 5525
rect 18512 5729 18535 5763
rect 18535 5729 18564 5763
rect 18512 5720 18564 5729
rect 20536 5720 20588 5772
rect 22100 5720 22152 5772
rect 23296 5763 23348 5772
rect 23296 5729 23305 5763
rect 23305 5729 23339 5763
rect 23339 5729 23348 5763
rect 23296 5720 23348 5729
rect 26424 5720 26476 5772
rect 27160 5720 27212 5772
rect 29000 5720 29052 5772
rect 32312 5720 32364 5772
rect 36268 5865 36277 5899
rect 36277 5865 36311 5899
rect 36311 5865 36320 5899
rect 36268 5856 36320 5865
rect 38200 5899 38252 5908
rect 38200 5865 38211 5899
rect 38211 5865 38245 5899
rect 38245 5865 38252 5899
rect 42064 5899 42116 5908
rect 38200 5856 38252 5865
rect 42064 5865 42073 5899
rect 42073 5865 42107 5899
rect 42107 5865 42116 5899
rect 42064 5856 42116 5865
rect 43812 5899 43864 5908
rect 43812 5865 43821 5899
rect 43821 5865 43855 5899
rect 43855 5865 43864 5899
rect 43812 5856 43864 5865
rect 44364 5856 44416 5908
rect 37740 5788 37792 5840
rect 35440 5720 35492 5772
rect 40684 5763 40736 5772
rect 18236 5695 18288 5704
rect 18236 5661 18245 5695
rect 18245 5661 18279 5695
rect 18279 5661 18288 5695
rect 18236 5652 18288 5661
rect 22560 5695 22612 5704
rect 20996 5627 21048 5636
rect 20996 5593 21005 5627
rect 21005 5593 21039 5627
rect 21039 5593 21048 5627
rect 20996 5584 21048 5593
rect 22560 5661 22569 5695
rect 22569 5661 22603 5695
rect 22603 5661 22612 5695
rect 22560 5652 22612 5661
rect 23020 5695 23072 5704
rect 23020 5661 23029 5695
rect 23029 5661 23063 5695
rect 23063 5661 23072 5695
rect 23020 5652 23072 5661
rect 31852 5652 31904 5704
rect 19984 5516 20036 5568
rect 20628 5516 20680 5568
rect 24032 5516 24084 5568
rect 27620 5516 27672 5568
rect 30748 5516 30800 5568
rect 34612 5652 34664 5704
rect 36544 5652 36596 5704
rect 37096 5652 37148 5704
rect 40684 5729 40693 5763
rect 40693 5729 40727 5763
rect 40727 5729 40736 5763
rect 40684 5720 40736 5729
rect 40960 5763 41012 5772
rect 40960 5729 40994 5763
rect 40994 5729 41012 5763
rect 40960 5720 41012 5729
rect 38476 5695 38528 5704
rect 38476 5661 38485 5695
rect 38485 5661 38519 5695
rect 38519 5661 38528 5695
rect 38476 5652 38528 5661
rect 33048 5516 33100 5568
rect 33600 5516 33652 5568
rect 34336 5559 34388 5568
rect 34336 5525 34345 5559
rect 34345 5525 34379 5559
rect 34379 5525 34388 5559
rect 34336 5516 34388 5525
rect 39948 5516 40000 5568
rect 40684 5516 40736 5568
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 34966 5414 35018 5466
rect 35030 5414 35082 5466
rect 35094 5414 35146 5466
rect 35158 5414 35210 5466
rect 3332 5312 3384 5364
rect 4620 5312 4672 5364
rect 6184 5312 6236 5364
rect 8208 5312 8260 5364
rect 9220 5355 9272 5364
rect 9220 5321 9229 5355
rect 9229 5321 9263 5355
rect 9263 5321 9272 5355
rect 9220 5312 9272 5321
rect 11336 5312 11388 5364
rect 11520 5312 11572 5364
rect 12440 5312 12492 5364
rect 15752 5355 15804 5364
rect 9588 5244 9640 5296
rect 15752 5321 15761 5355
rect 15761 5321 15795 5355
rect 15795 5321 15804 5355
rect 15752 5312 15804 5321
rect 17408 5355 17460 5364
rect 17408 5321 17417 5355
rect 17417 5321 17451 5355
rect 17451 5321 17460 5355
rect 17408 5312 17460 5321
rect 18052 5312 18104 5364
rect 18236 5312 18288 5364
rect 20536 5355 20588 5364
rect 13544 5176 13596 5228
rect 19432 5244 19484 5296
rect 20536 5321 20545 5355
rect 20545 5321 20579 5355
rect 20579 5321 20588 5355
rect 20536 5312 20588 5321
rect 23112 5355 23164 5364
rect 23112 5321 23121 5355
rect 23121 5321 23155 5355
rect 23155 5321 23164 5355
rect 23112 5312 23164 5321
rect 23480 5355 23532 5364
rect 23480 5321 23489 5355
rect 23489 5321 23523 5355
rect 23523 5321 23532 5355
rect 23480 5312 23532 5321
rect 23756 5355 23808 5364
rect 23756 5321 23765 5355
rect 23765 5321 23799 5355
rect 23799 5321 23808 5355
rect 23756 5312 23808 5321
rect 26884 5312 26936 5364
rect 27160 5355 27212 5364
rect 27160 5321 27169 5355
rect 27169 5321 27203 5355
rect 27203 5321 27212 5355
rect 27160 5312 27212 5321
rect 28448 5312 28500 5364
rect 29092 5312 29144 5364
rect 33048 5312 33100 5364
rect 34612 5312 34664 5364
rect 35440 5355 35492 5364
rect 35440 5321 35449 5355
rect 35449 5321 35483 5355
rect 35483 5321 35492 5355
rect 35440 5312 35492 5321
rect 3332 5040 3384 5092
rect 4068 5040 4120 5092
rect 6828 5151 6880 5160
rect 6828 5117 6837 5151
rect 6837 5117 6871 5151
rect 6871 5117 6880 5151
rect 6828 5108 6880 5117
rect 11244 5151 11296 5160
rect 11244 5117 11253 5151
rect 11253 5117 11287 5151
rect 11287 5117 11296 5151
rect 11244 5108 11296 5117
rect 8852 5083 8904 5092
rect 8852 5049 8861 5083
rect 8861 5049 8895 5083
rect 8895 5049 8904 5083
rect 8852 5040 8904 5049
rect 4160 4972 4212 5024
rect 4804 4972 4856 5024
rect 5540 5015 5592 5024
rect 5540 4981 5549 5015
rect 5549 4981 5583 5015
rect 5583 4981 5592 5015
rect 5540 4972 5592 4981
rect 5816 5015 5868 5024
rect 5816 4981 5825 5015
rect 5825 4981 5859 5015
rect 5859 4981 5868 5015
rect 5816 4972 5868 4981
rect 6276 5015 6328 5024
rect 6276 4981 6285 5015
rect 6285 4981 6319 5015
rect 6319 4981 6328 5015
rect 6276 4972 6328 4981
rect 8760 5015 8812 5024
rect 8760 4981 8769 5015
rect 8769 4981 8803 5015
rect 8803 4981 8812 5015
rect 8760 4972 8812 4981
rect 11612 4972 11664 5024
rect 11704 4972 11756 5024
rect 14004 5151 14056 5160
rect 14004 5117 14038 5151
rect 14038 5117 14056 5151
rect 14004 5108 14056 5117
rect 18512 5040 18564 5092
rect 15108 5015 15160 5024
rect 15108 4981 15117 5015
rect 15117 4981 15151 5015
rect 15151 4981 15160 5015
rect 15108 4972 15160 4981
rect 16120 5015 16172 5024
rect 16120 4981 16129 5015
rect 16129 4981 16163 5015
rect 16163 4981 16172 5015
rect 16120 4972 16172 4981
rect 17408 4972 17460 5024
rect 19340 4972 19392 5024
rect 25964 5244 26016 5296
rect 26608 5244 26660 5296
rect 24216 5176 24268 5228
rect 24768 5176 24820 5228
rect 29000 5219 29052 5228
rect 21088 5151 21140 5160
rect 21088 5117 21097 5151
rect 21097 5117 21131 5151
rect 21131 5117 21140 5151
rect 21088 5108 21140 5117
rect 26608 5108 26660 5160
rect 21548 5040 21600 5092
rect 19984 5015 20036 5024
rect 19984 4981 19993 5015
rect 19993 4981 20027 5015
rect 20027 4981 20036 5015
rect 19984 4972 20036 4981
rect 22744 5040 22796 5092
rect 23664 5040 23716 5092
rect 23572 4972 23624 5024
rect 25964 5015 26016 5024
rect 25964 4981 25973 5015
rect 25973 4981 26007 5015
rect 26007 4981 26016 5015
rect 25964 4972 26016 4981
rect 26056 4972 26108 5024
rect 29000 5185 29009 5219
rect 29009 5185 29043 5219
rect 29043 5185 29052 5219
rect 29000 5176 29052 5185
rect 29920 5219 29972 5228
rect 29920 5185 29929 5219
rect 29929 5185 29963 5219
rect 29963 5185 29972 5219
rect 29920 5176 29972 5185
rect 37188 5312 37240 5364
rect 38660 5355 38712 5364
rect 38660 5321 38669 5355
rect 38669 5321 38703 5355
rect 38703 5321 38712 5355
rect 38660 5312 38712 5321
rect 31852 5108 31904 5160
rect 30748 5083 30800 5092
rect 30748 5049 30757 5083
rect 30757 5049 30791 5083
rect 30791 5049 30800 5083
rect 30748 5040 30800 5049
rect 31392 5040 31444 5092
rect 29092 4972 29144 5024
rect 32312 4972 32364 5024
rect 34612 4972 34664 5024
rect 40592 5108 40644 5160
rect 36268 5040 36320 5092
rect 37372 5040 37424 5092
rect 38476 5040 38528 5092
rect 37464 5015 37516 5024
rect 37464 4981 37473 5015
rect 37473 4981 37507 5015
rect 37507 4981 37516 5015
rect 37464 4972 37516 4981
rect 38200 4972 38252 5024
rect 39120 5015 39172 5024
rect 39120 4981 39129 5015
rect 39129 4981 39163 5015
rect 39163 4981 39172 5015
rect 39120 4972 39172 4981
rect 40684 5040 40736 5092
rect 40960 4972 41012 5024
rect 19606 4870 19658 4922
rect 19670 4870 19722 4922
rect 19734 4870 19786 4922
rect 19798 4870 19850 4922
rect 3332 4768 3384 4820
rect 4620 4768 4672 4820
rect 5632 4768 5684 4820
rect 6184 4768 6236 4820
rect 7840 4811 7892 4820
rect 7840 4777 7849 4811
rect 7849 4777 7883 4811
rect 7883 4777 7892 4811
rect 7840 4768 7892 4777
rect 11704 4811 11756 4820
rect 11704 4777 11713 4811
rect 11713 4777 11747 4811
rect 11747 4777 11756 4811
rect 11704 4768 11756 4777
rect 12900 4768 12952 4820
rect 13820 4768 13872 4820
rect 15844 4811 15896 4820
rect 15844 4777 15853 4811
rect 15853 4777 15887 4811
rect 15887 4777 15896 4811
rect 15844 4768 15896 4777
rect 18512 4768 18564 4820
rect 21548 4768 21600 4820
rect 22560 4811 22612 4820
rect 22560 4777 22569 4811
rect 22569 4777 22603 4811
rect 22603 4777 22612 4811
rect 22560 4768 22612 4777
rect 23020 4768 23072 4820
rect 5724 4700 5776 4752
rect 23756 4768 23808 4820
rect 24032 4768 24084 4820
rect 24216 4768 24268 4820
rect 24952 4811 25004 4820
rect 24952 4777 24961 4811
rect 24961 4777 24995 4811
rect 24995 4777 25004 4811
rect 24952 4768 25004 4777
rect 26056 4768 26108 4820
rect 6092 4632 6144 4684
rect 8300 4700 8352 4752
rect 16672 4700 16724 4752
rect 21456 4743 21508 4752
rect 21456 4709 21465 4743
rect 21465 4709 21499 4743
rect 21499 4709 21508 4743
rect 21456 4700 21508 4709
rect 22008 4700 22060 4752
rect 23388 4743 23440 4752
rect 23388 4709 23397 4743
rect 23397 4709 23431 4743
rect 23431 4709 23440 4743
rect 23388 4700 23440 4709
rect 23664 4743 23716 4752
rect 23664 4709 23673 4743
rect 23673 4709 23707 4743
rect 23707 4709 23716 4743
rect 27528 4768 27580 4820
rect 30564 4811 30616 4820
rect 30564 4777 30573 4811
rect 30573 4777 30607 4811
rect 30607 4777 30616 4811
rect 30564 4768 30616 4777
rect 31392 4811 31444 4820
rect 31392 4777 31401 4811
rect 31401 4777 31435 4811
rect 31435 4777 31444 4811
rect 31392 4768 31444 4777
rect 32496 4811 32548 4820
rect 32496 4777 32505 4811
rect 32505 4777 32539 4811
rect 32539 4777 32548 4811
rect 32496 4768 32548 4777
rect 33600 4811 33652 4820
rect 33600 4777 33609 4811
rect 33609 4777 33643 4811
rect 33643 4777 33652 4811
rect 33600 4768 33652 4777
rect 36268 4768 36320 4820
rect 37096 4811 37148 4820
rect 37096 4777 37105 4811
rect 37105 4777 37139 4811
rect 37139 4777 37148 4811
rect 37096 4768 37148 4777
rect 39120 4768 39172 4820
rect 40592 4811 40644 4820
rect 40592 4777 40601 4811
rect 40601 4777 40635 4811
rect 40635 4777 40644 4811
rect 40592 4768 40644 4777
rect 40960 4811 41012 4820
rect 40960 4777 40969 4811
rect 40969 4777 41003 4811
rect 41003 4777 41012 4811
rect 40960 4768 41012 4777
rect 23664 4700 23716 4709
rect 27068 4743 27120 4752
rect 27068 4709 27077 4743
rect 27077 4709 27111 4743
rect 27111 4709 27120 4743
rect 27068 4700 27120 4709
rect 38108 4743 38160 4752
rect 6828 4496 6880 4548
rect 2688 4471 2740 4480
rect 2688 4437 2697 4471
rect 2697 4437 2731 4471
rect 2731 4437 2740 4471
rect 2688 4428 2740 4437
rect 4712 4471 4764 4480
rect 4712 4437 4721 4471
rect 4721 4437 4755 4471
rect 4755 4437 4764 4471
rect 4712 4428 4764 4437
rect 5356 4428 5408 4480
rect 7104 4428 7156 4480
rect 8852 4632 8904 4684
rect 10324 4632 10376 4684
rect 11520 4675 11572 4684
rect 11520 4641 11529 4675
rect 11529 4641 11563 4675
rect 11563 4641 11572 4675
rect 11520 4632 11572 4641
rect 8576 4607 8628 4616
rect 8576 4573 8585 4607
rect 8585 4573 8619 4607
rect 8619 4573 8628 4607
rect 8576 4564 8628 4573
rect 11796 4607 11848 4616
rect 11796 4573 11805 4607
rect 11805 4573 11839 4607
rect 11839 4573 11848 4607
rect 11796 4564 11848 4573
rect 8208 4496 8260 4548
rect 11244 4539 11296 4548
rect 11244 4505 11253 4539
rect 11253 4505 11287 4539
rect 11287 4505 11296 4539
rect 11244 4496 11296 4505
rect 15016 4564 15068 4616
rect 16948 4632 17000 4684
rect 17224 4675 17276 4684
rect 17224 4641 17233 4675
rect 17233 4641 17267 4675
rect 17267 4641 17276 4675
rect 17224 4632 17276 4641
rect 18696 4632 18748 4684
rect 19708 4675 19760 4684
rect 19708 4641 19717 4675
rect 19717 4641 19751 4675
rect 19751 4641 19760 4675
rect 19708 4632 19760 4641
rect 20720 4632 20772 4684
rect 24584 4632 24636 4684
rect 26976 4632 27028 4684
rect 38108 4709 38117 4743
rect 38117 4709 38151 4743
rect 38151 4709 38160 4743
rect 38108 4700 38160 4709
rect 38292 4743 38344 4752
rect 38292 4709 38301 4743
rect 38301 4709 38335 4743
rect 38335 4709 38344 4743
rect 38292 4700 38344 4709
rect 29460 4675 29512 4684
rect 17132 4607 17184 4616
rect 17132 4573 17141 4607
rect 17141 4573 17175 4607
rect 17175 4573 17184 4607
rect 17132 4564 17184 4573
rect 20628 4564 20680 4616
rect 21364 4607 21416 4616
rect 21364 4573 21373 4607
rect 21373 4573 21407 4607
rect 21407 4573 21416 4607
rect 21364 4564 21416 4573
rect 21548 4607 21600 4616
rect 21548 4573 21557 4607
rect 21557 4573 21591 4607
rect 21591 4573 21600 4607
rect 21548 4564 21600 4573
rect 25596 4607 25648 4616
rect 25596 4573 25605 4607
rect 25605 4573 25639 4607
rect 25639 4573 25648 4607
rect 25596 4564 25648 4573
rect 16212 4496 16264 4548
rect 20720 4496 20772 4548
rect 20904 4496 20956 4548
rect 23572 4496 23624 4548
rect 26608 4539 26660 4548
rect 26608 4505 26617 4539
rect 26617 4505 26651 4539
rect 26651 4505 26660 4539
rect 26608 4496 26660 4505
rect 10232 4471 10284 4480
rect 10232 4437 10241 4471
rect 10241 4437 10275 4471
rect 10275 4437 10284 4471
rect 10232 4428 10284 4437
rect 11060 4471 11112 4480
rect 11060 4437 11069 4471
rect 11069 4437 11103 4471
rect 11103 4437 11112 4471
rect 11060 4428 11112 4437
rect 12808 4471 12860 4480
rect 12808 4437 12817 4471
rect 12817 4437 12851 4471
rect 12851 4437 12860 4471
rect 12808 4428 12860 4437
rect 13176 4471 13228 4480
rect 13176 4437 13185 4471
rect 13185 4437 13219 4471
rect 13219 4437 13228 4471
rect 13176 4428 13228 4437
rect 13452 4471 13504 4480
rect 13452 4437 13461 4471
rect 13461 4437 13495 4471
rect 13495 4437 13504 4471
rect 13452 4428 13504 4437
rect 13820 4428 13872 4480
rect 14096 4428 14148 4480
rect 15016 4471 15068 4480
rect 15016 4437 15025 4471
rect 15025 4437 15059 4471
rect 15059 4437 15068 4471
rect 15016 4428 15068 4437
rect 15476 4471 15528 4480
rect 15476 4437 15485 4471
rect 15485 4437 15519 4471
rect 15519 4437 15528 4471
rect 15476 4428 15528 4437
rect 17960 4428 18012 4480
rect 20536 4428 20588 4480
rect 24400 4471 24452 4480
rect 24400 4437 24409 4471
rect 24409 4437 24443 4471
rect 24443 4437 24452 4471
rect 24400 4428 24452 4437
rect 25872 4471 25924 4480
rect 25872 4437 25881 4471
rect 25881 4437 25915 4471
rect 25915 4437 25924 4471
rect 29460 4641 29494 4675
rect 29494 4641 29512 4675
rect 29460 4632 29512 4641
rect 32128 4675 32180 4684
rect 32128 4641 32137 4675
rect 32137 4641 32171 4675
rect 32171 4641 32180 4675
rect 32128 4632 32180 4641
rect 32312 4675 32364 4684
rect 32312 4641 32321 4675
rect 32321 4641 32355 4675
rect 32355 4641 32364 4675
rect 32312 4632 32364 4641
rect 33140 4632 33192 4684
rect 37464 4632 37516 4684
rect 29000 4564 29052 4616
rect 31852 4539 31904 4548
rect 31852 4505 31861 4539
rect 31861 4505 31895 4539
rect 31895 4505 31904 4539
rect 31852 4496 31904 4505
rect 37372 4496 37424 4548
rect 27712 4471 27764 4480
rect 25872 4428 25924 4437
rect 27712 4437 27721 4471
rect 27721 4437 27755 4471
rect 27755 4437 27764 4471
rect 27712 4428 27764 4437
rect 28356 4428 28408 4480
rect 33048 4428 33100 4480
rect 33232 4471 33284 4480
rect 33232 4437 33241 4471
rect 33241 4437 33275 4471
rect 33275 4437 33284 4471
rect 33232 4428 33284 4437
rect 37832 4471 37884 4480
rect 37832 4437 37841 4471
rect 37841 4437 37875 4471
rect 37875 4437 37884 4471
rect 37832 4428 37884 4437
rect 40500 4428 40552 4480
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 34966 4326 35018 4378
rect 35030 4326 35082 4378
rect 35094 4326 35146 4378
rect 35158 4326 35210 4378
rect 6184 4267 6236 4276
rect 6184 4233 6193 4267
rect 6193 4233 6227 4267
rect 6227 4233 6236 4267
rect 6184 4224 6236 4233
rect 7840 4224 7892 4276
rect 8300 4224 8352 4276
rect 8576 4224 8628 4276
rect 11796 4224 11848 4276
rect 13452 4224 13504 4276
rect 16212 4267 16264 4276
rect 16212 4233 16221 4267
rect 16221 4233 16255 4267
rect 16255 4233 16264 4267
rect 16212 4224 16264 4233
rect 16672 4267 16724 4276
rect 16672 4233 16681 4267
rect 16681 4233 16715 4267
rect 16715 4233 16724 4267
rect 16672 4224 16724 4233
rect 17132 4224 17184 4276
rect 21456 4224 21508 4276
rect 22744 4267 22796 4276
rect 22744 4233 22753 4267
rect 22753 4233 22787 4267
rect 22787 4233 22796 4267
rect 22744 4224 22796 4233
rect 23388 4267 23440 4276
rect 23388 4233 23397 4267
rect 23397 4233 23431 4267
rect 23431 4233 23440 4267
rect 23388 4224 23440 4233
rect 25872 4224 25924 4276
rect 29000 4267 29052 4276
rect 29000 4233 29009 4267
rect 29009 4233 29043 4267
rect 29043 4233 29052 4267
rect 29000 4224 29052 4233
rect 33140 4224 33192 4276
rect 37464 4224 37516 4276
rect 38108 4224 38160 4276
rect 5172 4156 5224 4208
rect 5356 4156 5408 4208
rect 5816 4156 5868 4208
rect 5632 4131 5684 4140
rect 5632 4097 5641 4131
rect 5641 4097 5675 4131
rect 5675 4097 5684 4131
rect 5632 4088 5684 4097
rect 8116 4088 8168 4140
rect 11520 4156 11572 4208
rect 11980 4199 12032 4208
rect 11980 4165 11989 4199
rect 11989 4165 12023 4199
rect 12023 4165 12032 4199
rect 11980 4156 12032 4165
rect 11704 4131 11756 4140
rect 11704 4097 11713 4131
rect 11713 4097 11747 4131
rect 11747 4097 11756 4131
rect 11704 4088 11756 4097
rect 13176 4131 13228 4140
rect 13176 4097 13185 4131
rect 13185 4097 13219 4131
rect 13219 4097 13228 4131
rect 13176 4088 13228 4097
rect 13360 4131 13412 4140
rect 13360 4097 13369 4131
rect 13369 4097 13403 4131
rect 13403 4097 13412 4131
rect 13360 4088 13412 4097
rect 2780 3952 2832 4004
rect 4068 3952 4120 4004
rect 4712 3995 4764 4004
rect 4712 3961 4721 3995
rect 4721 3961 4755 3995
rect 4755 3961 4764 3995
rect 5816 3995 5868 4004
rect 4712 3952 4764 3961
rect 5816 3961 5825 3995
rect 5825 3961 5859 3995
rect 5859 3961 5868 3995
rect 5816 3952 5868 3961
rect 2596 3884 2648 3936
rect 2964 3884 3016 3936
rect 5080 3927 5132 3936
rect 5080 3893 5089 3927
rect 5089 3893 5123 3927
rect 5123 3893 5132 3927
rect 8760 3995 8812 4004
rect 8760 3961 8769 3995
rect 8769 3961 8803 3995
rect 8803 3961 8812 3995
rect 8760 3952 8812 3961
rect 11060 4063 11112 4072
rect 11060 4029 11069 4063
rect 11069 4029 11103 4063
rect 11103 4029 11112 4063
rect 11060 4020 11112 4029
rect 12348 4020 12400 4072
rect 12808 4020 12860 4072
rect 13544 3952 13596 4004
rect 19432 4088 19484 4140
rect 19524 4088 19576 4140
rect 21364 4156 21416 4208
rect 20720 4088 20772 4140
rect 25964 4088 26016 4140
rect 27712 4088 27764 4140
rect 29552 4088 29604 4140
rect 32312 4156 32364 4208
rect 33600 4131 33652 4140
rect 15108 4020 15160 4072
rect 16856 4020 16908 4072
rect 17776 4020 17828 4072
rect 18696 4063 18748 4072
rect 18696 4029 18705 4063
rect 18705 4029 18739 4063
rect 18739 4029 18748 4063
rect 18696 4020 18748 4029
rect 19340 4020 19392 4072
rect 19708 4063 19760 4072
rect 19708 4029 19717 4063
rect 19717 4029 19751 4063
rect 19751 4029 19760 4063
rect 19708 4020 19760 4029
rect 20260 4020 20312 4072
rect 23572 4020 23624 4072
rect 24768 4063 24820 4072
rect 24768 4029 24777 4063
rect 24777 4029 24811 4063
rect 24811 4029 24820 4063
rect 24768 4020 24820 4029
rect 5080 3884 5132 3893
rect 7748 3884 7800 3936
rect 8300 3884 8352 3936
rect 9220 3927 9272 3936
rect 9220 3893 9229 3927
rect 9229 3893 9263 3927
rect 9263 3893 9272 3927
rect 9220 3884 9272 3893
rect 10324 3927 10376 3936
rect 10324 3893 10333 3927
rect 10333 3893 10367 3927
rect 10367 3893 10376 3927
rect 10324 3884 10376 3893
rect 15660 3927 15712 3936
rect 15660 3893 15669 3927
rect 15669 3893 15703 3927
rect 15703 3893 15712 3927
rect 15660 3884 15712 3893
rect 16948 3927 17000 3936
rect 16948 3893 16957 3927
rect 16957 3893 16991 3927
rect 16991 3893 17000 3927
rect 16948 3884 17000 3893
rect 17868 3927 17920 3936
rect 17868 3893 17877 3927
rect 17877 3893 17911 3927
rect 17911 3893 17920 3927
rect 18604 3927 18656 3936
rect 17868 3884 17920 3893
rect 18604 3893 18613 3927
rect 18613 3893 18647 3927
rect 18647 3893 18656 3927
rect 18604 3884 18656 3893
rect 20168 3927 20220 3936
rect 20168 3893 20177 3927
rect 20177 3893 20211 3927
rect 20211 3893 20220 3927
rect 20168 3884 20220 3893
rect 20812 3952 20864 4004
rect 23112 3927 23164 3936
rect 23112 3893 23121 3927
rect 23121 3893 23155 3927
rect 23155 3893 23164 3927
rect 23112 3884 23164 3893
rect 24952 3952 25004 4004
rect 26240 3995 26292 4004
rect 26240 3961 26249 3995
rect 26249 3961 26283 3995
rect 26283 3961 26292 3995
rect 26240 3952 26292 3961
rect 27620 3952 27672 4004
rect 29000 4020 29052 4072
rect 29276 4063 29328 4072
rect 29276 4029 29285 4063
rect 29285 4029 29319 4063
rect 29319 4029 29328 4063
rect 29276 4020 29328 4029
rect 30380 4063 30432 4072
rect 30380 4029 30389 4063
rect 30389 4029 30423 4063
rect 30423 4029 30432 4063
rect 30380 4020 30432 4029
rect 24584 3927 24636 3936
rect 24584 3893 24593 3927
rect 24593 3893 24627 3927
rect 24627 3893 24636 3927
rect 24584 3884 24636 3893
rect 26332 3927 26384 3936
rect 26332 3893 26341 3927
rect 26341 3893 26375 3927
rect 26375 3893 26384 3927
rect 26332 3884 26384 3893
rect 26608 3884 26660 3936
rect 28080 3884 28132 3936
rect 28172 3927 28224 3936
rect 28172 3893 28181 3927
rect 28181 3893 28215 3927
rect 28215 3893 28224 3927
rect 28632 3927 28684 3936
rect 28172 3884 28224 3893
rect 28632 3893 28641 3927
rect 28641 3893 28675 3927
rect 28675 3893 28684 3927
rect 28632 3884 28684 3893
rect 30288 3952 30340 4004
rect 32588 3952 32640 4004
rect 33600 4097 33609 4131
rect 33609 4097 33643 4131
rect 33643 4097 33652 4131
rect 33600 4088 33652 4097
rect 38292 4088 38344 4140
rect 39856 4131 39908 4140
rect 39856 4097 39865 4131
rect 39865 4097 39899 4131
rect 39899 4097 39908 4131
rect 39856 4088 39908 4097
rect 40408 4088 40460 4140
rect 40500 4063 40552 4072
rect 40500 4029 40509 4063
rect 40509 4029 40543 4063
rect 40543 4029 40552 4063
rect 40500 4020 40552 4029
rect 33232 3995 33284 4004
rect 33232 3961 33241 3995
rect 33241 3961 33275 3995
rect 33275 3961 33284 3995
rect 33232 3952 33284 3961
rect 40040 3952 40092 4004
rect 40776 4020 40828 4072
rect 31484 3927 31536 3936
rect 31484 3893 31493 3927
rect 31493 3893 31527 3927
rect 31527 3893 31536 3927
rect 31484 3884 31536 3893
rect 32128 3927 32180 3936
rect 32128 3893 32137 3927
rect 32137 3893 32171 3927
rect 32171 3893 32180 3927
rect 32128 3884 32180 3893
rect 33048 3884 33100 3936
rect 33140 3927 33192 3936
rect 33140 3893 33149 3927
rect 33149 3893 33183 3927
rect 33183 3893 33192 3927
rect 33140 3884 33192 3893
rect 33968 3884 34020 3936
rect 34888 3927 34940 3936
rect 34888 3893 34897 3927
rect 34897 3893 34931 3927
rect 34931 3893 34940 3927
rect 34888 3884 34940 3893
rect 37372 3884 37424 3936
rect 39396 3927 39448 3936
rect 39396 3893 39405 3927
rect 39405 3893 39439 3927
rect 39439 3893 39448 3927
rect 39396 3884 39448 3893
rect 41052 3884 41104 3936
rect 42340 3927 42392 3936
rect 42340 3893 42349 3927
rect 42349 3893 42383 3927
rect 42383 3893 42392 3927
rect 42340 3884 42392 3893
rect 19606 3782 19658 3834
rect 19670 3782 19722 3834
rect 19734 3782 19786 3834
rect 19798 3782 19850 3834
rect 2320 3723 2372 3732
rect 2320 3689 2329 3723
rect 2329 3689 2363 3723
rect 2363 3689 2372 3723
rect 2964 3723 3016 3732
rect 2320 3680 2372 3689
rect 2964 3689 2973 3723
rect 2973 3689 3007 3723
rect 3007 3689 3016 3723
rect 2964 3680 3016 3689
rect 4620 3680 4672 3732
rect 5724 3723 5776 3732
rect 5724 3689 5733 3723
rect 5733 3689 5767 3723
rect 5767 3689 5776 3723
rect 5724 3680 5776 3689
rect 6092 3723 6144 3732
rect 6092 3689 6101 3723
rect 6101 3689 6135 3723
rect 6135 3689 6144 3723
rect 6092 3680 6144 3689
rect 8208 3723 8260 3732
rect 8208 3689 8217 3723
rect 8217 3689 8251 3723
rect 8251 3689 8260 3723
rect 8208 3680 8260 3689
rect 13636 3723 13688 3732
rect 13636 3689 13645 3723
rect 13645 3689 13679 3723
rect 13679 3689 13688 3723
rect 13636 3680 13688 3689
rect 15476 3680 15528 3732
rect 16764 3680 16816 3732
rect 17224 3723 17276 3732
rect 17224 3689 17233 3723
rect 17233 3689 17267 3723
rect 17267 3689 17276 3723
rect 17224 3680 17276 3689
rect 18604 3680 18656 3732
rect 19432 3680 19484 3732
rect 20076 3680 20128 3732
rect 20260 3723 20312 3732
rect 20260 3689 20269 3723
rect 20269 3689 20303 3723
rect 20303 3689 20312 3723
rect 20260 3680 20312 3689
rect 20720 3680 20772 3732
rect 21548 3723 21600 3732
rect 21548 3689 21557 3723
rect 21557 3689 21591 3723
rect 21591 3689 21600 3723
rect 21548 3680 21600 3689
rect 24400 3680 24452 3732
rect 26148 3680 26200 3732
rect 26240 3680 26292 3732
rect 26976 3680 27028 3732
rect 29460 3723 29512 3732
rect 29460 3689 29469 3723
rect 29469 3689 29503 3723
rect 29503 3689 29512 3723
rect 29460 3680 29512 3689
rect 30472 3723 30524 3732
rect 30472 3689 30481 3723
rect 30481 3689 30515 3723
rect 30515 3689 30524 3723
rect 30472 3680 30524 3689
rect 32680 3680 32732 3732
rect 33968 3723 34020 3732
rect 33968 3689 33977 3723
rect 33977 3689 34011 3723
rect 34011 3689 34020 3723
rect 33968 3680 34020 3689
rect 34520 3723 34572 3732
rect 34520 3689 34529 3723
rect 34529 3689 34563 3723
rect 34563 3689 34572 3723
rect 34520 3680 34572 3689
rect 37832 3680 37884 3732
rect 40776 3723 40828 3732
rect 40776 3689 40785 3723
rect 40785 3689 40819 3723
rect 40819 3689 40828 3723
rect 40776 3680 40828 3689
rect 4712 3612 4764 3664
rect 5632 3612 5684 3664
rect 9496 3612 9548 3664
rect 13176 3612 13228 3664
rect 15660 3612 15712 3664
rect 15844 3612 15896 3664
rect 17132 3612 17184 3664
rect 20168 3612 20220 3664
rect 23940 3612 23992 3664
rect 26332 3612 26384 3664
rect 6092 3544 6144 3596
rect 11244 3544 11296 3596
rect 13820 3587 13872 3596
rect 13820 3553 13829 3587
rect 13829 3553 13863 3587
rect 13863 3553 13872 3587
rect 13820 3544 13872 3553
rect 16948 3544 17000 3596
rect 17684 3544 17736 3596
rect 20720 3544 20772 3596
rect 22100 3544 22152 3596
rect 22376 3587 22428 3596
rect 22376 3553 22385 3587
rect 22385 3553 22419 3587
rect 22419 3553 22428 3587
rect 22376 3544 22428 3553
rect 23480 3544 23532 3596
rect 25596 3544 25648 3596
rect 28632 3612 28684 3664
rect 34888 3612 34940 3664
rect 35256 3612 35308 3664
rect 37464 3655 37516 3664
rect 37464 3621 37473 3655
rect 37473 3621 37507 3655
rect 37507 3621 37516 3655
rect 37464 3612 37516 3621
rect 39396 3612 39448 3664
rect 40224 3655 40276 3664
rect 40224 3621 40233 3655
rect 40233 3621 40267 3655
rect 40267 3621 40276 3655
rect 40224 3612 40276 3621
rect 27712 3544 27764 3596
rect 28356 3587 28408 3596
rect 28356 3553 28390 3587
rect 28390 3553 28408 3587
rect 28356 3544 28408 3553
rect 29092 3544 29144 3596
rect 30932 3587 30984 3596
rect 30932 3553 30941 3587
rect 30941 3553 30975 3587
rect 30975 3553 30984 3587
rect 30932 3544 30984 3553
rect 31944 3587 31996 3596
rect 31944 3553 31953 3587
rect 31953 3553 31987 3587
rect 31987 3553 31996 3587
rect 31944 3544 31996 3553
rect 37372 3544 37424 3596
rect 5172 3519 5224 3528
rect 2504 3451 2556 3460
rect 2504 3417 2513 3451
rect 2513 3417 2547 3451
rect 2547 3417 2556 3451
rect 2504 3408 2556 3417
rect 5172 3485 5181 3519
rect 5181 3485 5215 3519
rect 5215 3485 5224 3519
rect 5172 3476 5224 3485
rect 6184 3519 6236 3528
rect 6184 3485 6193 3519
rect 6193 3485 6227 3519
rect 6227 3485 6236 3519
rect 6184 3476 6236 3485
rect 9588 3476 9640 3528
rect 11336 3519 11388 3528
rect 11336 3485 11345 3519
rect 11345 3485 11379 3519
rect 11379 3485 11388 3519
rect 11336 3476 11388 3485
rect 15108 3476 15160 3528
rect 15844 3476 15896 3528
rect 22836 3476 22888 3528
rect 23756 3476 23808 3528
rect 26424 3476 26476 3528
rect 5448 3408 5500 3460
rect 9220 3408 9272 3460
rect 15476 3451 15528 3460
rect 15476 3417 15485 3451
rect 15485 3417 15519 3451
rect 15519 3417 15528 3451
rect 15476 3408 15528 3417
rect 20720 3451 20772 3460
rect 20720 3417 20729 3451
rect 20729 3417 20763 3451
rect 20763 3417 20772 3451
rect 20720 3408 20772 3417
rect 23848 3451 23900 3460
rect 23848 3417 23857 3451
rect 23857 3417 23891 3451
rect 23891 3417 23900 3451
rect 23848 3408 23900 3417
rect 26608 3451 26660 3460
rect 26608 3417 26617 3451
rect 26617 3417 26651 3451
rect 26651 3417 26660 3451
rect 26608 3408 26660 3417
rect 27620 3451 27672 3460
rect 27620 3417 27629 3451
rect 27629 3417 27663 3451
rect 27663 3417 27672 3451
rect 27620 3408 27672 3417
rect 1676 3383 1728 3392
rect 1676 3349 1685 3383
rect 1685 3349 1719 3383
rect 1719 3349 1728 3383
rect 1676 3340 1728 3349
rect 3516 3383 3568 3392
rect 3516 3349 3525 3383
rect 3525 3349 3559 3383
rect 3559 3349 3568 3383
rect 3516 3340 3568 3349
rect 7656 3340 7708 3392
rect 8300 3340 8352 3392
rect 9496 3383 9548 3392
rect 9496 3349 9505 3383
rect 9505 3349 9539 3383
rect 9539 3349 9548 3383
rect 9496 3340 9548 3349
rect 12716 3383 12768 3392
rect 12716 3349 12725 3383
rect 12725 3349 12759 3383
rect 12759 3349 12768 3383
rect 12716 3340 12768 3349
rect 15016 3340 15068 3392
rect 16488 3383 16540 3392
rect 16488 3349 16497 3383
rect 16497 3349 16531 3383
rect 16531 3349 16540 3383
rect 16488 3340 16540 3349
rect 16856 3383 16908 3392
rect 16856 3349 16865 3383
rect 16865 3349 16899 3383
rect 16899 3349 16908 3383
rect 16856 3340 16908 3349
rect 17776 3383 17828 3392
rect 17776 3349 17785 3383
rect 17785 3349 17819 3383
rect 17819 3349 17828 3383
rect 17776 3340 17828 3349
rect 23480 3340 23532 3392
rect 24860 3383 24912 3392
rect 24860 3349 24869 3383
rect 24869 3349 24903 3383
rect 24903 3349 24912 3383
rect 24860 3340 24912 3349
rect 31852 3476 31904 3528
rect 32588 3519 32640 3528
rect 32588 3485 32597 3519
rect 32597 3485 32631 3519
rect 32631 3485 32640 3519
rect 32588 3476 32640 3485
rect 35348 3476 35400 3528
rect 38568 3476 38620 3528
rect 40684 3476 40736 3528
rect 28816 3340 28868 3392
rect 30380 3340 30432 3392
rect 31116 3383 31168 3392
rect 31116 3349 31125 3383
rect 31125 3349 31159 3383
rect 31159 3349 31168 3383
rect 31116 3340 31168 3349
rect 34520 3340 34572 3392
rect 37832 3383 37884 3392
rect 37832 3349 37841 3383
rect 37841 3349 37875 3383
rect 37875 3349 37884 3383
rect 37832 3340 37884 3349
rect 39764 3383 39816 3392
rect 39764 3349 39773 3383
rect 39773 3349 39807 3383
rect 39807 3349 39816 3383
rect 39764 3340 39816 3349
rect 41052 3383 41104 3392
rect 41052 3349 41061 3383
rect 41061 3349 41095 3383
rect 41095 3349 41104 3383
rect 41052 3340 41104 3349
rect 41144 3340 41196 3392
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 34966 3238 35018 3290
rect 35030 3238 35082 3290
rect 35094 3238 35146 3290
rect 35158 3238 35210 3290
rect 2320 3179 2372 3188
rect 2320 3145 2329 3179
rect 2329 3145 2363 3179
rect 2363 3145 2372 3179
rect 2320 3136 2372 3145
rect 3516 3136 3568 3188
rect 4712 3179 4764 3188
rect 4712 3145 4721 3179
rect 4721 3145 4755 3179
rect 4755 3145 4764 3179
rect 4712 3136 4764 3145
rect 5172 3179 5224 3188
rect 5172 3145 5181 3179
rect 5181 3145 5215 3179
rect 5215 3145 5224 3179
rect 5172 3136 5224 3145
rect 5816 3179 5868 3188
rect 5816 3145 5825 3179
rect 5825 3145 5859 3179
rect 5859 3145 5868 3179
rect 5816 3136 5868 3145
rect 8484 3136 8536 3188
rect 11244 3179 11296 3188
rect 11244 3145 11253 3179
rect 11253 3145 11287 3179
rect 11287 3145 11296 3179
rect 11244 3136 11296 3145
rect 13820 3136 13872 3188
rect 14096 3136 14148 3188
rect 16396 3179 16448 3188
rect 16396 3145 16405 3179
rect 16405 3145 16439 3179
rect 16439 3145 16448 3179
rect 16396 3136 16448 3145
rect 16672 3136 16724 3188
rect 16856 3136 16908 3188
rect 20720 3136 20772 3188
rect 22376 3136 22428 3188
rect 23664 3136 23716 3188
rect 26056 3179 26108 3188
rect 26056 3145 26065 3179
rect 26065 3145 26099 3179
rect 26099 3145 26108 3179
rect 26056 3136 26108 3145
rect 16764 3068 16816 3120
rect 17132 3068 17184 3120
rect 17316 3068 17368 3120
rect 17684 3068 17736 3120
rect 18052 3068 18104 3120
rect 16488 3000 16540 3052
rect 18696 3043 18748 3052
rect 18696 3009 18705 3043
rect 18705 3009 18739 3043
rect 18739 3009 18748 3043
rect 18696 3000 18748 3009
rect 22100 3068 22152 3120
rect 26516 3136 26568 3188
rect 28172 3136 28224 3188
rect 28908 3136 28960 3188
rect 29368 3136 29420 3188
rect 29552 3179 29604 3188
rect 29552 3145 29561 3179
rect 29561 3145 29595 3179
rect 29595 3145 29604 3179
rect 29552 3136 29604 3145
rect 30932 3136 30984 3188
rect 31668 3136 31720 3188
rect 33600 3179 33652 3188
rect 33600 3145 33609 3179
rect 33609 3145 33643 3179
rect 33643 3145 33652 3179
rect 33600 3136 33652 3145
rect 34612 3179 34664 3188
rect 34612 3145 34621 3179
rect 34621 3145 34655 3179
rect 34655 3145 34664 3179
rect 34612 3136 34664 3145
rect 37372 3136 37424 3188
rect 39396 3136 39448 3188
rect 40500 3136 40552 3188
rect 40684 3136 40736 3188
rect 29092 3111 29144 3120
rect 29092 3077 29101 3111
rect 29101 3077 29135 3111
rect 29135 3077 29144 3111
rect 29092 3068 29144 3077
rect 30196 3111 30248 3120
rect 30196 3077 30205 3111
rect 30205 3077 30239 3111
rect 30239 3077 30248 3111
rect 30196 3068 30248 3077
rect 2596 2932 2648 2984
rect 7196 2932 7248 2984
rect 7656 2975 7708 2984
rect 7656 2941 7690 2975
rect 7690 2941 7708 2975
rect 1492 2796 1544 2848
rect 2964 2864 3016 2916
rect 5356 2796 5408 2848
rect 6184 2796 6236 2848
rect 7656 2932 7708 2941
rect 9772 2932 9824 2984
rect 11336 2932 11388 2984
rect 12716 2975 12768 2984
rect 12716 2941 12750 2975
rect 12750 2941 12768 2975
rect 9496 2864 9548 2916
rect 11152 2864 11204 2916
rect 12716 2932 12768 2941
rect 13544 2864 13596 2916
rect 15660 2932 15712 2984
rect 17776 2932 17828 2984
rect 17960 2864 18012 2916
rect 26424 3000 26476 3052
rect 26608 3000 26660 3052
rect 30380 3000 30432 3052
rect 36268 3111 36320 3120
rect 36268 3077 36277 3111
rect 36277 3077 36311 3111
rect 36311 3077 36320 3111
rect 36268 3068 36320 3077
rect 20076 2975 20128 2984
rect 20076 2941 20110 2975
rect 20110 2941 20128 2975
rect 20076 2932 20128 2941
rect 20720 2864 20772 2916
rect 23756 2932 23808 2984
rect 24860 2932 24912 2984
rect 27252 2932 27304 2984
rect 31484 2932 31536 2984
rect 22284 2907 22336 2916
rect 22284 2873 22293 2907
rect 22293 2873 22327 2907
rect 22327 2873 22336 2907
rect 22284 2864 22336 2873
rect 29368 2864 29420 2916
rect 31760 2864 31812 2916
rect 34244 2864 34296 2916
rect 35348 2864 35400 2916
rect 37464 2932 37516 2984
rect 37280 2907 37332 2916
rect 37280 2873 37289 2907
rect 37289 2873 37323 2907
rect 37323 2873 37332 2907
rect 37280 2864 37332 2873
rect 40040 2864 40092 2916
rect 41052 2864 41104 2916
rect 41328 2864 41380 2916
rect 8760 2839 8812 2848
rect 8760 2805 8769 2839
rect 8769 2805 8803 2839
rect 8803 2805 8812 2839
rect 8760 2796 8812 2805
rect 9772 2839 9824 2848
rect 9772 2805 9781 2839
rect 9781 2805 9815 2839
rect 9815 2805 9824 2839
rect 9772 2796 9824 2805
rect 13912 2796 13964 2848
rect 21180 2839 21232 2848
rect 21180 2805 21189 2839
rect 21189 2805 21223 2839
rect 21223 2805 21232 2839
rect 21180 2796 21232 2805
rect 24768 2796 24820 2848
rect 25596 2839 25648 2848
rect 25596 2805 25605 2839
rect 25605 2805 25639 2839
rect 25639 2805 25648 2839
rect 25596 2796 25648 2805
rect 26056 2796 26108 2848
rect 26792 2796 26844 2848
rect 30472 2796 30524 2848
rect 33140 2796 33192 2848
rect 38568 2796 38620 2848
rect 19606 2694 19658 2746
rect 19670 2694 19722 2746
rect 19734 2694 19786 2746
rect 19798 2694 19850 2746
rect 1676 2524 1728 2576
rect 5632 2592 5684 2644
rect 7104 2635 7156 2644
rect 7104 2601 7113 2635
rect 7113 2601 7147 2635
rect 7147 2601 7156 2635
rect 7104 2592 7156 2601
rect 7564 2635 7616 2644
rect 7564 2601 7573 2635
rect 7573 2601 7607 2635
rect 7607 2601 7616 2635
rect 7564 2592 7616 2601
rect 7656 2592 7708 2644
rect 11152 2635 11204 2644
rect 11152 2601 11161 2635
rect 11161 2601 11195 2635
rect 11195 2601 11204 2635
rect 11152 2592 11204 2601
rect 12532 2592 12584 2644
rect 15108 2592 15160 2644
rect 17316 2592 17368 2644
rect 17868 2592 17920 2644
rect 18052 2635 18104 2644
rect 18052 2601 18061 2635
rect 18061 2601 18095 2635
rect 18095 2601 18104 2635
rect 18052 2592 18104 2601
rect 20076 2592 20128 2644
rect 21180 2592 21232 2644
rect 22836 2635 22888 2644
rect 22836 2601 22845 2635
rect 22845 2601 22879 2635
rect 22879 2601 22888 2635
rect 22836 2592 22888 2601
rect 23480 2635 23532 2644
rect 23480 2601 23489 2635
rect 23489 2601 23523 2635
rect 23523 2601 23532 2635
rect 23480 2592 23532 2601
rect 23664 2592 23716 2644
rect 25688 2635 25740 2644
rect 25688 2601 25697 2635
rect 25697 2601 25731 2635
rect 25731 2601 25740 2635
rect 25688 2592 25740 2601
rect 26332 2592 26384 2644
rect 5080 2524 5132 2576
rect 1492 2499 1544 2508
rect 1492 2465 1501 2499
rect 1501 2465 1535 2499
rect 1535 2465 1544 2499
rect 1492 2456 1544 2465
rect 2596 2456 2648 2508
rect 5356 2456 5408 2508
rect 8760 2524 8812 2576
rect 12716 2524 12768 2576
rect 8484 2456 8536 2508
rect 9588 2456 9640 2508
rect 11428 2456 11480 2508
rect 9772 2431 9824 2440
rect 9772 2397 9781 2431
rect 9781 2397 9815 2431
rect 9815 2397 9824 2431
rect 9772 2388 9824 2397
rect 8208 2320 8260 2372
rect 7748 2252 7800 2304
rect 8760 2252 8812 2304
rect 16488 2524 16540 2576
rect 20720 2524 20772 2576
rect 29368 2592 29420 2644
rect 16396 2456 16448 2508
rect 18052 2456 18104 2508
rect 24768 2524 24820 2576
rect 27252 2567 27304 2576
rect 27252 2533 27261 2567
rect 27261 2533 27295 2567
rect 27295 2533 27304 2567
rect 27252 2524 27304 2533
rect 27620 2524 27672 2576
rect 23664 2456 23716 2508
rect 27712 2456 27764 2508
rect 28448 2499 28500 2508
rect 28448 2465 28457 2499
rect 28457 2465 28491 2499
rect 28491 2465 28500 2499
rect 28448 2456 28500 2465
rect 30380 2592 30432 2644
rect 31760 2635 31812 2644
rect 31760 2601 31769 2635
rect 31769 2601 31803 2635
rect 31803 2601 31812 2635
rect 31760 2592 31812 2601
rect 32680 2592 32732 2644
rect 34244 2635 34296 2644
rect 34244 2601 34253 2635
rect 34253 2601 34287 2635
rect 34287 2601 34296 2635
rect 34244 2592 34296 2601
rect 35256 2592 35308 2644
rect 37280 2592 37332 2644
rect 40040 2592 40092 2644
rect 40408 2592 40460 2644
rect 29552 2524 29604 2576
rect 33140 2567 33192 2576
rect 33140 2533 33174 2567
rect 33174 2533 33192 2567
rect 33140 2524 33192 2533
rect 38568 2567 38620 2576
rect 38568 2533 38580 2567
rect 38580 2533 38620 2567
rect 38568 2524 38620 2533
rect 34520 2456 34572 2508
rect 36636 2499 36688 2508
rect 36636 2465 36645 2499
rect 36645 2465 36679 2499
rect 36679 2465 36688 2499
rect 36636 2456 36688 2465
rect 37096 2456 37148 2508
rect 42340 2524 42392 2576
rect 41420 2456 41472 2508
rect 42432 2456 42484 2508
rect 42708 2499 42760 2508
rect 42708 2465 42717 2499
rect 42717 2465 42751 2499
rect 42751 2465 42760 2499
rect 42708 2456 42760 2465
rect 45192 2456 45244 2508
rect 26976 2363 27028 2372
rect 26976 2329 26985 2363
rect 26985 2329 27019 2363
rect 27019 2329 27028 2363
rect 26976 2320 27028 2329
rect 27620 2320 27672 2372
rect 38200 2320 38252 2372
rect 40224 2320 40276 2372
rect 43812 2320 43864 2372
rect 46480 2320 46532 2372
rect 15476 2252 15528 2304
rect 35716 2252 35768 2304
rect 45192 2252 45244 2304
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 34966 2150 35018 2202
rect 35030 2150 35082 2202
rect 35094 2150 35146 2202
rect 35158 2150 35210 2202
rect 4712 552 4764 604
rect 4988 552 5040 604
<< metal2 >>
rect 8298 49520 8354 50000
rect 24950 49520 25006 50000
rect 41602 49520 41658 50000
rect 4220 46812 4516 46832
rect 4276 46810 4300 46812
rect 4356 46810 4380 46812
rect 4436 46810 4460 46812
rect 4298 46758 4300 46810
rect 4362 46758 4374 46810
rect 4436 46758 4438 46810
rect 4276 46756 4300 46758
rect 4356 46756 4380 46758
rect 4436 46756 4460 46758
rect 4220 46736 4516 46756
rect 4220 45724 4516 45744
rect 4276 45722 4300 45724
rect 4356 45722 4380 45724
rect 4436 45722 4460 45724
rect 4298 45670 4300 45722
rect 4362 45670 4374 45722
rect 4436 45670 4438 45722
rect 4276 45668 4300 45670
rect 4356 45668 4380 45670
rect 4436 45668 4460 45670
rect 4220 45648 4516 45668
rect 4220 44636 4516 44656
rect 4276 44634 4300 44636
rect 4356 44634 4380 44636
rect 4436 44634 4460 44636
rect 4298 44582 4300 44634
rect 4362 44582 4374 44634
rect 4436 44582 4438 44634
rect 4276 44580 4300 44582
rect 4356 44580 4380 44582
rect 4436 44580 4460 44582
rect 4220 44560 4516 44580
rect 4220 43548 4516 43568
rect 4276 43546 4300 43548
rect 4356 43546 4380 43548
rect 4436 43546 4460 43548
rect 4298 43494 4300 43546
rect 4362 43494 4374 43546
rect 4436 43494 4438 43546
rect 4276 43492 4300 43494
rect 4356 43492 4380 43494
rect 4436 43492 4460 43494
rect 4220 43472 4516 43492
rect 4220 42460 4516 42480
rect 4276 42458 4300 42460
rect 4356 42458 4380 42460
rect 4436 42458 4460 42460
rect 4298 42406 4300 42458
rect 4362 42406 4374 42458
rect 4436 42406 4438 42458
rect 4276 42404 4300 42406
rect 4356 42404 4380 42406
rect 4436 42404 4460 42406
rect 4220 42384 4516 42404
rect 4220 41372 4516 41392
rect 4276 41370 4300 41372
rect 4356 41370 4380 41372
rect 4436 41370 4460 41372
rect 4298 41318 4300 41370
rect 4362 41318 4374 41370
rect 4436 41318 4438 41370
rect 4276 41316 4300 41318
rect 4356 41316 4380 41318
rect 4436 41316 4460 41318
rect 4220 41296 4516 41316
rect 4220 40284 4516 40304
rect 4276 40282 4300 40284
rect 4356 40282 4380 40284
rect 4436 40282 4460 40284
rect 4298 40230 4300 40282
rect 4362 40230 4374 40282
rect 4436 40230 4438 40282
rect 4276 40228 4300 40230
rect 4356 40228 4380 40230
rect 4436 40228 4460 40230
rect 4220 40208 4516 40228
rect 4220 39196 4516 39216
rect 4276 39194 4300 39196
rect 4356 39194 4380 39196
rect 4436 39194 4460 39196
rect 4298 39142 4300 39194
rect 4362 39142 4374 39194
rect 4436 39142 4438 39194
rect 4276 39140 4300 39142
rect 4356 39140 4380 39142
rect 4436 39140 4460 39142
rect 4220 39120 4516 39140
rect 4220 38108 4516 38128
rect 4276 38106 4300 38108
rect 4356 38106 4380 38108
rect 4436 38106 4460 38108
rect 4298 38054 4300 38106
rect 4362 38054 4374 38106
rect 4436 38054 4438 38106
rect 4276 38052 4300 38054
rect 4356 38052 4380 38054
rect 4436 38052 4460 38054
rect 4220 38032 4516 38052
rect 3422 37632 3478 37641
rect 3422 37567 3478 37576
rect 3436 17105 3464 37567
rect 4220 37020 4516 37040
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4298 36966 4300 37018
rect 4362 36966 4374 37018
rect 4436 36966 4438 37018
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4220 36944 4516 36964
rect 4220 35932 4516 35952
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4298 35878 4300 35930
rect 4362 35878 4374 35930
rect 4436 35878 4438 35930
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4220 35856 4516 35876
rect 4220 34844 4516 34864
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4298 34790 4300 34842
rect 4362 34790 4374 34842
rect 4436 34790 4438 34842
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 4220 34768 4516 34788
rect 4220 33756 4516 33776
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4298 33702 4300 33754
rect 4362 33702 4374 33754
rect 4436 33702 4438 33754
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 4220 33680 4516 33700
rect 4220 32668 4516 32688
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4298 32614 4300 32666
rect 4362 32614 4374 32666
rect 4436 32614 4438 32666
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4220 32592 4516 32612
rect 4220 31580 4516 31600
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4298 31526 4300 31578
rect 4362 31526 4374 31578
rect 4436 31526 4438 31578
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4220 31504 4516 31524
rect 4220 30492 4516 30512
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4298 30438 4300 30490
rect 4362 30438 4374 30490
rect 4436 30438 4438 30490
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4220 30416 4516 30436
rect 4220 29404 4516 29424
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4298 29350 4300 29402
rect 4362 29350 4374 29402
rect 4436 29350 4438 29402
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4220 29328 4516 29348
rect 4220 28316 4516 28336
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4298 28262 4300 28314
rect 4362 28262 4374 28314
rect 4436 28262 4438 28314
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4220 28240 4516 28260
rect 4220 27228 4516 27248
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4298 27174 4300 27226
rect 4362 27174 4374 27226
rect 4436 27174 4438 27226
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4220 27152 4516 27172
rect 4220 26140 4516 26160
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4298 26086 4300 26138
rect 4362 26086 4374 26138
rect 4436 26086 4438 26138
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4220 26064 4516 26084
rect 4220 25052 4516 25072
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4220 23888 4516 23908
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4220 22800 4516 22820
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 8312 21457 8340 49520
rect 19580 47356 19876 47376
rect 19636 47354 19660 47356
rect 19716 47354 19740 47356
rect 19796 47354 19820 47356
rect 19658 47302 19660 47354
rect 19722 47302 19734 47354
rect 19796 47302 19798 47354
rect 19636 47300 19660 47302
rect 19716 47300 19740 47302
rect 19796 47300 19820 47302
rect 19580 47280 19876 47300
rect 19580 46268 19876 46288
rect 19636 46266 19660 46268
rect 19716 46266 19740 46268
rect 19796 46266 19820 46268
rect 19658 46214 19660 46266
rect 19722 46214 19734 46266
rect 19796 46214 19798 46266
rect 19636 46212 19660 46214
rect 19716 46212 19740 46214
rect 19796 46212 19820 46214
rect 19580 46192 19876 46212
rect 24964 45665 24992 49520
rect 41616 49450 41644 49520
rect 41616 49422 42104 49450
rect 34940 46812 35236 46832
rect 34996 46810 35020 46812
rect 35076 46810 35100 46812
rect 35156 46810 35180 46812
rect 35018 46758 35020 46810
rect 35082 46758 35094 46810
rect 35156 46758 35158 46810
rect 34996 46756 35020 46758
rect 35076 46756 35100 46758
rect 35156 46756 35180 46758
rect 34940 46736 35236 46756
rect 34940 45724 35236 45744
rect 34996 45722 35020 45724
rect 35076 45722 35100 45724
rect 35156 45722 35180 45724
rect 35018 45670 35020 45722
rect 35082 45670 35094 45722
rect 35156 45670 35158 45722
rect 34996 45668 35020 45670
rect 35076 45668 35100 45670
rect 35156 45668 35180 45670
rect 24950 45656 25006 45665
rect 24950 45591 25006 45600
rect 28078 45656 28134 45665
rect 34940 45648 35236 45668
rect 28078 45591 28134 45600
rect 19580 45180 19876 45200
rect 19636 45178 19660 45180
rect 19716 45178 19740 45180
rect 19796 45178 19820 45180
rect 19658 45126 19660 45178
rect 19722 45126 19734 45178
rect 19796 45126 19798 45178
rect 19636 45124 19660 45126
rect 19716 45124 19740 45126
rect 19796 45124 19820 45126
rect 19580 45104 19876 45124
rect 19580 44092 19876 44112
rect 19636 44090 19660 44092
rect 19716 44090 19740 44092
rect 19796 44090 19820 44092
rect 19658 44038 19660 44090
rect 19722 44038 19734 44090
rect 19796 44038 19798 44090
rect 19636 44036 19660 44038
rect 19716 44036 19740 44038
rect 19796 44036 19820 44038
rect 19580 44016 19876 44036
rect 19580 43004 19876 43024
rect 19636 43002 19660 43004
rect 19716 43002 19740 43004
rect 19796 43002 19820 43004
rect 19658 42950 19660 43002
rect 19722 42950 19734 43002
rect 19796 42950 19798 43002
rect 19636 42948 19660 42950
rect 19716 42948 19740 42950
rect 19796 42948 19820 42950
rect 19580 42928 19876 42948
rect 19580 41916 19876 41936
rect 19636 41914 19660 41916
rect 19716 41914 19740 41916
rect 19796 41914 19820 41916
rect 19658 41862 19660 41914
rect 19722 41862 19734 41914
rect 19796 41862 19798 41914
rect 19636 41860 19660 41862
rect 19716 41860 19740 41862
rect 19796 41860 19820 41862
rect 19580 41840 19876 41860
rect 19580 40828 19876 40848
rect 19636 40826 19660 40828
rect 19716 40826 19740 40828
rect 19796 40826 19820 40828
rect 19658 40774 19660 40826
rect 19722 40774 19734 40826
rect 19796 40774 19798 40826
rect 19636 40772 19660 40774
rect 19716 40772 19740 40774
rect 19796 40772 19820 40774
rect 19580 40752 19876 40772
rect 19580 39740 19876 39760
rect 19636 39738 19660 39740
rect 19716 39738 19740 39740
rect 19796 39738 19820 39740
rect 19658 39686 19660 39738
rect 19722 39686 19734 39738
rect 19796 39686 19798 39738
rect 19636 39684 19660 39686
rect 19716 39684 19740 39686
rect 19796 39684 19820 39686
rect 19580 39664 19876 39684
rect 19580 38652 19876 38672
rect 19636 38650 19660 38652
rect 19716 38650 19740 38652
rect 19796 38650 19820 38652
rect 19658 38598 19660 38650
rect 19722 38598 19734 38650
rect 19796 38598 19798 38650
rect 19636 38596 19660 38598
rect 19716 38596 19740 38598
rect 19796 38596 19820 38598
rect 19580 38576 19876 38596
rect 19580 37564 19876 37584
rect 19636 37562 19660 37564
rect 19716 37562 19740 37564
rect 19796 37562 19820 37564
rect 19658 37510 19660 37562
rect 19722 37510 19734 37562
rect 19796 37510 19798 37562
rect 19636 37508 19660 37510
rect 19716 37508 19740 37510
rect 19796 37508 19820 37510
rect 19580 37488 19876 37508
rect 19580 36476 19876 36496
rect 19636 36474 19660 36476
rect 19716 36474 19740 36476
rect 19796 36474 19820 36476
rect 19658 36422 19660 36474
rect 19722 36422 19734 36474
rect 19796 36422 19798 36474
rect 19636 36420 19660 36422
rect 19716 36420 19740 36422
rect 19796 36420 19820 36422
rect 19580 36400 19876 36420
rect 19580 35388 19876 35408
rect 19636 35386 19660 35388
rect 19716 35386 19740 35388
rect 19796 35386 19820 35388
rect 19658 35334 19660 35386
rect 19722 35334 19734 35386
rect 19796 35334 19798 35386
rect 19636 35332 19660 35334
rect 19716 35332 19740 35334
rect 19796 35332 19820 35334
rect 19580 35312 19876 35332
rect 19580 34300 19876 34320
rect 19636 34298 19660 34300
rect 19716 34298 19740 34300
rect 19796 34298 19820 34300
rect 19658 34246 19660 34298
rect 19722 34246 19734 34298
rect 19796 34246 19798 34298
rect 19636 34244 19660 34246
rect 19716 34244 19740 34246
rect 19796 34244 19820 34246
rect 19580 34224 19876 34244
rect 19580 33212 19876 33232
rect 19636 33210 19660 33212
rect 19716 33210 19740 33212
rect 19796 33210 19820 33212
rect 19658 33158 19660 33210
rect 19722 33158 19734 33210
rect 19796 33158 19798 33210
rect 19636 33156 19660 33158
rect 19716 33156 19740 33158
rect 19796 33156 19820 33158
rect 19580 33136 19876 33156
rect 19580 32124 19876 32144
rect 19636 32122 19660 32124
rect 19716 32122 19740 32124
rect 19796 32122 19820 32124
rect 19658 32070 19660 32122
rect 19722 32070 19734 32122
rect 19796 32070 19798 32122
rect 19636 32068 19660 32070
rect 19716 32068 19740 32070
rect 19796 32068 19820 32070
rect 19580 32048 19876 32068
rect 19580 31036 19876 31056
rect 19636 31034 19660 31036
rect 19716 31034 19740 31036
rect 19796 31034 19820 31036
rect 19658 30982 19660 31034
rect 19722 30982 19734 31034
rect 19796 30982 19798 31034
rect 19636 30980 19660 30982
rect 19716 30980 19740 30982
rect 19796 30980 19820 30982
rect 19580 30960 19876 30980
rect 19580 29948 19876 29968
rect 19636 29946 19660 29948
rect 19716 29946 19740 29948
rect 19796 29946 19820 29948
rect 19658 29894 19660 29946
rect 19722 29894 19734 29946
rect 19796 29894 19798 29946
rect 19636 29892 19660 29894
rect 19716 29892 19740 29894
rect 19796 29892 19820 29894
rect 19580 29872 19876 29892
rect 19580 28860 19876 28880
rect 19636 28858 19660 28860
rect 19716 28858 19740 28860
rect 19796 28858 19820 28860
rect 19658 28806 19660 28858
rect 19722 28806 19734 28858
rect 19796 28806 19798 28858
rect 19636 28804 19660 28806
rect 19716 28804 19740 28806
rect 19796 28804 19820 28806
rect 19580 28784 19876 28804
rect 19580 27772 19876 27792
rect 19636 27770 19660 27772
rect 19716 27770 19740 27772
rect 19796 27770 19820 27772
rect 19658 27718 19660 27770
rect 19722 27718 19734 27770
rect 19796 27718 19798 27770
rect 19636 27716 19660 27718
rect 19716 27716 19740 27718
rect 19796 27716 19820 27718
rect 19580 27696 19876 27716
rect 19580 26684 19876 26704
rect 19636 26682 19660 26684
rect 19716 26682 19740 26684
rect 19796 26682 19820 26684
rect 19658 26630 19660 26682
rect 19722 26630 19734 26682
rect 19796 26630 19798 26682
rect 19636 26628 19660 26630
rect 19716 26628 19740 26630
rect 19796 26628 19820 26630
rect 19580 26608 19876 26628
rect 19580 25596 19876 25616
rect 19636 25594 19660 25596
rect 19716 25594 19740 25596
rect 19796 25594 19820 25596
rect 19658 25542 19660 25594
rect 19722 25542 19734 25594
rect 19796 25542 19798 25594
rect 19636 25540 19660 25542
rect 19716 25540 19740 25542
rect 19796 25540 19820 25542
rect 19580 25520 19876 25540
rect 19580 24508 19876 24528
rect 19636 24506 19660 24508
rect 19716 24506 19740 24508
rect 19796 24506 19820 24508
rect 19658 24454 19660 24506
rect 19722 24454 19734 24506
rect 19796 24454 19798 24506
rect 19636 24452 19660 24454
rect 19716 24452 19740 24454
rect 19796 24452 19820 24454
rect 19580 24432 19876 24452
rect 19580 23420 19876 23440
rect 19636 23418 19660 23420
rect 19716 23418 19740 23420
rect 19796 23418 19820 23420
rect 19658 23366 19660 23418
rect 19722 23366 19734 23418
rect 19796 23366 19798 23418
rect 19636 23364 19660 23366
rect 19716 23364 19740 23366
rect 19796 23364 19820 23366
rect 19580 23344 19876 23364
rect 19580 22332 19876 22352
rect 19636 22330 19660 22332
rect 19716 22330 19740 22332
rect 19796 22330 19820 22332
rect 19658 22278 19660 22330
rect 19722 22278 19734 22330
rect 19796 22278 19798 22330
rect 19636 22276 19660 22278
rect 19716 22276 19740 22278
rect 19796 22276 19820 22278
rect 19580 22256 19876 22276
rect 27988 22024 28040 22030
rect 27988 21966 28040 21972
rect 27896 21616 27948 21622
rect 27896 21558 27948 21564
rect 8298 21448 8354 21457
rect 8298 21383 8354 21392
rect 19580 21244 19876 21264
rect 19636 21242 19660 21244
rect 19716 21242 19740 21244
rect 19796 21242 19820 21244
rect 19658 21190 19660 21242
rect 19722 21190 19734 21242
rect 19796 21190 19798 21242
rect 19636 21188 19660 21190
rect 19716 21188 19740 21190
rect 19796 21188 19820 21190
rect 19580 21168 19876 21188
rect 27908 20942 27936 21558
rect 28000 21486 28028 21966
rect 27988 21480 28040 21486
rect 27988 21422 28040 21428
rect 28092 21010 28120 45591
rect 34940 44636 35236 44656
rect 34996 44634 35020 44636
rect 35076 44634 35100 44636
rect 35156 44634 35180 44636
rect 35018 44582 35020 44634
rect 35082 44582 35094 44634
rect 35156 44582 35158 44634
rect 34996 44580 35020 44582
rect 35076 44580 35100 44582
rect 35156 44580 35180 44582
rect 34940 44560 35236 44580
rect 34940 43548 35236 43568
rect 34996 43546 35020 43548
rect 35076 43546 35100 43548
rect 35156 43546 35180 43548
rect 35018 43494 35020 43546
rect 35082 43494 35094 43546
rect 35156 43494 35158 43546
rect 34996 43492 35020 43494
rect 35076 43492 35100 43494
rect 35156 43492 35180 43494
rect 34940 43472 35236 43492
rect 34940 42460 35236 42480
rect 34996 42458 35020 42460
rect 35076 42458 35100 42460
rect 35156 42458 35180 42460
rect 35018 42406 35020 42458
rect 35082 42406 35094 42458
rect 35156 42406 35158 42458
rect 34996 42404 35020 42406
rect 35076 42404 35100 42406
rect 35156 42404 35180 42406
rect 34940 42384 35236 42404
rect 34940 41372 35236 41392
rect 34996 41370 35020 41372
rect 35076 41370 35100 41372
rect 35156 41370 35180 41372
rect 35018 41318 35020 41370
rect 35082 41318 35094 41370
rect 35156 41318 35158 41370
rect 34996 41316 35020 41318
rect 35076 41316 35100 41318
rect 35156 41316 35180 41318
rect 34940 41296 35236 41316
rect 42076 41290 42104 49422
rect 46938 49192 46994 49201
rect 46938 49127 46994 49136
rect 46754 47696 46810 47705
rect 46754 47631 46810 47640
rect 46768 45422 46796 47631
rect 46846 46064 46902 46073
rect 46846 45999 46902 46008
rect 46756 45416 46808 45422
rect 46756 45358 46808 45364
rect 46768 44962 46796 45358
rect 46860 45098 46888 45999
rect 46952 45558 46980 49127
rect 46940 45552 46992 45558
rect 46940 45494 46992 45500
rect 46860 45070 46980 45098
rect 46676 44934 46796 44962
rect 46112 44328 46164 44334
rect 46112 44270 46164 44276
rect 42076 41262 42196 41290
rect 34940 40284 35236 40304
rect 34996 40282 35020 40284
rect 35076 40282 35100 40284
rect 35156 40282 35180 40284
rect 35018 40230 35020 40282
rect 35082 40230 35094 40282
rect 35156 40230 35158 40282
rect 34996 40228 35020 40230
rect 35076 40228 35100 40230
rect 35156 40228 35180 40230
rect 34940 40208 35236 40228
rect 34940 39196 35236 39216
rect 34996 39194 35020 39196
rect 35076 39194 35100 39196
rect 35156 39194 35180 39196
rect 35018 39142 35020 39194
rect 35082 39142 35094 39194
rect 35156 39142 35158 39194
rect 34996 39140 35020 39142
rect 35076 39140 35100 39142
rect 35156 39140 35180 39142
rect 34940 39120 35236 39140
rect 34940 38108 35236 38128
rect 34996 38106 35020 38108
rect 35076 38106 35100 38108
rect 35156 38106 35180 38108
rect 35018 38054 35020 38106
rect 35082 38054 35094 38106
rect 35156 38054 35158 38106
rect 34996 38052 35020 38054
rect 35076 38052 35100 38054
rect 35156 38052 35180 38054
rect 34940 38032 35236 38052
rect 34940 37020 35236 37040
rect 34996 37018 35020 37020
rect 35076 37018 35100 37020
rect 35156 37018 35180 37020
rect 35018 36966 35020 37018
rect 35082 36966 35094 37018
rect 35156 36966 35158 37018
rect 34996 36964 35020 36966
rect 35076 36964 35100 36966
rect 35156 36964 35180 36966
rect 34940 36944 35236 36964
rect 34940 35932 35236 35952
rect 34996 35930 35020 35932
rect 35076 35930 35100 35932
rect 35156 35930 35180 35932
rect 35018 35878 35020 35930
rect 35082 35878 35094 35930
rect 35156 35878 35158 35930
rect 34996 35876 35020 35878
rect 35076 35876 35100 35878
rect 35156 35876 35180 35878
rect 34940 35856 35236 35876
rect 34940 34844 35236 34864
rect 34996 34842 35020 34844
rect 35076 34842 35100 34844
rect 35156 34842 35180 34844
rect 35018 34790 35020 34842
rect 35082 34790 35094 34842
rect 35156 34790 35158 34842
rect 34996 34788 35020 34790
rect 35076 34788 35100 34790
rect 35156 34788 35180 34790
rect 34940 34768 35236 34788
rect 34940 33756 35236 33776
rect 34996 33754 35020 33756
rect 35076 33754 35100 33756
rect 35156 33754 35180 33756
rect 35018 33702 35020 33754
rect 35082 33702 35094 33754
rect 35156 33702 35158 33754
rect 34996 33700 35020 33702
rect 35076 33700 35100 33702
rect 35156 33700 35180 33702
rect 34940 33680 35236 33700
rect 34940 32668 35236 32688
rect 34996 32666 35020 32668
rect 35076 32666 35100 32668
rect 35156 32666 35180 32668
rect 35018 32614 35020 32666
rect 35082 32614 35094 32666
rect 35156 32614 35158 32666
rect 34996 32612 35020 32614
rect 35076 32612 35100 32614
rect 35156 32612 35180 32614
rect 34940 32592 35236 32612
rect 34940 31580 35236 31600
rect 34996 31578 35020 31580
rect 35076 31578 35100 31580
rect 35156 31578 35180 31580
rect 35018 31526 35020 31578
rect 35082 31526 35094 31578
rect 35156 31526 35158 31578
rect 34996 31524 35020 31526
rect 35076 31524 35100 31526
rect 35156 31524 35180 31526
rect 34940 31504 35236 31524
rect 42064 30864 42116 30870
rect 42064 30806 42116 30812
rect 41880 30796 41932 30802
rect 41880 30738 41932 30744
rect 41788 30592 41840 30598
rect 41788 30534 41840 30540
rect 34940 30492 35236 30512
rect 34996 30490 35020 30492
rect 35076 30490 35100 30492
rect 35156 30490 35180 30492
rect 35018 30438 35020 30490
rect 35082 30438 35094 30490
rect 35156 30438 35158 30490
rect 34996 30436 35020 30438
rect 35076 30436 35100 30438
rect 35156 30436 35180 30438
rect 34940 30416 35236 30436
rect 41696 30252 41748 30258
rect 41696 30194 41748 30200
rect 41420 30048 41472 30054
rect 41420 29990 41472 29996
rect 39580 29776 39632 29782
rect 39580 29718 39632 29724
rect 39028 29640 39080 29646
rect 39028 29582 39080 29588
rect 34940 29404 35236 29424
rect 34996 29402 35020 29404
rect 35076 29402 35100 29404
rect 35156 29402 35180 29404
rect 35018 29350 35020 29402
rect 35082 29350 35094 29402
rect 35156 29350 35158 29402
rect 34996 29348 35020 29350
rect 35076 29348 35100 29350
rect 35156 29348 35180 29350
rect 34940 29328 35236 29348
rect 39040 28966 39068 29582
rect 39592 29345 39620 29718
rect 41432 29646 41460 29990
rect 41420 29640 41472 29646
rect 41420 29582 41472 29588
rect 40224 29504 40276 29510
rect 40224 29446 40276 29452
rect 39578 29336 39634 29345
rect 39578 29271 39580 29280
rect 39632 29271 39634 29280
rect 39580 29242 39632 29248
rect 40236 29102 40264 29446
rect 41328 29232 41380 29238
rect 41156 29170 41276 29186
rect 41328 29174 41380 29180
rect 41156 29164 41288 29170
rect 41156 29158 41236 29164
rect 40224 29096 40276 29102
rect 40224 29038 40276 29044
rect 39396 29028 39448 29034
rect 39396 28970 39448 28976
rect 39028 28960 39080 28966
rect 39028 28902 39080 28908
rect 39212 28960 39264 28966
rect 39212 28902 39264 28908
rect 39040 28626 39068 28902
rect 39224 28626 39252 28902
rect 39028 28620 39080 28626
rect 39028 28562 39080 28568
rect 39212 28620 39264 28626
rect 39212 28562 39264 28568
rect 39040 28506 39068 28562
rect 39040 28478 39160 28506
rect 34940 28316 35236 28336
rect 34996 28314 35020 28316
rect 35076 28314 35100 28316
rect 35156 28314 35180 28316
rect 35018 28262 35020 28314
rect 35082 28262 35094 28314
rect 35156 28262 35158 28314
rect 34996 28260 35020 28262
rect 35076 28260 35100 28262
rect 35156 28260 35180 28262
rect 34940 28240 35236 28260
rect 39132 28014 39160 28478
rect 39224 28218 39252 28562
rect 39212 28212 39264 28218
rect 39212 28154 39264 28160
rect 39120 28008 39172 28014
rect 39120 27950 39172 27956
rect 39132 27878 39160 27950
rect 39120 27872 39172 27878
rect 39120 27814 39172 27820
rect 39132 27470 39160 27814
rect 39408 27606 39436 28970
rect 40236 28966 40264 29038
rect 40316 29028 40368 29034
rect 40316 28970 40368 28976
rect 40224 28960 40276 28966
rect 40224 28902 40276 28908
rect 40328 28762 40356 28970
rect 40316 28756 40368 28762
rect 40316 28698 40368 28704
rect 40316 28484 40368 28490
rect 40316 28426 40368 28432
rect 39948 27872 40000 27878
rect 39948 27814 40000 27820
rect 39960 27674 39988 27814
rect 39948 27668 40000 27674
rect 39948 27610 40000 27616
rect 39396 27600 39448 27606
rect 39396 27542 39448 27548
rect 38108 27464 38160 27470
rect 38108 27406 38160 27412
rect 39120 27464 39172 27470
rect 39120 27406 39172 27412
rect 34940 27228 35236 27248
rect 34996 27226 35020 27228
rect 35076 27226 35100 27228
rect 35156 27226 35180 27228
rect 35018 27174 35020 27226
rect 35082 27174 35094 27226
rect 35156 27174 35158 27226
rect 34996 27172 35020 27174
rect 35076 27172 35100 27174
rect 35156 27172 35180 27174
rect 34940 27152 35236 27172
rect 38120 27130 38148 27406
rect 38292 27328 38344 27334
rect 38292 27270 38344 27276
rect 38108 27124 38160 27130
rect 38108 27066 38160 27072
rect 35900 26852 35952 26858
rect 35900 26794 35952 26800
rect 35912 26586 35940 26794
rect 38304 26790 38332 27270
rect 38382 27160 38438 27169
rect 38382 27095 38384 27104
rect 38436 27095 38438 27104
rect 38384 27066 38436 27072
rect 39132 26926 39160 27406
rect 39408 27130 39436 27542
rect 39396 27124 39448 27130
rect 39396 27066 39448 27072
rect 38660 26920 38712 26926
rect 38660 26862 38712 26868
rect 39120 26920 39172 26926
rect 39120 26862 39172 26868
rect 38384 26852 38436 26858
rect 38384 26794 38436 26800
rect 35992 26784 36044 26790
rect 35992 26726 36044 26732
rect 37188 26784 37240 26790
rect 37188 26726 37240 26732
rect 38292 26784 38344 26790
rect 38292 26726 38344 26732
rect 35900 26580 35952 26586
rect 35900 26522 35952 26528
rect 34940 26140 35236 26160
rect 34996 26138 35020 26140
rect 35076 26138 35100 26140
rect 35156 26138 35180 26140
rect 35018 26086 35020 26138
rect 35082 26086 35094 26138
rect 35156 26086 35158 26138
rect 34996 26084 35020 26086
rect 35076 26084 35100 26086
rect 35156 26084 35180 26086
rect 34940 26064 35236 26084
rect 36004 25838 36032 26726
rect 36728 26240 36780 26246
rect 36728 26182 36780 26188
rect 37096 26240 37148 26246
rect 37096 26182 37148 26188
rect 36740 25838 36768 26182
rect 35992 25832 36044 25838
rect 35992 25774 36044 25780
rect 36728 25832 36780 25838
rect 36728 25774 36780 25780
rect 37108 25770 37136 26182
rect 37096 25764 37148 25770
rect 37096 25706 37148 25712
rect 35992 25696 36044 25702
rect 35992 25638 36044 25644
rect 36360 25696 36412 25702
rect 36360 25638 36412 25644
rect 36004 25498 36032 25638
rect 35992 25492 36044 25498
rect 35992 25434 36044 25440
rect 36176 25492 36228 25498
rect 36176 25434 36228 25440
rect 35990 25256 36046 25265
rect 35990 25191 35992 25200
rect 36044 25191 36046 25200
rect 35992 25162 36044 25168
rect 34940 25052 35236 25072
rect 34996 25050 35020 25052
rect 35076 25050 35100 25052
rect 35156 25050 35180 25052
rect 35018 24998 35020 25050
rect 35082 24998 35094 25050
rect 35156 24998 35158 25050
rect 34996 24996 35020 24998
rect 35076 24996 35100 24998
rect 35156 24996 35180 24998
rect 34940 24976 35236 24996
rect 35808 24676 35860 24682
rect 35808 24618 35860 24624
rect 35440 24608 35492 24614
rect 35440 24550 35492 24556
rect 31298 24168 31354 24177
rect 31298 24103 31354 24112
rect 30472 24064 30524 24070
rect 30472 24006 30524 24012
rect 30484 23526 30512 24006
rect 31312 23866 31340 24103
rect 34940 23964 35236 23984
rect 34996 23962 35020 23964
rect 35076 23962 35100 23964
rect 35156 23962 35180 23964
rect 35018 23910 35020 23962
rect 35082 23910 35094 23962
rect 35156 23910 35158 23962
rect 34996 23908 35020 23910
rect 35076 23908 35100 23910
rect 35156 23908 35180 23910
rect 34940 23888 35236 23908
rect 31300 23860 31352 23866
rect 31300 23802 31352 23808
rect 35452 23662 35480 24550
rect 35820 24274 35848 24618
rect 35808 24268 35860 24274
rect 35808 24210 35860 24216
rect 35716 24200 35768 24206
rect 35716 24142 35768 24148
rect 35728 23798 35756 24142
rect 35820 23866 35848 24210
rect 36188 24138 36216 25434
rect 36268 25356 36320 25362
rect 36268 25298 36320 25304
rect 36280 24410 36308 25298
rect 36372 24750 36400 25638
rect 36912 25288 36964 25294
rect 36912 25230 36964 25236
rect 36924 24954 36952 25230
rect 36912 24948 36964 24954
rect 36912 24890 36964 24896
rect 36360 24744 36412 24750
rect 36360 24686 36412 24692
rect 36268 24404 36320 24410
rect 36268 24346 36320 24352
rect 36636 24336 36688 24342
rect 36636 24278 36688 24284
rect 36176 24132 36228 24138
rect 36176 24074 36228 24080
rect 35808 23860 35860 23866
rect 35808 23802 35860 23808
rect 35716 23792 35768 23798
rect 35716 23734 35768 23740
rect 35440 23656 35492 23662
rect 35440 23598 35492 23604
rect 31668 23588 31720 23594
rect 31668 23530 31720 23536
rect 31852 23588 31904 23594
rect 31852 23530 31904 23536
rect 30472 23520 30524 23526
rect 30472 23462 30524 23468
rect 31680 23474 31708 23530
rect 29552 22432 29604 22438
rect 29552 22374 29604 22380
rect 29564 22234 29592 22374
rect 29552 22228 29604 22234
rect 29552 22170 29604 22176
rect 29920 22228 29972 22234
rect 29920 22170 29972 22176
rect 28908 22024 28960 22030
rect 28908 21966 28960 21972
rect 28264 21888 28316 21894
rect 28264 21830 28316 21836
rect 28276 21554 28304 21830
rect 28920 21690 28948 21966
rect 28908 21684 28960 21690
rect 28908 21626 28960 21632
rect 29736 21684 29788 21690
rect 29736 21626 29788 21632
rect 28264 21548 28316 21554
rect 28264 21490 28316 21496
rect 28080 21004 28132 21010
rect 28080 20946 28132 20952
rect 27252 20936 27304 20942
rect 27252 20878 27304 20884
rect 27620 20936 27672 20942
rect 27620 20878 27672 20884
rect 27896 20936 27948 20942
rect 27896 20878 27948 20884
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 27264 20262 27292 20878
rect 27632 20641 27660 20878
rect 27618 20632 27674 20641
rect 27448 20590 27618 20618
rect 27448 20262 27476 20590
rect 27908 20602 27936 20878
rect 27618 20567 27674 20576
rect 27896 20596 27948 20602
rect 27632 20507 27660 20567
rect 27896 20538 27948 20544
rect 28092 20466 28120 20946
rect 28276 20777 28304 21490
rect 29642 21448 29698 21457
rect 29748 21418 29776 21626
rect 29932 21554 29960 22170
rect 30288 22092 30340 22098
rect 30288 22034 30340 22040
rect 30300 22001 30328 22034
rect 30286 21992 30342 22001
rect 30286 21927 30342 21936
rect 29920 21548 29972 21554
rect 29920 21490 29972 21496
rect 29642 21383 29644 21392
rect 29696 21383 29698 21392
rect 29736 21412 29788 21418
rect 29644 21354 29696 21360
rect 29736 21354 29788 21360
rect 28262 20768 28318 20777
rect 28262 20703 28318 20712
rect 28080 20460 28132 20466
rect 28080 20402 28132 20408
rect 29748 20398 29776 21354
rect 29828 21344 29880 21350
rect 29828 21286 29880 21292
rect 29840 20806 29868 21286
rect 29828 20800 29880 20806
rect 29828 20742 29880 20748
rect 29932 20398 29960 21490
rect 30484 20874 30512 23462
rect 31680 23446 31800 23474
rect 31772 23322 31800 23446
rect 31760 23316 31812 23322
rect 31760 23258 31812 23264
rect 31864 23254 31892 23530
rect 35808 23520 35860 23526
rect 35808 23462 35860 23468
rect 31852 23248 31904 23254
rect 31852 23190 31904 23196
rect 33232 23248 33284 23254
rect 33232 23190 33284 23196
rect 31864 22642 31892 23190
rect 31852 22636 31904 22642
rect 31852 22578 31904 22584
rect 32404 22568 32456 22574
rect 32404 22510 32456 22516
rect 32220 22432 32272 22438
rect 32220 22374 32272 22380
rect 32232 22234 32260 22374
rect 31760 22228 31812 22234
rect 31760 22170 31812 22176
rect 32220 22228 32272 22234
rect 32220 22170 32272 22176
rect 31208 21888 31260 21894
rect 31208 21830 31260 21836
rect 31220 21486 31248 21830
rect 31208 21480 31260 21486
rect 31772 21434 31800 22170
rect 32416 22166 32444 22510
rect 33048 22228 33100 22234
rect 33048 22170 33100 22176
rect 32404 22160 32456 22166
rect 32404 22102 32456 22108
rect 32416 21690 32444 22102
rect 33060 22030 33088 22170
rect 33048 22024 33100 22030
rect 33048 21966 33100 21972
rect 33244 21894 33272 23190
rect 34060 23112 34112 23118
rect 33598 23080 33654 23089
rect 34060 23054 34112 23060
rect 34612 23112 34664 23118
rect 34612 23054 34664 23060
rect 33598 23015 33600 23024
rect 33652 23015 33654 23024
rect 33600 22986 33652 22992
rect 34072 22778 34100 23054
rect 34060 22772 34112 22778
rect 34060 22714 34112 22720
rect 34624 22710 34652 23054
rect 34940 22876 35236 22896
rect 34996 22874 35020 22876
rect 35076 22874 35100 22876
rect 35156 22874 35180 22876
rect 35018 22822 35020 22874
rect 35082 22822 35094 22874
rect 35156 22822 35158 22874
rect 34996 22820 35020 22822
rect 35076 22820 35100 22822
rect 35156 22820 35180 22822
rect 34940 22800 35236 22820
rect 34612 22704 34664 22710
rect 34612 22646 34664 22652
rect 33600 22432 33652 22438
rect 33600 22374 33652 22380
rect 33612 22166 33640 22374
rect 34624 22234 34652 22646
rect 35820 22438 35848 23462
rect 36176 22976 36228 22982
rect 36174 22944 36176 22953
rect 36648 22953 36676 24278
rect 36924 23662 36952 24890
rect 37200 24342 37228 26726
rect 38198 25664 38254 25673
rect 38198 25599 38254 25608
rect 37832 25424 37884 25430
rect 37832 25366 37884 25372
rect 37844 24954 37872 25366
rect 38212 25294 38240 25599
rect 38200 25288 38252 25294
rect 38200 25230 38252 25236
rect 38212 24954 38240 25230
rect 38304 25226 38332 26726
rect 38396 26586 38424 26794
rect 38384 26580 38436 26586
rect 38384 26522 38436 26528
rect 38568 26580 38620 26586
rect 38568 26522 38620 26528
rect 38396 26042 38424 26522
rect 38384 26036 38436 26042
rect 38384 25978 38436 25984
rect 38580 25838 38608 26522
rect 38672 26246 38700 26862
rect 38752 26444 38804 26450
rect 38752 26386 38804 26392
rect 38660 26240 38712 26246
rect 38660 26182 38712 26188
rect 38672 26042 38700 26182
rect 38764 26042 38792 26386
rect 38660 26036 38712 26042
rect 38660 25978 38712 25984
rect 38752 26036 38804 26042
rect 38752 25978 38804 25984
rect 38568 25832 38620 25838
rect 38568 25774 38620 25780
rect 38580 25430 38608 25774
rect 38568 25424 38620 25430
rect 38568 25366 38620 25372
rect 38292 25220 38344 25226
rect 38292 25162 38344 25168
rect 37832 24948 37884 24954
rect 37832 24890 37884 24896
rect 38200 24948 38252 24954
rect 38200 24890 38252 24896
rect 37188 24336 37240 24342
rect 37188 24278 37240 24284
rect 37188 24200 37240 24206
rect 37240 24148 37412 24154
rect 37188 24142 37412 24148
rect 37200 24126 37412 24142
rect 36912 23656 36964 23662
rect 36912 23598 36964 23604
rect 36924 23322 36952 23598
rect 37280 23520 37332 23526
rect 37280 23462 37332 23468
rect 36912 23316 36964 23322
rect 36912 23258 36964 23264
rect 36228 22944 36230 22953
rect 36174 22879 36230 22888
rect 36634 22944 36690 22953
rect 36634 22879 36690 22888
rect 35808 22432 35860 22438
rect 35808 22374 35860 22380
rect 34612 22228 34664 22234
rect 34612 22170 34664 22176
rect 33600 22160 33652 22166
rect 33600 22102 33652 22108
rect 33508 22024 33560 22030
rect 33508 21966 33560 21972
rect 33232 21888 33284 21894
rect 33232 21830 33284 21836
rect 32404 21684 32456 21690
rect 32404 21626 32456 21632
rect 31208 21422 31260 21428
rect 31220 21078 31248 21422
rect 31680 21418 31800 21434
rect 31668 21412 31800 21418
rect 31720 21406 31800 21412
rect 31668 21354 31720 21360
rect 30932 21072 30984 21078
rect 30932 21014 30984 21020
rect 31208 21072 31260 21078
rect 31208 21014 31260 21020
rect 30472 20868 30524 20874
rect 30472 20810 30524 20816
rect 30380 20800 30432 20806
rect 30380 20742 30432 20748
rect 29736 20392 29788 20398
rect 29736 20334 29788 20340
rect 29920 20392 29972 20398
rect 29920 20334 29972 20340
rect 27252 20256 27304 20262
rect 27252 20198 27304 20204
rect 27436 20256 27488 20262
rect 27436 20198 27488 20204
rect 19580 20156 19876 20176
rect 19636 20154 19660 20156
rect 19716 20154 19740 20156
rect 19796 20154 19820 20156
rect 19658 20102 19660 20154
rect 19722 20102 19734 20154
rect 19796 20102 19798 20154
rect 19636 20100 19660 20102
rect 19716 20100 19740 20102
rect 19796 20100 19820 20102
rect 19580 20080 19876 20100
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 19580 19068 19876 19088
rect 19636 19066 19660 19068
rect 19716 19066 19740 19068
rect 19796 19066 19820 19068
rect 19658 19014 19660 19066
rect 19722 19014 19734 19066
rect 19796 19014 19798 19066
rect 19636 19012 19660 19014
rect 19716 19012 19740 19014
rect 19796 19012 19820 19014
rect 19580 18992 19876 19012
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4220 18448 4516 18468
rect 19580 17980 19876 18000
rect 19636 17978 19660 17980
rect 19716 17978 19740 17980
rect 19796 17978 19820 17980
rect 19658 17926 19660 17978
rect 19722 17926 19734 17978
rect 19796 17926 19798 17978
rect 19636 17924 19660 17926
rect 19716 17924 19740 17926
rect 19796 17924 19820 17926
rect 19580 17904 19876 17924
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 26516 17264 26568 17270
rect 26516 17206 26568 17212
rect 23756 17128 23808 17134
rect 3422 17096 3478 17105
rect 3422 17031 3478 17040
rect 23478 17096 23534 17105
rect 23756 17070 23808 17076
rect 23478 17031 23480 17040
rect 23532 17031 23534 17040
rect 23480 17002 23532 17008
rect 19580 16892 19876 16912
rect 19636 16890 19660 16892
rect 19716 16890 19740 16892
rect 19796 16890 19820 16892
rect 19658 16838 19660 16890
rect 19722 16838 19734 16890
rect 19796 16838 19798 16890
rect 19636 16836 19660 16838
rect 19716 16836 19740 16838
rect 19796 16836 19820 16838
rect 19580 16816 19876 16836
rect 23768 16658 23796 17070
rect 25780 16992 25832 16998
rect 25780 16934 25832 16940
rect 23756 16652 23808 16658
rect 23756 16594 23808 16600
rect 25320 16584 25372 16590
rect 25320 16526 25372 16532
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 25332 16250 25360 16526
rect 25320 16244 25372 16250
rect 25320 16186 25372 16192
rect 25792 16046 25820 16934
rect 26528 16833 26556 17206
rect 26792 17128 26844 17134
rect 26792 17070 26844 17076
rect 27160 17128 27212 17134
rect 27160 17070 27212 17076
rect 26514 16824 26570 16833
rect 26514 16759 26570 16768
rect 26804 16250 26832 17070
rect 26884 17060 26936 17066
rect 26884 17002 26936 17008
rect 26896 16726 26924 17002
rect 27172 16726 27200 17070
rect 26884 16720 26936 16726
rect 26884 16662 26936 16668
rect 27160 16720 27212 16726
rect 27160 16662 27212 16668
rect 26884 16584 26936 16590
rect 26884 16526 26936 16532
rect 26792 16244 26844 16250
rect 26792 16186 26844 16192
rect 25780 16040 25832 16046
rect 25780 15982 25832 15988
rect 19580 15804 19876 15824
rect 19636 15802 19660 15804
rect 19716 15802 19740 15804
rect 19796 15802 19820 15804
rect 19658 15750 19660 15802
rect 19722 15750 19734 15802
rect 19796 15750 19798 15802
rect 19636 15748 19660 15750
rect 19716 15748 19740 15750
rect 19796 15748 19820 15750
rect 19580 15728 19876 15748
rect 25792 15706 25820 15982
rect 26608 15904 26660 15910
rect 26608 15846 26660 15852
rect 25780 15700 25832 15706
rect 25780 15642 25832 15648
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 19580 14716 19876 14736
rect 19636 14714 19660 14716
rect 19716 14714 19740 14716
rect 19796 14714 19820 14716
rect 19658 14662 19660 14714
rect 19722 14662 19734 14714
rect 19796 14662 19798 14714
rect 19636 14660 19660 14662
rect 19716 14660 19740 14662
rect 19796 14660 19820 14662
rect 19580 14640 19876 14660
rect 20258 14512 20314 14521
rect 26620 14482 26648 15846
rect 26804 15706 26832 16186
rect 26896 15910 26924 16526
rect 26884 15904 26936 15910
rect 26884 15846 26936 15852
rect 26792 15700 26844 15706
rect 26792 15642 26844 15648
rect 20258 14447 20314 14456
rect 26608 14476 26660 14482
rect 8390 14376 8446 14385
rect 8390 14311 8392 14320
rect 8444 14311 8446 14320
rect 8392 14282 8444 14288
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 8404 13870 8432 14282
rect 19800 14272 19852 14278
rect 19800 14214 19852 14220
rect 19340 14000 19392 14006
rect 19340 13942 19392 13948
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 8392 13864 8444 13870
rect 8392 13806 8444 13812
rect 4712 13728 4764 13734
rect 4712 13670 4764 13676
rect 4724 13462 4752 13670
rect 4804 13524 4856 13530
rect 4804 13466 4856 13472
rect 5632 13524 5684 13530
rect 5632 13466 5684 13472
rect 4712 13456 4764 13462
rect 4712 13398 4764 13404
rect 2044 13320 2096 13326
rect 2044 13262 2096 13268
rect 4620 13320 4672 13326
rect 4620 13262 4672 13268
rect 1492 13184 1544 13190
rect 1492 13126 1544 13132
rect 1504 12782 1532 13126
rect 2056 12782 2084 13262
rect 4068 13184 4120 13190
rect 4068 13126 4120 13132
rect 1492 12776 1544 12782
rect 1492 12718 1544 12724
rect 2044 12776 2096 12782
rect 2044 12718 2096 12724
rect 1504 12306 1532 12718
rect 2688 12640 2740 12646
rect 2688 12582 2740 12588
rect 2700 12374 2728 12582
rect 2320 12368 2372 12374
rect 2320 12310 2372 12316
rect 2688 12368 2740 12374
rect 2688 12310 2740 12316
rect 1492 12300 1544 12306
rect 1492 12242 1544 12248
rect 1504 11898 1532 12242
rect 1492 11892 1544 11898
rect 1492 11834 1544 11840
rect 1504 10674 1532 11834
rect 2332 11626 2360 12310
rect 3976 12232 4028 12238
rect 3976 12174 4028 12180
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 2884 11898 2912 12038
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 2780 11824 2832 11830
rect 2780 11766 2832 11772
rect 3424 11824 3476 11830
rect 3424 11766 3476 11772
rect 2412 11756 2464 11762
rect 2412 11698 2464 11704
rect 2320 11620 2372 11626
rect 2320 11562 2372 11568
rect 2332 11286 2360 11562
rect 2424 11354 2452 11698
rect 2792 11626 2820 11766
rect 2688 11620 2740 11626
rect 2688 11562 2740 11568
rect 2780 11620 2832 11626
rect 2780 11562 2832 11568
rect 2700 11354 2728 11562
rect 2792 11354 2820 11562
rect 2412 11348 2464 11354
rect 2412 11290 2464 11296
rect 2688 11348 2740 11354
rect 2688 11290 2740 11296
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2320 11280 2372 11286
rect 2320 11222 2372 11228
rect 1492 10668 1544 10674
rect 1492 10610 1544 10616
rect 1504 10266 1532 10610
rect 2424 10606 2452 11290
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2504 10464 2556 10470
rect 2504 10406 2556 10412
rect 2516 10266 2544 10406
rect 1492 10260 1544 10266
rect 1492 10202 1544 10208
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 1504 9518 1532 10202
rect 2044 10192 2096 10198
rect 2516 10146 2544 10202
rect 2700 10198 2728 11290
rect 3436 11218 3464 11766
rect 3896 11608 3924 12038
rect 3988 11898 4016 12174
rect 3976 11892 4028 11898
rect 3976 11834 4028 11840
rect 3976 11620 4028 11626
rect 3896 11580 3976 11608
rect 3976 11562 4028 11568
rect 3424 11212 3476 11218
rect 3424 11154 3476 11160
rect 2044 10134 2096 10140
rect 1492 9512 1544 9518
rect 1492 9454 1544 9460
rect 1504 9178 1532 9454
rect 1492 9172 1544 9178
rect 1492 9114 1544 9120
rect 1504 8566 1532 9114
rect 2056 9042 2084 10134
rect 2424 10118 2544 10146
rect 2688 10192 2740 10198
rect 2688 10134 2740 10140
rect 2424 9518 2452 10118
rect 2504 10056 2556 10062
rect 2504 9998 2556 10004
rect 2516 9722 2544 9998
rect 2688 9920 2740 9926
rect 2688 9862 2740 9868
rect 2504 9716 2556 9722
rect 2504 9658 2556 9664
rect 2700 9586 2728 9862
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 2424 9178 2452 9454
rect 2792 9178 2820 9590
rect 3988 9382 4016 11562
rect 4080 11558 4108 13126
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 4172 12306 4200 12718
rect 4632 12442 4660 13262
rect 4620 12436 4672 12442
rect 4620 12378 4672 12384
rect 4816 12374 4844 13466
rect 5644 12986 5672 13466
rect 6736 13388 6788 13394
rect 6736 13330 6788 13336
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 6472 12986 6500 13262
rect 5632 12980 5684 12986
rect 5632 12922 5684 12928
rect 6460 12980 6512 12986
rect 6460 12922 6512 12928
rect 6472 12782 6500 12922
rect 6460 12776 6512 12782
rect 6460 12718 6512 12724
rect 5540 12708 5592 12714
rect 5540 12650 5592 12656
rect 5552 12442 5580 12650
rect 6748 12646 6776 13330
rect 7196 13184 7248 13190
rect 7196 13126 7248 13132
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 6920 12912 6972 12918
rect 6920 12854 6972 12860
rect 6828 12844 6880 12850
rect 6828 12786 6880 12792
rect 6736 12640 6788 12646
rect 6736 12582 6788 12588
rect 6840 12442 6868 12786
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 4804 12368 4856 12374
rect 4804 12310 4856 12316
rect 4160 12300 4212 12306
rect 4160 12242 4212 12248
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 4816 11898 4844 12310
rect 6932 12306 6960 12854
rect 7208 12782 7236 13126
rect 7392 12850 7420 13126
rect 7656 12980 7708 12986
rect 7656 12922 7708 12928
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 7012 12776 7064 12782
rect 7010 12744 7012 12753
rect 7196 12776 7248 12782
rect 7064 12744 7066 12753
rect 7196 12718 7248 12724
rect 7010 12679 7066 12688
rect 7104 12368 7156 12374
rect 7104 12310 7156 12316
rect 6920 12300 6972 12306
rect 6920 12242 6972 12248
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 5552 11898 5580 12038
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 5446 11656 5502 11665
rect 5446 11591 5502 11600
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 5460 11354 5488 11591
rect 5816 11552 5868 11558
rect 5816 11494 5868 11500
rect 5828 11354 5856 11494
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 4632 10810 4660 11154
rect 5540 11076 5592 11082
rect 5540 11018 5592 11024
rect 4988 11008 5040 11014
rect 4988 10950 5040 10956
rect 5448 11008 5500 11014
rect 5448 10950 5500 10956
rect 5000 10810 5028 10950
rect 5262 10840 5318 10849
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4988 10804 5040 10810
rect 5262 10775 5264 10784
rect 4988 10746 5040 10752
rect 5316 10775 5318 10784
rect 5264 10746 5316 10752
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 5276 10266 5304 10406
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 5354 10160 5410 10169
rect 4620 10124 4672 10130
rect 5354 10095 5356 10104
rect 4620 10066 4672 10072
rect 5408 10095 5410 10104
rect 5356 10066 5408 10072
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 4632 9654 4660 10066
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4620 9648 4672 9654
rect 4620 9590 4672 9596
rect 4724 9450 4752 9862
rect 5368 9722 5396 10066
rect 5460 9926 5488 10950
rect 5552 10606 5580 11018
rect 5828 10810 5856 11290
rect 5908 11144 5960 11150
rect 5908 11086 5960 11092
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 5540 10600 5592 10606
rect 5540 10542 5592 10548
rect 5552 10266 5580 10542
rect 5920 10538 5948 11086
rect 6472 11082 6500 12174
rect 6932 11898 6960 12242
rect 6920 11892 6972 11898
rect 6920 11834 6972 11840
rect 7116 11830 7144 12310
rect 7104 11824 7156 11830
rect 7104 11766 7156 11772
rect 7208 11626 7236 12718
rect 7668 12646 7696 12922
rect 8312 12782 8340 13806
rect 8300 12776 8352 12782
rect 8298 12744 8300 12753
rect 8352 12744 8354 12753
rect 8298 12679 8354 12688
rect 7656 12640 7708 12646
rect 7656 12582 7708 12588
rect 7668 12442 7696 12582
rect 7656 12436 7708 12442
rect 7656 12378 7708 12384
rect 7656 11756 7708 11762
rect 7656 11698 7708 11704
rect 7196 11620 7248 11626
rect 7196 11562 7248 11568
rect 7668 11354 7696 11698
rect 7840 11620 7892 11626
rect 7840 11562 7892 11568
rect 7656 11348 7708 11354
rect 7656 11290 7708 11296
rect 6460 11076 6512 11082
rect 6460 11018 6512 11024
rect 7472 11076 7524 11082
rect 7472 11018 7524 11024
rect 7196 11008 7248 11014
rect 7196 10950 7248 10956
rect 6920 10736 6972 10742
rect 6920 10678 6972 10684
rect 5908 10532 5960 10538
rect 5908 10474 5960 10480
rect 5920 10266 5948 10474
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5908 10260 5960 10266
rect 5908 10202 5960 10208
rect 5448 9920 5500 9926
rect 5448 9862 5500 9868
rect 5920 9722 5948 10202
rect 6564 9994 6592 10406
rect 6932 10169 6960 10678
rect 7208 10606 7236 10950
rect 7484 10674 7512 11018
rect 7852 11014 7880 11562
rect 8404 11558 8432 13806
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 8772 12782 8800 13670
rect 19352 13462 19380 13942
rect 19812 13818 19840 14214
rect 20272 13938 20300 14447
rect 26608 14418 26660 14424
rect 26884 14476 26936 14482
rect 26884 14418 26936 14424
rect 26620 14074 26648 14418
rect 26896 14074 26924 14418
rect 26608 14068 26660 14074
rect 26608 14010 26660 14016
rect 26884 14068 26936 14074
rect 26884 14010 26936 14016
rect 20260 13932 20312 13938
rect 20260 13874 20312 13880
rect 19812 13802 19932 13818
rect 19800 13796 19932 13802
rect 19852 13790 19932 13796
rect 19800 13738 19852 13744
rect 19580 13628 19876 13648
rect 19636 13626 19660 13628
rect 19716 13626 19740 13628
rect 19796 13626 19820 13628
rect 19658 13574 19660 13626
rect 19722 13574 19734 13626
rect 19796 13574 19798 13626
rect 19636 13572 19660 13574
rect 19716 13572 19740 13574
rect 19796 13572 19820 13574
rect 19580 13552 19876 13572
rect 19340 13456 19392 13462
rect 19340 13398 19392 13404
rect 18880 13320 18932 13326
rect 18880 13262 18932 13268
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 8772 12442 8800 12718
rect 18892 12646 18920 13262
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 8760 12436 8812 12442
rect 8760 12378 8812 12384
rect 8772 11762 8800 12378
rect 9600 12322 9628 12582
rect 18236 12368 18288 12374
rect 9954 12336 10010 12345
rect 9600 12294 9720 12322
rect 9692 12238 9720 12294
rect 18892 12345 18920 12582
rect 19352 12442 19380 13398
rect 19616 13388 19668 13394
rect 19616 13330 19668 13336
rect 19628 12986 19656 13330
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19616 12980 19668 12986
rect 19616 12922 19668 12928
rect 19444 12442 19472 12922
rect 19580 12540 19876 12560
rect 19636 12538 19660 12540
rect 19716 12538 19740 12540
rect 19796 12538 19820 12540
rect 19658 12486 19660 12538
rect 19722 12486 19734 12538
rect 19796 12486 19798 12538
rect 19636 12484 19660 12486
rect 19716 12484 19740 12486
rect 19796 12484 19820 12486
rect 19580 12464 19876 12484
rect 19340 12436 19392 12442
rect 19340 12378 19392 12384
rect 19432 12436 19484 12442
rect 19432 12378 19484 12384
rect 18236 12310 18288 12316
rect 18878 12336 18934 12345
rect 9954 12271 9956 12280
rect 10008 12271 10010 12280
rect 17868 12300 17920 12306
rect 9956 12242 10008 12248
rect 17868 12242 17920 12248
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9692 11762 9720 12174
rect 9968 11898 9996 12242
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 13636 12096 13688 12102
rect 13636 12038 13688 12044
rect 16028 12096 16080 12102
rect 16028 12038 16080 12044
rect 9956 11892 10008 11898
rect 9956 11834 10008 11840
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 7840 11008 7892 11014
rect 7840 10950 7892 10956
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 7104 10192 7156 10198
rect 6918 10160 6974 10169
rect 7104 10134 7156 10140
rect 6918 10095 6974 10104
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 6552 9988 6604 9994
rect 6552 9930 6604 9936
rect 7024 9722 7052 9998
rect 5356 9716 5408 9722
rect 5356 9658 5408 9664
rect 5908 9716 5960 9722
rect 5908 9658 5960 9664
rect 7012 9716 7064 9722
rect 7012 9658 7064 9664
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 4160 9444 4212 9450
rect 4160 9386 4212 9392
rect 4712 9444 4764 9450
rect 4712 9386 4764 9392
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 2780 9172 2832 9178
rect 2780 9114 2832 9120
rect 2044 9036 2096 9042
rect 2044 8978 2096 8984
rect 2056 8634 2084 8978
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 1492 8560 1544 8566
rect 1492 8502 1544 8508
rect 2056 8090 2084 8570
rect 2792 8514 2820 9114
rect 2700 8486 2820 8514
rect 2700 8090 2728 8486
rect 2792 8430 2820 8486
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 1952 7948 2004 7954
rect 1952 7890 2004 7896
rect 1964 7206 1992 7890
rect 1952 7200 2004 7206
rect 1952 7142 2004 7148
rect 1676 3392 1728 3398
rect 1676 3334 1728 3340
rect 662 3088 718 3097
rect 662 3023 718 3032
rect 676 480 704 3023
rect 1492 2848 1544 2854
rect 1492 2790 1544 2796
rect 1504 2514 1532 2790
rect 1688 2582 1716 3334
rect 1676 2576 1728 2582
rect 1676 2518 1728 2524
rect 1492 2508 1544 2514
rect 1492 2450 1544 2456
rect 1964 480 1992 7142
rect 3332 6928 3384 6934
rect 3332 6870 3384 6876
rect 3240 6860 3292 6866
rect 3240 6802 3292 6808
rect 3252 6118 3280 6802
rect 3344 6458 3372 6870
rect 3988 6730 4016 9318
rect 4172 8906 4200 9386
rect 4620 9104 4672 9110
rect 4620 9046 4672 9052
rect 4160 8900 4212 8906
rect 4160 8842 4212 8848
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4220 8656 4516 8676
rect 4632 8634 4660 9046
rect 4804 8900 4856 8906
rect 4804 8842 4856 8848
rect 4816 8634 4844 8842
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 4080 7886 4108 8230
rect 4632 8022 4660 8570
rect 4816 8090 4844 8570
rect 4804 8084 4856 8090
rect 4804 8026 4856 8032
rect 4620 8016 4672 8022
rect 4620 7958 4672 7964
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 4080 7188 4108 7822
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 4632 7546 4660 7958
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 4160 7200 4212 7206
rect 4080 7160 4160 7188
rect 4160 7142 4212 7148
rect 4172 6934 4200 7142
rect 4160 6928 4212 6934
rect 4160 6870 4212 6876
rect 4080 6730 4200 6746
rect 3976 6724 4028 6730
rect 3976 6666 4028 6672
rect 4080 6724 4212 6730
rect 4080 6718 4160 6724
rect 3332 6452 3384 6458
rect 3332 6394 3384 6400
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 3252 4706 3280 6054
rect 3344 5914 3372 6394
rect 3332 5908 3384 5914
rect 3332 5850 3384 5856
rect 3344 5370 3372 5850
rect 3332 5364 3384 5370
rect 3332 5306 3384 5312
rect 4080 5098 4108 6718
rect 4160 6666 4212 6672
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 4620 6180 4672 6186
rect 4620 6122 4672 6128
rect 4632 5914 4660 6122
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 4632 5370 4660 5850
rect 4724 5710 4752 6598
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 3332 5092 3384 5098
rect 3332 5034 3384 5040
rect 4068 5092 4120 5098
rect 4068 5034 4120 5040
rect 3344 4826 3372 5034
rect 4160 5024 4212 5030
rect 4080 4972 4160 4978
rect 4080 4966 4212 4972
rect 4080 4950 4200 4966
rect 3332 4820 3384 4826
rect 3332 4762 3384 4768
rect 3252 4678 3372 4706
rect 2688 4480 2740 4486
rect 2740 4440 2820 4468
rect 2688 4422 2740 4428
rect 2792 4010 2820 4440
rect 2780 4004 2832 4010
rect 2780 3946 2832 3952
rect 2596 3936 2648 3942
rect 2596 3878 2648 3884
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 2332 3194 2360 3674
rect 2502 3496 2558 3505
rect 2502 3431 2504 3440
rect 2556 3431 2558 3440
rect 2504 3402 2556 3408
rect 2320 3188 2372 3194
rect 2320 3130 2372 3136
rect 2608 2990 2636 3878
rect 2976 3738 3004 3878
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 2596 2984 2648 2990
rect 2596 2926 2648 2932
rect 2608 2514 2636 2926
rect 2976 2922 3004 3674
rect 2964 2916 3016 2922
rect 2964 2858 3016 2864
rect 2596 2508 2648 2514
rect 2596 2450 2648 2456
rect 3344 480 3372 4678
rect 4080 4010 4108 4950
rect 4632 4826 4660 5306
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 4724 4486 4752 5646
rect 4816 5642 4844 6054
rect 4804 5636 4856 5642
rect 4804 5578 4856 5584
rect 4816 5030 4844 5578
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 4712 4480 4764 4486
rect 4712 4422 4764 4428
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 4724 4010 4752 4422
rect 4068 4004 4120 4010
rect 4068 3946 4120 3952
rect 4712 4004 4764 4010
rect 4712 3946 4764 3952
rect 4724 3754 4752 3946
rect 4632 3738 4752 3754
rect 4620 3732 4752 3738
rect 4672 3726 4752 3732
rect 4620 3674 4672 3680
rect 4712 3664 4764 3670
rect 4712 3606 4764 3612
rect 4724 3505 4752 3606
rect 4710 3496 4766 3505
rect 4710 3431 4766 3440
rect 3516 3392 3568 3398
rect 3516 3334 3568 3340
rect 3528 3194 3556 3334
rect 4220 3292 4516 3312
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 4724 3194 4752 3431
rect 3516 3188 3568 3194
rect 3516 3130 3568 3136
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4220 2128 4516 2148
rect 5000 610 5028 9454
rect 6460 9444 6512 9450
rect 6460 9386 6512 9392
rect 5172 9036 5224 9042
rect 5172 8978 5224 8984
rect 5184 8566 5212 8978
rect 6472 8974 6500 9386
rect 7116 9382 7144 10134
rect 7208 9926 7236 10542
rect 7852 10062 7880 10950
rect 8496 10606 8524 10950
rect 8484 10600 8536 10606
rect 8484 10542 8536 10548
rect 8496 10266 8524 10542
rect 9692 10538 9720 11698
rect 11152 11688 11204 11694
rect 11150 11656 11152 11665
rect 11204 11656 11206 11665
rect 11150 11591 11206 11600
rect 10692 11212 10744 11218
rect 10692 11154 10744 11160
rect 10414 11112 10470 11121
rect 10414 11047 10416 11056
rect 10468 11047 10470 11056
rect 10416 11018 10468 11024
rect 9680 10532 9732 10538
rect 9680 10474 9732 10480
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 7288 10056 7340 10062
rect 7288 9998 7340 10004
rect 7840 10056 7892 10062
rect 7840 9998 7892 10004
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 6564 9042 6592 9318
rect 7300 9110 7328 9998
rect 8496 9722 8524 10202
rect 9692 10062 9720 10474
rect 10704 10470 10732 11154
rect 11058 10840 11114 10849
rect 11114 10784 11192 10792
rect 11058 10775 11060 10784
rect 11112 10764 11192 10784
rect 11060 10746 11112 10752
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 9784 10130 9812 10406
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 8484 9716 8536 9722
rect 8484 9658 8536 9664
rect 7840 9512 7892 9518
rect 7840 9454 7892 9460
rect 7852 9178 7880 9454
rect 8496 9178 8524 9658
rect 9956 9444 10008 9450
rect 9956 9386 10008 9392
rect 10140 9444 10192 9450
rect 10140 9386 10192 9392
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 7840 9172 7892 9178
rect 7840 9114 7892 9120
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 7288 9104 7340 9110
rect 7288 9046 7340 9052
rect 6552 9036 6604 9042
rect 6552 8978 6604 8984
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 5172 8560 5224 8566
rect 5172 8502 5224 8508
rect 6472 8362 6500 8910
rect 6564 8634 6592 8978
rect 6552 8628 6604 8634
rect 6552 8570 6604 8576
rect 6460 8356 6512 8362
rect 6460 8298 6512 8304
rect 6564 8090 6592 8570
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 6932 7750 6960 8298
rect 9692 8294 9720 9318
rect 9680 8288 9732 8294
rect 9680 8230 9732 8236
rect 9692 7886 9720 8230
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 5448 7472 5500 7478
rect 5448 7414 5500 7420
rect 5460 5114 5488 7414
rect 5540 7268 5592 7274
rect 5540 7210 5592 7216
rect 5632 7268 5684 7274
rect 5632 7210 5684 7216
rect 5552 6934 5580 7210
rect 5540 6928 5592 6934
rect 5540 6870 5592 6876
rect 5552 6798 5580 6870
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5644 6662 5672 7210
rect 6932 7206 6960 7686
rect 9324 7342 9352 7822
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 9586 7304 9642 7313
rect 5724 7200 5776 7206
rect 5724 7142 5776 7148
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 5736 6662 5764 7142
rect 6932 7018 6960 7142
rect 6748 6990 6960 7018
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 6196 6746 6224 6802
rect 6274 6760 6330 6769
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5920 6118 5948 6734
rect 6196 6718 6274 6746
rect 6274 6695 6330 6704
rect 6184 6656 6236 6662
rect 6184 6598 6236 6604
rect 5908 6112 5960 6118
rect 5908 6054 5960 6060
rect 5920 5710 5948 6054
rect 6196 5846 6224 6598
rect 6288 6458 6316 6695
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6748 6118 6776 6990
rect 6828 6928 6880 6934
rect 6828 6870 6880 6876
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6840 5930 6868 6870
rect 9324 6458 9352 7278
rect 9586 7239 9588 7248
rect 9640 7239 9642 7248
rect 9588 7210 9640 7216
rect 9600 7002 9628 7210
rect 9588 6996 9640 7002
rect 9588 6938 9640 6944
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 8208 6384 8260 6390
rect 8208 6326 8260 6332
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 6840 5914 6960 5930
rect 6840 5908 6972 5914
rect 6840 5902 6920 5908
rect 6920 5850 6972 5856
rect 6184 5840 6236 5846
rect 6184 5782 6236 5788
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 5460 5086 5672 5114
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5356 4480 5408 4486
rect 5552 4468 5580 4966
rect 5644 4826 5672 5086
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5736 4758 5764 5510
rect 6196 5370 6224 5782
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 6184 5364 6236 5370
rect 6184 5306 6236 5312
rect 6288 5030 6316 5510
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 5724 4752 5776 4758
rect 5724 4694 5776 4700
rect 5356 4422 5408 4428
rect 5460 4440 5580 4468
rect 5368 4214 5396 4422
rect 5172 4208 5224 4214
rect 5172 4150 5224 4156
rect 5356 4208 5408 4214
rect 5356 4150 5408 4156
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 5092 2582 5120 3878
rect 5184 3534 5212 4150
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 5184 3194 5212 3470
rect 5460 3466 5488 4440
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5644 3670 5672 4082
rect 5736 3738 5764 4694
rect 5828 4214 5856 4966
rect 6184 4820 6236 4826
rect 6184 4762 6236 4768
rect 6092 4684 6144 4690
rect 6092 4626 6144 4632
rect 5816 4208 5868 4214
rect 5816 4150 5868 4156
rect 5816 4004 5868 4010
rect 5816 3946 5868 3952
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5632 3664 5684 3670
rect 5632 3606 5684 3612
rect 5448 3460 5500 3466
rect 5448 3402 5500 3408
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5356 2848 5408 2854
rect 5356 2790 5408 2796
rect 5080 2576 5132 2582
rect 5080 2518 5132 2524
rect 5368 2514 5396 2790
rect 5644 2650 5672 3606
rect 5828 3194 5856 3946
rect 5998 3904 6054 3913
rect 5998 3839 6054 3848
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5356 2508 5408 2514
rect 5356 2450 5408 2456
rect 4712 604 4764 610
rect 4712 546 4764 552
rect 4988 604 5040 610
rect 4988 546 5040 552
rect 4724 480 4752 546
rect 6012 480 6040 3839
rect 6104 3738 6132 4626
rect 6196 4282 6224 4762
rect 6184 4276 6236 4282
rect 6184 4218 6236 4224
rect 6288 4162 6316 4966
rect 6840 4554 6868 5102
rect 7852 4826 7880 6190
rect 8220 5778 8248 6326
rect 9416 6322 9444 6598
rect 9404 6316 9456 6322
rect 9404 6258 9456 6264
rect 8666 6216 8722 6225
rect 8666 6151 8668 6160
rect 8720 6151 8722 6160
rect 8668 6122 8720 6128
rect 8208 5772 8260 5778
rect 8208 5714 8260 5720
rect 9220 5772 9272 5778
rect 9220 5714 9272 5720
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8760 5568 8812 5574
rect 8760 5510 8812 5516
rect 8852 5568 8904 5574
rect 8852 5510 8904 5516
rect 8208 5364 8260 5370
rect 8312 5352 8340 5510
rect 8260 5324 8340 5352
rect 8208 5306 8260 5312
rect 8772 5030 8800 5510
rect 8864 5098 8892 5510
rect 9232 5370 9260 5714
rect 9508 5574 9536 6734
rect 9496 5568 9548 5574
rect 9496 5510 9548 5516
rect 9220 5364 9272 5370
rect 9220 5306 9272 5312
rect 8852 5092 8904 5098
rect 8852 5034 8904 5040
rect 8760 5024 8812 5030
rect 8760 4966 8812 4972
rect 7840 4820 7892 4826
rect 7840 4762 7892 4768
rect 6828 4548 6880 4554
rect 6828 4490 6880 4496
rect 7104 4480 7156 4486
rect 7104 4422 7156 4428
rect 6196 4134 6316 4162
rect 6092 3732 6144 3738
rect 6092 3674 6144 3680
rect 6104 3602 6132 3674
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 6196 3534 6224 4134
rect 6184 3528 6236 3534
rect 6184 3470 6236 3476
rect 6196 2854 6224 3470
rect 6184 2848 6236 2854
rect 6184 2790 6236 2796
rect 7116 2650 7144 4422
rect 7852 4282 7880 4762
rect 8300 4752 8352 4758
rect 8128 4700 8300 4706
rect 8128 4694 8352 4700
rect 8128 4678 8340 4694
rect 8864 4690 8892 5034
rect 9508 4706 9536 5510
rect 9588 5296 9640 5302
rect 9588 5238 9640 5244
rect 9600 4865 9628 5238
rect 9586 4856 9642 4865
rect 9586 4791 9642 4800
rect 8852 4684 8904 4690
rect 7840 4276 7892 4282
rect 7840 4218 7892 4224
rect 7852 4049 7880 4218
rect 8128 4146 8156 4678
rect 9508 4678 9628 4706
rect 8852 4626 8904 4632
rect 8576 4616 8628 4622
rect 8206 4584 8262 4593
rect 8576 4558 8628 4564
rect 8206 4519 8208 4528
rect 8260 4519 8262 4528
rect 8208 4490 8260 4496
rect 8588 4282 8616 4558
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 8576 4276 8628 4282
rect 8576 4218 8628 4224
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 7838 4040 7894 4049
rect 8312 4026 8340 4218
rect 7838 3975 7894 3984
rect 8220 3998 8340 4026
rect 8758 4040 8814 4049
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7656 3392 7708 3398
rect 7656 3334 7708 3340
rect 7668 2990 7696 3334
rect 7196 2984 7248 2990
rect 7196 2926 7248 2932
rect 7656 2984 7708 2990
rect 7656 2926 7708 2932
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 7208 592 7236 2926
rect 7562 2816 7618 2825
rect 7562 2751 7618 2760
rect 7576 2650 7604 2751
rect 7668 2650 7696 2926
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 7656 2644 7708 2650
rect 7656 2586 7708 2592
rect 7760 2310 7788 3878
rect 8220 3738 8248 3998
rect 8758 3975 8760 3984
rect 8812 3975 8814 3984
rect 8760 3946 8812 3952
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 8312 3398 8340 3878
rect 9232 3466 9260 3878
rect 9496 3664 9548 3670
rect 9496 3606 9548 3612
rect 9220 3460 9272 3466
rect 9220 3402 9272 3408
rect 9508 3398 9536 3606
rect 9600 3534 9628 4678
rect 9968 3913 9996 9386
rect 10152 9110 10180 9386
rect 10428 9178 10456 10066
rect 10704 9994 10732 10406
rect 10692 9988 10744 9994
rect 10692 9930 10744 9936
rect 11072 9926 11100 10610
rect 11164 10606 11192 10764
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 11164 10198 11192 10542
rect 11152 10192 11204 10198
rect 11152 10134 11204 10140
rect 11060 9920 11112 9926
rect 10980 9880 11060 9908
rect 10980 9450 11008 9880
rect 11060 9862 11112 9868
rect 10968 9444 11020 9450
rect 10968 9386 11020 9392
rect 10416 9172 10468 9178
rect 10416 9114 10468 9120
rect 10140 9104 10192 9110
rect 10140 9046 10192 9052
rect 11256 8022 11284 12038
rect 12440 11824 12492 11830
rect 12440 11766 12492 11772
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11900 11286 11928 11698
rect 12348 11688 12400 11694
rect 12348 11630 12400 11636
rect 11888 11280 11940 11286
rect 11888 11222 11940 11228
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 11428 10736 11480 10742
rect 11426 10704 11428 10713
rect 11480 10704 11482 10713
rect 11624 10674 11652 11154
rect 11900 10810 11928 11222
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 11426 10639 11482 10648
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 12360 10266 12388 11630
rect 12452 10606 12480 11766
rect 13544 11756 13596 11762
rect 13544 11698 13596 11704
rect 12530 11520 12586 11529
rect 12530 11455 12586 11464
rect 12544 10810 12572 11455
rect 13084 11348 13136 11354
rect 13084 11290 13136 11296
rect 12990 11112 13046 11121
rect 12990 11047 13046 11056
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 13004 10538 13032 11047
rect 13096 10674 13124 11290
rect 13556 11218 13584 11698
rect 13648 11694 13676 12038
rect 16040 11762 16068 12038
rect 17880 11898 17908 12242
rect 18248 11898 18276 12310
rect 19904 12306 19932 13790
rect 20272 12782 20300 13874
rect 20628 13864 20680 13870
rect 20680 13812 20760 13818
rect 20628 13806 20760 13812
rect 20640 13790 20760 13806
rect 20732 13682 20760 13790
rect 20732 13654 20852 13682
rect 20352 13184 20404 13190
rect 20352 13126 20404 13132
rect 20364 12850 20392 13126
rect 20442 12880 20498 12889
rect 20352 12844 20404 12850
rect 20442 12815 20498 12824
rect 20352 12786 20404 12792
rect 19984 12776 20036 12782
rect 19984 12718 20036 12724
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 18878 12271 18934 12280
rect 19892 12300 19944 12306
rect 19892 12242 19944 12248
rect 18512 12232 18564 12238
rect 18432 12180 18512 12186
rect 18432 12174 18564 12180
rect 18432 12158 18552 12174
rect 17868 11892 17920 11898
rect 17868 11834 17920 11840
rect 18236 11892 18288 11898
rect 18236 11834 18288 11840
rect 16028 11756 16080 11762
rect 16028 11698 16080 11704
rect 13636 11688 13688 11694
rect 13636 11630 13688 11636
rect 13648 11354 13676 11630
rect 14924 11552 14976 11558
rect 15476 11552 15528 11558
rect 14924 11494 14976 11500
rect 15474 11520 15476 11529
rect 15844 11552 15896 11558
rect 15528 11520 15530 11529
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 14936 11286 14964 11494
rect 15844 11494 15896 11500
rect 15474 11455 15530 11464
rect 15856 11354 15884 11494
rect 15844 11348 15896 11354
rect 15844 11290 15896 11296
rect 16040 11286 16068 11698
rect 18144 11552 18196 11558
rect 18144 11494 18196 11500
rect 14924 11280 14976 11286
rect 14924 11222 14976 11228
rect 16028 11280 16080 11286
rect 16028 11222 16080 11228
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 15672 10810 15700 11154
rect 16040 10810 16068 11222
rect 18156 11150 18184 11494
rect 18432 11218 18460 12158
rect 19996 12102 20024 12718
rect 20272 12442 20300 12718
rect 20456 12646 20484 12815
rect 20444 12640 20496 12646
rect 20444 12582 20496 12588
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20260 12436 20312 12442
rect 20260 12378 20312 12384
rect 20628 12368 20680 12374
rect 20732 12322 20760 12582
rect 20824 12374 20852 13654
rect 26620 13394 26648 14010
rect 26608 13388 26660 13394
rect 26608 13330 26660 13336
rect 27160 13388 27212 13394
rect 27160 13330 27212 13336
rect 27172 12986 27200 13330
rect 27160 12980 27212 12986
rect 27160 12922 27212 12928
rect 20994 12880 21050 12889
rect 20994 12815 21050 12824
rect 20680 12316 20760 12322
rect 20628 12310 20760 12316
rect 20812 12368 20864 12374
rect 20812 12310 20864 12316
rect 20640 12294 20760 12310
rect 18604 12096 18656 12102
rect 18604 12038 18656 12044
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 19984 12096 20036 12102
rect 19984 12038 20036 12044
rect 20444 12096 20496 12102
rect 20444 12038 20496 12044
rect 18420 11212 18472 11218
rect 18420 11154 18472 11160
rect 18144 11144 18196 11150
rect 18144 11086 18196 11092
rect 17776 11008 17828 11014
rect 17776 10950 17828 10956
rect 15660 10804 15712 10810
rect 15580 10764 15660 10792
rect 13084 10668 13136 10674
rect 13084 10610 13136 10616
rect 12992 10532 13044 10538
rect 12992 10474 13044 10480
rect 13004 10266 13032 10474
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 12254 9616 12310 9625
rect 12360 9586 12388 10202
rect 12532 10192 12584 10198
rect 12532 10134 12584 10140
rect 12544 9722 12572 10134
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 15200 10056 15252 10062
rect 15200 9998 15252 10004
rect 12820 9722 12848 9998
rect 12532 9716 12584 9722
rect 12532 9658 12584 9664
rect 12808 9716 12860 9722
rect 12808 9658 12860 9664
rect 15212 9602 15240 9998
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 12254 9551 12310 9560
rect 12348 9580 12400 9586
rect 12268 9110 12296 9551
rect 12348 9522 12400 9528
rect 15120 9574 15240 9602
rect 14648 9444 14700 9450
rect 14648 9386 14700 9392
rect 12256 9104 12308 9110
rect 12256 9046 12308 9052
rect 11980 8968 12032 8974
rect 11980 8910 12032 8916
rect 11992 8430 12020 8910
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 11992 8294 12020 8366
rect 11980 8288 12032 8294
rect 11980 8230 12032 8236
rect 11244 8016 11296 8022
rect 11244 7958 11296 7964
rect 11256 7546 11284 7958
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 10232 7200 10284 7206
rect 10232 7142 10284 7148
rect 10244 7002 10272 7142
rect 11256 7002 11284 7482
rect 11808 7313 11836 7686
rect 11992 7546 12020 8230
rect 12268 8090 12296 9046
rect 13820 8900 13872 8906
rect 13820 8842 13872 8848
rect 12624 8832 12676 8838
rect 12544 8780 12624 8786
rect 12544 8774 12676 8780
rect 12544 8758 12664 8774
rect 12544 8362 12572 8758
rect 12532 8356 12584 8362
rect 12532 8298 12584 8304
rect 12256 8084 12308 8090
rect 12256 8026 12308 8032
rect 12544 8022 12572 8298
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 12532 8016 12584 8022
rect 12532 7958 12584 7964
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 11992 7342 12020 7482
rect 11980 7336 12032 7342
rect 11794 7304 11850 7313
rect 11980 7278 12032 7284
rect 12348 7336 12400 7342
rect 12348 7278 12400 7284
rect 11794 7239 11850 7248
rect 10232 6996 10284 7002
rect 10232 6938 10284 6944
rect 11244 6996 11296 7002
rect 11244 6938 11296 6944
rect 11612 6996 11664 7002
rect 11612 6938 11664 6944
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 10060 6769 10088 6802
rect 10046 6760 10102 6769
rect 10046 6695 10102 6704
rect 10060 6458 10088 6695
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10060 5778 10088 6394
rect 10244 6254 10272 6938
rect 11336 6656 11388 6662
rect 11336 6598 11388 6604
rect 10232 6248 10284 6254
rect 11348 6225 11376 6598
rect 11624 6458 11652 6938
rect 11808 6798 11836 7239
rect 12360 7206 12388 7278
rect 12348 7200 12400 7206
rect 12348 7142 12400 7148
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 11980 6860 12032 6866
rect 11980 6802 12032 6808
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 11808 6458 11836 6734
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 10232 6190 10284 6196
rect 11334 6216 11390 6225
rect 10244 5914 10272 6190
rect 11334 6151 11390 6160
rect 11992 5914 12020 6802
rect 10232 5908 10284 5914
rect 10232 5850 10284 5856
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 11520 5840 11572 5846
rect 11520 5782 11572 5788
rect 10048 5772 10100 5778
rect 10048 5714 10100 5720
rect 11336 5772 11388 5778
rect 11336 5714 11388 5720
rect 11058 5672 11114 5681
rect 11058 5607 11060 5616
rect 11112 5607 11114 5616
rect 11060 5578 11112 5584
rect 11348 5370 11376 5714
rect 11532 5370 11560 5782
rect 12452 5778 12480 7142
rect 12544 7002 12572 7958
rect 12912 7886 12940 8230
rect 13832 7954 13860 8842
rect 14660 8838 14688 9386
rect 15016 9036 15068 9042
rect 15016 8978 15068 8984
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14660 8498 14688 8774
rect 15028 8634 15056 8978
rect 15120 8906 15148 9574
rect 15292 9512 15344 9518
rect 15292 9454 15344 9460
rect 15304 8974 15332 9454
rect 15292 8968 15344 8974
rect 15292 8910 15344 8916
rect 15108 8900 15160 8906
rect 15108 8842 15160 8848
rect 15016 8628 15068 8634
rect 15016 8570 15068 8576
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 15120 8401 15148 8842
rect 15304 8634 15332 8910
rect 15292 8628 15344 8634
rect 15292 8570 15344 8576
rect 15106 8392 15162 8401
rect 15106 8327 15162 8336
rect 13820 7948 13872 7954
rect 13820 7890 13872 7896
rect 12900 7880 12952 7886
rect 12900 7822 12952 7828
rect 13084 7880 13136 7886
rect 13084 7822 13136 7828
rect 12808 7540 12860 7546
rect 12912 7528 12940 7822
rect 12860 7500 12940 7528
rect 12808 7482 12860 7488
rect 12912 7274 12940 7500
rect 12900 7268 12952 7274
rect 12900 7210 12952 7216
rect 12912 7002 12940 7210
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 13096 6186 13124 7822
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 13832 6866 13860 7686
rect 15028 7206 15056 7686
rect 15108 7472 15160 7478
rect 15160 7420 15240 7426
rect 15108 7414 15240 7420
rect 15120 7398 15240 7414
rect 13912 7200 13964 7206
rect 13912 7142 13964 7148
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 13820 6860 13872 6866
rect 13820 6802 13872 6808
rect 13360 6656 13412 6662
rect 13360 6598 13412 6604
rect 13372 6254 13400 6598
rect 13636 6384 13688 6390
rect 13636 6326 13688 6332
rect 13360 6248 13412 6254
rect 13360 6190 13412 6196
rect 13084 6180 13136 6186
rect 13084 6122 13136 6128
rect 12900 6112 12952 6118
rect 12900 6054 12952 6060
rect 12912 5846 12940 6054
rect 13372 5914 13400 6190
rect 13360 5908 13412 5914
rect 13360 5850 13412 5856
rect 12900 5840 12952 5846
rect 12900 5782 12952 5788
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 11612 5704 11664 5710
rect 11612 5646 11664 5652
rect 11336 5364 11388 5370
rect 11336 5306 11388 5312
rect 11520 5364 11572 5370
rect 11520 5306 11572 5312
rect 11244 5160 11296 5166
rect 11244 5102 11296 5108
rect 10324 4684 10376 4690
rect 10324 4626 10376 4632
rect 10232 4480 10284 4486
rect 10232 4422 10284 4428
rect 10244 4321 10272 4422
rect 10230 4312 10286 4321
rect 10230 4247 10286 4256
rect 10336 3942 10364 4626
rect 11256 4554 11284 5102
rect 11624 5030 11652 5646
rect 12452 5370 12480 5714
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 11612 5024 11664 5030
rect 11612 4966 11664 4972
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 11532 4593 11560 4626
rect 11518 4584 11574 4593
rect 11244 4548 11296 4554
rect 11518 4519 11574 4528
rect 11244 4490 11296 4496
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 11072 4078 11100 4422
rect 11532 4214 11560 4519
rect 11624 4457 11652 4966
rect 11716 4865 11744 4966
rect 11702 4856 11758 4865
rect 12912 4826 12940 5782
rect 13544 5228 13596 5234
rect 13544 5170 13596 5176
rect 11702 4791 11704 4800
rect 11756 4791 11758 4800
rect 12900 4820 12952 4826
rect 11704 4762 11756 4768
rect 12900 4762 12952 4768
rect 11610 4448 11666 4457
rect 11610 4383 11666 4392
rect 11520 4208 11572 4214
rect 11520 4150 11572 4156
rect 11716 4146 11744 4762
rect 11796 4616 11848 4622
rect 11796 4558 11848 4564
rect 11808 4282 11836 4558
rect 12808 4480 12860 4486
rect 12808 4422 12860 4428
rect 13176 4480 13228 4486
rect 13176 4422 13228 4428
rect 13452 4480 13504 4486
rect 13452 4422 13504 4428
rect 11796 4276 11848 4282
rect 11796 4218 11848 4224
rect 11980 4208 12032 4214
rect 11978 4176 11980 4185
rect 12032 4176 12034 4185
rect 11704 4140 11756 4146
rect 11978 4111 12034 4120
rect 11704 4082 11756 4088
rect 12820 4078 12848 4422
rect 13188 4146 13216 4422
rect 13358 4312 13414 4321
rect 13464 4282 13492 4422
rect 13358 4247 13414 4256
rect 13452 4276 13504 4282
rect 13372 4146 13400 4247
rect 13452 4218 13504 4224
rect 13176 4140 13228 4146
rect 13176 4082 13228 4088
rect 13360 4140 13412 4146
rect 13360 4082 13412 4088
rect 11060 4072 11112 4078
rect 11060 4014 11112 4020
rect 12348 4072 12400 4078
rect 12808 4072 12860 4078
rect 12400 4020 12572 4026
rect 12348 4014 12572 4020
rect 12808 4014 12860 4020
rect 12360 3998 12572 4014
rect 10324 3936 10376 3942
rect 9954 3904 10010 3913
rect 9954 3839 10010 3848
rect 10322 3904 10324 3913
rect 10376 3904 10378 3913
rect 10322 3839 10378 3848
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 8300 3392 8352 3398
rect 8220 3352 8300 3380
rect 8220 2378 8248 3352
rect 8300 3334 8352 3340
rect 9496 3392 9548 3398
rect 9496 3334 9548 3340
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8496 2514 8524 3130
rect 9508 2922 9536 3334
rect 9496 2916 9548 2922
rect 9496 2858 9548 2864
rect 8760 2848 8812 2854
rect 8760 2790 8812 2796
rect 8772 2582 8800 2790
rect 8760 2576 8812 2582
rect 8760 2518 8812 2524
rect 9600 2514 9628 3470
rect 11256 3194 11284 3538
rect 11336 3528 11388 3534
rect 11336 3470 11388 3476
rect 11244 3188 11296 3194
rect 11244 3130 11296 3136
rect 11348 2990 11376 3470
rect 9772 2984 9824 2990
rect 9772 2926 9824 2932
rect 11336 2984 11388 2990
rect 11336 2926 11388 2932
rect 9784 2854 9812 2926
rect 11152 2916 11204 2922
rect 11152 2858 11204 2864
rect 9772 2848 9824 2854
rect 9772 2790 9824 2796
rect 10046 2816 10102 2825
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 9588 2508 9640 2514
rect 9588 2450 9640 2456
rect 9784 2446 9812 2790
rect 10046 2751 10102 2760
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 8208 2372 8260 2378
rect 8208 2314 8260 2320
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 8760 2304 8812 2310
rect 8760 2246 8812 2252
rect 7208 564 7420 592
rect 7392 480 7420 564
rect 8772 480 8800 2246
rect 10060 480 10088 2751
rect 11164 2650 11192 2858
rect 12544 2650 12572 3998
rect 12806 3904 12862 3913
rect 12806 3839 12862 3848
rect 12716 3392 12768 3398
rect 12716 3334 12768 3340
rect 12728 2990 12756 3334
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 12532 2644 12584 2650
rect 12532 2586 12584 2592
rect 12728 2582 12756 2926
rect 12716 2576 12768 2582
rect 12716 2518 12768 2524
rect 11428 2508 11480 2514
rect 11428 2450 11480 2456
rect 11440 480 11468 2450
rect 12820 480 12848 3839
rect 13188 3670 13216 4082
rect 13556 4010 13584 5170
rect 13648 4842 13676 6326
rect 13924 6202 13952 7142
rect 13740 6174 13952 6202
rect 13740 6118 13768 6174
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 14096 6112 14148 6118
rect 14096 6054 14148 6060
rect 14004 5908 14056 5914
rect 14004 5850 14056 5856
rect 14016 5166 14044 5850
rect 14004 5160 14056 5166
rect 14004 5102 14056 5108
rect 13648 4826 13860 4842
rect 13648 4820 13872 4826
rect 13648 4814 13820 4820
rect 13544 4004 13596 4010
rect 13544 3946 13596 3952
rect 13176 3664 13228 3670
rect 13176 3606 13228 3612
rect 13556 2922 13584 3946
rect 13648 3738 13676 4814
rect 13820 4762 13872 4768
rect 14108 4486 14136 6054
rect 15028 4622 15056 7142
rect 15212 6866 15240 7398
rect 15396 7274 15424 9862
rect 15580 9518 15608 10764
rect 15660 10746 15712 10752
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 17788 10470 17816 10950
rect 18432 10810 18460 11154
rect 18512 11008 18564 11014
rect 18512 10950 18564 10956
rect 18420 10804 18472 10810
rect 18420 10746 18472 10752
rect 18524 10606 18552 10950
rect 18512 10600 18564 10606
rect 18512 10542 18564 10548
rect 17868 10532 17920 10538
rect 17868 10474 17920 10480
rect 17776 10464 17828 10470
rect 17776 10406 17828 10412
rect 15936 10192 15988 10198
rect 15936 10134 15988 10140
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 15672 9722 15700 10066
rect 15660 9716 15712 9722
rect 15660 9658 15712 9664
rect 15672 9625 15700 9658
rect 15658 9616 15714 9625
rect 15658 9551 15714 9560
rect 15568 9512 15620 9518
rect 15568 9454 15620 9460
rect 15948 9382 15976 10134
rect 16672 9648 16724 9654
rect 16672 9590 16724 9596
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 15948 9042 15976 9318
rect 16684 9178 16712 9590
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 15936 9036 15988 9042
rect 15936 8978 15988 8984
rect 17788 8974 17816 10406
rect 17880 10266 17908 10474
rect 18524 10266 18552 10542
rect 18616 10538 18644 12038
rect 19260 11626 19288 12038
rect 19248 11620 19300 11626
rect 19248 11562 19300 11568
rect 19260 11082 19288 11562
rect 19580 11452 19876 11472
rect 19636 11450 19660 11452
rect 19716 11450 19740 11452
rect 19796 11450 19820 11452
rect 19658 11398 19660 11450
rect 19722 11398 19734 11450
rect 19796 11398 19798 11450
rect 19636 11396 19660 11398
rect 19716 11396 19740 11398
rect 19796 11396 19820 11398
rect 19580 11376 19876 11396
rect 19248 11076 19300 11082
rect 19248 11018 19300 11024
rect 19248 10736 19300 10742
rect 20456 10713 20484 12038
rect 20732 11642 20760 12294
rect 20904 12232 20956 12238
rect 20904 12174 20956 12180
rect 20916 11830 20944 12174
rect 20904 11824 20956 11830
rect 20904 11766 20956 11772
rect 20732 11614 20944 11642
rect 20628 11552 20680 11558
rect 20628 11494 20680 11500
rect 20640 10996 20668 11494
rect 20916 11082 20944 11614
rect 20904 11076 20956 11082
rect 20904 11018 20956 11024
rect 20720 11008 20772 11014
rect 20640 10968 20720 10996
rect 20720 10950 20772 10956
rect 19248 10678 19300 10684
rect 20258 10704 20314 10713
rect 18604 10532 18656 10538
rect 18604 10474 18656 10480
rect 18616 10266 18644 10474
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 18512 10260 18564 10266
rect 18512 10202 18564 10208
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 18052 9036 18104 9042
rect 18052 8978 18104 8984
rect 17776 8968 17828 8974
rect 17776 8910 17828 8916
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 17684 8832 17736 8838
rect 17684 8774 17736 8780
rect 16396 8560 16448 8566
rect 16396 8502 16448 8508
rect 16408 8022 16436 8502
rect 16946 8392 17002 8401
rect 17604 8362 17632 8774
rect 17696 8498 17724 8774
rect 17788 8634 17816 8910
rect 17776 8628 17828 8634
rect 17776 8570 17828 8576
rect 17684 8492 17736 8498
rect 17684 8434 17736 8440
rect 16946 8327 16948 8336
rect 17000 8327 17002 8336
rect 17592 8356 17644 8362
rect 16948 8298 17000 8304
rect 17592 8298 17644 8304
rect 16856 8288 16908 8294
rect 16856 8230 16908 8236
rect 16868 8090 16896 8230
rect 16856 8084 16908 8090
rect 16856 8026 16908 8032
rect 16960 8022 16988 8298
rect 16396 8016 16448 8022
rect 16396 7958 16448 7964
rect 16488 8016 16540 8022
rect 16488 7958 16540 7964
rect 16948 8016 17000 8022
rect 16948 7958 17000 7964
rect 16028 7744 16080 7750
rect 16028 7686 16080 7692
rect 15292 7268 15344 7274
rect 15292 7210 15344 7216
rect 15384 7268 15436 7274
rect 15384 7210 15436 7216
rect 15304 7002 15332 7210
rect 15292 6996 15344 7002
rect 15292 6938 15344 6944
rect 16040 6866 16068 7686
rect 16408 7546 16436 7958
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16500 7478 16528 7958
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 16488 7472 16540 7478
rect 16488 7414 16540 7420
rect 16592 7206 16620 7822
rect 16960 7342 16988 7958
rect 17788 7954 17816 8570
rect 18064 8090 18092 8978
rect 18512 8356 18564 8362
rect 18512 8298 18564 8304
rect 18052 8084 18104 8090
rect 18052 8026 18104 8032
rect 17776 7948 17828 7954
rect 17776 7890 17828 7896
rect 17788 7546 17816 7890
rect 17776 7540 17828 7546
rect 17828 7500 17908 7528
rect 17776 7482 17828 7488
rect 16948 7336 17000 7342
rect 16948 7278 17000 7284
rect 16580 7200 16632 7206
rect 16580 7142 16632 7148
rect 15200 6860 15252 6866
rect 15200 6802 15252 6808
rect 15476 6860 15528 6866
rect 15476 6802 15528 6808
rect 16028 6860 16080 6866
rect 16028 6802 16080 6808
rect 16396 6860 16448 6866
rect 16396 6802 16448 6808
rect 15488 5914 15516 6802
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15936 6656 15988 6662
rect 15936 6598 15988 6604
rect 15764 6254 15792 6598
rect 15844 6316 15896 6322
rect 15844 6258 15896 6264
rect 15752 6248 15804 6254
rect 15752 6190 15804 6196
rect 15476 5908 15528 5914
rect 15476 5850 15528 5856
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 15764 5370 15792 5714
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 15108 5024 15160 5030
rect 15108 4966 15160 4972
rect 15016 4616 15068 4622
rect 15016 4558 15068 4564
rect 15028 4486 15056 4558
rect 13820 4480 13872 4486
rect 14096 4480 14148 4486
rect 13820 4422 13872 4428
rect 13910 4448 13966 4457
rect 13832 4321 13860 4422
rect 14096 4422 14148 4428
rect 15016 4480 15068 4486
rect 15016 4422 15068 4428
rect 13910 4383 13966 4392
rect 13818 4312 13874 4321
rect 13818 4247 13874 4256
rect 13636 3732 13688 3738
rect 13636 3674 13688 3680
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 13832 3194 13860 3538
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 13544 2916 13596 2922
rect 13544 2858 13596 2864
rect 13924 2854 13952 4383
rect 15028 3398 15056 4422
rect 15120 4078 15148 4966
rect 15856 4826 15884 6258
rect 15948 6186 15976 6598
rect 16408 6458 16436 6802
rect 16396 6452 16448 6458
rect 16396 6394 16448 6400
rect 16488 6384 16540 6390
rect 16488 6326 16540 6332
rect 15936 6180 15988 6186
rect 15936 6122 15988 6128
rect 16120 5840 16172 5846
rect 16120 5782 16172 5788
rect 16132 5030 16160 5782
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 15844 4820 15896 4826
rect 15844 4762 15896 4768
rect 15476 4480 15528 4486
rect 15476 4422 15528 4428
rect 15108 4072 15160 4078
rect 15108 4014 15160 4020
rect 15488 3738 15516 4422
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 15476 3732 15528 3738
rect 15476 3674 15528 3680
rect 15672 3670 15700 3878
rect 15856 3670 15884 4762
rect 16132 4457 16160 4966
rect 16212 4548 16264 4554
rect 16212 4490 16264 4496
rect 16118 4448 16174 4457
rect 16118 4383 16174 4392
rect 16224 4282 16252 4490
rect 16212 4276 16264 4282
rect 16212 4218 16264 4224
rect 16500 3913 16528 6326
rect 16672 4752 16724 4758
rect 16672 4694 16724 4700
rect 16684 4282 16712 4694
rect 16960 4690 16988 7278
rect 17880 6882 17908 7500
rect 18524 7274 18552 8298
rect 18604 8288 18656 8294
rect 18604 8230 18656 8236
rect 18616 8022 18644 8230
rect 18604 8016 18656 8022
rect 18604 7958 18656 7964
rect 18616 7410 18644 7958
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18512 7268 18564 7274
rect 18512 7210 18564 7216
rect 17880 6854 18000 6882
rect 18524 6866 18552 7210
rect 18616 7002 18644 7346
rect 18604 6996 18656 7002
rect 18604 6938 18656 6944
rect 17972 6458 18000 6854
rect 18512 6860 18564 6866
rect 18512 6802 18564 6808
rect 17960 6452 18012 6458
rect 17960 6394 18012 6400
rect 18236 6452 18288 6458
rect 18236 6394 18288 6400
rect 18052 6112 18104 6118
rect 18052 6054 18104 6060
rect 17684 5772 17736 5778
rect 17684 5714 17736 5720
rect 17406 5672 17462 5681
rect 17406 5607 17462 5616
rect 17420 5370 17448 5607
rect 17408 5364 17460 5370
rect 17408 5306 17460 5312
rect 17420 5030 17448 5306
rect 17408 5024 17460 5030
rect 17408 4966 17460 4972
rect 16948 4684 17000 4690
rect 16948 4626 17000 4632
rect 17224 4684 17276 4690
rect 17224 4626 17276 4632
rect 17132 4616 17184 4622
rect 17132 4558 17184 4564
rect 17144 4282 17172 4558
rect 16672 4276 16724 4282
rect 16672 4218 16724 4224
rect 17132 4276 17184 4282
rect 17132 4218 17184 4224
rect 16486 3904 16542 3913
rect 16486 3839 16542 3848
rect 15660 3664 15712 3670
rect 15660 3606 15712 3612
rect 15844 3664 15896 3670
rect 15844 3606 15896 3612
rect 15108 3528 15160 3534
rect 15108 3470 15160 3476
rect 15474 3496 15530 3505
rect 15016 3392 15068 3398
rect 15016 3334 15068 3340
rect 14096 3188 14148 3194
rect 14096 3130 14148 3136
rect 13912 2848 13964 2854
rect 13912 2790 13964 2796
rect 14108 480 14136 3130
rect 15120 2650 15148 3470
rect 15474 3431 15476 3440
rect 15528 3431 15530 3440
rect 15476 3402 15528 3408
rect 15672 2990 15700 3606
rect 15856 3534 15884 3606
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 16488 3392 16540 3398
rect 16486 3360 16488 3369
rect 16540 3360 16542 3369
rect 16486 3295 16542 3304
rect 16684 3194 16712 4218
rect 16856 4072 16908 4078
rect 16856 4014 16908 4020
rect 16764 3732 16816 3738
rect 16764 3674 16816 3680
rect 16396 3188 16448 3194
rect 16396 3130 16448 3136
rect 16672 3188 16724 3194
rect 16672 3130 16724 3136
rect 15660 2984 15712 2990
rect 15660 2926 15712 2932
rect 15108 2644 15160 2650
rect 15108 2586 15160 2592
rect 16408 2514 16436 3130
rect 16776 3126 16804 3674
rect 16868 3398 16896 4014
rect 16948 3936 17000 3942
rect 16948 3878 17000 3884
rect 16960 3602 16988 3878
rect 17144 3670 17172 4218
rect 17236 3738 17264 4626
rect 17224 3732 17276 3738
rect 17224 3674 17276 3680
rect 17132 3664 17184 3670
rect 17132 3606 17184 3612
rect 16948 3596 17000 3602
rect 16948 3538 17000 3544
rect 16856 3392 16908 3398
rect 16856 3334 16908 3340
rect 16868 3194 16896 3334
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 17144 3126 17172 3606
rect 17696 3602 17724 5714
rect 18064 5370 18092 6054
rect 18248 5846 18276 6394
rect 18236 5840 18288 5846
rect 18236 5782 18288 5788
rect 18248 5710 18276 5782
rect 18512 5772 18564 5778
rect 18512 5714 18564 5720
rect 18236 5704 18288 5710
rect 18236 5646 18288 5652
rect 18248 5370 18276 5646
rect 18052 5364 18104 5370
rect 18052 5306 18104 5312
rect 18236 5364 18288 5370
rect 18236 5306 18288 5312
rect 18524 5098 18552 5714
rect 18512 5092 18564 5098
rect 18512 5034 18564 5040
rect 18524 4826 18552 5034
rect 18512 4820 18564 4826
rect 18512 4762 18564 4768
rect 18696 4684 18748 4690
rect 18696 4626 18748 4632
rect 17960 4480 18012 4486
rect 17960 4422 18012 4428
rect 17776 4072 17828 4078
rect 17776 4014 17828 4020
rect 17684 3596 17736 3602
rect 17684 3538 17736 3544
rect 17696 3126 17724 3538
rect 17788 3398 17816 4014
rect 17868 3936 17920 3942
rect 17868 3878 17920 3884
rect 17776 3392 17828 3398
rect 17776 3334 17828 3340
rect 16764 3120 16816 3126
rect 16764 3062 16816 3068
rect 17132 3120 17184 3126
rect 17132 3062 17184 3068
rect 17316 3120 17368 3126
rect 17316 3062 17368 3068
rect 17684 3120 17736 3126
rect 17684 3062 17736 3068
rect 16488 3052 16540 3058
rect 16488 2994 16540 3000
rect 16500 2582 16528 2994
rect 16854 2952 16910 2961
rect 16854 2887 16910 2896
rect 16488 2576 16540 2582
rect 16488 2518 16540 2524
rect 16396 2508 16448 2514
rect 16396 2450 16448 2456
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 15488 480 15516 2246
rect 16868 480 16896 2887
rect 17328 2650 17356 3062
rect 17788 2990 17816 3334
rect 17776 2984 17828 2990
rect 17776 2926 17828 2932
rect 17880 2650 17908 3878
rect 17972 2922 18000 4422
rect 18708 4078 18736 4626
rect 18696 4072 18748 4078
rect 18142 4040 18198 4049
rect 18696 4014 18748 4020
rect 18142 3975 18198 3984
rect 18052 3120 18104 3126
rect 18052 3062 18104 3068
rect 17960 2916 18012 2922
rect 17960 2858 18012 2864
rect 18064 2650 18092 3062
rect 17316 2644 17368 2650
rect 17316 2586 17368 2592
rect 17868 2644 17920 2650
rect 17868 2586 17920 2592
rect 18052 2644 18104 2650
rect 18052 2586 18104 2592
rect 18064 2514 18092 2586
rect 18052 2508 18104 2514
rect 18052 2450 18104 2456
rect 18156 480 18184 3975
rect 18604 3936 18656 3942
rect 18604 3878 18656 3884
rect 18616 3738 18644 3878
rect 18604 3732 18656 3738
rect 18604 3674 18656 3680
rect 18694 3360 18750 3369
rect 18694 3295 18750 3304
rect 18708 3058 18736 3295
rect 19260 3233 19288 10678
rect 20258 10639 20260 10648
rect 20312 10639 20314 10648
rect 20442 10704 20498 10713
rect 20916 10674 20944 11018
rect 20442 10639 20498 10648
rect 20904 10668 20956 10674
rect 20260 10610 20312 10616
rect 19580 10364 19876 10384
rect 19636 10362 19660 10364
rect 19716 10362 19740 10364
rect 19796 10362 19820 10364
rect 19658 10310 19660 10362
rect 19722 10310 19734 10362
rect 19796 10310 19798 10362
rect 19636 10308 19660 10310
rect 19716 10308 19740 10310
rect 19796 10308 19820 10310
rect 19580 10288 19876 10308
rect 20272 10266 20300 10610
rect 20456 10606 20484 10639
rect 20904 10610 20956 10616
rect 20444 10600 20496 10606
rect 20444 10542 20496 10548
rect 21008 10470 21036 12815
rect 22284 12436 22336 12442
rect 22284 12378 22336 12384
rect 21364 12368 21416 12374
rect 22296 12345 22324 12378
rect 21364 12310 21416 12316
rect 22282 12336 22338 12345
rect 21376 11937 21404 12310
rect 27172 12306 27200 12922
rect 22282 12271 22338 12280
rect 27160 12300 27212 12306
rect 27160 12242 27212 12248
rect 23572 12096 23624 12102
rect 23572 12038 23624 12044
rect 21362 11928 21418 11937
rect 21362 11863 21364 11872
rect 21416 11863 21418 11872
rect 21364 11834 21416 11840
rect 22192 11824 22244 11830
rect 22192 11766 22244 11772
rect 22204 11150 22232 11766
rect 23584 11626 23612 12038
rect 25042 11928 25098 11937
rect 25042 11863 25044 11872
rect 25096 11863 25098 11872
rect 25044 11834 25096 11840
rect 23664 11756 23716 11762
rect 23664 11698 23716 11704
rect 23572 11620 23624 11626
rect 23572 11562 23624 11568
rect 22192 11144 22244 11150
rect 22244 11092 22324 11098
rect 22192 11086 22324 11092
rect 22204 11070 22324 11086
rect 23584 11082 23612 11562
rect 23676 11257 23704 11698
rect 26240 11280 26292 11286
rect 23662 11248 23718 11257
rect 26240 11222 26292 11228
rect 26606 11248 26662 11257
rect 23662 11183 23718 11192
rect 22192 11008 22244 11014
rect 22192 10950 22244 10956
rect 22098 10704 22154 10713
rect 22098 10639 22154 10648
rect 20996 10464 21048 10470
rect 20996 10406 21048 10412
rect 21456 10464 21508 10470
rect 21456 10406 21508 10412
rect 20260 10260 20312 10266
rect 20260 10202 20312 10208
rect 19580 9276 19876 9296
rect 19636 9274 19660 9276
rect 19716 9274 19740 9276
rect 19796 9274 19820 9276
rect 19658 9222 19660 9274
rect 19722 9222 19734 9274
rect 19796 9222 19798 9274
rect 19636 9220 19660 9222
rect 19716 9220 19740 9222
rect 19796 9220 19820 9222
rect 19580 9200 19876 9220
rect 20904 8968 20956 8974
rect 20904 8910 20956 8916
rect 20812 8832 20864 8838
rect 20812 8774 20864 8780
rect 20824 8430 20852 8774
rect 20812 8424 20864 8430
rect 20812 8366 20864 8372
rect 19580 8188 19876 8208
rect 19636 8186 19660 8188
rect 19716 8186 19740 8188
rect 19796 8186 19820 8188
rect 19658 8134 19660 8186
rect 19722 8134 19734 8186
rect 19796 8134 19798 8186
rect 19636 8132 19660 8134
rect 19716 8132 19740 8134
rect 19796 8132 19820 8134
rect 19580 8112 19876 8132
rect 20824 8090 20852 8366
rect 20260 8084 20312 8090
rect 20260 8026 20312 8032
rect 20812 8084 20864 8090
rect 20812 8026 20864 8032
rect 20272 7546 20300 8026
rect 20812 7744 20864 7750
rect 20812 7686 20864 7692
rect 20260 7540 20312 7546
rect 20260 7482 20312 7488
rect 20824 7478 20852 7686
rect 20916 7546 20944 8910
rect 21008 7886 21036 10406
rect 21468 10198 21496 10406
rect 21272 10192 21324 10198
rect 21272 10134 21324 10140
rect 21456 10192 21508 10198
rect 21456 10134 21508 10140
rect 21732 10192 21784 10198
rect 21732 10134 21784 10140
rect 21284 9654 21312 10134
rect 21468 9722 21496 10134
rect 21744 9722 21772 10134
rect 21456 9716 21508 9722
rect 21456 9658 21508 9664
rect 21732 9716 21784 9722
rect 21732 9658 21784 9664
rect 21272 9648 21324 9654
rect 21272 9590 21324 9596
rect 21916 9648 21968 9654
rect 21916 9590 21968 9596
rect 21180 8084 21232 8090
rect 21180 8026 21232 8032
rect 20996 7880 21048 7886
rect 20996 7822 21048 7828
rect 20904 7540 20956 7546
rect 20904 7482 20956 7488
rect 21192 7478 21220 8026
rect 21928 7886 21956 9590
rect 22008 8084 22060 8090
rect 22008 8026 22060 8032
rect 22020 7886 22048 8026
rect 22112 7886 22140 10639
rect 22204 10198 22232 10950
rect 22296 10810 22324 11070
rect 23572 11076 23624 11082
rect 23572 11018 23624 11024
rect 23112 11008 23164 11014
rect 23112 10950 23164 10956
rect 22284 10804 22336 10810
rect 22284 10746 22336 10752
rect 22192 10192 22244 10198
rect 22192 10134 22244 10140
rect 22296 9042 22324 10746
rect 23020 10464 23072 10470
rect 23020 10406 23072 10412
rect 23032 10062 23060 10406
rect 23124 10062 23152 10950
rect 26252 10826 26280 11222
rect 27172 11218 27200 12242
rect 26606 11183 26608 11192
rect 26660 11183 26662 11192
rect 27160 11212 27212 11218
rect 26608 11154 26660 11160
rect 27160 11154 27212 11160
rect 26160 10810 26280 10826
rect 26148 10804 26280 10810
rect 26200 10798 26280 10804
rect 26148 10746 26200 10752
rect 26056 10532 26108 10538
rect 26056 10474 26108 10480
rect 25410 10296 25466 10305
rect 23204 10260 23256 10266
rect 25410 10231 25412 10240
rect 23204 10202 23256 10208
rect 25464 10231 25466 10240
rect 25412 10202 25464 10208
rect 23020 10056 23072 10062
rect 23020 9998 23072 10004
rect 23112 10056 23164 10062
rect 23112 9998 23164 10004
rect 23032 9722 23060 9998
rect 23020 9716 23072 9722
rect 23020 9658 23072 9664
rect 23124 9654 23152 9998
rect 23216 9722 23244 10202
rect 25320 10056 25372 10062
rect 25320 9998 25372 10004
rect 23572 9920 23624 9926
rect 23572 9862 23624 9868
rect 24952 9920 25004 9926
rect 24952 9862 25004 9868
rect 23204 9716 23256 9722
rect 23204 9658 23256 9664
rect 23112 9648 23164 9654
rect 23112 9590 23164 9596
rect 22284 9036 22336 9042
rect 22284 8978 22336 8984
rect 22928 9036 22980 9042
rect 22928 8978 22980 8984
rect 22296 8634 22324 8978
rect 22940 8634 22968 8978
rect 22284 8628 22336 8634
rect 22284 8570 22336 8576
rect 22928 8628 22980 8634
rect 22928 8570 22980 8576
rect 21456 7880 21508 7886
rect 21456 7822 21508 7828
rect 21640 7880 21692 7886
rect 21640 7822 21692 7828
rect 21916 7880 21968 7886
rect 21916 7822 21968 7828
rect 22008 7880 22060 7886
rect 22008 7822 22060 7828
rect 22100 7880 22152 7886
rect 22100 7822 22152 7828
rect 21468 7478 21496 7822
rect 21652 7750 21680 7822
rect 21640 7744 21692 7750
rect 21640 7686 21692 7692
rect 21652 7546 21680 7686
rect 21640 7540 21692 7546
rect 21640 7482 21692 7488
rect 21928 7478 21956 7822
rect 20812 7472 20864 7478
rect 20812 7414 20864 7420
rect 21180 7472 21232 7478
rect 21180 7414 21232 7420
rect 21456 7472 21508 7478
rect 21456 7414 21508 7420
rect 21916 7472 21968 7478
rect 21916 7414 21968 7420
rect 21180 7336 21232 7342
rect 21180 7278 21232 7284
rect 19580 7100 19876 7120
rect 19636 7098 19660 7100
rect 19716 7098 19740 7100
rect 19796 7098 19820 7100
rect 19658 7046 19660 7098
rect 19722 7046 19734 7098
rect 19796 7046 19798 7098
rect 19636 7044 19660 7046
rect 19716 7044 19740 7046
rect 19796 7044 19820 7046
rect 19580 7024 19876 7044
rect 20536 6792 20588 6798
rect 20536 6734 20588 6740
rect 19984 6180 20036 6186
rect 19984 6122 20036 6128
rect 19580 6012 19876 6032
rect 19636 6010 19660 6012
rect 19716 6010 19740 6012
rect 19796 6010 19820 6012
rect 19658 5958 19660 6010
rect 19722 5958 19734 6010
rect 19796 5958 19798 6010
rect 19636 5956 19660 5958
rect 19716 5956 19740 5958
rect 19796 5956 19820 5958
rect 19580 5936 19876 5956
rect 19996 5574 20024 6122
rect 20548 5778 20576 6734
rect 21192 6730 21220 7278
rect 21928 6866 21956 7414
rect 22008 7404 22060 7410
rect 22008 7346 22060 7352
rect 22020 7188 22048 7346
rect 22112 7342 22140 7822
rect 22100 7336 22152 7342
rect 22100 7278 22152 7284
rect 22560 7336 22612 7342
rect 22560 7278 22612 7284
rect 22020 7160 22140 7188
rect 21364 6860 21416 6866
rect 21364 6802 21416 6808
rect 21916 6860 21968 6866
rect 21916 6802 21968 6808
rect 21180 6724 21232 6730
rect 21180 6666 21232 6672
rect 21376 6186 21404 6802
rect 21928 6458 21956 6802
rect 21916 6452 21968 6458
rect 21916 6394 21968 6400
rect 21364 6180 21416 6186
rect 21364 6122 21416 6128
rect 20994 5944 21050 5953
rect 20994 5879 21050 5888
rect 20904 5840 20956 5846
rect 20904 5782 20956 5788
rect 20536 5772 20588 5778
rect 20536 5714 20588 5720
rect 19984 5568 20036 5574
rect 19984 5510 20036 5516
rect 20548 5370 20576 5714
rect 20628 5568 20680 5574
rect 20680 5516 20760 5522
rect 20628 5510 20760 5516
rect 20640 5494 20760 5510
rect 20536 5364 20588 5370
rect 20536 5306 20588 5312
rect 19432 5296 19484 5302
rect 19432 5238 19484 5244
rect 19340 5024 19392 5030
rect 19340 4966 19392 4972
rect 19352 4185 19380 4966
rect 19444 4298 19472 5238
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 19580 4924 19876 4944
rect 19636 4922 19660 4924
rect 19716 4922 19740 4924
rect 19796 4922 19820 4924
rect 19658 4870 19660 4922
rect 19722 4870 19734 4922
rect 19796 4870 19798 4922
rect 19636 4868 19660 4870
rect 19716 4868 19740 4870
rect 19796 4868 19820 4870
rect 19580 4848 19876 4868
rect 19996 4865 20024 4966
rect 19982 4856 20038 4865
rect 19982 4791 20038 4800
rect 20732 4690 20760 5494
rect 19708 4684 19760 4690
rect 19708 4626 19760 4632
rect 20720 4684 20772 4690
rect 20720 4626 20772 4632
rect 19444 4270 19564 4298
rect 19338 4176 19394 4185
rect 19536 4146 19564 4270
rect 19338 4111 19394 4120
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 19524 4140 19576 4146
rect 19524 4082 19576 4088
rect 19340 4072 19392 4078
rect 19340 4014 19392 4020
rect 19352 3913 19380 4014
rect 19338 3904 19394 3913
rect 19338 3839 19394 3848
rect 19444 3738 19472 4082
rect 19720 4078 19748 4626
rect 20628 4616 20680 4622
rect 20628 4558 20680 4564
rect 20536 4480 20588 4486
rect 20536 4422 20588 4428
rect 19708 4072 19760 4078
rect 19708 4014 19760 4020
rect 20260 4072 20312 4078
rect 20260 4014 20312 4020
rect 20168 3936 20220 3942
rect 20168 3878 20220 3884
rect 19580 3836 19876 3856
rect 19636 3834 19660 3836
rect 19716 3834 19740 3836
rect 19796 3834 19820 3836
rect 19658 3782 19660 3834
rect 19722 3782 19734 3834
rect 19796 3782 19798 3834
rect 19636 3780 19660 3782
rect 19716 3780 19740 3782
rect 19796 3780 19820 3782
rect 19580 3760 19876 3780
rect 19432 3732 19484 3738
rect 19432 3674 19484 3680
rect 20076 3732 20128 3738
rect 20076 3674 20128 3680
rect 19430 3632 19486 3641
rect 19430 3567 19486 3576
rect 19246 3224 19302 3233
rect 19246 3159 19302 3168
rect 18696 3052 18748 3058
rect 18696 2994 18748 3000
rect 19444 2632 19472 3567
rect 20088 2990 20116 3674
rect 20180 3670 20208 3878
rect 20272 3738 20300 4014
rect 20260 3732 20312 3738
rect 20260 3674 20312 3680
rect 20168 3664 20220 3670
rect 20168 3606 20220 3612
rect 20548 3210 20576 4422
rect 20640 3584 20668 4558
rect 20916 4554 20944 5782
rect 21008 5642 21036 5879
rect 20996 5636 21048 5642
rect 20996 5578 21048 5584
rect 21086 5536 21142 5545
rect 21086 5471 21142 5480
rect 21100 5166 21128 5471
rect 21088 5160 21140 5166
rect 21088 5102 21140 5108
rect 21376 4622 21404 6122
rect 21548 6112 21600 6118
rect 21548 6054 21600 6060
rect 21560 5846 21588 6054
rect 22112 5914 22140 7160
rect 22100 5908 22152 5914
rect 22100 5850 22152 5856
rect 21548 5840 21600 5846
rect 21548 5782 21600 5788
rect 21560 5098 21588 5782
rect 22100 5772 22152 5778
rect 22100 5714 22152 5720
rect 21548 5092 21600 5098
rect 21548 5034 21600 5040
rect 21560 4826 21588 5034
rect 22112 4842 22140 5714
rect 22572 5710 22600 7278
rect 22940 6798 22968 8570
rect 23296 7744 23348 7750
rect 23296 7686 23348 7692
rect 22928 6792 22980 6798
rect 22928 6734 22980 6740
rect 22940 6458 22968 6734
rect 22928 6452 22980 6458
rect 22928 6394 22980 6400
rect 23112 5908 23164 5914
rect 23112 5850 23164 5856
rect 22560 5704 22612 5710
rect 22558 5672 22560 5681
rect 23020 5704 23072 5710
rect 22612 5672 22614 5681
rect 23020 5646 23072 5652
rect 22558 5607 22614 5616
rect 22744 5092 22796 5098
rect 22744 5034 22796 5040
rect 21548 4820 21600 4826
rect 21548 4762 21600 4768
rect 22020 4814 22140 4842
rect 22558 4856 22614 4865
rect 22020 4758 22048 4814
rect 22558 4791 22560 4800
rect 22612 4791 22614 4800
rect 22560 4762 22612 4768
rect 21456 4752 21508 4758
rect 21456 4694 21508 4700
rect 22008 4752 22060 4758
rect 22008 4694 22060 4700
rect 21364 4616 21416 4622
rect 21364 4558 21416 4564
rect 20720 4548 20772 4554
rect 20720 4490 20772 4496
rect 20904 4548 20956 4554
rect 20904 4490 20956 4496
rect 20732 4146 20760 4490
rect 21376 4214 21404 4558
rect 21468 4282 21496 4694
rect 21548 4616 21600 4622
rect 21548 4558 21600 4564
rect 21456 4276 21508 4282
rect 21456 4218 21508 4224
rect 21364 4208 21416 4214
rect 21364 4150 21416 4156
rect 20720 4140 20772 4146
rect 20720 4082 20772 4088
rect 20732 3738 20760 4082
rect 20812 4004 20864 4010
rect 20812 3946 20864 3952
rect 20720 3732 20772 3738
rect 20720 3674 20772 3680
rect 20720 3596 20772 3602
rect 20640 3556 20720 3584
rect 20720 3538 20772 3544
rect 20718 3496 20774 3505
rect 20824 3482 20852 3946
rect 21560 3738 21588 4558
rect 22756 4282 22784 5034
rect 23032 4826 23060 5646
rect 23124 5370 23152 5850
rect 23308 5778 23336 7686
rect 23480 7200 23532 7206
rect 23480 7142 23532 7148
rect 23296 5772 23348 5778
rect 23296 5714 23348 5720
rect 23492 5370 23520 7142
rect 23112 5364 23164 5370
rect 23112 5306 23164 5312
rect 23480 5364 23532 5370
rect 23480 5306 23532 5312
rect 23020 4820 23072 4826
rect 23020 4762 23072 4768
rect 22744 4276 22796 4282
rect 22744 4218 22796 4224
rect 23124 4185 23152 5306
rect 23584 5114 23612 9862
rect 24584 9648 24636 9654
rect 24584 9590 24636 9596
rect 24596 9110 24624 9590
rect 24676 9376 24728 9382
rect 24676 9318 24728 9324
rect 24584 9104 24636 9110
rect 24584 9046 24636 9052
rect 24688 8974 24716 9318
rect 24676 8968 24728 8974
rect 24676 8910 24728 8916
rect 24688 8430 24716 8910
rect 24676 8424 24728 8430
rect 24676 8366 24728 8372
rect 23940 8356 23992 8362
rect 23940 8298 23992 8304
rect 23848 8288 23900 8294
rect 23848 8230 23900 8236
rect 23756 6656 23808 6662
rect 23756 6598 23808 6604
rect 23768 6254 23796 6598
rect 23860 6458 23888 8230
rect 23952 7818 23980 8298
rect 24688 8090 24716 8366
rect 24964 8106 24992 9862
rect 25332 9450 25360 9998
rect 25424 9722 25452 10202
rect 26068 10198 26096 10474
rect 26620 10266 26648 11154
rect 27264 10810 27292 20198
rect 27448 13818 27476 20198
rect 29748 19378 29776 20334
rect 29932 20058 29960 20334
rect 29920 20052 29972 20058
rect 29920 19994 29972 20000
rect 30392 19854 30420 20742
rect 30944 20602 30972 21014
rect 31022 20768 31078 20777
rect 31022 20703 31078 20712
rect 30932 20596 30984 20602
rect 30932 20538 30984 20544
rect 30944 20058 30972 20538
rect 31036 20534 31064 20703
rect 31024 20528 31076 20534
rect 31024 20470 31076 20476
rect 30932 20052 30984 20058
rect 30932 19994 30984 20000
rect 29920 19848 29972 19854
rect 29920 19790 29972 19796
rect 30380 19848 30432 19854
rect 30380 19790 30432 19796
rect 29736 19372 29788 19378
rect 29736 19314 29788 19320
rect 29368 18896 29420 18902
rect 29368 18838 29420 18844
rect 29380 18086 29408 18838
rect 29748 18222 29776 19314
rect 29932 18834 29960 19790
rect 30392 19700 30420 19790
rect 30300 19672 30420 19700
rect 30196 19236 30248 19242
rect 30196 19178 30248 19184
rect 30208 18902 30236 19178
rect 30196 18896 30248 18902
rect 30196 18838 30248 18844
rect 29920 18828 29972 18834
rect 29920 18770 29972 18776
rect 29932 18426 29960 18770
rect 30104 18624 30156 18630
rect 30104 18566 30156 18572
rect 29920 18420 29972 18426
rect 29920 18362 29972 18368
rect 29736 18216 29788 18222
rect 29736 18158 29788 18164
rect 30116 18154 30144 18566
rect 30104 18148 30156 18154
rect 30104 18090 30156 18096
rect 29368 18080 29420 18086
rect 29368 18022 29420 18028
rect 29092 17740 29144 17746
rect 29092 17682 29144 17688
rect 29104 16998 29132 17682
rect 29380 17610 29408 18022
rect 30116 17746 30144 18090
rect 30208 18086 30236 18838
rect 30300 18698 30328 19672
rect 31036 19446 31064 20470
rect 31220 20058 31248 21014
rect 32496 21004 32548 21010
rect 32496 20946 32548 20952
rect 32402 20632 32458 20641
rect 32508 20618 32536 20946
rect 32864 20936 32916 20942
rect 32864 20878 32916 20884
rect 33048 20936 33100 20942
rect 33048 20878 33100 20884
rect 32772 20800 32824 20806
rect 32772 20742 32824 20748
rect 32458 20590 32536 20618
rect 32402 20567 32458 20576
rect 32416 20534 32444 20567
rect 32404 20528 32456 20534
rect 32404 20470 32456 20476
rect 31208 20052 31260 20058
rect 31208 19994 31260 20000
rect 31220 19514 31248 19994
rect 32128 19916 32180 19922
rect 32128 19858 32180 19864
rect 31208 19508 31260 19514
rect 31208 19450 31260 19456
rect 31024 19440 31076 19446
rect 31024 19382 31076 19388
rect 30288 18692 30340 18698
rect 30288 18634 30340 18640
rect 32140 18630 32168 19858
rect 32416 19417 32444 20470
rect 32784 20097 32812 20742
rect 32876 20330 32904 20878
rect 33060 20602 33088 20878
rect 33244 20602 33272 21830
rect 33520 21418 33548 21966
rect 33612 21486 33640 22102
rect 34624 22001 34652 22170
rect 34610 21992 34666 22001
rect 34610 21927 34666 21936
rect 34940 21788 35236 21808
rect 34996 21786 35020 21788
rect 35076 21786 35100 21788
rect 35156 21786 35180 21788
rect 35018 21734 35020 21786
rect 35082 21734 35094 21786
rect 35156 21734 35158 21786
rect 34996 21732 35020 21734
rect 35076 21732 35100 21734
rect 35156 21732 35180 21734
rect 34940 21712 35236 21732
rect 35820 21486 35848 22374
rect 33600 21480 33652 21486
rect 33600 21422 33652 21428
rect 35808 21480 35860 21486
rect 35808 21422 35860 21428
rect 33508 21412 33560 21418
rect 33508 21354 33560 21360
rect 33048 20596 33100 20602
rect 33048 20538 33100 20544
rect 33232 20596 33284 20602
rect 33232 20538 33284 20544
rect 33612 20330 33640 21422
rect 35532 21412 35584 21418
rect 35532 21354 35584 21360
rect 35544 21078 35572 21354
rect 35532 21072 35584 21078
rect 35532 21014 35584 21020
rect 34244 20800 34296 20806
rect 34244 20742 34296 20748
rect 32864 20324 32916 20330
rect 32864 20266 32916 20272
rect 33232 20324 33284 20330
rect 33232 20266 33284 20272
rect 33600 20324 33652 20330
rect 33600 20266 33652 20272
rect 32770 20088 32826 20097
rect 33244 20058 33272 20266
rect 33612 20058 33640 20266
rect 34256 20262 34284 20742
rect 34940 20700 35236 20720
rect 34996 20698 35020 20700
rect 35076 20698 35100 20700
rect 35156 20698 35180 20700
rect 35018 20646 35020 20698
rect 35082 20646 35094 20698
rect 35156 20646 35158 20698
rect 34996 20644 35020 20646
rect 35076 20644 35100 20646
rect 35156 20644 35180 20646
rect 34940 20624 35236 20644
rect 35622 20632 35678 20641
rect 34704 20596 34756 20602
rect 35820 20602 35848 21422
rect 35622 20567 35678 20576
rect 35808 20596 35860 20602
rect 34704 20538 34756 20544
rect 34244 20256 34296 20262
rect 34244 20198 34296 20204
rect 34520 20256 34572 20262
rect 34520 20198 34572 20204
rect 32770 20023 32826 20032
rect 33232 20052 33284 20058
rect 32784 19990 32812 20023
rect 33232 19994 33284 20000
rect 33600 20052 33652 20058
rect 33600 19994 33652 20000
rect 32772 19984 32824 19990
rect 32772 19926 32824 19932
rect 34428 19848 34480 19854
rect 34428 19790 34480 19796
rect 32402 19408 32458 19417
rect 32402 19343 32458 19352
rect 34440 19310 34468 19790
rect 32220 19304 32272 19310
rect 32220 19246 32272 19252
rect 34428 19304 34480 19310
rect 34428 19246 34480 19252
rect 31760 18624 31812 18630
rect 31760 18566 31812 18572
rect 32128 18624 32180 18630
rect 32128 18566 32180 18572
rect 30196 18080 30248 18086
rect 30196 18022 30248 18028
rect 30208 17814 30236 18022
rect 30196 17808 30248 17814
rect 30196 17750 30248 17756
rect 30564 17808 30616 17814
rect 30564 17750 30616 17756
rect 30748 17808 30800 17814
rect 30748 17750 30800 17756
rect 30104 17740 30156 17746
rect 30104 17682 30156 17688
rect 29368 17604 29420 17610
rect 29368 17546 29420 17552
rect 30576 17270 30604 17750
rect 30760 17338 30788 17750
rect 30748 17332 30800 17338
rect 30748 17274 30800 17280
rect 30564 17264 30616 17270
rect 30564 17206 30616 17212
rect 30472 17128 30524 17134
rect 30472 17070 30524 17076
rect 29092 16992 29144 16998
rect 29092 16934 29144 16940
rect 29918 16824 29974 16833
rect 29918 16759 29974 16768
rect 30378 16824 30434 16833
rect 30378 16759 30434 16768
rect 29932 16726 29960 16759
rect 29920 16720 29972 16726
rect 29920 16662 29972 16668
rect 28816 16652 28868 16658
rect 28816 16594 28868 16600
rect 30012 16652 30064 16658
rect 30012 16594 30064 16600
rect 28828 16046 28856 16594
rect 29368 16584 29420 16590
rect 29368 16526 29420 16532
rect 29000 16448 29052 16454
rect 29000 16390 29052 16396
rect 29012 16250 29040 16390
rect 29380 16250 29408 16526
rect 29000 16244 29052 16250
rect 29000 16186 29052 16192
rect 29368 16244 29420 16250
rect 29368 16186 29420 16192
rect 28816 16040 28868 16046
rect 28816 15982 28868 15988
rect 27620 15972 27672 15978
rect 27620 15914 27672 15920
rect 27632 15858 27660 15914
rect 29012 15910 29040 16186
rect 29552 15972 29604 15978
rect 29552 15914 29604 15920
rect 27540 15830 27660 15858
rect 28172 15904 28224 15910
rect 28172 15846 28224 15852
rect 28356 15904 28408 15910
rect 28356 15846 28408 15852
rect 29000 15904 29052 15910
rect 29000 15846 29052 15852
rect 27540 14550 27568 15830
rect 28184 15570 28212 15846
rect 28172 15564 28224 15570
rect 28172 15506 28224 15512
rect 28184 15162 28212 15506
rect 28172 15156 28224 15162
rect 28172 15098 28224 15104
rect 27620 14816 27672 14822
rect 27620 14758 27672 14764
rect 27528 14544 27580 14550
rect 27528 14486 27580 14492
rect 27632 13870 27660 14758
rect 28368 14618 28396 15846
rect 29012 15638 29040 15846
rect 29564 15706 29592 15914
rect 29552 15700 29604 15706
rect 29552 15642 29604 15648
rect 28632 15632 28684 15638
rect 28632 15574 28684 15580
rect 29000 15632 29052 15638
rect 29000 15574 29052 15580
rect 28644 15162 28672 15574
rect 28632 15156 28684 15162
rect 28632 15098 28684 15104
rect 28356 14612 28408 14618
rect 28356 14554 28408 14560
rect 30024 14550 30052 16594
rect 30392 16250 30420 16759
rect 30484 16454 30512 17070
rect 30564 16992 30616 16998
rect 30564 16934 30616 16940
rect 30472 16448 30524 16454
rect 30472 16390 30524 16396
rect 30484 16250 30512 16390
rect 30380 16244 30432 16250
rect 30380 16186 30432 16192
rect 30472 16244 30524 16250
rect 30472 16186 30524 16192
rect 30288 15972 30340 15978
rect 30288 15914 30340 15920
rect 30300 14822 30328 15914
rect 30576 15910 30604 16934
rect 30656 16584 30708 16590
rect 30656 16526 30708 16532
rect 30380 15904 30432 15910
rect 30380 15846 30432 15852
rect 30564 15904 30616 15910
rect 30564 15846 30616 15852
rect 30392 15162 30420 15846
rect 30668 15570 30696 16526
rect 31484 16448 31536 16454
rect 31484 16390 31536 16396
rect 31496 16114 31524 16390
rect 31772 16182 31800 18566
rect 32232 17746 32260 19246
rect 33600 19168 33652 19174
rect 33600 19110 33652 19116
rect 32220 17740 32272 17746
rect 32220 17682 32272 17688
rect 32312 17740 32364 17746
rect 32312 17682 32364 17688
rect 31944 17536 31996 17542
rect 31944 17478 31996 17484
rect 31852 17196 31904 17202
rect 31852 17138 31904 17144
rect 31864 16794 31892 17138
rect 31956 17134 31984 17478
rect 32232 17338 32260 17682
rect 32220 17332 32272 17338
rect 32220 17274 32272 17280
rect 31944 17128 31996 17134
rect 31944 17070 31996 17076
rect 31956 16794 31984 17070
rect 32324 16998 32352 17682
rect 32312 16992 32364 16998
rect 32312 16934 32364 16940
rect 31852 16788 31904 16794
rect 31852 16730 31904 16736
rect 31944 16788 31996 16794
rect 31944 16730 31996 16736
rect 32324 16658 32352 16934
rect 32128 16652 32180 16658
rect 32128 16594 32180 16600
rect 32312 16652 32364 16658
rect 32312 16594 32364 16600
rect 31760 16176 31812 16182
rect 31760 16118 31812 16124
rect 31300 16108 31352 16114
rect 31300 16050 31352 16056
rect 31484 16108 31536 16114
rect 31484 16050 31536 16056
rect 31312 15706 31340 16050
rect 31300 15700 31352 15706
rect 31300 15642 31352 15648
rect 30656 15564 30708 15570
rect 30656 15506 30708 15512
rect 31300 15564 31352 15570
rect 31300 15506 31352 15512
rect 30656 15360 30708 15366
rect 30656 15302 30708 15308
rect 30840 15360 30892 15366
rect 30840 15302 30892 15308
rect 30380 15156 30432 15162
rect 30380 15098 30432 15104
rect 30668 14958 30696 15302
rect 30656 14952 30708 14958
rect 30656 14894 30708 14900
rect 30288 14816 30340 14822
rect 30288 14758 30340 14764
rect 29368 14544 29420 14550
rect 29368 14486 29420 14492
rect 30012 14544 30064 14550
rect 30012 14486 30064 14492
rect 27988 14272 28040 14278
rect 27988 14214 28040 14220
rect 27620 13864 27672 13870
rect 27448 13790 27568 13818
rect 27620 13806 27672 13812
rect 28000 13802 28028 14214
rect 29380 14006 29408 14486
rect 29736 14476 29788 14482
rect 29736 14418 29788 14424
rect 29748 14074 29776 14418
rect 29736 14068 29788 14074
rect 29736 14010 29788 14016
rect 29368 14000 29420 14006
rect 29368 13942 29420 13948
rect 28632 13932 28684 13938
rect 28632 13874 28684 13880
rect 27436 13728 27488 13734
rect 27436 13670 27488 13676
rect 27448 13462 27476 13670
rect 27436 13456 27488 13462
rect 27436 13398 27488 13404
rect 27448 12986 27476 13398
rect 27436 12980 27488 12986
rect 27436 12922 27488 12928
rect 27540 12889 27568 13790
rect 27988 13796 28040 13802
rect 27988 13738 28040 13744
rect 28644 13734 28672 13874
rect 28632 13728 28684 13734
rect 28632 13670 28684 13676
rect 28644 13190 28672 13670
rect 29380 13530 29408 13942
rect 30300 13938 30328 14758
rect 30668 14618 30696 14894
rect 30852 14890 30880 15302
rect 31312 15162 31340 15506
rect 31772 15162 31800 16118
rect 32140 15910 32168 16594
rect 32324 16250 32352 16594
rect 32312 16244 32364 16250
rect 32312 16186 32364 16192
rect 33508 16176 33560 16182
rect 33508 16118 33560 16124
rect 32128 15904 32180 15910
rect 32128 15846 32180 15852
rect 32956 15904 33008 15910
rect 32956 15846 33008 15852
rect 32312 15360 32364 15366
rect 32312 15302 32364 15308
rect 31300 15156 31352 15162
rect 31300 15098 31352 15104
rect 31760 15156 31812 15162
rect 31760 15098 31812 15104
rect 32324 15026 32352 15302
rect 32312 15020 32364 15026
rect 32312 14962 32364 14968
rect 31944 14952 31996 14958
rect 31944 14894 31996 14900
rect 30840 14884 30892 14890
rect 30840 14826 30892 14832
rect 31668 14816 31720 14822
rect 31668 14758 31720 14764
rect 31680 14618 31708 14758
rect 31956 14618 31984 14894
rect 32324 14618 32352 14962
rect 30656 14612 30708 14618
rect 30656 14554 30708 14560
rect 31668 14612 31720 14618
rect 31668 14554 31720 14560
rect 31944 14612 31996 14618
rect 31944 14554 31996 14560
rect 32312 14612 32364 14618
rect 32312 14554 32364 14560
rect 30932 14476 30984 14482
rect 30932 14418 30984 14424
rect 32128 14476 32180 14482
rect 32128 14418 32180 14424
rect 30944 14074 30972 14418
rect 31576 14272 31628 14278
rect 31576 14214 31628 14220
rect 30932 14068 30984 14074
rect 30932 14010 30984 14016
rect 30288 13932 30340 13938
rect 30288 13874 30340 13880
rect 30300 13841 30328 13874
rect 31588 13870 31616 14214
rect 32140 13870 32168 14418
rect 32312 14340 32364 14346
rect 32312 14282 32364 14288
rect 32324 13938 32352 14282
rect 32312 13932 32364 13938
rect 32312 13874 32364 13880
rect 32864 13932 32916 13938
rect 32864 13874 32916 13880
rect 31576 13864 31628 13870
rect 30286 13832 30342 13841
rect 32128 13864 32180 13870
rect 31576 13806 31628 13812
rect 31758 13832 31814 13841
rect 30286 13767 30342 13776
rect 31024 13796 31076 13802
rect 31758 13767 31814 13776
rect 32048 13812 32128 13818
rect 32048 13806 32180 13812
rect 32048 13790 32168 13806
rect 31024 13738 31076 13744
rect 29920 13728 29972 13734
rect 29920 13670 29972 13676
rect 29368 13524 29420 13530
rect 29368 13466 29420 13472
rect 29932 13462 29960 13670
rect 31036 13530 31064 13738
rect 31024 13524 31076 13530
rect 31024 13466 31076 13472
rect 29920 13456 29972 13462
rect 29920 13398 29972 13404
rect 29644 13320 29696 13326
rect 29644 13262 29696 13268
rect 28632 13184 28684 13190
rect 28632 13126 28684 13132
rect 27526 12880 27582 12889
rect 27526 12815 27582 12824
rect 28644 12306 28672 13126
rect 29656 12646 29684 13262
rect 29932 12986 29960 13398
rect 29920 12980 29972 12986
rect 29920 12922 29972 12928
rect 29644 12640 29696 12646
rect 29644 12582 29696 12588
rect 29656 12374 29684 12582
rect 29932 12442 29960 12922
rect 31772 12918 31800 13767
rect 31760 12912 31812 12918
rect 31760 12854 31812 12860
rect 31024 12640 31076 12646
rect 31022 12608 31024 12617
rect 31076 12608 31078 12617
rect 31022 12543 31078 12552
rect 31772 12458 31800 12854
rect 31680 12442 31800 12458
rect 29920 12436 29972 12442
rect 29920 12378 29972 12384
rect 31668 12436 31800 12442
rect 31720 12430 31800 12436
rect 31668 12378 31720 12384
rect 29644 12368 29696 12374
rect 29644 12310 29696 12316
rect 28356 12300 28408 12306
rect 28356 12242 28408 12248
rect 28632 12300 28684 12306
rect 28632 12242 28684 12248
rect 28368 11898 28396 12242
rect 28644 11898 28672 12242
rect 29656 11937 29684 12310
rect 29642 11928 29698 11937
rect 28356 11892 28408 11898
rect 28356 11834 28408 11840
rect 28632 11892 28684 11898
rect 29642 11863 29698 11872
rect 28632 11834 28684 11840
rect 27528 11280 27580 11286
rect 27528 11222 27580 11228
rect 27252 10804 27304 10810
rect 27252 10746 27304 10752
rect 27264 10713 27292 10746
rect 27250 10704 27306 10713
rect 27250 10639 27306 10648
rect 26608 10260 26660 10266
rect 26608 10202 26660 10208
rect 27540 10198 27568 11222
rect 28368 11218 28396 11834
rect 28356 11212 28408 11218
rect 28356 11154 28408 11160
rect 29644 11212 29696 11218
rect 29644 11154 29696 11160
rect 27988 11076 28040 11082
rect 27988 11018 28040 11024
rect 28000 10305 28028 11018
rect 28368 10674 28396 11154
rect 29656 10810 29684 11154
rect 30472 11076 30524 11082
rect 30472 11018 30524 11024
rect 29644 10804 29696 10810
rect 29644 10746 29696 10752
rect 28356 10668 28408 10674
rect 28356 10610 28408 10616
rect 29276 10668 29328 10674
rect 29276 10610 29328 10616
rect 27986 10296 28042 10305
rect 28814 10296 28870 10305
rect 27986 10231 28042 10240
rect 28724 10260 28776 10266
rect 28814 10231 28870 10240
rect 28724 10202 28776 10208
rect 26056 10192 26108 10198
rect 26054 10160 26056 10169
rect 27528 10192 27580 10198
rect 26108 10160 26110 10169
rect 27528 10134 27580 10140
rect 26054 10095 26110 10104
rect 25504 10056 25556 10062
rect 25502 10024 25504 10033
rect 25556 10024 25558 10033
rect 25502 9959 25558 9968
rect 27158 10024 27214 10033
rect 27158 9959 27214 9968
rect 25412 9716 25464 9722
rect 25412 9658 25464 9664
rect 27172 9654 27200 9959
rect 28540 9920 28592 9926
rect 28540 9862 28592 9868
rect 28552 9722 28580 9862
rect 28736 9722 28764 10202
rect 28828 10198 28856 10231
rect 28816 10192 28868 10198
rect 28816 10134 28868 10140
rect 28828 9722 28856 10134
rect 29000 10056 29052 10062
rect 29000 9998 29052 10004
rect 27804 9716 27856 9722
rect 27804 9658 27856 9664
rect 28540 9716 28592 9722
rect 28540 9658 28592 9664
rect 28724 9716 28776 9722
rect 28724 9658 28776 9664
rect 28816 9716 28868 9722
rect 28816 9658 28868 9664
rect 27160 9648 27212 9654
rect 27160 9590 27212 9596
rect 25320 9444 25372 9450
rect 25320 9386 25372 9392
rect 26056 9444 26108 9450
rect 26056 9386 26108 9392
rect 26068 9178 26096 9386
rect 26608 9376 26660 9382
rect 26608 9318 26660 9324
rect 26620 9178 26648 9318
rect 26056 9172 26108 9178
rect 26608 9172 26660 9178
rect 26056 9114 26108 9120
rect 26528 9132 26608 9160
rect 26240 8832 26292 8838
rect 26240 8774 26292 8780
rect 26252 8106 26280 8774
rect 26528 8362 26556 9132
rect 26608 9114 26660 9120
rect 27172 9110 27200 9590
rect 27816 9110 27844 9658
rect 27896 9376 27948 9382
rect 27896 9318 27948 9324
rect 28264 9376 28316 9382
rect 28264 9318 28316 9324
rect 27160 9104 27212 9110
rect 27160 9046 27212 9052
rect 27804 9104 27856 9110
rect 27804 9046 27856 9052
rect 27068 8968 27120 8974
rect 27068 8910 27120 8916
rect 27080 8634 27108 8910
rect 27068 8628 27120 8634
rect 27068 8570 27120 8576
rect 26516 8356 26568 8362
rect 26516 8298 26568 8304
rect 24872 8090 24992 8106
rect 24676 8084 24728 8090
rect 24676 8026 24728 8032
rect 24872 8084 25004 8090
rect 24872 8078 24952 8084
rect 24584 7880 24636 7886
rect 24584 7822 24636 7828
rect 23940 7812 23992 7818
rect 23940 7754 23992 7760
rect 24596 7546 24624 7822
rect 24768 7812 24820 7818
rect 24768 7754 24820 7760
rect 24584 7540 24636 7546
rect 24584 7482 24636 7488
rect 23940 6792 23992 6798
rect 23940 6734 23992 6740
rect 23848 6452 23900 6458
rect 23848 6394 23900 6400
rect 23756 6248 23808 6254
rect 23492 5086 23612 5114
rect 23676 6208 23756 6236
rect 23676 5098 23704 6208
rect 23756 6190 23808 6196
rect 23860 5545 23888 6394
rect 23846 5536 23902 5545
rect 23846 5471 23902 5480
rect 23754 5400 23810 5409
rect 23754 5335 23756 5344
rect 23808 5335 23810 5344
rect 23756 5306 23808 5312
rect 23664 5092 23716 5098
rect 23388 4752 23440 4758
rect 23388 4694 23440 4700
rect 23400 4282 23428 4694
rect 23492 4434 23520 5086
rect 23664 5034 23716 5040
rect 23572 5024 23624 5030
rect 23572 4966 23624 4972
rect 23584 4554 23612 4966
rect 23676 4758 23704 5034
rect 23756 4820 23808 4826
rect 23756 4762 23808 4768
rect 23664 4752 23716 4758
rect 23664 4694 23716 4700
rect 23572 4548 23624 4554
rect 23572 4490 23624 4496
rect 23492 4406 23612 4434
rect 23388 4276 23440 4282
rect 23388 4218 23440 4224
rect 23110 4176 23166 4185
rect 23110 4111 23166 4120
rect 23584 4078 23612 4406
rect 23572 4072 23624 4078
rect 23572 4014 23624 4020
rect 23112 3936 23164 3942
rect 23110 3904 23112 3913
rect 23164 3904 23166 3913
rect 23110 3839 23166 3848
rect 21548 3732 21600 3738
rect 21548 3674 21600 3680
rect 22100 3596 22152 3602
rect 22100 3538 22152 3544
rect 22376 3596 22428 3602
rect 22376 3538 22428 3544
rect 23480 3596 23532 3602
rect 23480 3538 23532 3544
rect 20774 3454 20852 3482
rect 20718 3431 20720 3440
rect 20772 3431 20774 3440
rect 20720 3402 20772 3408
rect 20548 3194 20760 3210
rect 20548 3188 20772 3194
rect 20548 3182 20720 3188
rect 20720 3130 20772 3136
rect 22112 3126 22140 3538
rect 22190 3360 22246 3369
rect 22190 3295 22246 3304
rect 22100 3120 22152 3126
rect 22100 3062 22152 3068
rect 20076 2984 20128 2990
rect 20076 2926 20128 2932
rect 19580 2748 19876 2768
rect 19636 2746 19660 2748
rect 19716 2746 19740 2748
rect 19796 2746 19820 2748
rect 19658 2694 19660 2746
rect 19722 2694 19734 2746
rect 19796 2694 19798 2746
rect 19636 2692 19660 2694
rect 19716 2692 19740 2694
rect 19796 2692 19820 2694
rect 19580 2672 19876 2692
rect 20088 2650 20116 2926
rect 20720 2916 20772 2922
rect 20720 2858 20772 2864
rect 20076 2644 20128 2650
rect 19444 2604 19564 2632
rect 19536 480 19564 2604
rect 20076 2586 20128 2592
rect 20732 2582 20760 2858
rect 21180 2848 21232 2854
rect 20902 2816 20958 2825
rect 21180 2790 21232 2796
rect 20902 2751 20958 2760
rect 20720 2576 20772 2582
rect 20720 2518 20772 2524
rect 20916 480 20944 2751
rect 21192 2650 21220 2790
rect 21180 2644 21232 2650
rect 21180 2586 21232 2592
rect 22204 480 22232 3295
rect 22388 3194 22416 3538
rect 22836 3528 22888 3534
rect 22836 3470 22888 3476
rect 22376 3188 22428 3194
rect 22376 3130 22428 3136
rect 22282 2952 22338 2961
rect 22282 2887 22284 2896
rect 22336 2887 22338 2896
rect 22284 2858 22336 2864
rect 22848 2650 22876 3470
rect 23492 3398 23520 3538
rect 23480 3392 23532 3398
rect 23480 3334 23532 3340
rect 23492 2650 23520 3334
rect 22836 2644 22888 2650
rect 22836 2586 22888 2592
rect 23480 2644 23532 2650
rect 23480 2586 23532 2592
rect 23584 480 23612 4014
rect 23768 3913 23796 4762
rect 23754 3904 23810 3913
rect 23754 3839 23810 3848
rect 23860 3618 23888 5471
rect 23952 3670 23980 6734
rect 24780 6440 24808 7754
rect 24872 7546 24900 8078
rect 24952 8026 25004 8032
rect 26160 8078 26280 8106
rect 26528 8090 26556 8298
rect 26608 8288 26660 8294
rect 26608 8230 26660 8236
rect 26516 8084 26568 8090
rect 24952 7948 25004 7954
rect 24952 7890 25004 7896
rect 24860 7540 24912 7546
rect 24860 7482 24912 7488
rect 24964 6866 24992 7890
rect 26160 7886 26188 8078
rect 26516 8026 26568 8032
rect 26620 7954 26648 8230
rect 27080 8022 27108 8570
rect 27068 8016 27120 8022
rect 27068 7958 27120 7964
rect 26608 7948 26660 7954
rect 26608 7890 26660 7896
rect 26148 7880 26200 7886
rect 26148 7822 26200 7828
rect 25320 7744 25372 7750
rect 25320 7686 25372 7692
rect 25332 7342 25360 7686
rect 25320 7336 25372 7342
rect 25320 7278 25372 7284
rect 26620 7206 26648 7890
rect 27080 7546 27108 7958
rect 27068 7540 27120 7546
rect 27068 7482 27120 7488
rect 25504 7200 25556 7206
rect 25504 7142 25556 7148
rect 26608 7200 26660 7206
rect 26608 7142 26660 7148
rect 24952 6860 25004 6866
rect 24952 6802 25004 6808
rect 24860 6452 24912 6458
rect 24780 6412 24860 6440
rect 24032 5568 24084 5574
rect 24032 5510 24084 5516
rect 24044 4826 24072 5510
rect 24780 5234 24808 6412
rect 24860 6394 24912 6400
rect 24216 5228 24268 5234
rect 24216 5170 24268 5176
rect 24768 5228 24820 5234
rect 24768 5170 24820 5176
rect 24228 4826 24256 5170
rect 24964 4826 24992 6802
rect 25516 6458 25544 7142
rect 26240 6656 26292 6662
rect 26160 6604 26240 6610
rect 26160 6598 26292 6604
rect 26516 6656 26568 6662
rect 26516 6598 26568 6604
rect 26160 6582 26280 6598
rect 25504 6452 25556 6458
rect 25504 6394 25556 6400
rect 26160 6202 26188 6582
rect 26424 6452 26476 6458
rect 26424 6394 26476 6400
rect 26240 6384 26292 6390
rect 26238 6352 26240 6361
rect 26292 6352 26294 6361
rect 26238 6287 26294 6296
rect 26240 6248 26292 6254
rect 26160 6196 26240 6202
rect 26160 6190 26292 6196
rect 26160 6174 26280 6190
rect 25594 5672 25650 5681
rect 25594 5607 25650 5616
rect 24032 4820 24084 4826
rect 24032 4762 24084 4768
rect 24216 4820 24268 4826
rect 24216 4762 24268 4768
rect 24952 4820 25004 4826
rect 24952 4762 25004 4768
rect 24584 4684 24636 4690
rect 24584 4626 24636 4632
rect 24400 4480 24452 4486
rect 24400 4422 24452 4428
rect 24412 3738 24440 4422
rect 24596 3942 24624 4626
rect 25608 4622 25636 5607
rect 25964 5296 26016 5302
rect 25964 5238 26016 5244
rect 25976 5030 26004 5238
rect 25964 5024 26016 5030
rect 25964 4966 26016 4972
rect 26056 5024 26108 5030
rect 26056 4966 26108 4972
rect 25596 4616 25648 4622
rect 25594 4584 25596 4593
rect 25648 4584 25650 4593
rect 25594 4519 25650 4528
rect 25872 4480 25924 4486
rect 25872 4422 25924 4428
rect 25884 4282 25912 4422
rect 25872 4276 25924 4282
rect 25872 4218 25924 4224
rect 25976 4146 26004 4966
rect 26068 4826 26096 4966
rect 26056 4820 26108 4826
rect 26056 4762 26108 4768
rect 26054 4176 26110 4185
rect 25964 4140 26016 4146
rect 26054 4111 26110 4120
rect 25964 4082 26016 4088
rect 24768 4072 24820 4078
rect 24766 4040 24768 4049
rect 24820 4040 24822 4049
rect 25686 4040 25742 4049
rect 24766 3975 24822 3984
rect 24952 4004 25004 4010
rect 25686 3975 25742 3984
rect 24952 3946 25004 3952
rect 24584 3936 24636 3942
rect 24584 3878 24636 3884
rect 24400 3732 24452 3738
rect 24400 3674 24452 3680
rect 23676 3590 23888 3618
rect 23940 3664 23992 3670
rect 24596 3641 24624 3878
rect 23940 3606 23992 3612
rect 24582 3632 24638 3641
rect 23676 3194 23704 3590
rect 24582 3567 24638 3576
rect 23756 3528 23808 3534
rect 23756 3470 23808 3476
rect 23846 3496 23902 3505
rect 23664 3188 23716 3194
rect 23664 3130 23716 3136
rect 23676 2650 23704 3130
rect 23768 2990 23796 3470
rect 23846 3431 23848 3440
rect 23900 3431 23902 3440
rect 23848 3402 23900 3408
rect 24860 3392 24912 3398
rect 24860 3334 24912 3340
rect 24872 2990 24900 3334
rect 23756 2984 23808 2990
rect 23756 2926 23808 2932
rect 24860 2984 24912 2990
rect 24860 2926 24912 2932
rect 24768 2848 24820 2854
rect 24768 2790 24820 2796
rect 23664 2644 23716 2650
rect 23664 2586 23716 2592
rect 23676 2514 23704 2586
rect 24780 2582 24808 2790
rect 24768 2576 24820 2582
rect 24768 2518 24820 2524
rect 23664 2508 23716 2514
rect 23664 2450 23716 2456
rect 24964 480 24992 3946
rect 25596 3596 25648 3602
rect 25596 3538 25648 3544
rect 25608 2854 25636 3538
rect 25596 2848 25648 2854
rect 25594 2816 25596 2825
rect 25648 2816 25650 2825
rect 25594 2751 25650 2760
rect 25700 2650 25728 3975
rect 26068 3194 26096 4111
rect 26160 3738 26188 6174
rect 26436 5778 26464 6394
rect 26528 6186 26556 6598
rect 26620 6458 26648 7142
rect 27172 6882 27200 9046
rect 27908 8906 27936 9318
rect 28080 9104 28132 9110
rect 28080 9046 28132 9052
rect 27896 8900 27948 8906
rect 27896 8842 27948 8848
rect 28092 8634 28120 9046
rect 28172 8968 28224 8974
rect 28172 8910 28224 8916
rect 28080 8628 28132 8634
rect 28080 8570 28132 8576
rect 28184 8090 28212 8910
rect 28172 8084 28224 8090
rect 28172 8026 28224 8032
rect 27620 7744 27672 7750
rect 27620 7686 27672 7692
rect 27632 7018 27660 7686
rect 27712 7472 27764 7478
rect 27710 7440 27712 7449
rect 27764 7440 27766 7449
rect 28276 7410 28304 9318
rect 29012 9042 29040 9998
rect 29288 9722 29316 10610
rect 29552 10532 29604 10538
rect 29552 10474 29604 10480
rect 29564 9926 29592 10474
rect 29656 10266 29684 10746
rect 30484 10305 30512 11018
rect 30470 10296 30526 10305
rect 29644 10260 29696 10266
rect 30470 10231 30526 10240
rect 29644 10202 29696 10208
rect 29552 9920 29604 9926
rect 29552 9862 29604 9868
rect 30012 9920 30064 9926
rect 30012 9862 30064 9868
rect 29276 9716 29328 9722
rect 29276 9658 29328 9664
rect 30024 9382 30052 9862
rect 30104 9580 30156 9586
rect 30104 9522 30156 9528
rect 30012 9376 30064 9382
rect 30012 9318 30064 9324
rect 29552 9172 29604 9178
rect 29552 9114 29604 9120
rect 29092 9104 29144 9110
rect 29092 9046 29144 9052
rect 29000 9036 29052 9042
rect 29000 8978 29052 8984
rect 29104 8566 29132 9046
rect 29184 8832 29236 8838
rect 29184 8774 29236 8780
rect 29196 8634 29224 8774
rect 29564 8634 29592 9114
rect 30024 9110 30052 9318
rect 30012 9104 30064 9110
rect 30012 9046 30064 9052
rect 30116 8974 30144 9522
rect 30380 9444 30432 9450
rect 30380 9386 30432 9392
rect 30392 9178 30420 9386
rect 30380 9172 30432 9178
rect 30380 9114 30432 9120
rect 30196 9036 30248 9042
rect 30196 8978 30248 8984
rect 30840 9036 30892 9042
rect 30840 8978 30892 8984
rect 31852 9036 31904 9042
rect 31852 8978 31904 8984
rect 30104 8968 30156 8974
rect 30104 8910 30156 8916
rect 29184 8628 29236 8634
rect 29184 8570 29236 8576
rect 29552 8628 29604 8634
rect 29552 8570 29604 8576
rect 29092 8560 29144 8566
rect 29092 8502 29144 8508
rect 29368 8560 29420 8566
rect 29368 8502 29420 8508
rect 28448 8084 28500 8090
rect 28448 8026 28500 8032
rect 27710 7375 27766 7384
rect 28264 7404 28316 7410
rect 28264 7346 28316 7352
rect 28170 7304 28226 7313
rect 28170 7239 28226 7248
rect 28264 7268 28316 7274
rect 28184 7206 28212 7239
rect 28264 7210 28316 7216
rect 28172 7200 28224 7206
rect 28172 7142 28224 7148
rect 26884 6860 26936 6866
rect 26884 6802 26936 6808
rect 26988 6854 27200 6882
rect 27540 6990 27660 7018
rect 26608 6452 26660 6458
rect 26608 6394 26660 6400
rect 26516 6180 26568 6186
rect 26516 6122 26568 6128
rect 26528 5914 26556 6122
rect 26896 6118 26924 6802
rect 26884 6112 26936 6118
rect 26884 6054 26936 6060
rect 26516 5908 26568 5914
rect 26516 5850 26568 5856
rect 26608 5840 26660 5846
rect 26608 5782 26660 5788
rect 26424 5772 26476 5778
rect 26424 5714 26476 5720
rect 26620 5302 26648 5782
rect 26896 5370 26924 6054
rect 26884 5364 26936 5370
rect 26884 5306 26936 5312
rect 26608 5296 26660 5302
rect 26608 5238 26660 5244
rect 26608 5160 26660 5166
rect 26608 5102 26660 5108
rect 26514 4584 26570 4593
rect 26620 4554 26648 5102
rect 26988 4690 27016 6854
rect 27540 5846 27568 6990
rect 28276 6934 28304 7210
rect 28460 6934 28488 8026
rect 29380 8022 29408 8502
rect 29368 8016 29420 8022
rect 29368 7958 29420 7964
rect 29552 8016 29604 8022
rect 29552 7958 29604 7964
rect 29564 7546 29592 7958
rect 29552 7540 29604 7546
rect 29552 7482 29604 7488
rect 30208 7410 30236 8978
rect 30748 8832 30800 8838
rect 30748 8774 30800 8780
rect 30760 8498 30788 8774
rect 30852 8498 30880 8978
rect 31576 8968 31628 8974
rect 31576 8910 31628 8916
rect 31588 8634 31616 8910
rect 31576 8628 31628 8634
rect 31576 8570 31628 8576
rect 31864 8616 31892 8978
rect 31944 8628 31996 8634
rect 31864 8588 31944 8616
rect 30748 8492 30800 8498
rect 30748 8434 30800 8440
rect 30840 8492 30892 8498
rect 30840 8434 30892 8440
rect 30760 8362 30788 8434
rect 30748 8356 30800 8362
rect 30748 8298 30800 8304
rect 30288 8288 30340 8294
rect 30288 8230 30340 8236
rect 30300 8090 30328 8230
rect 31588 8090 31616 8570
rect 31864 8362 31892 8588
rect 31944 8570 31996 8576
rect 31852 8356 31904 8362
rect 31852 8298 31904 8304
rect 31864 8090 31892 8298
rect 30288 8084 30340 8090
rect 30288 8026 30340 8032
rect 31576 8084 31628 8090
rect 31576 8026 31628 8032
rect 31852 8084 31904 8090
rect 31852 8026 31904 8032
rect 30656 7812 30708 7818
rect 30656 7754 30708 7760
rect 29644 7404 29696 7410
rect 29644 7346 29696 7352
rect 30196 7404 30248 7410
rect 30196 7346 30248 7352
rect 28264 6928 28316 6934
rect 28264 6870 28316 6876
rect 28448 6928 28500 6934
rect 28448 6870 28500 6876
rect 29184 6928 29236 6934
rect 29184 6870 29236 6876
rect 27620 6860 27672 6866
rect 27620 6802 27672 6808
rect 27632 6186 27660 6802
rect 27712 6792 27764 6798
rect 27712 6734 27764 6740
rect 27724 6458 27752 6734
rect 27712 6452 27764 6458
rect 27712 6394 27764 6400
rect 27620 6180 27672 6186
rect 27620 6122 27672 6128
rect 27068 5840 27120 5846
rect 27068 5782 27120 5788
rect 27528 5840 27580 5846
rect 27528 5782 27580 5788
rect 27080 4758 27108 5782
rect 27160 5772 27212 5778
rect 27160 5714 27212 5720
rect 27172 5370 27200 5714
rect 27632 5574 27660 6122
rect 27620 5568 27672 5574
rect 27540 5516 27620 5522
rect 27540 5510 27672 5516
rect 27540 5494 27660 5510
rect 27160 5364 27212 5370
rect 27160 5306 27212 5312
rect 27540 4826 27568 5494
rect 28460 5370 28488 6870
rect 29092 6656 29144 6662
rect 29092 6598 29144 6604
rect 29000 6180 29052 6186
rect 29000 6122 29052 6128
rect 29012 5778 29040 6122
rect 29104 5846 29132 6598
rect 29196 6458 29224 6870
rect 29184 6452 29236 6458
rect 29184 6394 29236 6400
rect 29656 6118 29684 7346
rect 29736 7336 29788 7342
rect 29736 7278 29788 7284
rect 29748 7002 29776 7278
rect 30472 7200 30524 7206
rect 30472 7142 30524 7148
rect 29736 6996 29788 7002
rect 29736 6938 29788 6944
rect 30484 6746 30512 7142
rect 30668 7002 30696 7754
rect 30748 7744 30800 7750
rect 30748 7686 30800 7692
rect 30760 7313 30788 7686
rect 31588 7562 31616 8026
rect 31496 7546 31616 7562
rect 31484 7540 31616 7546
rect 31536 7534 31616 7540
rect 31484 7482 31536 7488
rect 30746 7304 30802 7313
rect 30746 7239 30802 7248
rect 31208 7268 31260 7274
rect 31208 7210 31260 7216
rect 30656 6996 30708 7002
rect 30656 6938 30708 6944
rect 30484 6718 30604 6746
rect 30576 6662 30604 6718
rect 31220 6662 31248 7210
rect 30564 6656 30616 6662
rect 30564 6598 30616 6604
rect 31208 6656 31260 6662
rect 31208 6598 31260 6604
rect 30576 6186 30604 6598
rect 31220 6458 31248 6598
rect 31208 6452 31260 6458
rect 31208 6394 31260 6400
rect 30564 6180 30616 6186
rect 30564 6122 30616 6128
rect 29644 6112 29696 6118
rect 29644 6054 29696 6060
rect 29920 6112 29972 6118
rect 29920 6054 29972 6060
rect 29092 5840 29144 5846
rect 29092 5782 29144 5788
rect 29000 5772 29052 5778
rect 29000 5714 29052 5720
rect 28448 5364 28500 5370
rect 28448 5306 28500 5312
rect 29012 5234 29040 5714
rect 29104 5370 29132 5782
rect 29274 5400 29330 5409
rect 29092 5364 29144 5370
rect 29274 5335 29330 5344
rect 29092 5306 29144 5312
rect 29000 5228 29052 5234
rect 29000 5170 29052 5176
rect 27528 4820 27580 4826
rect 27528 4762 27580 4768
rect 27068 4752 27120 4758
rect 27068 4694 27120 4700
rect 26976 4684 27028 4690
rect 26976 4626 27028 4632
rect 29012 4622 29040 5170
rect 29104 5030 29132 5306
rect 29092 5024 29144 5030
rect 29092 4966 29144 4972
rect 29000 4616 29052 4622
rect 29000 4558 29052 4564
rect 26514 4519 26570 4528
rect 26608 4548 26660 4554
rect 26240 4004 26292 4010
rect 26240 3946 26292 3952
rect 26252 3738 26280 3946
rect 26332 3936 26384 3942
rect 26332 3878 26384 3884
rect 26422 3904 26478 3913
rect 26148 3732 26200 3738
rect 26148 3674 26200 3680
rect 26240 3732 26292 3738
rect 26240 3674 26292 3680
rect 26344 3670 26372 3878
rect 26422 3839 26478 3848
rect 26332 3664 26384 3670
rect 26332 3606 26384 3612
rect 26238 3224 26294 3233
rect 26056 3188 26108 3194
rect 26238 3159 26294 3168
rect 26056 3130 26108 3136
rect 26068 2854 26096 3130
rect 26056 2848 26108 2854
rect 26056 2790 26108 2796
rect 25688 2644 25740 2650
rect 25688 2586 25740 2592
rect 26252 480 26280 3159
rect 26344 2650 26372 3606
rect 26436 3534 26464 3839
rect 26424 3528 26476 3534
rect 26424 3470 26476 3476
rect 26436 3058 26464 3470
rect 26528 3194 26556 4519
rect 26608 4490 26660 4496
rect 27712 4480 27764 4486
rect 27712 4422 27764 4428
rect 28356 4480 28408 4486
rect 28356 4422 28408 4428
rect 27724 4146 27752 4422
rect 27712 4140 27764 4146
rect 27712 4082 27764 4088
rect 27724 4049 27752 4082
rect 27710 4040 27766 4049
rect 27620 4004 27672 4010
rect 27710 3975 27766 3984
rect 27620 3946 27672 3952
rect 26608 3936 26660 3942
rect 26608 3878 26660 3884
rect 26620 3466 26648 3878
rect 26976 3732 27028 3738
rect 26976 3674 27028 3680
rect 26608 3460 26660 3466
rect 26608 3402 26660 3408
rect 26516 3188 26568 3194
rect 26516 3130 26568 3136
rect 26620 3058 26648 3402
rect 26790 3088 26846 3097
rect 26424 3052 26476 3058
rect 26424 2994 26476 3000
rect 26608 3052 26660 3058
rect 26790 3023 26846 3032
rect 26608 2994 26660 3000
rect 26804 2854 26832 3023
rect 26792 2848 26844 2854
rect 26792 2790 26844 2796
rect 26332 2644 26384 2650
rect 26332 2586 26384 2592
rect 26988 2378 27016 3674
rect 27632 3505 27660 3946
rect 28080 3936 28132 3942
rect 28078 3904 28080 3913
rect 28172 3936 28224 3942
rect 28132 3904 28134 3913
rect 28172 3878 28224 3884
rect 28078 3839 28134 3848
rect 28184 3641 28212 3878
rect 28170 3632 28226 3641
rect 27712 3596 27764 3602
rect 28368 3602 28396 4422
rect 29012 4282 29040 4558
rect 29000 4276 29052 4282
rect 29000 4218 29052 4224
rect 29012 4162 29040 4218
rect 28920 4134 29040 4162
rect 28632 3936 28684 3942
rect 28632 3878 28684 3884
rect 28644 3670 28672 3878
rect 28632 3664 28684 3670
rect 28632 3606 28684 3612
rect 28170 3567 28226 3576
rect 28356 3596 28408 3602
rect 27712 3538 27764 3544
rect 27618 3496 27674 3505
rect 27618 3431 27620 3440
rect 27672 3431 27674 3440
rect 27620 3402 27672 3408
rect 27252 2984 27304 2990
rect 27252 2926 27304 2932
rect 27264 2582 27292 2926
rect 27632 2582 27660 3402
rect 27252 2576 27304 2582
rect 27252 2518 27304 2524
rect 27620 2576 27672 2582
rect 27620 2518 27672 2524
rect 27724 2514 27752 3538
rect 28184 3194 28212 3567
rect 28356 3538 28408 3544
rect 28816 3392 28868 3398
rect 28920 3346 28948 4134
rect 29288 4078 29316 5335
rect 29932 5234 29960 6054
rect 29920 5228 29972 5234
rect 29920 5170 29972 5176
rect 30576 4826 30604 6122
rect 30930 5944 30986 5953
rect 30930 5879 30986 5888
rect 30748 5568 30800 5574
rect 30748 5510 30800 5516
rect 30760 5098 30788 5510
rect 30748 5092 30800 5098
rect 30748 5034 30800 5040
rect 30564 4820 30616 4826
rect 30564 4762 30616 4768
rect 29460 4684 29512 4690
rect 29460 4626 29512 4632
rect 29000 4072 29052 4078
rect 29000 4014 29052 4020
rect 29276 4072 29328 4078
rect 29276 4014 29328 4020
rect 28868 3340 28948 3346
rect 28816 3334 28948 3340
rect 28828 3318 28948 3334
rect 28446 3224 28502 3233
rect 28172 3188 28224 3194
rect 28920 3194 28948 3318
rect 28446 3159 28502 3168
rect 28908 3188 28960 3194
rect 28172 3130 28224 3136
rect 28460 2514 28488 3159
rect 28908 3130 28960 3136
rect 27712 2508 27764 2514
rect 27712 2450 27764 2456
rect 28448 2508 28500 2514
rect 28448 2450 28500 2456
rect 26976 2372 27028 2378
rect 26976 2314 27028 2320
rect 27620 2372 27672 2378
rect 27620 2314 27672 2320
rect 27632 480 27660 2314
rect 29012 480 29040 4014
rect 29472 3738 29500 4626
rect 29552 4140 29604 4146
rect 29552 4082 29604 4088
rect 29460 3732 29512 3738
rect 29460 3674 29512 3680
rect 29092 3596 29144 3602
rect 29092 3538 29144 3544
rect 29104 3126 29132 3538
rect 29564 3194 29592 4082
rect 30380 4072 30432 4078
rect 30380 4014 30432 4020
rect 30288 4004 30340 4010
rect 30288 3946 30340 3952
rect 29368 3188 29420 3194
rect 29368 3130 29420 3136
rect 29552 3188 29604 3194
rect 29552 3130 29604 3136
rect 29092 3120 29144 3126
rect 29090 3088 29092 3097
rect 29144 3088 29146 3097
rect 29090 3023 29146 3032
rect 29380 2922 29408 3130
rect 29368 2916 29420 2922
rect 29368 2858 29420 2864
rect 29380 2650 29408 2858
rect 29368 2644 29420 2650
rect 29368 2586 29420 2592
rect 29564 2582 29592 3130
rect 30196 3120 30248 3126
rect 30196 3062 30248 3068
rect 30208 2961 30236 3062
rect 30194 2952 30250 2961
rect 30194 2887 30250 2896
rect 29552 2576 29604 2582
rect 29552 2518 29604 2524
rect 30300 480 30328 3946
rect 30392 3777 30420 4014
rect 30470 3904 30526 3913
rect 30470 3839 30526 3848
rect 30378 3768 30434 3777
rect 30484 3738 30512 3839
rect 30378 3703 30434 3712
rect 30472 3732 30524 3738
rect 30472 3674 30524 3680
rect 30380 3392 30432 3398
rect 30380 3334 30432 3340
rect 30392 3058 30420 3334
rect 30380 3052 30432 3058
rect 30380 2994 30432 3000
rect 30392 2650 30420 2994
rect 30484 2854 30512 3674
rect 30944 3602 30972 5879
rect 31852 5704 31904 5710
rect 31852 5646 31904 5652
rect 31864 5166 31892 5646
rect 31852 5160 31904 5166
rect 31852 5102 31904 5108
rect 31392 5092 31444 5098
rect 31392 5034 31444 5040
rect 31404 4826 31432 5034
rect 31392 4820 31444 4826
rect 31392 4762 31444 4768
rect 31850 4584 31906 4593
rect 31850 4519 31852 4528
rect 31904 4519 31906 4528
rect 31852 4490 31904 4496
rect 31484 3936 31536 3942
rect 31484 3878 31536 3884
rect 30932 3596 30984 3602
rect 30932 3538 30984 3544
rect 30944 3194 30972 3538
rect 31116 3392 31168 3398
rect 31116 3334 31168 3340
rect 30932 3188 30984 3194
rect 30932 3130 30984 3136
rect 30472 2848 30524 2854
rect 31128 2825 31156 3334
rect 31496 2990 31524 3878
rect 31864 3534 31892 4490
rect 32048 3913 32076 13790
rect 32220 13728 32272 13734
rect 32220 13670 32272 13676
rect 32232 13258 32260 13670
rect 32876 13462 32904 13874
rect 32680 13456 32732 13462
rect 32680 13398 32732 13404
rect 32864 13456 32916 13462
rect 32864 13398 32916 13404
rect 32220 13252 32272 13258
rect 32220 13194 32272 13200
rect 32692 12986 32720 13398
rect 32772 13184 32824 13190
rect 32772 13126 32824 13132
rect 32680 12980 32732 12986
rect 32680 12922 32732 12928
rect 32128 12776 32180 12782
rect 32128 12718 32180 12724
rect 32140 12238 32168 12718
rect 32692 12374 32720 12922
rect 32784 12782 32812 13126
rect 32876 12918 32904 13398
rect 32864 12912 32916 12918
rect 32864 12854 32916 12860
rect 32772 12776 32824 12782
rect 32772 12718 32824 12724
rect 32680 12368 32732 12374
rect 32680 12310 32732 12316
rect 32128 12232 32180 12238
rect 32128 12174 32180 12180
rect 32140 11937 32168 12174
rect 32126 11928 32182 11937
rect 32692 11898 32720 12310
rect 32126 11863 32128 11872
rect 32180 11863 32182 11872
rect 32680 11892 32732 11898
rect 32128 11834 32180 11840
rect 32680 11834 32732 11840
rect 32496 8832 32548 8838
rect 32496 8774 32548 8780
rect 32508 8362 32536 8774
rect 32496 8356 32548 8362
rect 32496 8298 32548 8304
rect 32508 7546 32536 8298
rect 32496 7540 32548 7546
rect 32496 7482 32548 7488
rect 32496 6860 32548 6866
rect 32496 6802 32548 6808
rect 32508 6662 32536 6802
rect 32496 6656 32548 6662
rect 32496 6598 32548 6604
rect 32402 6352 32458 6361
rect 32402 6287 32404 6296
rect 32456 6287 32458 6296
rect 32404 6258 32456 6264
rect 32312 5772 32364 5778
rect 32312 5714 32364 5720
rect 32324 5030 32352 5714
rect 32312 5024 32364 5030
rect 32312 4966 32364 4972
rect 32324 4690 32352 4966
rect 32508 4826 32536 6598
rect 32496 4820 32548 4826
rect 32496 4762 32548 4768
rect 32128 4684 32180 4690
rect 32128 4626 32180 4632
rect 32312 4684 32364 4690
rect 32312 4626 32364 4632
rect 32140 3942 32168 4626
rect 32324 4214 32352 4626
rect 32312 4208 32364 4214
rect 32968 4185 32996 15846
rect 33048 15632 33100 15638
rect 33048 15574 33100 15580
rect 33060 15162 33088 15574
rect 33520 15502 33548 16118
rect 33508 15496 33560 15502
rect 33508 15438 33560 15444
rect 33140 15360 33192 15366
rect 33140 15302 33192 15308
rect 33152 15162 33180 15302
rect 33048 15156 33100 15162
rect 33048 15098 33100 15104
rect 33140 15156 33192 15162
rect 33140 15098 33192 15104
rect 33520 14618 33548 15438
rect 33508 14612 33560 14618
rect 33508 14554 33560 14560
rect 33612 14362 33640 19110
rect 34440 18290 34468 19246
rect 34532 18902 34560 20198
rect 34612 19916 34664 19922
rect 34612 19858 34664 19864
rect 34624 18970 34652 19858
rect 34716 19854 34744 20538
rect 35440 20256 35492 20262
rect 35440 20198 35492 20204
rect 34794 20088 34850 20097
rect 34794 20023 34850 20032
rect 34704 19848 34756 19854
rect 34704 19790 34756 19796
rect 34704 19712 34756 19718
rect 34808 19700 34836 20023
rect 34978 19952 35034 19961
rect 34978 19887 34980 19896
rect 35032 19887 35034 19896
rect 34980 19858 35032 19864
rect 34756 19672 34836 19700
rect 34704 19654 34756 19660
rect 34702 19408 34758 19417
rect 34702 19343 34758 19352
rect 34716 19310 34744 19343
rect 34808 19310 34836 19672
rect 34940 19612 35236 19632
rect 34996 19610 35020 19612
rect 35076 19610 35100 19612
rect 35156 19610 35180 19612
rect 35018 19558 35020 19610
rect 35082 19558 35094 19610
rect 35156 19558 35158 19610
rect 34996 19556 35020 19558
rect 35076 19556 35100 19558
rect 35156 19556 35180 19558
rect 34940 19536 35236 19556
rect 35452 19378 35480 20198
rect 35440 19372 35492 19378
rect 35440 19314 35492 19320
rect 34704 19304 34756 19310
rect 34704 19246 34756 19252
rect 34796 19304 34848 19310
rect 34796 19246 34848 19252
rect 35348 19304 35400 19310
rect 35348 19246 35400 19252
rect 34612 18964 34664 18970
rect 34612 18906 34664 18912
rect 34520 18896 34572 18902
rect 34520 18838 34572 18844
rect 34520 18760 34572 18766
rect 34520 18702 34572 18708
rect 34428 18284 34480 18290
rect 34428 18226 34480 18232
rect 33692 16788 33744 16794
rect 33692 16730 33744 16736
rect 33704 16114 33732 16730
rect 34440 16726 34468 18226
rect 34532 17678 34560 18702
rect 34808 18222 34836 19246
rect 35360 18902 35388 19246
rect 35348 18896 35400 18902
rect 35348 18838 35400 18844
rect 35256 18624 35308 18630
rect 35256 18566 35308 18572
rect 34940 18524 35236 18544
rect 34996 18522 35020 18524
rect 35076 18522 35100 18524
rect 35156 18522 35180 18524
rect 35018 18470 35020 18522
rect 35082 18470 35094 18522
rect 35156 18470 35158 18522
rect 34996 18468 35020 18470
rect 35076 18468 35100 18470
rect 35156 18468 35180 18470
rect 34940 18448 35236 18468
rect 34796 18216 34848 18222
rect 34796 18158 34848 18164
rect 35268 17814 35296 18566
rect 35360 18358 35388 18838
rect 35348 18352 35400 18358
rect 35348 18294 35400 18300
rect 35348 18216 35400 18222
rect 35348 18158 35400 18164
rect 34704 17808 34756 17814
rect 34704 17750 34756 17756
rect 35256 17808 35308 17814
rect 35256 17750 35308 17756
rect 34520 17672 34572 17678
rect 34520 17614 34572 17620
rect 34716 17338 34744 17750
rect 35256 17672 35308 17678
rect 35256 17614 35308 17620
rect 34940 17436 35236 17456
rect 34996 17434 35020 17436
rect 35076 17434 35100 17436
rect 35156 17434 35180 17436
rect 35018 17382 35020 17434
rect 35082 17382 35094 17434
rect 35156 17382 35158 17434
rect 34996 17380 35020 17382
rect 35076 17380 35100 17382
rect 35156 17380 35180 17382
rect 34940 17360 35236 17380
rect 35268 17338 35296 17614
rect 34704 17332 34756 17338
rect 34704 17274 34756 17280
rect 35256 17332 35308 17338
rect 35256 17274 35308 17280
rect 34428 16720 34480 16726
rect 34428 16662 34480 16668
rect 33784 16652 33836 16658
rect 33784 16594 33836 16600
rect 34060 16652 34112 16658
rect 34060 16594 34112 16600
rect 33796 16250 33824 16594
rect 33968 16448 34020 16454
rect 33968 16390 34020 16396
rect 33784 16244 33836 16250
rect 33784 16186 33836 16192
rect 33692 16108 33744 16114
rect 33692 16050 33744 16056
rect 33796 15314 33824 16186
rect 33980 15978 34008 16390
rect 34072 16182 34100 16594
rect 34940 16348 35236 16368
rect 34996 16346 35020 16348
rect 35076 16346 35100 16348
rect 35156 16346 35180 16348
rect 35018 16294 35020 16346
rect 35082 16294 35094 16346
rect 35156 16294 35158 16346
rect 34996 16292 35020 16294
rect 35076 16292 35100 16294
rect 35156 16292 35180 16294
rect 34940 16272 35236 16292
rect 34060 16176 34112 16182
rect 34060 16118 34112 16124
rect 33968 15972 34020 15978
rect 33968 15914 34020 15920
rect 34336 15972 34388 15978
rect 34336 15914 34388 15920
rect 34348 15314 34376 15914
rect 35256 15632 35308 15638
rect 35256 15574 35308 15580
rect 34796 15564 34848 15570
rect 34796 15506 34848 15512
rect 34428 15496 34480 15502
rect 34480 15444 34560 15450
rect 34428 15438 34560 15444
rect 34440 15422 34560 15438
rect 34428 15360 34480 15366
rect 33796 15286 33916 15314
rect 34348 15308 34428 15314
rect 34348 15302 34480 15308
rect 34348 15286 34468 15302
rect 33612 14334 33732 14362
rect 33600 14272 33652 14278
rect 33600 14214 33652 14220
rect 33612 13870 33640 14214
rect 33600 13864 33652 13870
rect 33600 13806 33652 13812
rect 33232 13524 33284 13530
rect 33232 13466 33284 13472
rect 33048 13388 33100 13394
rect 33048 13330 33100 13336
rect 33060 12458 33088 13330
rect 33244 12782 33272 13466
rect 33324 13388 33376 13394
rect 33324 13330 33376 13336
rect 33232 12776 33284 12782
rect 33232 12718 33284 12724
rect 33232 12640 33284 12646
rect 33336 12594 33364 13330
rect 33284 12588 33364 12594
rect 33232 12582 33364 12588
rect 33244 12566 33364 12582
rect 33060 12442 33180 12458
rect 33060 12436 33192 12442
rect 33060 12430 33140 12436
rect 33140 12378 33192 12384
rect 33244 12102 33272 12566
rect 33232 12096 33284 12102
rect 33232 12038 33284 12044
rect 33244 10169 33272 12038
rect 33704 11286 33732 14334
rect 33888 13802 33916 15286
rect 33968 14272 34020 14278
rect 33968 14214 34020 14220
rect 33980 14006 34008 14214
rect 34440 14006 34468 15286
rect 34532 14346 34560 15422
rect 34808 15162 34836 15506
rect 34940 15260 35236 15280
rect 34996 15258 35020 15260
rect 35076 15258 35100 15260
rect 35156 15258 35180 15260
rect 35018 15206 35020 15258
rect 35082 15206 35094 15258
rect 35156 15206 35158 15258
rect 34996 15204 35020 15206
rect 35076 15204 35100 15206
rect 35156 15204 35180 15206
rect 34940 15184 35236 15204
rect 34796 15156 34848 15162
rect 34796 15098 34848 15104
rect 34808 14618 34836 15098
rect 35164 14952 35216 14958
rect 35164 14894 35216 14900
rect 34796 14612 34848 14618
rect 34796 14554 34848 14560
rect 35176 14362 35204 14894
rect 35268 14890 35296 15574
rect 35256 14884 35308 14890
rect 35256 14826 35308 14832
rect 34520 14340 34572 14346
rect 35176 14334 35296 14362
rect 34520 14282 34572 14288
rect 33968 14000 34020 14006
rect 33968 13942 34020 13948
rect 34428 14000 34480 14006
rect 34428 13942 34480 13948
rect 33876 13796 33928 13802
rect 33876 13738 33928 13744
rect 33784 13728 33836 13734
rect 33784 13670 33836 13676
rect 33796 12714 33824 13670
rect 33888 13190 33916 13738
rect 34440 13410 34468 13942
rect 34532 13530 34560 14282
rect 35268 14278 35296 14334
rect 35256 14272 35308 14278
rect 35256 14214 35308 14220
rect 34940 14172 35236 14192
rect 34996 14170 35020 14172
rect 35076 14170 35100 14172
rect 35156 14170 35180 14172
rect 35018 14118 35020 14170
rect 35082 14118 35094 14170
rect 35156 14118 35158 14170
rect 34996 14116 35020 14118
rect 35076 14116 35100 14118
rect 35156 14116 35180 14118
rect 34940 14096 35236 14116
rect 34796 13864 34848 13870
rect 35164 13864 35216 13870
rect 35162 13832 35164 13841
rect 35216 13832 35218 13841
rect 34848 13812 35162 13818
rect 34796 13806 35162 13812
rect 34808 13790 35162 13806
rect 35268 13802 35296 14214
rect 35162 13767 35218 13776
rect 35256 13796 35308 13802
rect 35176 13707 35204 13767
rect 35256 13738 35308 13744
rect 34520 13524 34572 13530
rect 34520 13466 34572 13472
rect 35360 13462 35388 18158
rect 35452 17610 35480 19314
rect 35636 19174 35664 20567
rect 35808 20538 35860 20544
rect 36084 19712 36136 19718
rect 36084 19654 36136 19660
rect 35624 19168 35676 19174
rect 35624 19110 35676 19116
rect 36096 18902 36124 19654
rect 35624 18896 35676 18902
rect 35622 18864 35624 18873
rect 36084 18896 36136 18902
rect 35676 18864 35678 18873
rect 35622 18799 35678 18808
rect 36004 18856 36084 18884
rect 35636 18426 35664 18799
rect 35624 18420 35676 18426
rect 35624 18362 35676 18368
rect 36004 18222 36032 18856
rect 36084 18838 36136 18844
rect 35808 18216 35860 18222
rect 35808 18158 35860 18164
rect 35992 18216 36044 18222
rect 35992 18158 36044 18164
rect 35820 18086 35848 18158
rect 35808 18080 35860 18086
rect 35808 18022 35860 18028
rect 36004 17882 36032 18158
rect 35992 17876 36044 17882
rect 35992 17818 36044 17824
rect 35532 17672 35584 17678
rect 35532 17614 35584 17620
rect 35440 17604 35492 17610
rect 35440 17546 35492 17552
rect 35544 17270 35572 17614
rect 35532 17264 35584 17270
rect 35530 17232 35532 17241
rect 35584 17232 35586 17241
rect 35530 17167 35586 17176
rect 35716 15972 35768 15978
rect 35716 15914 35768 15920
rect 35728 15570 35756 15914
rect 35716 15564 35768 15570
rect 35716 15506 35768 15512
rect 36188 14521 36216 22879
rect 37292 22658 37320 23462
rect 37384 22778 37412 24126
rect 38212 23322 38240 24890
rect 38580 24410 38608 25366
rect 38672 25362 38700 25978
rect 39578 25528 39634 25537
rect 39578 25463 39634 25472
rect 39592 25430 39620 25463
rect 39580 25424 39632 25430
rect 39580 25366 39632 25372
rect 38660 25356 38712 25362
rect 38660 25298 38712 25304
rect 38672 24954 38700 25298
rect 39592 24954 39620 25366
rect 38660 24948 38712 24954
rect 38660 24890 38712 24896
rect 39580 24948 39632 24954
rect 39580 24890 39632 24896
rect 38752 24812 38804 24818
rect 38752 24754 38804 24760
rect 38660 24744 38712 24750
rect 38658 24712 38660 24721
rect 38712 24712 38714 24721
rect 38658 24647 38714 24656
rect 38568 24404 38620 24410
rect 38568 24346 38620 24352
rect 38476 23520 38528 23526
rect 38476 23462 38528 23468
rect 38660 23520 38712 23526
rect 38660 23462 38712 23468
rect 38200 23316 38252 23322
rect 38200 23258 38252 23264
rect 37372 22772 37424 22778
rect 37372 22714 37424 22720
rect 37200 22630 37320 22658
rect 38488 22642 38516 23462
rect 38672 23186 38700 23462
rect 38764 23186 38792 24754
rect 39120 24608 39172 24614
rect 39120 24550 39172 24556
rect 38936 23316 38988 23322
rect 38936 23258 38988 23264
rect 38660 23180 38712 23186
rect 38660 23122 38712 23128
rect 38752 23180 38804 23186
rect 38752 23122 38804 23128
rect 38568 22704 38620 22710
rect 38568 22646 38620 22652
rect 38672 22658 38700 23122
rect 38476 22636 38528 22642
rect 37200 22574 37228 22630
rect 38476 22578 38528 22584
rect 37188 22568 37240 22574
rect 37188 22510 37240 22516
rect 38200 22568 38252 22574
rect 38200 22510 38252 22516
rect 37280 22432 37332 22438
rect 37280 22374 37332 22380
rect 36452 22092 36504 22098
rect 36452 22034 36504 22040
rect 36544 22092 36596 22098
rect 36544 22034 36596 22040
rect 37188 22092 37240 22098
rect 37292 22080 37320 22374
rect 37372 22228 37424 22234
rect 37372 22170 37424 22176
rect 37240 22052 37320 22080
rect 37188 22034 37240 22040
rect 36464 21418 36492 22034
rect 36452 21412 36504 21418
rect 36452 21354 36504 21360
rect 36464 21146 36492 21354
rect 36556 21146 36584 22034
rect 37384 21690 37412 22170
rect 37556 22092 37608 22098
rect 37556 22034 37608 22040
rect 37568 21894 37596 22034
rect 38212 22030 38240 22510
rect 38580 22234 38608 22646
rect 38672 22630 38792 22658
rect 38660 22500 38712 22506
rect 38660 22442 38712 22448
rect 38568 22228 38620 22234
rect 38568 22170 38620 22176
rect 38672 22030 38700 22442
rect 38764 22234 38792 22630
rect 38948 22438 38976 23258
rect 39132 23118 39160 24550
rect 40328 24177 40356 28426
rect 41156 28014 41184 29158
rect 41236 29106 41288 29112
rect 41236 29028 41288 29034
rect 41236 28970 41288 28976
rect 41248 28937 41276 28970
rect 41234 28928 41290 28937
rect 41234 28863 41290 28872
rect 41248 28762 41276 28863
rect 41236 28756 41288 28762
rect 41236 28698 41288 28704
rect 41144 28008 41196 28014
rect 41144 27950 41196 27956
rect 41340 27554 41368 29174
rect 41708 29034 41736 30194
rect 41800 29034 41828 30534
rect 41892 30394 41920 30738
rect 42076 30394 42104 30806
rect 41880 30388 41932 30394
rect 41880 30330 41932 30336
rect 42064 30388 42116 30394
rect 42064 30330 42116 30336
rect 41880 29844 41932 29850
rect 41880 29786 41932 29792
rect 41892 29306 41920 29786
rect 42064 29640 42116 29646
rect 42064 29582 42116 29588
rect 42076 29306 42104 29582
rect 41880 29300 41932 29306
rect 41880 29242 41932 29248
rect 42064 29300 42116 29306
rect 42064 29242 42116 29248
rect 41696 29028 41748 29034
rect 41696 28970 41748 28976
rect 41788 29028 41840 29034
rect 41788 28970 41840 28976
rect 42076 28937 42104 29242
rect 42062 28928 42118 28937
rect 42062 28863 42118 28872
rect 41972 28688 42024 28694
rect 41972 28630 42024 28636
rect 41880 28552 41932 28558
rect 41880 28494 41932 28500
rect 41512 28416 41564 28422
rect 41512 28358 41564 28364
rect 41420 27600 41472 27606
rect 41340 27548 41420 27554
rect 41340 27542 41472 27548
rect 41340 27526 41460 27542
rect 41524 27538 41552 28358
rect 41694 27976 41750 27985
rect 41694 27911 41750 27920
rect 41512 27532 41564 27538
rect 41512 27474 41564 27480
rect 41420 26920 41472 26926
rect 41420 26862 41472 26868
rect 40684 26444 40736 26450
rect 40684 26386 40736 26392
rect 40592 25968 40644 25974
rect 40592 25910 40644 25916
rect 40604 25673 40632 25910
rect 40696 25906 40724 26386
rect 41328 26308 41380 26314
rect 41328 26250 41380 26256
rect 40684 25900 40736 25906
rect 40684 25842 40736 25848
rect 40590 25664 40646 25673
rect 40590 25599 40646 25608
rect 40696 25498 40724 25842
rect 41340 25770 41368 26250
rect 41432 25974 41460 26862
rect 41524 26586 41552 27474
rect 41708 27402 41736 27911
rect 41892 27878 41920 28494
rect 41880 27872 41932 27878
rect 41880 27814 41932 27820
rect 41696 27396 41748 27402
rect 41696 27338 41748 27344
rect 41892 26858 41920 27814
rect 41984 27674 42012 28630
rect 42076 28626 42104 28863
rect 42064 28620 42116 28626
rect 42064 28562 42116 28568
rect 41972 27668 42024 27674
rect 41972 27610 42024 27616
rect 41880 26852 41932 26858
rect 41880 26794 41932 26800
rect 41512 26580 41564 26586
rect 41512 26522 41564 26528
rect 41880 26512 41932 26518
rect 41880 26454 41932 26460
rect 41604 26308 41656 26314
rect 41604 26250 41656 26256
rect 41616 26042 41644 26250
rect 41604 26036 41656 26042
rect 41604 25978 41656 25984
rect 41420 25968 41472 25974
rect 41420 25910 41472 25916
rect 41328 25764 41380 25770
rect 41328 25706 41380 25712
rect 41892 25498 41920 26454
rect 41972 26376 42024 26382
rect 41972 26318 42024 26324
rect 41984 26042 42012 26318
rect 41972 26036 42024 26042
rect 41972 25978 42024 25984
rect 41984 25537 42012 25978
rect 41970 25528 42026 25537
rect 40684 25492 40736 25498
rect 40684 25434 40736 25440
rect 41880 25492 41932 25498
rect 41970 25463 42026 25472
rect 41880 25434 41932 25440
rect 41050 24848 41106 24857
rect 41050 24783 41106 24792
rect 40314 24168 40370 24177
rect 40314 24103 40370 24112
rect 41064 23866 41092 24783
rect 41892 24410 41920 25434
rect 41984 25430 42012 25463
rect 41972 25424 42024 25430
rect 41972 25366 42024 25372
rect 42064 24608 42116 24614
rect 42064 24550 42116 24556
rect 41880 24404 41932 24410
rect 41880 24346 41932 24352
rect 42076 24274 42104 24550
rect 42064 24268 42116 24274
rect 42064 24210 42116 24216
rect 41604 24064 41656 24070
rect 41604 24006 41656 24012
rect 41052 23860 41104 23866
rect 41052 23802 41104 23808
rect 41616 23730 41644 24006
rect 42076 23866 42104 24210
rect 42064 23860 42116 23866
rect 42064 23802 42116 23808
rect 42168 23746 42196 41262
rect 45652 37664 45704 37670
rect 45652 37606 45704 37612
rect 42340 31680 42392 31686
rect 42340 31622 42392 31628
rect 42352 31210 42380 31622
rect 42616 31272 42668 31278
rect 42616 31214 42668 31220
rect 42340 31204 42392 31210
rect 42340 31146 42392 31152
rect 42352 30938 42380 31146
rect 42340 30932 42392 30938
rect 42340 30874 42392 30880
rect 42628 30734 42656 31214
rect 43444 31136 43496 31142
rect 43444 31078 43496 31084
rect 42340 30728 42392 30734
rect 42340 30670 42392 30676
rect 42616 30728 42668 30734
rect 42616 30670 42668 30676
rect 43352 30728 43404 30734
rect 43352 30670 43404 30676
rect 42352 29646 42380 30670
rect 42628 30394 42656 30670
rect 42616 30388 42668 30394
rect 42616 30330 42668 30336
rect 42800 30184 42852 30190
rect 42800 30126 42852 30132
rect 42812 29850 42840 30126
rect 43364 29850 43392 30670
rect 43456 30190 43484 31078
rect 43628 30796 43680 30802
rect 43628 30738 43680 30744
rect 45560 30796 45612 30802
rect 45560 30738 45612 30744
rect 43640 30705 43668 30738
rect 43626 30696 43682 30705
rect 43626 30631 43682 30640
rect 43444 30184 43496 30190
rect 43444 30126 43496 30132
rect 43640 29850 43668 30631
rect 45572 30326 45600 30738
rect 45560 30320 45612 30326
rect 45560 30262 45612 30268
rect 44088 30048 44140 30054
rect 44088 29990 44140 29996
rect 45192 30048 45244 30054
rect 45192 29990 45244 29996
rect 42800 29844 42852 29850
rect 42800 29786 42852 29792
rect 43352 29844 43404 29850
rect 43352 29786 43404 29792
rect 43628 29844 43680 29850
rect 43628 29786 43680 29792
rect 42432 29776 42484 29782
rect 42432 29718 42484 29724
rect 42340 29640 42392 29646
rect 42340 29582 42392 29588
rect 42340 29504 42392 29510
rect 42340 29446 42392 29452
rect 42352 29102 42380 29446
rect 42444 29345 42472 29718
rect 43364 29714 43392 29786
rect 44100 29782 44128 29990
rect 45008 29844 45060 29850
rect 45008 29786 45060 29792
rect 44088 29776 44140 29782
rect 44088 29718 44140 29724
rect 43352 29708 43404 29714
rect 43352 29650 43404 29656
rect 42430 29336 42486 29345
rect 42430 29271 42486 29280
rect 42340 29096 42392 29102
rect 42340 29038 42392 29044
rect 42444 28762 42472 29271
rect 42892 29232 42944 29238
rect 42892 29174 42944 29180
rect 44916 29232 44968 29238
rect 44916 29174 44968 29180
rect 42800 29164 42852 29170
rect 42800 29106 42852 29112
rect 42812 28762 42840 29106
rect 42432 28756 42484 28762
rect 42432 28698 42484 28704
rect 42800 28756 42852 28762
rect 42800 28698 42852 28704
rect 42904 28626 42932 29174
rect 44928 28626 44956 29174
rect 45020 29170 45048 29786
rect 45204 29714 45232 29990
rect 45572 29850 45600 30262
rect 45560 29844 45612 29850
rect 45560 29786 45612 29792
rect 45192 29708 45244 29714
rect 45192 29650 45244 29656
rect 45204 29306 45232 29650
rect 45100 29300 45152 29306
rect 45100 29242 45152 29248
rect 45192 29300 45244 29306
rect 45192 29242 45244 29248
rect 45560 29300 45612 29306
rect 45560 29242 45612 29248
rect 45008 29164 45060 29170
rect 45008 29106 45060 29112
rect 45112 29034 45140 29242
rect 45100 29028 45152 29034
rect 45100 28970 45152 28976
rect 45468 29028 45520 29034
rect 45468 28970 45520 28976
rect 45192 28960 45244 28966
rect 45192 28902 45244 28908
rect 45100 28688 45152 28694
rect 45100 28630 45152 28636
rect 42892 28620 42944 28626
rect 42892 28562 42944 28568
rect 43996 28620 44048 28626
rect 43996 28562 44048 28568
rect 44916 28620 44968 28626
rect 44916 28562 44968 28568
rect 43536 28416 43588 28422
rect 43536 28358 43588 28364
rect 42892 28144 42944 28150
rect 42892 28086 42944 28092
rect 42800 27872 42852 27878
rect 42800 27814 42852 27820
rect 42812 27674 42840 27814
rect 42800 27668 42852 27674
rect 42800 27610 42852 27616
rect 42248 27464 42300 27470
rect 42246 27432 42248 27441
rect 42300 27432 42302 27441
rect 42246 27367 42302 27376
rect 42432 26784 42484 26790
rect 42432 26726 42484 26732
rect 42444 26246 42472 26726
rect 42432 26240 42484 26246
rect 42432 26182 42484 26188
rect 42248 25968 42300 25974
rect 42248 25910 42300 25916
rect 42260 23866 42288 25910
rect 42444 25770 42472 26182
rect 42432 25764 42484 25770
rect 42432 25706 42484 25712
rect 42616 25288 42668 25294
rect 42616 25230 42668 25236
rect 42340 25152 42392 25158
rect 42340 25094 42392 25100
rect 42352 24954 42380 25094
rect 42340 24948 42392 24954
rect 42340 24890 42392 24896
rect 42338 24712 42394 24721
rect 42338 24647 42394 24656
rect 42352 24614 42380 24647
rect 42340 24608 42392 24614
rect 42340 24550 42392 24556
rect 42352 24410 42380 24550
rect 42628 24410 42656 25230
rect 42904 24614 42932 28086
rect 43168 28076 43220 28082
rect 43168 28018 43220 28024
rect 43180 27674 43208 28018
rect 43548 27946 43576 28358
rect 44008 28218 44036 28562
rect 44640 28416 44692 28422
rect 44640 28358 44692 28364
rect 43996 28212 44048 28218
rect 43996 28154 44048 28160
rect 44548 28008 44600 28014
rect 44546 27976 44548 27985
rect 44600 27976 44602 27985
rect 43536 27940 43588 27946
rect 43536 27882 43588 27888
rect 44088 27940 44140 27946
rect 44546 27911 44602 27920
rect 44088 27882 44140 27888
rect 43168 27668 43220 27674
rect 43168 27610 43220 27616
rect 43260 27600 43312 27606
rect 43260 27542 43312 27548
rect 43272 27130 43300 27542
rect 43260 27124 43312 27130
rect 43260 27066 43312 27072
rect 43904 27056 43956 27062
rect 43904 26998 43956 27004
rect 43916 26450 43944 26998
rect 44100 26858 44128 27882
rect 44652 27538 44680 28358
rect 44928 27674 44956 28562
rect 45112 28218 45140 28630
rect 45204 28558 45232 28902
rect 45192 28552 45244 28558
rect 45192 28494 45244 28500
rect 45100 28212 45152 28218
rect 45100 28154 45152 28160
rect 44916 27668 44968 27674
rect 44916 27610 44968 27616
rect 44640 27532 44692 27538
rect 44640 27474 44692 27480
rect 44272 27328 44324 27334
rect 44272 27270 44324 27276
rect 44284 26994 44312 27270
rect 44652 27130 44680 27474
rect 45204 27441 45232 28494
rect 45480 27878 45508 28970
rect 45572 28626 45600 29242
rect 45560 28620 45612 28626
rect 45560 28562 45612 28568
rect 45572 28150 45600 28562
rect 45560 28144 45612 28150
rect 45560 28086 45612 28092
rect 45468 27872 45520 27878
rect 45468 27814 45520 27820
rect 45572 27538 45600 28086
rect 45560 27532 45612 27538
rect 45560 27474 45612 27480
rect 45190 27432 45246 27441
rect 45190 27367 45246 27376
rect 45204 27334 45232 27367
rect 45192 27328 45244 27334
rect 45192 27270 45244 27276
rect 44640 27124 44692 27130
rect 44640 27066 44692 27072
rect 44272 26988 44324 26994
rect 44272 26930 44324 26936
rect 44088 26852 44140 26858
rect 44088 26794 44140 26800
rect 45008 26784 45060 26790
rect 45008 26726 45060 26732
rect 44732 26512 44784 26518
rect 44732 26454 44784 26460
rect 43352 26444 43404 26450
rect 43352 26386 43404 26392
rect 43904 26444 43956 26450
rect 43904 26386 43956 26392
rect 44548 26444 44600 26450
rect 44548 26386 44600 26392
rect 43364 24750 43392 26386
rect 44560 25974 44588 26386
rect 44640 26240 44692 26246
rect 44640 26182 44692 26188
rect 44548 25968 44600 25974
rect 44548 25910 44600 25916
rect 43536 25764 43588 25770
rect 43536 25706 43588 25712
rect 43444 25424 43496 25430
rect 43444 25366 43496 25372
rect 43352 24744 43404 24750
rect 43352 24686 43404 24692
rect 43456 24614 43484 25366
rect 43548 25362 43576 25706
rect 44560 25498 44588 25910
rect 44652 25838 44680 26182
rect 44640 25832 44692 25838
rect 44640 25774 44692 25780
rect 44652 25498 44680 25774
rect 44744 25702 44772 26454
rect 45020 26042 45048 26726
rect 45204 26382 45232 27270
rect 45572 27130 45600 27474
rect 45560 27124 45612 27130
rect 45560 27066 45612 27072
rect 45284 26784 45336 26790
rect 45282 26752 45284 26761
rect 45336 26752 45338 26761
rect 45282 26687 45338 26696
rect 45572 26450 45600 27066
rect 45560 26444 45612 26450
rect 45560 26386 45612 26392
rect 45192 26376 45244 26382
rect 45190 26344 45192 26353
rect 45244 26344 45246 26353
rect 45190 26279 45246 26288
rect 45572 26042 45600 26386
rect 45008 26036 45060 26042
rect 45008 25978 45060 25984
rect 45560 26036 45612 26042
rect 45560 25978 45612 25984
rect 44732 25696 44784 25702
rect 44732 25638 44784 25644
rect 44548 25492 44600 25498
rect 44548 25434 44600 25440
rect 44640 25492 44692 25498
rect 44640 25434 44692 25440
rect 43536 25356 43588 25362
rect 43536 25298 43588 25304
rect 43548 24954 43576 25298
rect 44744 25226 44772 25638
rect 44732 25220 44784 25226
rect 44732 25162 44784 25168
rect 45572 24954 45600 25978
rect 43536 24948 43588 24954
rect 43536 24890 43588 24896
rect 45560 24948 45612 24954
rect 45560 24890 45612 24896
rect 45664 24857 45692 37606
rect 45836 30728 45888 30734
rect 45836 30670 45888 30676
rect 45848 30190 45876 30670
rect 45928 30388 45980 30394
rect 45928 30330 45980 30336
rect 45836 30184 45888 30190
rect 45836 30126 45888 30132
rect 45848 30054 45876 30126
rect 45836 30048 45888 30054
rect 45836 29990 45888 29996
rect 45836 29776 45888 29782
rect 45836 29718 45888 29724
rect 45848 29306 45876 29718
rect 45836 29300 45888 29306
rect 45836 29242 45888 29248
rect 45848 29102 45876 29242
rect 45836 29096 45888 29102
rect 45836 29038 45888 29044
rect 45744 29028 45796 29034
rect 45744 28970 45796 28976
rect 45756 28490 45784 28970
rect 45744 28484 45796 28490
rect 45744 28426 45796 28432
rect 45836 25288 45888 25294
rect 45836 25230 45888 25236
rect 45650 24848 45706 24857
rect 45650 24783 45706 24792
rect 42892 24608 42944 24614
rect 42892 24550 42944 24556
rect 43444 24608 43496 24614
rect 43444 24550 43496 24556
rect 42340 24404 42392 24410
rect 42340 24346 42392 24352
rect 42616 24404 42668 24410
rect 42616 24346 42668 24352
rect 43456 24177 43484 24550
rect 45848 24410 45876 25230
rect 45836 24404 45888 24410
rect 45836 24346 45888 24352
rect 45468 24200 45520 24206
rect 43442 24168 43498 24177
rect 45468 24142 45520 24148
rect 43442 24103 43498 24112
rect 42248 23860 42300 23866
rect 42248 23802 42300 23808
rect 41604 23724 41656 23730
rect 41604 23666 41656 23672
rect 41892 23718 42196 23746
rect 41420 23588 41472 23594
rect 41420 23530 41472 23536
rect 41052 23520 41104 23526
rect 41052 23462 41104 23468
rect 39856 23180 39908 23186
rect 39856 23122 39908 23128
rect 39028 23112 39080 23118
rect 39028 23054 39080 23060
rect 39120 23112 39172 23118
rect 39120 23054 39172 23060
rect 39040 22574 39068 23054
rect 39132 22778 39160 23054
rect 39868 22778 39896 23122
rect 40500 22976 40552 22982
rect 40498 22944 40500 22953
rect 40552 22944 40554 22953
rect 40498 22879 40554 22888
rect 39120 22772 39172 22778
rect 39120 22714 39172 22720
rect 39856 22772 39908 22778
rect 39856 22714 39908 22720
rect 39028 22568 39080 22574
rect 39028 22510 39080 22516
rect 38936 22432 38988 22438
rect 38936 22374 38988 22380
rect 39868 22234 39896 22714
rect 40408 22432 40460 22438
rect 40408 22374 40460 22380
rect 38752 22228 38804 22234
rect 38752 22170 38804 22176
rect 39856 22228 39908 22234
rect 39856 22170 39908 22176
rect 38200 22024 38252 22030
rect 38200 21966 38252 21972
rect 38660 22024 38712 22030
rect 38660 21966 38712 21972
rect 37556 21888 37608 21894
rect 37556 21830 37608 21836
rect 37568 21690 37596 21830
rect 37372 21684 37424 21690
rect 37372 21626 37424 21632
rect 37556 21684 37608 21690
rect 37556 21626 37608 21632
rect 38212 21350 38240 21966
rect 38292 21888 38344 21894
rect 38292 21830 38344 21836
rect 36636 21344 36688 21350
rect 36636 21286 36688 21292
rect 38200 21344 38252 21350
rect 38200 21286 38252 21292
rect 36452 21140 36504 21146
rect 36452 21082 36504 21088
rect 36544 21140 36596 21146
rect 36544 21082 36596 21088
rect 36268 14884 36320 14890
rect 36268 14826 36320 14832
rect 36174 14512 36230 14521
rect 36174 14447 36230 14456
rect 36280 14074 36308 14826
rect 36648 14385 36676 21286
rect 38016 20800 38068 20806
rect 38212 20777 38240 21286
rect 38304 20806 38332 21830
rect 38672 21690 38700 21966
rect 38764 21894 38792 22170
rect 38752 21888 38804 21894
rect 38752 21830 38804 21836
rect 38660 21684 38712 21690
rect 38660 21626 38712 21632
rect 40316 20936 40368 20942
rect 40316 20878 40368 20884
rect 38292 20800 38344 20806
rect 38016 20742 38068 20748
rect 38198 20768 38254 20777
rect 37740 20460 37792 20466
rect 37740 20402 37792 20408
rect 37188 20256 37240 20262
rect 37188 20198 37240 20204
rect 37200 19242 37228 20198
rect 37752 19922 37780 20402
rect 38028 20398 38056 20742
rect 38292 20742 38344 20748
rect 38198 20703 38254 20712
rect 38016 20392 38068 20398
rect 38016 20334 38068 20340
rect 38028 20058 38056 20334
rect 38304 20097 38332 20742
rect 40328 20602 40356 20878
rect 40316 20596 40368 20602
rect 40316 20538 40368 20544
rect 39304 20256 39356 20262
rect 39304 20198 39356 20204
rect 39856 20256 39908 20262
rect 39856 20198 39908 20204
rect 38290 20088 38346 20097
rect 38016 20052 38068 20058
rect 38290 20023 38346 20032
rect 38660 20052 38712 20058
rect 38016 19994 38068 20000
rect 38660 19994 38712 20000
rect 37740 19916 37792 19922
rect 37740 19858 37792 19864
rect 38384 19916 38436 19922
rect 38384 19858 38436 19864
rect 37752 19514 37780 19858
rect 37740 19508 37792 19514
rect 37740 19450 37792 19456
rect 37188 19236 37240 19242
rect 37188 19178 37240 19184
rect 36912 19168 36964 19174
rect 36912 19110 36964 19116
rect 36924 18902 36952 19110
rect 36912 18896 36964 18902
rect 36912 18838 36964 18844
rect 36924 18426 36952 18838
rect 36912 18420 36964 18426
rect 36912 18362 36964 18368
rect 37188 18080 37240 18086
rect 37188 18022 37240 18028
rect 37200 17218 37228 18022
rect 37278 17232 37334 17241
rect 37200 17190 37278 17218
rect 37278 17167 37334 17176
rect 37292 17134 37320 17167
rect 37280 17128 37332 17134
rect 37280 17070 37332 17076
rect 37292 16794 37320 17070
rect 37752 17066 37780 19450
rect 37832 19168 37884 19174
rect 37832 19110 37884 19116
rect 37844 18698 37872 19110
rect 38106 18864 38162 18873
rect 38106 18799 38108 18808
rect 38160 18799 38162 18808
rect 38108 18770 38160 18776
rect 37832 18692 37884 18698
rect 37832 18634 37884 18640
rect 38120 18426 38148 18770
rect 38396 18766 38424 19858
rect 38672 19378 38700 19994
rect 39316 19990 39344 20198
rect 39304 19984 39356 19990
rect 39868 19961 39896 20198
rect 40224 19984 40276 19990
rect 39304 19926 39356 19932
rect 39854 19952 39910 19961
rect 40224 19926 40276 19932
rect 39854 19887 39910 19896
rect 40236 19378 40264 19926
rect 40420 19718 40448 22374
rect 40776 22092 40828 22098
rect 40776 22034 40828 22040
rect 40788 21486 40816 22034
rect 41064 21962 41092 23462
rect 41432 23322 41460 23530
rect 41420 23316 41472 23322
rect 41420 23258 41472 23264
rect 41328 22976 41380 22982
rect 41328 22918 41380 22924
rect 41340 22506 41368 22918
rect 41328 22500 41380 22506
rect 41328 22442 41380 22448
rect 41604 22500 41656 22506
rect 41604 22442 41656 22448
rect 41512 22160 41564 22166
rect 41512 22102 41564 22108
rect 41328 22092 41380 22098
rect 41328 22034 41380 22040
rect 41052 21956 41104 21962
rect 41052 21898 41104 21904
rect 41340 21554 41368 22034
rect 41524 21706 41552 22102
rect 41616 22030 41644 22442
rect 41604 22024 41656 22030
rect 41602 21992 41604 22001
rect 41656 21992 41658 22001
rect 41602 21927 41658 21936
rect 41432 21690 41552 21706
rect 41420 21684 41552 21690
rect 41472 21678 41552 21684
rect 41420 21626 41472 21632
rect 41328 21548 41380 21554
rect 41328 21490 41380 21496
rect 40776 21480 40828 21486
rect 40696 21440 40776 21468
rect 40590 20632 40646 20641
rect 40590 20567 40592 20576
rect 40644 20567 40646 20576
rect 40592 20538 40644 20544
rect 40696 20398 40724 21440
rect 40776 21422 40828 21428
rect 40776 21344 40828 21350
rect 40776 21286 40828 21292
rect 40788 20806 40816 21286
rect 41432 21146 41460 21626
rect 41616 21146 41644 21927
rect 41420 21140 41472 21146
rect 41420 21082 41472 21088
rect 41604 21140 41656 21146
rect 41604 21082 41656 21088
rect 40776 20800 40828 20806
rect 40774 20768 40776 20777
rect 41328 20800 41380 20806
rect 40828 20768 40830 20777
rect 41328 20742 41380 20748
rect 40774 20703 40830 20712
rect 40684 20392 40736 20398
rect 40684 20334 40736 20340
rect 40592 20256 40644 20262
rect 40592 20198 40644 20204
rect 40408 19712 40460 19718
rect 40408 19654 40460 19660
rect 38660 19372 38712 19378
rect 38660 19314 38712 19320
rect 40224 19372 40276 19378
rect 40224 19314 40276 19320
rect 38568 19304 38620 19310
rect 38566 19272 38568 19281
rect 38620 19272 38622 19281
rect 38566 19207 38622 19216
rect 38672 18970 38700 19314
rect 39120 19168 39172 19174
rect 39120 19110 39172 19116
rect 38660 18964 38712 18970
rect 38660 18906 38712 18912
rect 38384 18760 38436 18766
rect 38384 18702 38436 18708
rect 37832 18420 37884 18426
rect 37832 18362 37884 18368
rect 38108 18420 38160 18426
rect 38108 18362 38160 18368
rect 37740 17060 37792 17066
rect 37740 17002 37792 17008
rect 37280 16788 37332 16794
rect 37280 16730 37332 16736
rect 37648 14816 37700 14822
rect 37648 14758 37700 14764
rect 37660 14414 37688 14758
rect 37648 14408 37700 14414
rect 36634 14376 36690 14385
rect 37648 14350 37700 14356
rect 36634 14311 36690 14320
rect 36268 14068 36320 14074
rect 36268 14010 36320 14016
rect 37660 13870 37688 14350
rect 35716 13864 35768 13870
rect 35714 13832 35716 13841
rect 37648 13864 37700 13870
rect 35768 13832 35770 13841
rect 37648 13806 37700 13812
rect 35714 13767 35770 13776
rect 36268 13796 36320 13802
rect 36268 13738 36320 13744
rect 35348 13456 35400 13462
rect 34440 13382 34560 13410
rect 35348 13398 35400 13404
rect 33876 13184 33928 13190
rect 33876 13126 33928 13132
rect 33784 12708 33836 12714
rect 33784 12650 33836 12656
rect 33888 12238 33916 13126
rect 34244 12436 34296 12442
rect 34244 12378 34296 12384
rect 33876 12232 33928 12238
rect 33876 12174 33928 12180
rect 33692 11280 33744 11286
rect 33692 11222 33744 11228
rect 33888 11234 33916 12174
rect 34256 11898 34284 12378
rect 34244 11892 34296 11898
rect 34244 11834 34296 11840
rect 34532 11830 34560 13382
rect 36176 13388 36228 13394
rect 36176 13330 36228 13336
rect 36188 13190 36216 13330
rect 36176 13184 36228 13190
rect 36176 13126 36228 13132
rect 34940 13084 35236 13104
rect 34996 13082 35020 13084
rect 35076 13082 35100 13084
rect 35156 13082 35180 13084
rect 35018 13030 35020 13082
rect 35082 13030 35094 13082
rect 35156 13030 35158 13082
rect 34996 13028 35020 13030
rect 35076 13028 35100 13030
rect 35156 13028 35180 13030
rect 34940 13008 35236 13028
rect 34612 12776 34664 12782
rect 34612 12718 34664 12724
rect 34624 12238 34652 12718
rect 35256 12708 35308 12714
rect 35256 12650 35308 12656
rect 35268 12442 35296 12650
rect 35256 12436 35308 12442
rect 35256 12378 35308 12384
rect 34612 12232 34664 12238
rect 34612 12174 34664 12180
rect 34624 11898 34652 12174
rect 34940 11996 35236 12016
rect 34996 11994 35020 11996
rect 35076 11994 35100 11996
rect 35156 11994 35180 11996
rect 35018 11942 35020 11994
rect 35082 11942 35094 11994
rect 35156 11942 35158 11994
rect 34996 11940 35020 11942
rect 35076 11940 35100 11942
rect 35156 11940 35180 11942
rect 34940 11920 35236 11940
rect 35268 11898 35296 12378
rect 34612 11892 34664 11898
rect 34612 11834 34664 11840
rect 35256 11892 35308 11898
rect 35256 11834 35308 11840
rect 34520 11824 34572 11830
rect 34520 11766 34572 11772
rect 36084 11552 36136 11558
rect 36084 11494 36136 11500
rect 34244 11280 34296 11286
rect 33888 11218 34008 11234
rect 34244 11222 34296 11228
rect 33888 11212 34020 11218
rect 33888 11206 33968 11212
rect 33888 10810 33916 11206
rect 33968 11154 34020 11160
rect 34256 10810 34284 11222
rect 35348 11008 35400 11014
rect 35348 10950 35400 10956
rect 34940 10908 35236 10928
rect 34996 10906 35020 10908
rect 35076 10906 35100 10908
rect 35156 10906 35180 10908
rect 35018 10854 35020 10906
rect 35082 10854 35094 10906
rect 35156 10854 35158 10906
rect 34996 10852 35020 10854
rect 35076 10852 35100 10854
rect 35156 10852 35180 10854
rect 34940 10832 35236 10852
rect 33876 10804 33928 10810
rect 33876 10746 33928 10752
rect 34244 10804 34296 10810
rect 34244 10746 34296 10752
rect 34256 10266 34284 10746
rect 34796 10736 34848 10742
rect 34796 10678 34848 10684
rect 34244 10260 34296 10266
rect 34244 10202 34296 10208
rect 33230 10160 33286 10169
rect 33230 10095 33286 10104
rect 34256 9722 34284 10202
rect 34520 10124 34572 10130
rect 34520 10066 34572 10072
rect 34244 9716 34296 9722
rect 34244 9658 34296 9664
rect 34532 9654 34560 10066
rect 34808 9722 34836 10678
rect 35360 10538 35388 10950
rect 35348 10532 35400 10538
rect 35348 10474 35400 10480
rect 35360 10062 35388 10474
rect 35808 10124 35860 10130
rect 35808 10066 35860 10072
rect 35348 10056 35400 10062
rect 35348 9998 35400 10004
rect 34940 9820 35236 9840
rect 34996 9818 35020 9820
rect 35076 9818 35100 9820
rect 35156 9818 35180 9820
rect 35018 9766 35020 9818
rect 35082 9766 35094 9818
rect 35156 9766 35158 9818
rect 34996 9764 35020 9766
rect 35076 9764 35100 9766
rect 35156 9764 35180 9766
rect 34940 9744 35236 9764
rect 34796 9716 34848 9722
rect 34796 9658 34848 9664
rect 34520 9648 34572 9654
rect 34520 9590 34572 9596
rect 35360 9178 35388 9998
rect 35440 9920 35492 9926
rect 35440 9862 35492 9868
rect 35452 9761 35480 9862
rect 35438 9752 35494 9761
rect 35438 9687 35494 9696
rect 35532 9580 35584 9586
rect 35532 9522 35584 9528
rect 35348 9172 35400 9178
rect 35348 9114 35400 9120
rect 34940 8732 35236 8752
rect 34996 8730 35020 8732
rect 35076 8730 35100 8732
rect 35156 8730 35180 8732
rect 35018 8678 35020 8730
rect 35082 8678 35094 8730
rect 35156 8678 35158 8730
rect 34996 8676 35020 8678
rect 35076 8676 35100 8678
rect 35156 8676 35180 8678
rect 34940 8656 35236 8676
rect 35544 8430 35572 9522
rect 35820 9110 35848 10066
rect 35992 9172 36044 9178
rect 35992 9114 36044 9120
rect 35808 9104 35860 9110
rect 35808 9046 35860 9052
rect 36004 8634 36032 9114
rect 35992 8628 36044 8634
rect 35992 8570 36044 8576
rect 35532 8424 35584 8430
rect 35532 8366 35584 8372
rect 34940 7644 35236 7664
rect 34996 7642 35020 7644
rect 35076 7642 35100 7644
rect 35156 7642 35180 7644
rect 35018 7590 35020 7642
rect 35082 7590 35094 7642
rect 35156 7590 35158 7642
rect 34996 7588 35020 7590
rect 35076 7588 35100 7590
rect 35156 7588 35180 7590
rect 34940 7568 35236 7588
rect 33598 7440 33654 7449
rect 33598 7375 33654 7384
rect 33612 7342 33640 7375
rect 33600 7336 33652 7342
rect 33600 7278 33652 7284
rect 33324 6656 33376 6662
rect 33324 6598 33376 6604
rect 33140 6384 33192 6390
rect 33140 6326 33192 6332
rect 33048 5568 33100 5574
rect 33048 5510 33100 5516
rect 33060 5370 33088 5510
rect 33048 5364 33100 5370
rect 33048 5306 33100 5312
rect 33152 4690 33180 6326
rect 33336 6322 33364 6598
rect 33324 6316 33376 6322
rect 33324 6258 33376 6264
rect 33322 6216 33378 6225
rect 33612 6186 33640 7278
rect 33784 7200 33836 7206
rect 33784 7142 33836 7148
rect 33796 6934 33824 7142
rect 33784 6928 33836 6934
rect 33784 6870 33836 6876
rect 34336 6928 34388 6934
rect 34336 6870 34388 6876
rect 33692 6656 33744 6662
rect 33692 6598 33744 6604
rect 33322 6151 33324 6160
rect 33376 6151 33378 6160
rect 33600 6180 33652 6186
rect 33324 6122 33376 6128
rect 33600 6122 33652 6128
rect 33704 5914 33732 6598
rect 33796 6458 33824 6870
rect 33876 6656 33928 6662
rect 33876 6598 33928 6604
rect 33784 6452 33836 6458
rect 33784 6394 33836 6400
rect 33888 6118 33916 6598
rect 33876 6112 33928 6118
rect 33876 6054 33928 6060
rect 33692 5908 33744 5914
rect 33692 5850 33744 5856
rect 34348 5574 34376 6870
rect 35256 6656 35308 6662
rect 35256 6598 35308 6604
rect 34940 6556 35236 6576
rect 34996 6554 35020 6556
rect 35076 6554 35100 6556
rect 35156 6554 35180 6556
rect 35018 6502 35020 6554
rect 35082 6502 35094 6554
rect 35156 6502 35158 6554
rect 34996 6500 35020 6502
rect 35076 6500 35100 6502
rect 35156 6500 35180 6502
rect 34940 6480 35236 6500
rect 35268 6254 35296 6598
rect 35532 6384 35584 6390
rect 35532 6326 35584 6332
rect 35256 6248 35308 6254
rect 35256 6190 35308 6196
rect 35440 5772 35492 5778
rect 35440 5714 35492 5720
rect 34612 5704 34664 5710
rect 34612 5646 34664 5652
rect 33600 5568 33652 5574
rect 33600 5510 33652 5516
rect 34336 5568 34388 5574
rect 34336 5510 34388 5516
rect 33612 4826 33640 5510
rect 34624 5370 34652 5646
rect 34940 5468 35236 5488
rect 34996 5466 35020 5468
rect 35076 5466 35100 5468
rect 35156 5466 35180 5468
rect 35018 5414 35020 5466
rect 35082 5414 35094 5466
rect 35156 5414 35158 5466
rect 34996 5412 35020 5414
rect 35076 5412 35100 5414
rect 35156 5412 35180 5414
rect 34940 5392 35236 5412
rect 35452 5370 35480 5714
rect 35544 5681 35572 6326
rect 35530 5672 35586 5681
rect 35530 5607 35586 5616
rect 34612 5364 34664 5370
rect 34612 5306 34664 5312
rect 35440 5364 35492 5370
rect 35440 5306 35492 5312
rect 34624 5030 34652 5306
rect 34612 5024 34664 5030
rect 34612 4966 34664 4972
rect 33600 4820 33652 4826
rect 33600 4762 33652 4768
rect 33140 4684 33192 4690
rect 33140 4626 33192 4632
rect 33048 4480 33100 4486
rect 33048 4422 33100 4428
rect 32312 4150 32364 4156
rect 32954 4176 33010 4185
rect 33060 4162 33088 4422
rect 33152 4282 33180 4626
rect 33966 4584 34022 4593
rect 33966 4519 34022 4528
rect 33232 4480 33284 4486
rect 33232 4422 33284 4428
rect 33140 4276 33192 4282
rect 33140 4218 33192 4224
rect 33060 4134 33180 4162
rect 32954 4111 33010 4120
rect 32678 4040 32734 4049
rect 32588 4004 32640 4010
rect 32678 3975 32734 3984
rect 32588 3946 32640 3952
rect 32128 3936 32180 3942
rect 32034 3904 32090 3913
rect 32128 3878 32180 3884
rect 32034 3839 32090 3848
rect 31942 3632 31998 3641
rect 31942 3567 31944 3576
rect 31996 3567 31998 3576
rect 31944 3538 31996 3544
rect 31852 3528 31904 3534
rect 31852 3470 31904 3476
rect 32140 3369 32168 3878
rect 32600 3534 32628 3946
rect 32692 3738 32720 3975
rect 33152 3942 33180 4134
rect 33244 4010 33272 4422
rect 33600 4140 33652 4146
rect 33600 4082 33652 4088
rect 33232 4004 33284 4010
rect 33232 3946 33284 3952
rect 33048 3936 33100 3942
rect 33048 3878 33100 3884
rect 33140 3936 33192 3942
rect 33140 3878 33192 3884
rect 33060 3777 33088 3878
rect 33046 3768 33102 3777
rect 32680 3732 32732 3738
rect 33046 3703 33102 3712
rect 32680 3674 32732 3680
rect 32588 3528 32640 3534
rect 32588 3470 32640 3476
rect 32126 3360 32182 3369
rect 32126 3295 32182 3304
rect 32692 3233 32720 3674
rect 32678 3224 32734 3233
rect 31668 3188 31720 3194
rect 32678 3159 32734 3168
rect 31668 3130 31720 3136
rect 31484 2984 31536 2990
rect 31484 2926 31536 2932
rect 30472 2790 30524 2796
rect 31114 2816 31170 2825
rect 31114 2751 31170 2760
rect 30380 2644 30432 2650
rect 30380 2586 30432 2592
rect 31680 480 31708 3130
rect 31760 2916 31812 2922
rect 31760 2858 31812 2864
rect 31772 2650 31800 2858
rect 32692 2650 32720 3159
rect 33140 2848 33192 2854
rect 33046 2816 33102 2825
rect 33244 2836 33272 3946
rect 33612 3194 33640 4082
rect 33980 3942 34008 4519
rect 33968 3936 34020 3942
rect 33968 3878 34020 3884
rect 33980 3738 34008 3878
rect 34518 3768 34574 3777
rect 33968 3732 34020 3738
rect 34518 3703 34520 3712
rect 33968 3674 34020 3680
rect 34572 3703 34574 3712
rect 34520 3674 34572 3680
rect 34520 3392 34572 3398
rect 34520 3334 34572 3340
rect 33600 3188 33652 3194
rect 33600 3130 33652 3136
rect 34244 2916 34296 2922
rect 34244 2858 34296 2864
rect 33192 2808 33272 2836
rect 33140 2790 33192 2796
rect 33046 2751 33102 2760
rect 31760 2644 31812 2650
rect 31760 2586 31812 2592
rect 32680 2644 32732 2650
rect 32680 2586 32732 2592
rect 33060 480 33088 2751
rect 33152 2582 33180 2790
rect 34256 2650 34284 2858
rect 34244 2644 34296 2650
rect 34244 2586 34296 2592
rect 33140 2576 33192 2582
rect 33140 2518 33192 2524
rect 34532 2514 34560 3334
rect 34624 3194 34652 4966
rect 34940 4380 35236 4400
rect 34996 4378 35020 4380
rect 35076 4378 35100 4380
rect 35156 4378 35180 4380
rect 35018 4326 35020 4378
rect 35082 4326 35094 4378
rect 35156 4326 35158 4378
rect 34996 4324 35020 4326
rect 35076 4324 35100 4326
rect 35156 4324 35180 4326
rect 34940 4304 35236 4324
rect 34888 3936 34940 3942
rect 34888 3878 34940 3884
rect 34900 3670 34928 3878
rect 34888 3664 34940 3670
rect 34888 3606 34940 3612
rect 35256 3664 35308 3670
rect 35256 3606 35308 3612
rect 34940 3292 35236 3312
rect 34996 3290 35020 3292
rect 35076 3290 35100 3292
rect 35156 3290 35180 3292
rect 35018 3238 35020 3290
rect 35082 3238 35094 3290
rect 35156 3238 35158 3290
rect 34996 3236 35020 3238
rect 35076 3236 35100 3238
rect 35156 3236 35180 3238
rect 34940 3216 35236 3236
rect 34612 3188 34664 3194
rect 34612 3130 34664 3136
rect 35268 2650 35296 3606
rect 35348 3528 35400 3534
rect 35348 3470 35400 3476
rect 35360 2922 35388 3470
rect 35348 2916 35400 2922
rect 35348 2858 35400 2864
rect 35256 2644 35308 2650
rect 35256 2586 35308 2592
rect 34520 2508 34572 2514
rect 34520 2450 34572 2456
rect 34532 2394 34560 2450
rect 34348 2366 34560 2394
rect 34348 480 34376 2366
rect 35716 2304 35768 2310
rect 35716 2246 35768 2252
rect 34940 2204 35236 2224
rect 34996 2202 35020 2204
rect 35076 2202 35100 2204
rect 35156 2202 35180 2204
rect 35018 2150 35020 2202
rect 35082 2150 35094 2202
rect 35156 2150 35158 2202
rect 34996 2148 35020 2150
rect 35076 2148 35100 2150
rect 35156 2148 35180 2150
rect 34940 2128 35236 2148
rect 35728 480 35756 2246
rect 662 0 718 480
rect 1950 0 2006 480
rect 3330 0 3386 480
rect 4710 0 4766 480
rect 5998 0 6054 480
rect 7378 0 7434 480
rect 8758 0 8814 480
rect 10046 0 10102 480
rect 11426 0 11482 480
rect 12806 0 12862 480
rect 14094 0 14150 480
rect 15474 0 15530 480
rect 16854 0 16910 480
rect 18142 0 18198 480
rect 19522 0 19578 480
rect 20902 0 20958 480
rect 22190 0 22246 480
rect 23570 0 23626 480
rect 24950 0 25006 480
rect 26238 0 26294 480
rect 27618 0 27674 480
rect 28998 0 29054 480
rect 30286 0 30342 480
rect 31666 0 31722 480
rect 33046 0 33102 480
rect 34334 0 34390 480
rect 35714 0 35770 480
rect 36096 105 36124 11494
rect 36188 1465 36216 13126
rect 36280 12986 36308 13738
rect 37372 13728 37424 13734
rect 37372 13670 37424 13676
rect 37384 13326 37412 13670
rect 36636 13320 36688 13326
rect 36636 13262 36688 13268
rect 37372 13320 37424 13326
rect 37372 13262 37424 13268
rect 36268 12980 36320 12986
rect 36268 12922 36320 12928
rect 36360 10464 36412 10470
rect 36360 10406 36412 10412
rect 36372 9450 36400 10406
rect 36360 9444 36412 9450
rect 36360 9386 36412 9392
rect 36372 9178 36400 9386
rect 36452 9376 36504 9382
rect 36452 9318 36504 9324
rect 36360 9172 36412 9178
rect 36360 9114 36412 9120
rect 36464 8974 36492 9318
rect 36452 8968 36504 8974
rect 36452 8910 36504 8916
rect 36464 8412 36492 8910
rect 36544 8424 36596 8430
rect 36464 8384 36544 8412
rect 36464 8090 36492 8384
rect 36544 8366 36596 8372
rect 36648 8276 36676 13262
rect 36912 13184 36964 13190
rect 36912 13126 36964 13132
rect 36924 12782 36952 13126
rect 36820 12776 36872 12782
rect 36820 12718 36872 12724
rect 36912 12776 36964 12782
rect 36912 12718 36964 12724
rect 36832 12374 36860 12718
rect 37188 12708 37240 12714
rect 37188 12650 37240 12656
rect 36820 12368 36872 12374
rect 36820 12310 36872 12316
rect 37200 12186 37228 12650
rect 37660 12374 37688 13806
rect 37844 13258 37872 18362
rect 38396 18086 38424 18702
rect 39132 18086 39160 19110
rect 40236 18970 40264 19314
rect 40420 19174 40448 19654
rect 40604 19514 40632 20198
rect 40592 19508 40644 19514
rect 40592 19450 40644 19456
rect 40408 19168 40460 19174
rect 40408 19110 40460 19116
rect 40224 18964 40276 18970
rect 40224 18906 40276 18912
rect 40224 18828 40276 18834
rect 40224 18770 40276 18776
rect 39948 18760 40000 18766
rect 39948 18702 40000 18708
rect 39960 18426 39988 18702
rect 39948 18420 40000 18426
rect 39948 18362 40000 18368
rect 40236 18358 40264 18770
rect 40420 18612 40448 19110
rect 40696 18766 40724 20334
rect 40788 18970 40816 20703
rect 41340 20584 41368 20742
rect 41420 20596 41472 20602
rect 41340 20556 41420 20584
rect 41420 20538 41472 20544
rect 41604 20324 41656 20330
rect 41604 20266 41656 20272
rect 41616 20058 41644 20266
rect 41604 20052 41656 20058
rect 41604 19994 41656 20000
rect 41892 19292 41920 23718
rect 42260 23662 42288 23802
rect 42248 23656 42300 23662
rect 42248 23598 42300 23604
rect 42616 23656 42668 23662
rect 42616 23598 42668 23604
rect 42628 23322 42656 23598
rect 45480 23526 45508 24142
rect 44088 23520 44140 23526
rect 44088 23462 44140 23468
rect 44640 23520 44692 23526
rect 44640 23462 44692 23468
rect 45468 23520 45520 23526
rect 45468 23462 45520 23468
rect 42616 23316 42668 23322
rect 42616 23258 42668 23264
rect 42628 22778 42656 23258
rect 44100 22982 44128 23462
rect 44652 23118 44680 23462
rect 44916 23180 44968 23186
rect 44916 23122 44968 23128
rect 44640 23112 44692 23118
rect 44640 23054 44692 23060
rect 44088 22976 44140 22982
rect 44088 22918 44140 22924
rect 42616 22772 42668 22778
rect 42616 22714 42668 22720
rect 44100 22506 44128 22918
rect 44652 22574 44680 23054
rect 44928 22778 44956 23122
rect 44916 22772 44968 22778
rect 44916 22714 44968 22720
rect 44640 22568 44692 22574
rect 44640 22510 44692 22516
rect 44088 22500 44140 22506
rect 44140 22460 44220 22488
rect 44088 22442 44140 22448
rect 43904 22160 43956 22166
rect 43904 22102 43956 22108
rect 43444 22092 43496 22098
rect 43444 22034 43496 22040
rect 42340 21888 42392 21894
rect 42340 21830 42392 21836
rect 41972 21548 42024 21554
rect 41972 21490 42024 21496
rect 41800 19264 41920 19292
rect 40960 19236 41012 19242
rect 40960 19178 41012 19184
rect 40776 18964 40828 18970
rect 40776 18906 40828 18912
rect 40684 18760 40736 18766
rect 40684 18702 40736 18708
rect 40500 18624 40552 18630
rect 40420 18584 40500 18612
rect 40224 18352 40276 18358
rect 40224 18294 40276 18300
rect 38384 18080 38436 18086
rect 38384 18022 38436 18028
rect 39120 18080 39172 18086
rect 39120 18022 39172 18028
rect 38660 16992 38712 16998
rect 38660 16934 38712 16940
rect 38568 16720 38620 16726
rect 38672 16708 38700 16934
rect 38620 16680 38700 16708
rect 38568 16662 38620 16668
rect 38292 16584 38344 16590
rect 38292 16526 38344 16532
rect 38304 15910 38332 16526
rect 38672 16250 38700 16680
rect 38660 16244 38712 16250
rect 38660 16186 38712 16192
rect 38672 15978 38700 16186
rect 38660 15972 38712 15978
rect 38660 15914 38712 15920
rect 37924 15904 37976 15910
rect 37924 15846 37976 15852
rect 38292 15904 38344 15910
rect 38292 15846 38344 15852
rect 37936 14958 37964 15846
rect 38672 15706 38700 15914
rect 38660 15700 38712 15706
rect 38660 15642 38712 15648
rect 38200 15632 38252 15638
rect 38200 15574 38252 15580
rect 38212 14958 38240 15574
rect 37924 14952 37976 14958
rect 37924 14894 37976 14900
rect 38200 14952 38252 14958
rect 38200 14894 38252 14900
rect 39132 14618 39160 18022
rect 40040 17060 40092 17066
rect 39960 17020 40040 17048
rect 39396 16788 39448 16794
rect 39396 16730 39448 16736
rect 39408 16114 39436 16730
rect 39960 16250 39988 17020
rect 40040 17002 40092 17008
rect 40420 16590 40448 18584
rect 40500 18566 40552 18572
rect 40788 18426 40816 18906
rect 40972 18766 41000 19178
rect 40960 18760 41012 18766
rect 41012 18720 41092 18748
rect 40960 18702 41012 18708
rect 40776 18420 40828 18426
rect 40776 18362 40828 18368
rect 41064 18086 41092 18720
rect 41142 18592 41198 18601
rect 41142 18527 41198 18536
rect 41052 18080 41104 18086
rect 41052 18022 41104 18028
rect 40408 16584 40460 16590
rect 40408 16526 40460 16532
rect 40776 16584 40828 16590
rect 40776 16526 40828 16532
rect 39948 16244 40000 16250
rect 39948 16186 40000 16192
rect 39396 16108 39448 16114
rect 39396 16050 39448 16056
rect 39408 15706 39436 16050
rect 40788 16046 40816 16526
rect 40776 16040 40828 16046
rect 40776 15982 40828 15988
rect 40868 15972 40920 15978
rect 40868 15914 40920 15920
rect 39396 15700 39448 15706
rect 39396 15642 39448 15648
rect 40776 15700 40828 15706
rect 40776 15642 40828 15648
rect 40788 15162 40816 15642
rect 40880 15502 40908 15914
rect 40868 15496 40920 15502
rect 40868 15438 40920 15444
rect 40776 15156 40828 15162
rect 40776 15098 40828 15104
rect 40880 15094 40908 15438
rect 40868 15088 40920 15094
rect 40868 15030 40920 15036
rect 39304 14816 39356 14822
rect 39304 14758 39356 14764
rect 39120 14612 39172 14618
rect 39120 14554 39172 14560
rect 39316 14550 39344 14758
rect 40880 14550 40908 15030
rect 39304 14544 39356 14550
rect 39304 14486 39356 14492
rect 40868 14544 40920 14550
rect 40868 14486 40920 14492
rect 38292 14476 38344 14482
rect 38292 14418 38344 14424
rect 38304 13734 38332 14418
rect 39316 14074 39344 14486
rect 40684 14408 40736 14414
rect 40684 14350 40736 14356
rect 39304 14068 39356 14074
rect 39304 14010 39356 14016
rect 39212 13796 39264 13802
rect 39212 13738 39264 13744
rect 38292 13728 38344 13734
rect 38292 13670 38344 13676
rect 38108 13456 38160 13462
rect 38108 13398 38160 13404
rect 37832 13252 37884 13258
rect 37832 13194 37884 13200
rect 37648 12368 37700 12374
rect 37648 12310 37700 12316
rect 37280 12232 37332 12238
rect 37200 12180 37280 12186
rect 37200 12174 37332 12180
rect 37200 12158 37320 12174
rect 37200 11370 37228 12158
rect 37660 11762 37688 12310
rect 38120 12170 38148 13398
rect 38304 13326 38332 13670
rect 39224 13326 39252 13738
rect 39316 13462 39344 14010
rect 40040 13932 40092 13938
rect 40040 13874 40092 13880
rect 39304 13456 39356 13462
rect 39304 13398 39356 13404
rect 38200 13320 38252 13326
rect 38200 13262 38252 13268
rect 38292 13320 38344 13326
rect 38292 13262 38344 13268
rect 39212 13320 39264 13326
rect 39212 13262 39264 13268
rect 38212 12986 38240 13262
rect 38200 12980 38252 12986
rect 38200 12922 38252 12928
rect 38200 12640 38252 12646
rect 38304 12628 38332 13262
rect 39224 12918 39252 13262
rect 39316 12986 39344 13398
rect 40052 13002 40080 13874
rect 40696 13802 40724 14350
rect 40684 13796 40736 13802
rect 40684 13738 40736 13744
rect 40696 13530 40724 13738
rect 40684 13524 40736 13530
rect 40684 13466 40736 13472
rect 39304 12980 39356 12986
rect 39304 12922 39356 12928
rect 39960 12974 40080 13002
rect 39960 12918 39988 12974
rect 39212 12912 39264 12918
rect 39212 12854 39264 12860
rect 39948 12912 40000 12918
rect 39948 12854 40000 12860
rect 38252 12600 38332 12628
rect 38200 12582 38252 12588
rect 38212 12442 38240 12582
rect 41064 12442 41092 18022
rect 41156 17882 41184 18527
rect 41144 17876 41196 17882
rect 41144 17818 41196 17824
rect 41604 17536 41656 17542
rect 41604 17478 41656 17484
rect 41616 17202 41644 17478
rect 41328 17196 41380 17202
rect 41328 17138 41380 17144
rect 41604 17196 41656 17202
rect 41604 17138 41656 17144
rect 41236 16040 41288 16046
rect 41236 15982 41288 15988
rect 41248 15706 41276 15982
rect 41236 15700 41288 15706
rect 41236 15642 41288 15648
rect 41144 15632 41196 15638
rect 41144 15574 41196 15580
rect 41156 15162 41184 15574
rect 41340 15366 41368 17138
rect 41420 16788 41472 16794
rect 41420 16730 41472 16736
rect 41432 16046 41460 16730
rect 41420 16040 41472 16046
rect 41420 15982 41472 15988
rect 41328 15360 41380 15366
rect 41328 15302 41380 15308
rect 41144 15156 41196 15162
rect 41144 15098 41196 15104
rect 41800 14958 41828 19264
rect 41984 18426 42012 21490
rect 42352 21146 42380 21830
rect 43456 21690 43484 22034
rect 43444 21684 43496 21690
rect 43444 21626 43496 21632
rect 43168 21616 43220 21622
rect 43168 21558 43220 21564
rect 42800 21480 42852 21486
rect 42800 21422 42852 21428
rect 42340 21140 42392 21146
rect 42340 21082 42392 21088
rect 42352 20482 42380 21082
rect 42812 20602 42840 21422
rect 43180 21146 43208 21558
rect 43456 21146 43484 21626
rect 43916 21622 43944 22102
rect 43904 21616 43956 21622
rect 43904 21558 43956 21564
rect 44192 21554 44220 22460
rect 44928 22166 44956 22714
rect 45100 22500 45152 22506
rect 45100 22442 45152 22448
rect 45112 22234 45140 22442
rect 45560 22432 45612 22438
rect 45480 22380 45560 22386
rect 45480 22374 45612 22380
rect 45480 22358 45600 22374
rect 45100 22228 45152 22234
rect 45100 22170 45152 22176
rect 44916 22160 44968 22166
rect 44916 22102 44968 22108
rect 44928 21690 44956 22102
rect 44916 21684 44968 21690
rect 44916 21626 44968 21632
rect 44180 21548 44232 21554
rect 44180 21490 44232 21496
rect 44088 21412 44140 21418
rect 44088 21354 44140 21360
rect 44100 21146 44128 21354
rect 44180 21344 44232 21350
rect 44180 21286 44232 21292
rect 43168 21140 43220 21146
rect 43168 21082 43220 21088
rect 43444 21140 43496 21146
rect 43444 21082 43496 21088
rect 44088 21140 44140 21146
rect 44088 21082 44140 21088
rect 44100 20754 44128 21082
rect 44192 21010 44220 21286
rect 44640 21072 44692 21078
rect 44640 21014 44692 21020
rect 44180 21004 44232 21010
rect 44180 20946 44232 20952
rect 44192 20806 44220 20946
rect 44008 20726 44128 20754
rect 44180 20800 44232 20806
rect 44180 20742 44232 20748
rect 42800 20596 42852 20602
rect 42800 20538 42852 20544
rect 42352 20466 42472 20482
rect 44008 20466 44036 20726
rect 44192 20618 44220 20742
rect 44100 20602 44220 20618
rect 44100 20596 44232 20602
rect 44100 20590 44180 20596
rect 42352 20460 42484 20466
rect 42352 20454 42432 20460
rect 42432 20402 42484 20408
rect 42984 20460 43036 20466
rect 42984 20402 43036 20408
rect 43996 20460 44048 20466
rect 43996 20402 44048 20408
rect 42248 20392 42300 20398
rect 42248 20334 42300 20340
rect 42260 20058 42288 20334
rect 42248 20052 42300 20058
rect 42248 19994 42300 20000
rect 42996 19990 43024 20402
rect 42156 19984 42208 19990
rect 42156 19926 42208 19932
rect 42984 19984 43036 19990
rect 42984 19926 43036 19932
rect 42168 19242 42196 19926
rect 43720 19848 43772 19854
rect 43720 19790 43772 19796
rect 43732 19514 43760 19790
rect 43720 19508 43772 19514
rect 43720 19450 43772 19456
rect 44100 19310 44128 20590
rect 44180 20538 44232 20544
rect 44192 20507 44220 20538
rect 44652 20534 44680 21014
rect 45100 20936 45152 20942
rect 45100 20878 45152 20884
rect 44640 20528 44692 20534
rect 44640 20470 44692 20476
rect 45112 20058 45140 20878
rect 45480 20874 45508 22358
rect 45560 22092 45612 22098
rect 45560 22034 45612 22040
rect 45572 21690 45600 22034
rect 45560 21684 45612 21690
rect 45560 21626 45612 21632
rect 45468 20868 45520 20874
rect 45468 20810 45520 20816
rect 45940 20641 45968 30330
rect 46020 25424 46072 25430
rect 46020 25366 46072 25372
rect 46032 24682 46060 25366
rect 46124 25265 46152 44270
rect 46296 40112 46348 40118
rect 46296 40054 46348 40060
rect 46204 30592 46256 30598
rect 46204 30534 46256 30540
rect 46216 30190 46244 30534
rect 46204 30184 46256 30190
rect 46204 30126 46256 30132
rect 46216 28082 46244 30126
rect 46204 28076 46256 28082
rect 46204 28018 46256 28024
rect 46204 27532 46256 27538
rect 46204 27474 46256 27480
rect 46216 27130 46244 27474
rect 46204 27124 46256 27130
rect 46204 27066 46256 27072
rect 46216 25838 46244 27066
rect 46204 25832 46256 25838
rect 46204 25774 46256 25780
rect 46110 25256 46166 25265
rect 46110 25191 46166 25200
rect 46020 24676 46072 24682
rect 46020 24618 46072 24624
rect 46032 24274 46060 24618
rect 46020 24268 46072 24274
rect 46020 24210 46072 24216
rect 46032 23526 46060 24210
rect 46020 23520 46072 23526
rect 46020 23462 46072 23468
rect 46032 23322 46060 23462
rect 46020 23316 46072 23322
rect 46020 23258 46072 23264
rect 46308 22778 46336 40054
rect 46388 28620 46440 28626
rect 46388 28562 46440 28568
rect 46400 28014 46428 28562
rect 46388 28008 46440 28014
rect 46388 27950 46440 27956
rect 46676 27169 46704 44934
rect 46952 44538 46980 45070
rect 47398 44568 47454 44577
rect 46940 44532 46992 44538
rect 47398 44503 47400 44512
rect 46940 44474 46992 44480
rect 47452 44503 47454 44512
rect 47400 44474 47452 44480
rect 47412 44334 47440 44474
rect 47400 44328 47452 44334
rect 47400 44270 47452 44276
rect 46938 42936 46994 42945
rect 46938 42871 46994 42880
rect 46952 41818 46980 42871
rect 46940 41812 46992 41818
rect 46940 41754 46992 41760
rect 46756 41676 46808 41682
rect 46756 41618 46808 41624
rect 46768 41449 46796 41618
rect 46754 41440 46810 41449
rect 46754 41375 46810 41384
rect 46768 40934 46796 41375
rect 46756 40928 46808 40934
rect 46756 40870 46808 40876
rect 46768 40118 46796 40870
rect 46756 40112 46808 40118
rect 46756 40054 46808 40060
rect 46938 39808 46994 39817
rect 46938 39743 46994 39752
rect 46952 38554 46980 39743
rect 46940 38548 46992 38554
rect 46940 38490 46992 38496
rect 46756 38412 46808 38418
rect 46756 38354 46808 38360
rect 46768 38321 46796 38354
rect 46754 38312 46810 38321
rect 46754 38247 46810 38256
rect 46768 37670 46796 38247
rect 46756 37664 46808 37670
rect 46756 37606 46808 37612
rect 46938 36680 46994 36689
rect 46938 36615 46994 36624
rect 46952 35290 46980 36615
rect 46940 35284 46992 35290
rect 46940 35226 46992 35232
rect 46754 35184 46810 35193
rect 46754 35119 46756 35128
rect 46808 35119 46810 35128
rect 46756 35090 46808 35096
rect 46768 34746 46796 35090
rect 46756 34740 46808 34746
rect 46756 34682 46808 34688
rect 46768 34082 46796 34682
rect 46768 34054 46888 34082
rect 46754 32056 46810 32065
rect 46754 31991 46810 32000
rect 46768 31890 46796 31991
rect 46756 31884 46808 31890
rect 46756 31826 46808 31832
rect 46768 31142 46796 31826
rect 46756 31136 46808 31142
rect 46756 31078 46808 31084
rect 46768 30394 46796 31078
rect 46756 30388 46808 30394
rect 46756 30330 46808 30336
rect 46662 27160 46718 27169
rect 46662 27095 46718 27104
rect 46860 26874 46888 34054
rect 46938 33552 46994 33561
rect 46938 33487 46994 33496
rect 46952 32026 46980 33487
rect 46940 32020 46992 32026
rect 46940 31962 46992 31968
rect 47214 30696 47270 30705
rect 47214 30631 47216 30640
rect 47268 30631 47270 30640
rect 47216 30602 47268 30608
rect 46938 30424 46994 30433
rect 46938 30359 46994 30368
rect 46952 29306 46980 30359
rect 47492 30048 47544 30054
rect 47492 29990 47544 29996
rect 47504 29782 47532 29990
rect 47492 29776 47544 29782
rect 47492 29718 47544 29724
rect 46940 29300 46992 29306
rect 46940 29242 46992 29248
rect 47308 29028 47360 29034
rect 47308 28970 47360 28976
rect 47320 28937 47348 28970
rect 47306 28928 47362 28937
rect 47306 28863 47362 28872
rect 47492 28416 47544 28422
rect 47492 28358 47544 28364
rect 47504 28082 47532 28358
rect 47492 28076 47544 28082
rect 47492 28018 47544 28024
rect 46940 28008 46992 28014
rect 46940 27950 46992 27956
rect 46952 27674 46980 27950
rect 47400 27940 47452 27946
rect 47400 27882 47452 27888
rect 46940 27668 46992 27674
rect 46940 27610 46992 27616
rect 46938 27296 46994 27305
rect 46938 27231 46994 27240
rect 46492 26846 46888 26874
rect 46388 25152 46440 25158
rect 46388 25094 46440 25100
rect 46400 24682 46428 25094
rect 46388 24676 46440 24682
rect 46388 24618 46440 24624
rect 46296 22772 46348 22778
rect 46296 22714 46348 22720
rect 46112 22568 46164 22574
rect 46112 22510 46164 22516
rect 46124 22030 46152 22510
rect 46112 22024 46164 22030
rect 46112 21966 46164 21972
rect 46124 21554 46152 21966
rect 46112 21548 46164 21554
rect 46112 21490 46164 21496
rect 46124 21146 46152 21490
rect 46388 21412 46440 21418
rect 46388 21354 46440 21360
rect 46112 21140 46164 21146
rect 46112 21082 46164 21088
rect 45926 20632 45982 20641
rect 45926 20567 45982 20576
rect 45100 20052 45152 20058
rect 45100 19994 45152 20000
rect 45008 19916 45060 19922
rect 45008 19858 45060 19864
rect 44732 19848 44784 19854
rect 44732 19790 44784 19796
rect 44180 19712 44232 19718
rect 44180 19654 44232 19660
rect 44192 19378 44220 19654
rect 44180 19372 44232 19378
rect 44180 19314 44232 19320
rect 44088 19304 44140 19310
rect 44088 19246 44140 19252
rect 42156 19236 42208 19242
rect 42156 19178 42208 19184
rect 42168 18970 42196 19178
rect 44744 19174 44772 19790
rect 45020 19378 45048 19858
rect 45008 19372 45060 19378
rect 45008 19314 45060 19320
rect 43444 19168 43496 19174
rect 43444 19110 43496 19116
rect 44732 19168 44784 19174
rect 44732 19110 44784 19116
rect 42156 18964 42208 18970
rect 42156 18906 42208 18912
rect 42892 18624 42944 18630
rect 42890 18592 42892 18601
rect 42944 18592 42946 18601
rect 42890 18527 42946 18536
rect 41972 18420 42024 18426
rect 41972 18362 42024 18368
rect 42904 18290 42932 18527
rect 42892 18284 42944 18290
rect 42892 18226 42944 18232
rect 43260 18148 43312 18154
rect 43260 18090 43312 18096
rect 42984 18080 43036 18086
rect 42984 18022 43036 18028
rect 42064 17740 42116 17746
rect 42064 17682 42116 17688
rect 42076 17338 42104 17682
rect 42616 17672 42668 17678
rect 42616 17614 42668 17620
rect 42248 17536 42300 17542
rect 42248 17478 42300 17484
rect 42064 17332 42116 17338
rect 42064 17274 42116 17280
rect 42260 16726 42288 17478
rect 42628 17377 42656 17614
rect 42614 17368 42670 17377
rect 42996 17338 43024 18022
rect 43168 17808 43220 17814
rect 43168 17750 43220 17756
rect 42614 17303 42616 17312
rect 42668 17303 42670 17312
rect 42984 17332 43036 17338
rect 42616 17274 42668 17280
rect 42984 17274 43036 17280
rect 42996 17134 43024 17274
rect 42708 17128 42760 17134
rect 42708 17070 42760 17076
rect 42984 17128 43036 17134
rect 42984 17070 43036 17076
rect 42248 16720 42300 16726
rect 42248 16662 42300 16668
rect 42064 15904 42116 15910
rect 42064 15846 42116 15852
rect 42246 15872 42302 15881
rect 42076 15638 42104 15846
rect 42246 15807 42302 15816
rect 42064 15632 42116 15638
rect 42064 15574 42116 15580
rect 41420 14952 41472 14958
rect 41420 14894 41472 14900
rect 41788 14952 41840 14958
rect 41788 14894 41840 14900
rect 41328 13864 41380 13870
rect 41328 13806 41380 13812
rect 41340 12646 41368 13806
rect 41328 12640 41380 12646
rect 41328 12582 41380 12588
rect 38200 12436 38252 12442
rect 38200 12378 38252 12384
rect 41052 12436 41104 12442
rect 41052 12378 41104 12384
rect 38568 12368 38620 12374
rect 38568 12310 38620 12316
rect 39764 12368 39816 12374
rect 39764 12310 39816 12316
rect 38384 12300 38436 12306
rect 38384 12242 38436 12248
rect 38108 12164 38160 12170
rect 38108 12106 38160 12112
rect 37648 11756 37700 11762
rect 37648 11698 37700 11704
rect 37200 11354 37320 11370
rect 38396 11354 38424 12242
rect 38580 11354 38608 12310
rect 39028 12232 39080 12238
rect 39028 12174 39080 12180
rect 39040 11898 39068 12174
rect 39672 12096 39724 12102
rect 39672 12038 39724 12044
rect 39028 11892 39080 11898
rect 39028 11834 39080 11840
rect 37200 11348 37332 11354
rect 37200 11342 37280 11348
rect 37280 11290 37332 11296
rect 38384 11348 38436 11354
rect 38384 11290 38436 11296
rect 38568 11348 38620 11354
rect 38568 11290 38620 11296
rect 39684 11218 39712 12038
rect 39776 11898 39804 12310
rect 40040 12232 40092 12238
rect 40040 12174 40092 12180
rect 40224 12232 40276 12238
rect 40224 12174 40276 12180
rect 40052 11898 40080 12174
rect 39764 11892 39816 11898
rect 39764 11834 39816 11840
rect 40040 11892 40092 11898
rect 40040 11834 40092 11840
rect 37740 11212 37792 11218
rect 37740 11154 37792 11160
rect 39672 11212 39724 11218
rect 39672 11154 39724 11160
rect 37752 10810 37780 11154
rect 39580 11008 39632 11014
rect 39580 10950 39632 10956
rect 37740 10804 37792 10810
rect 37740 10746 37792 10752
rect 37832 10600 37884 10606
rect 37832 10542 37884 10548
rect 37740 10192 37792 10198
rect 37740 10134 37792 10140
rect 37752 9761 37780 10134
rect 37844 9994 37872 10542
rect 39592 10538 39620 10950
rect 39684 10810 39712 11154
rect 39672 10804 39724 10810
rect 39672 10746 39724 10752
rect 39776 10742 39804 11834
rect 40236 11082 40264 12174
rect 40868 12096 40920 12102
rect 40868 12038 40920 12044
rect 40880 11626 40908 12038
rect 40868 11620 40920 11626
rect 40868 11562 40920 11568
rect 40880 11354 40908 11562
rect 41144 11552 41196 11558
rect 41144 11494 41196 11500
rect 40868 11348 40920 11354
rect 40868 11290 40920 11296
rect 40960 11212 41012 11218
rect 40960 11154 41012 11160
rect 40224 11076 40276 11082
rect 40224 11018 40276 11024
rect 40592 11076 40644 11082
rect 40592 11018 40644 11024
rect 39764 10736 39816 10742
rect 39764 10678 39816 10684
rect 39212 10532 39264 10538
rect 39212 10474 39264 10480
rect 39580 10532 39632 10538
rect 39580 10474 39632 10480
rect 39224 10266 39252 10474
rect 39212 10260 39264 10266
rect 39212 10202 39264 10208
rect 39592 10198 39620 10474
rect 40604 10266 40632 11018
rect 40972 10810 41000 11154
rect 40960 10804 41012 10810
rect 40960 10746 41012 10752
rect 40972 10305 41000 10746
rect 40958 10296 41014 10305
rect 40592 10260 40644 10266
rect 40958 10231 41014 10240
rect 40592 10202 40644 10208
rect 39580 10192 39632 10198
rect 39580 10134 39632 10140
rect 41156 10130 41184 11494
rect 41340 11286 41368 12582
rect 41328 11280 41380 11286
rect 41328 11222 41380 11228
rect 41340 10742 41368 11222
rect 41328 10736 41380 10742
rect 41328 10678 41380 10684
rect 38108 10124 38160 10130
rect 38108 10066 38160 10072
rect 39304 10124 39356 10130
rect 39304 10066 39356 10072
rect 40776 10124 40828 10130
rect 40776 10066 40828 10072
rect 41144 10124 41196 10130
rect 41144 10066 41196 10072
rect 37832 9988 37884 9994
rect 37832 9930 37884 9936
rect 37738 9752 37794 9761
rect 37738 9687 37740 9696
rect 37792 9687 37794 9696
rect 37740 9658 37792 9664
rect 38120 9382 38148 10066
rect 38568 10056 38620 10062
rect 38568 9998 38620 10004
rect 38580 9382 38608 9998
rect 39316 9382 39344 10066
rect 40788 9722 40816 10066
rect 41432 9722 41460 14894
rect 41972 14884 42024 14890
rect 41972 14826 42024 14832
rect 41788 14816 41840 14822
rect 41788 14758 41840 14764
rect 41800 14074 41828 14758
rect 41984 14618 42012 14826
rect 42260 14618 42288 15807
rect 42352 15366 42380 15397
rect 42340 15360 42392 15366
rect 42338 15328 42340 15337
rect 42392 15328 42394 15337
rect 42338 15263 42394 15272
rect 42352 14958 42380 15263
rect 42720 15178 42748 17070
rect 42996 16794 43024 17070
rect 42984 16788 43036 16794
rect 42984 16730 43036 16736
rect 43180 16658 43208 17750
rect 43272 17542 43300 18090
rect 43456 17610 43484 19110
rect 45020 18970 45048 19314
rect 46124 19174 46152 21082
rect 46400 20942 46428 21354
rect 46388 20936 46440 20942
rect 46388 20878 46440 20884
rect 46492 19281 46520 26846
rect 46848 26444 46900 26450
rect 46848 26386 46900 26392
rect 46860 25702 46888 26386
rect 46848 25696 46900 25702
rect 46848 25638 46900 25644
rect 46756 25356 46808 25362
rect 46756 25298 46808 25304
rect 46768 23089 46796 25298
rect 46860 25158 46888 25638
rect 46952 25498 46980 27231
rect 47030 26752 47086 26761
rect 47030 26687 47086 26696
rect 46940 25492 46992 25498
rect 46940 25434 46992 25440
rect 46848 25152 46900 25158
rect 46900 25100 46980 25106
rect 46848 25094 46980 25100
rect 46860 25078 46980 25094
rect 46848 24676 46900 24682
rect 46848 24618 46900 24624
rect 46860 24410 46888 24618
rect 46952 24614 46980 25078
rect 46940 24608 46992 24614
rect 46940 24550 46992 24556
rect 46848 24404 46900 24410
rect 46848 24346 46900 24352
rect 47044 23322 47072 26687
rect 47214 26344 47270 26353
rect 47214 26279 47270 26288
rect 47032 23316 47084 23322
rect 47032 23258 47084 23264
rect 46754 23080 46810 23089
rect 46754 23015 46810 23024
rect 46664 22976 46716 22982
rect 46664 22918 46716 22924
rect 46940 22976 46992 22982
rect 46940 22918 46992 22924
rect 46676 22642 46704 22918
rect 46664 22636 46716 22642
rect 46664 22578 46716 22584
rect 46848 22636 46900 22642
rect 46848 22578 46900 22584
rect 46860 22098 46888 22578
rect 46952 22438 46980 22918
rect 46940 22432 46992 22438
rect 46940 22374 46992 22380
rect 46848 22092 46900 22098
rect 46848 22034 46900 22040
rect 46860 21690 46888 22034
rect 46848 21684 46900 21690
rect 46848 21626 46900 21632
rect 47228 21146 47256 26279
rect 47306 25800 47362 25809
rect 47306 25735 47362 25744
rect 47320 25362 47348 25735
rect 47412 25702 47440 27882
rect 47492 26240 47544 26246
rect 47492 26182 47544 26188
rect 47504 25838 47532 26182
rect 47492 25832 47544 25838
rect 47492 25774 47544 25780
rect 47400 25696 47452 25702
rect 47400 25638 47452 25644
rect 47308 25356 47360 25362
rect 47308 25298 47360 25304
rect 47412 25294 47440 25638
rect 47400 25288 47452 25294
rect 47400 25230 47452 25236
rect 47308 23180 47360 23186
rect 47308 23122 47360 23128
rect 47320 22710 47348 23122
rect 47308 22704 47360 22710
rect 47306 22672 47308 22681
rect 47360 22672 47362 22681
rect 47306 22607 47362 22616
rect 47216 21140 47268 21146
rect 47216 21082 47268 21088
rect 46754 21040 46810 21049
rect 46754 20975 46756 20984
rect 46808 20975 46810 20984
rect 46756 20946 46808 20952
rect 46768 20602 46796 20946
rect 46756 20596 46808 20602
rect 46756 20538 46808 20544
rect 47412 20058 47440 25230
rect 47490 21992 47546 22001
rect 47490 21927 47492 21936
rect 47544 21927 47546 21936
rect 47492 21898 47544 21904
rect 47400 20052 47452 20058
rect 47400 19994 47452 20000
rect 47308 19916 47360 19922
rect 47308 19858 47360 19864
rect 47320 19553 47348 19858
rect 47306 19544 47362 19553
rect 47306 19479 47308 19488
rect 47360 19479 47362 19488
rect 47308 19450 47360 19456
rect 46478 19272 46534 19281
rect 46478 19207 46534 19216
rect 46112 19168 46164 19174
rect 46112 19110 46164 19116
rect 45008 18964 45060 18970
rect 45008 18906 45060 18912
rect 44364 18828 44416 18834
rect 44364 18770 44416 18776
rect 45560 18828 45612 18834
rect 45560 18770 45612 18776
rect 43628 18760 43680 18766
rect 43628 18702 43680 18708
rect 43640 18426 43668 18702
rect 44376 18465 44404 18770
rect 44362 18456 44418 18465
rect 43628 18420 43680 18426
rect 43628 18362 43680 18368
rect 43996 18420 44048 18426
rect 45572 18426 45600 18770
rect 46124 18766 46152 19110
rect 46940 18828 46992 18834
rect 46940 18770 46992 18776
rect 46112 18760 46164 18766
rect 46112 18702 46164 18708
rect 46124 18426 46152 18702
rect 44362 18391 44364 18400
rect 43996 18362 44048 18368
rect 44416 18391 44418 18400
rect 45560 18420 45612 18426
rect 44364 18362 44416 18368
rect 45560 18362 45612 18368
rect 46112 18420 46164 18426
rect 46112 18362 46164 18368
rect 44008 17814 44036 18362
rect 44088 18352 44140 18358
rect 44088 18294 44140 18300
rect 44100 17882 44128 18294
rect 46124 17882 46152 18362
rect 46388 18148 46440 18154
rect 46388 18090 46440 18096
rect 44088 17876 44140 17882
rect 44088 17818 44140 17824
rect 46112 17876 46164 17882
rect 46112 17818 46164 17824
rect 43996 17808 44048 17814
rect 43996 17750 44048 17756
rect 43720 17740 43772 17746
rect 43720 17682 43772 17688
rect 43444 17604 43496 17610
rect 43444 17546 43496 17552
rect 43260 17536 43312 17542
rect 43260 17478 43312 17484
rect 43168 16652 43220 16658
rect 43168 16594 43220 16600
rect 43168 15904 43220 15910
rect 43168 15846 43220 15852
rect 43076 15632 43128 15638
rect 43076 15574 43128 15580
rect 42720 15150 42840 15178
rect 43088 15162 43116 15574
rect 42524 15088 42576 15094
rect 42524 15030 42576 15036
rect 42340 14952 42392 14958
rect 42340 14894 42392 14900
rect 41972 14612 42024 14618
rect 41972 14554 42024 14560
rect 42248 14612 42300 14618
rect 42248 14554 42300 14560
rect 42536 14482 42564 15030
rect 42812 14958 42840 15150
rect 43076 15156 43128 15162
rect 43076 15098 43128 15104
rect 42800 14952 42852 14958
rect 42800 14894 42852 14900
rect 42616 14816 42668 14822
rect 42616 14758 42668 14764
rect 42524 14476 42576 14482
rect 42524 14418 42576 14424
rect 42536 14074 42564 14418
rect 42628 14346 42656 14758
rect 42800 14544 42852 14550
rect 42800 14486 42852 14492
rect 43076 14544 43128 14550
rect 43076 14486 43128 14492
rect 42616 14340 42668 14346
rect 42616 14282 42668 14288
rect 41788 14068 41840 14074
rect 41788 14010 41840 14016
rect 42524 14068 42576 14074
rect 42524 14010 42576 14016
rect 41512 12844 41564 12850
rect 41512 12786 41564 12792
rect 41524 12646 41552 12786
rect 41800 12782 41828 14010
rect 42812 13462 42840 14486
rect 43088 14074 43116 14486
rect 43180 14346 43208 15846
rect 43272 15434 43300 17478
rect 43732 17338 43760 17682
rect 44100 17338 44128 17818
rect 45744 17808 45796 17814
rect 45744 17750 45796 17756
rect 45560 17740 45612 17746
rect 45560 17682 45612 17688
rect 45284 17536 45336 17542
rect 45284 17478 45336 17484
rect 43720 17332 43772 17338
rect 43720 17274 43772 17280
rect 44088 17332 44140 17338
rect 44088 17274 44140 17280
rect 44548 17128 44600 17134
rect 44548 17070 44600 17076
rect 44180 16992 44232 16998
rect 44180 16934 44232 16940
rect 43812 16720 43864 16726
rect 43812 16662 43864 16668
rect 43720 16652 43772 16658
rect 43720 16594 43772 16600
rect 43444 15904 43496 15910
rect 43732 15881 43760 16594
rect 43824 16250 43852 16662
rect 43996 16584 44048 16590
rect 43996 16526 44048 16532
rect 43812 16244 43864 16250
rect 43812 16186 43864 16192
rect 44008 16114 44036 16526
rect 43996 16108 44048 16114
rect 43996 16050 44048 16056
rect 43444 15846 43496 15852
rect 43718 15872 43774 15881
rect 43456 15706 43484 15846
rect 43718 15807 43774 15816
rect 43444 15700 43496 15706
rect 43444 15642 43496 15648
rect 44008 15502 44036 16050
rect 44192 15858 44220 16934
rect 44560 16454 44588 17070
rect 45296 16794 45324 17478
rect 45572 17338 45600 17682
rect 45560 17332 45612 17338
rect 45560 17274 45612 17280
rect 45756 17066 45784 17750
rect 46124 17338 46152 17818
rect 46400 17746 46428 18090
rect 46952 18086 46980 18770
rect 47492 18624 47544 18630
rect 47492 18566 47544 18572
rect 47504 18465 47532 18566
rect 47490 18456 47546 18465
rect 47490 18391 47546 18400
rect 46940 18080 46992 18086
rect 46940 18022 46992 18028
rect 46754 17912 46810 17921
rect 46754 17847 46810 17856
rect 46768 17814 46796 17847
rect 46952 17814 46980 18022
rect 46756 17808 46808 17814
rect 46756 17750 46808 17756
rect 46940 17808 46992 17814
rect 46940 17750 46992 17756
rect 46388 17740 46440 17746
rect 46388 17682 46440 17688
rect 46400 17338 46428 17682
rect 46480 17604 46532 17610
rect 46480 17546 46532 17552
rect 46112 17332 46164 17338
rect 46112 17274 46164 17280
rect 46388 17332 46440 17338
rect 46388 17274 46440 17280
rect 45744 17060 45796 17066
rect 45744 17002 45796 17008
rect 45284 16788 45336 16794
rect 45284 16730 45336 16736
rect 44548 16448 44600 16454
rect 44548 16390 44600 16396
rect 44560 16250 44588 16390
rect 44548 16244 44600 16250
rect 44548 16186 44600 16192
rect 45296 16114 45324 16730
rect 46124 16726 46152 17274
rect 45560 16720 45612 16726
rect 45560 16662 45612 16668
rect 46112 16720 46164 16726
rect 46112 16662 46164 16668
rect 46492 16674 46520 17546
rect 46572 17060 46624 17066
rect 46572 17002 46624 17008
rect 46584 16794 46612 17002
rect 46768 16794 46796 17750
rect 47124 17536 47176 17542
rect 47124 17478 47176 17484
rect 47136 17377 47164 17478
rect 47122 17368 47178 17377
rect 47122 17303 47178 17312
rect 46572 16788 46624 16794
rect 46572 16730 46624 16736
rect 46756 16788 46808 16794
rect 46756 16730 46808 16736
rect 45468 16652 45520 16658
rect 45468 16594 45520 16600
rect 45284 16108 45336 16114
rect 45284 16050 45336 16056
rect 45480 15994 45508 16594
rect 45572 16250 45600 16662
rect 45560 16244 45612 16250
rect 45560 16186 45612 16192
rect 45480 15978 45600 15994
rect 44548 15972 44600 15978
rect 44548 15914 44600 15920
rect 45480 15972 45612 15978
rect 45480 15966 45560 15972
rect 44272 15904 44324 15910
rect 44100 15830 44220 15858
rect 44270 15872 44272 15881
rect 44324 15872 44326 15881
rect 44100 15638 44128 15830
rect 44270 15807 44326 15816
rect 44560 15706 44588 15914
rect 44824 15904 44876 15910
rect 44824 15846 44876 15852
rect 44180 15700 44232 15706
rect 44180 15642 44232 15648
rect 44548 15700 44600 15706
rect 44548 15642 44600 15648
rect 44088 15632 44140 15638
rect 44088 15574 44140 15580
rect 43996 15496 44048 15502
rect 43996 15438 44048 15444
rect 43260 15428 43312 15434
rect 43260 15370 43312 15376
rect 44008 15201 44036 15438
rect 43994 15192 44050 15201
rect 44192 15162 44220 15642
rect 44836 15366 44864 15846
rect 45480 15706 45508 15966
rect 45560 15914 45612 15920
rect 45468 15700 45520 15706
rect 45468 15642 45520 15648
rect 46124 15570 46152 16662
rect 46492 16646 46612 16674
rect 46584 15978 46612 16646
rect 46846 16416 46902 16425
rect 46846 16351 46902 16360
rect 46572 15972 46624 15978
rect 46572 15914 46624 15920
rect 46388 15904 46440 15910
rect 46388 15846 46440 15852
rect 46400 15570 46428 15846
rect 46112 15564 46164 15570
rect 46112 15506 46164 15512
rect 46388 15564 46440 15570
rect 46388 15506 46440 15512
rect 44824 15360 44876 15366
rect 44824 15302 44876 15308
rect 43994 15127 44050 15136
rect 44180 15156 44232 15162
rect 43260 14952 43312 14958
rect 43260 14894 43312 14900
rect 43168 14340 43220 14346
rect 43168 14282 43220 14288
rect 43076 14068 43128 14074
rect 43076 14010 43128 14016
rect 43272 13530 43300 14894
rect 44008 14618 44036 15127
rect 44180 15098 44232 15104
rect 44836 14958 44864 15302
rect 46124 15162 46152 15506
rect 46112 15156 46164 15162
rect 46112 15098 46164 15104
rect 44456 14952 44508 14958
rect 44456 14894 44508 14900
rect 44824 14952 44876 14958
rect 44824 14894 44876 14900
rect 43996 14612 44048 14618
rect 43996 14554 44048 14560
rect 44468 14550 44496 14894
rect 46400 14890 46428 15506
rect 46584 15337 46612 15914
rect 46570 15328 46626 15337
rect 46570 15263 46626 15272
rect 46388 14884 46440 14890
rect 46388 14826 46440 14832
rect 44088 14544 44140 14550
rect 44088 14486 44140 14492
rect 44456 14544 44508 14550
rect 44456 14486 44508 14492
rect 43628 14272 43680 14278
rect 43628 14214 43680 14220
rect 43640 13870 43668 14214
rect 43628 13864 43680 13870
rect 43628 13806 43680 13812
rect 43352 13728 43404 13734
rect 43352 13670 43404 13676
rect 43260 13524 43312 13530
rect 43260 13466 43312 13472
rect 42800 13456 42852 13462
rect 42800 13398 42852 13404
rect 42812 12918 42840 13398
rect 43364 13326 43392 13670
rect 43352 13320 43404 13326
rect 43352 13262 43404 13268
rect 43364 12986 43392 13262
rect 44100 12986 44128 14486
rect 44272 14408 44324 14414
rect 44272 14350 44324 14356
rect 44284 14074 44312 14350
rect 46584 14278 46612 15263
rect 46860 15162 46888 16351
rect 47492 16040 47544 16046
rect 47492 15982 47544 15988
rect 47504 15706 47532 15982
rect 47492 15700 47544 15706
rect 47492 15642 47544 15648
rect 46938 15192 46994 15201
rect 46848 15156 46900 15162
rect 46938 15127 46994 15136
rect 46848 15098 46900 15104
rect 46860 14958 46888 15098
rect 46952 15094 46980 15127
rect 46940 15088 46992 15094
rect 46940 15030 46992 15036
rect 46848 14952 46900 14958
rect 46848 14894 46900 14900
rect 46848 14816 46900 14822
rect 47214 14784 47270 14793
rect 46900 14764 46980 14770
rect 46848 14758 46980 14764
rect 46860 14742 46980 14758
rect 46756 14340 46808 14346
rect 46756 14282 46808 14288
rect 46572 14272 46624 14278
rect 46572 14214 46624 14220
rect 44272 14068 44324 14074
rect 44272 14010 44324 14016
rect 46584 13870 46612 14214
rect 46768 13938 46796 14282
rect 46756 13932 46808 13938
rect 46756 13874 46808 13880
rect 45468 13864 45520 13870
rect 45468 13806 45520 13812
rect 46572 13864 46624 13870
rect 46572 13806 46624 13812
rect 44732 13796 44784 13802
rect 44732 13738 44784 13744
rect 44744 13530 44772 13738
rect 44916 13728 44968 13734
rect 44916 13670 44968 13676
rect 44732 13524 44784 13530
rect 44732 13466 44784 13472
rect 43352 12980 43404 12986
rect 43352 12922 43404 12928
rect 44088 12980 44140 12986
rect 44088 12922 44140 12928
rect 42800 12912 42852 12918
rect 42800 12854 42852 12860
rect 43364 12782 43392 12922
rect 44548 12844 44600 12850
rect 44548 12786 44600 12792
rect 41788 12776 41840 12782
rect 41788 12718 41840 12724
rect 43352 12776 43404 12782
rect 43352 12718 43404 12724
rect 44088 12776 44140 12782
rect 44140 12724 44220 12730
rect 44088 12718 44220 12724
rect 44100 12702 44220 12718
rect 41512 12640 41564 12646
rect 41512 12582 41564 12588
rect 44088 12640 44140 12646
rect 44088 12582 44140 12588
rect 44100 12442 44128 12582
rect 44088 12436 44140 12442
rect 44088 12378 44140 12384
rect 41512 12300 41564 12306
rect 41512 12242 41564 12248
rect 41524 11558 41552 12242
rect 42708 11688 42760 11694
rect 42706 11656 42708 11665
rect 42760 11656 42762 11665
rect 42706 11591 42762 11600
rect 44192 11558 44220 12702
rect 44560 12306 44588 12786
rect 44744 12646 44772 13466
rect 44928 12850 44956 13670
rect 45480 12986 45508 13806
rect 46388 13728 46440 13734
rect 46388 13670 46440 13676
rect 46112 13320 46164 13326
rect 46112 13262 46164 13268
rect 45468 12980 45520 12986
rect 45468 12922 45520 12928
rect 44916 12844 44968 12850
rect 44916 12786 44968 12792
rect 46124 12782 46152 13262
rect 46400 12782 46428 13670
rect 46768 13394 46796 13874
rect 46952 13530 46980 14742
rect 47214 14719 47270 14728
rect 47228 14482 47256 14719
rect 47216 14476 47268 14482
rect 47216 14418 47268 14424
rect 47228 14074 47256 14418
rect 47216 14068 47268 14074
rect 47216 14010 47268 14016
rect 47032 13796 47084 13802
rect 47032 13738 47084 13744
rect 46940 13524 46992 13530
rect 46940 13466 46992 13472
rect 46756 13388 46808 13394
rect 46756 13330 46808 13336
rect 46768 12986 46796 13330
rect 46756 12980 46808 12986
rect 46756 12922 46808 12928
rect 46112 12776 46164 12782
rect 46112 12718 46164 12724
rect 46388 12776 46440 12782
rect 46388 12718 46440 12724
rect 44732 12640 44784 12646
rect 45560 12640 45612 12646
rect 44732 12582 44784 12588
rect 45480 12600 45560 12628
rect 45480 12374 45508 12600
rect 45560 12582 45612 12588
rect 45008 12368 45060 12374
rect 45008 12310 45060 12316
rect 45468 12368 45520 12374
rect 45468 12310 45520 12316
rect 44548 12300 44600 12306
rect 44548 12242 44600 12248
rect 45020 12238 45048 12310
rect 45284 12300 45336 12306
rect 45284 12242 45336 12248
rect 45008 12232 45060 12238
rect 45008 12174 45060 12180
rect 45020 11558 45048 12174
rect 45296 11898 45324 12242
rect 46400 12170 46428 12718
rect 47044 12442 47072 13738
rect 47490 13288 47546 13297
rect 47490 13223 47546 13232
rect 47032 12436 47084 12442
rect 47032 12378 47084 12384
rect 47504 12306 47532 13223
rect 47492 12300 47544 12306
rect 47492 12242 47544 12248
rect 46388 12164 46440 12170
rect 46388 12106 46440 12112
rect 47504 11898 47532 12242
rect 45284 11892 45336 11898
rect 45284 11834 45336 11840
rect 47492 11892 47544 11898
rect 47492 11834 47544 11840
rect 41512 11552 41564 11558
rect 41512 11494 41564 11500
rect 44180 11552 44232 11558
rect 44180 11494 44232 11500
rect 45008 11552 45060 11558
rect 45008 11494 45060 11500
rect 41524 10810 41552 11494
rect 43628 11280 43680 11286
rect 43628 11222 43680 11228
rect 43076 11212 43128 11218
rect 43076 11154 43128 11160
rect 43088 10810 43116 11154
rect 43168 11076 43220 11082
rect 43168 11018 43220 11024
rect 41512 10804 41564 10810
rect 41512 10746 41564 10752
rect 43076 10804 43128 10810
rect 43076 10746 43128 10752
rect 41788 10532 41840 10538
rect 41788 10474 41840 10480
rect 42064 10532 42116 10538
rect 42064 10474 42116 10480
rect 41800 10266 41828 10474
rect 41972 10464 42024 10470
rect 41972 10406 42024 10412
rect 41788 10260 41840 10266
rect 41788 10202 41840 10208
rect 41984 9926 42012 10406
rect 42076 10198 42104 10474
rect 43088 10305 43116 10746
rect 43074 10296 43130 10305
rect 43074 10231 43076 10240
rect 43128 10231 43130 10240
rect 43076 10202 43128 10208
rect 42064 10192 42116 10198
rect 42062 10160 42064 10169
rect 42116 10160 42118 10169
rect 42062 10095 42118 10104
rect 42432 10124 42484 10130
rect 42076 10069 42104 10095
rect 42432 10066 42484 10072
rect 41972 9920 42024 9926
rect 41972 9862 42024 9868
rect 40776 9716 40828 9722
rect 40776 9658 40828 9664
rect 41420 9716 41472 9722
rect 41420 9658 41472 9664
rect 41696 9716 41748 9722
rect 41696 9658 41748 9664
rect 41708 9586 41736 9658
rect 41696 9580 41748 9586
rect 41696 9522 41748 9528
rect 40776 9512 40828 9518
rect 40776 9454 40828 9460
rect 38108 9376 38160 9382
rect 38108 9318 38160 9324
rect 38568 9376 38620 9382
rect 38568 9318 38620 9324
rect 38660 9376 38712 9382
rect 38660 9318 38712 9324
rect 39304 9376 39356 9382
rect 39304 9318 39356 9324
rect 36728 8968 36780 8974
rect 36728 8910 36780 8916
rect 36556 8248 36676 8276
rect 36452 8084 36504 8090
rect 36452 8026 36504 8032
rect 36268 6316 36320 6322
rect 36268 6258 36320 6264
rect 36280 5914 36308 6258
rect 36268 5908 36320 5914
rect 36268 5850 36320 5856
rect 36280 5098 36308 5850
rect 36556 5710 36584 8248
rect 36740 8022 36768 8910
rect 38120 8906 38148 9318
rect 38580 9042 38608 9318
rect 38568 9036 38620 9042
rect 38568 8978 38620 8984
rect 38672 8906 38700 9318
rect 40040 9172 40092 9178
rect 40040 9114 40092 9120
rect 38936 9104 38988 9110
rect 38936 9046 38988 9052
rect 39120 9104 39172 9110
rect 39120 9046 39172 9052
rect 38108 8900 38160 8906
rect 38108 8842 38160 8848
rect 38660 8900 38712 8906
rect 38660 8842 38712 8848
rect 38948 8634 38976 9046
rect 38936 8628 38988 8634
rect 38936 8570 38988 8576
rect 39132 8362 39160 9046
rect 39212 8968 39264 8974
rect 39212 8910 39264 8916
rect 39224 8537 39252 8910
rect 39210 8528 39266 8537
rect 39210 8463 39266 8472
rect 39120 8356 39172 8362
rect 39120 8298 39172 8304
rect 37832 8288 37884 8294
rect 37832 8230 37884 8236
rect 37924 8288 37976 8294
rect 37924 8230 37976 8236
rect 37844 8022 37872 8230
rect 36728 8016 36780 8022
rect 36728 7958 36780 7964
rect 37832 8016 37884 8022
rect 37832 7958 37884 7964
rect 36740 7478 36768 7958
rect 37740 7880 37792 7886
rect 37740 7822 37792 7828
rect 36728 7472 36780 7478
rect 36728 7414 36780 7420
rect 37752 7206 37780 7822
rect 37844 7546 37872 7958
rect 37936 7546 37964 8230
rect 39948 7948 40000 7954
rect 39948 7890 40000 7896
rect 39960 7750 39988 7890
rect 38384 7744 38436 7750
rect 38384 7686 38436 7692
rect 39948 7744 40000 7750
rect 39948 7686 40000 7692
rect 37832 7540 37884 7546
rect 37832 7482 37884 7488
rect 37924 7540 37976 7546
rect 37924 7482 37976 7488
rect 37844 7206 37872 7482
rect 38396 7410 38424 7686
rect 39960 7546 39988 7686
rect 39948 7540 40000 7546
rect 39948 7482 40000 7488
rect 40052 7426 40080 9114
rect 40788 9110 40816 9454
rect 41984 9178 42012 9862
rect 42064 9580 42116 9586
rect 42064 9522 42116 9528
rect 41972 9172 42024 9178
rect 41972 9114 42024 9120
rect 40684 9104 40736 9110
rect 40684 9046 40736 9052
rect 40776 9104 40828 9110
rect 40776 9046 40828 9052
rect 40500 9036 40552 9042
rect 40500 8978 40552 8984
rect 40512 8634 40540 8978
rect 40500 8628 40552 8634
rect 40500 8570 40552 8576
rect 40316 8424 40368 8430
rect 40316 8366 40368 8372
rect 40328 8294 40356 8366
rect 40316 8288 40368 8294
rect 40316 8230 40368 8236
rect 40224 7880 40276 7886
rect 40328 7834 40356 8230
rect 40512 8090 40540 8570
rect 40696 8294 40724 9046
rect 41604 8356 41656 8362
rect 41604 8298 41656 8304
rect 40684 8288 40736 8294
rect 40684 8230 40736 8236
rect 41616 8090 41644 8298
rect 40500 8084 40552 8090
rect 40500 8026 40552 8032
rect 41604 8084 41656 8090
rect 41604 8026 41656 8032
rect 40276 7828 40356 7834
rect 40224 7822 40356 7828
rect 40236 7806 40356 7822
rect 39960 7410 40080 7426
rect 38384 7404 38436 7410
rect 38384 7346 38436 7352
rect 39948 7404 40080 7410
rect 40000 7398 40080 7404
rect 39948 7346 40000 7352
rect 37280 7200 37332 7206
rect 37280 7142 37332 7148
rect 37740 7200 37792 7206
rect 37740 7142 37792 7148
rect 37832 7200 37884 7206
rect 37832 7142 37884 7148
rect 36544 5704 36596 5710
rect 36544 5646 36596 5652
rect 37096 5704 37148 5710
rect 37096 5646 37148 5652
rect 36268 5092 36320 5098
rect 36268 5034 36320 5040
rect 36280 4826 36308 5034
rect 37108 4826 37136 5646
rect 37188 5364 37240 5370
rect 37292 5352 37320 7142
rect 38396 7002 38424 7346
rect 40328 7342 40356 7806
rect 40316 7336 40368 7342
rect 40316 7278 40368 7284
rect 40512 7274 40540 8026
rect 40684 7336 40736 7342
rect 40684 7278 40736 7284
rect 40500 7268 40552 7274
rect 40500 7210 40552 7216
rect 38384 6996 38436 7002
rect 38384 6938 38436 6944
rect 37832 6792 37884 6798
rect 37832 6734 37884 6740
rect 37740 6384 37792 6390
rect 37740 6326 37792 6332
rect 37752 5846 37780 6326
rect 37844 6254 37872 6734
rect 37832 6248 37884 6254
rect 39304 6248 39356 6254
rect 37832 6190 37884 6196
rect 39302 6216 39304 6225
rect 39356 6216 39358 6225
rect 38292 6180 38344 6186
rect 39302 6151 39358 6160
rect 38292 6122 38344 6128
rect 38304 6089 38332 6122
rect 38660 6112 38712 6118
rect 38290 6080 38346 6089
rect 38660 6054 38712 6060
rect 39856 6112 39908 6118
rect 39856 6054 39908 6060
rect 38290 6015 38346 6024
rect 38200 5908 38252 5914
rect 38200 5850 38252 5856
rect 37740 5840 37792 5846
rect 37740 5782 37792 5788
rect 38106 5672 38162 5681
rect 38106 5607 38162 5616
rect 37240 5324 37320 5352
rect 37188 5306 37240 5312
rect 37372 5092 37424 5098
rect 37372 5034 37424 5040
rect 36268 4820 36320 4826
rect 36268 4762 36320 4768
rect 37096 4820 37148 4826
rect 37096 4762 37148 4768
rect 37108 4321 37136 4762
rect 37384 4593 37412 5034
rect 37464 5024 37516 5030
rect 37464 4966 37516 4972
rect 37476 4690 37504 4966
rect 38120 4758 38148 5607
rect 38212 5030 38240 5850
rect 38476 5704 38528 5710
rect 38476 5646 38528 5652
rect 38488 5098 38516 5646
rect 38672 5370 38700 6054
rect 38660 5364 38712 5370
rect 38660 5306 38712 5312
rect 38476 5092 38528 5098
rect 38476 5034 38528 5040
rect 38200 5024 38252 5030
rect 38200 4966 38252 4972
rect 39120 5024 39172 5030
rect 39120 4966 39172 4972
rect 38108 4752 38160 4758
rect 38108 4694 38160 4700
rect 37464 4684 37516 4690
rect 37464 4626 37516 4632
rect 37370 4584 37426 4593
rect 37370 4519 37372 4528
rect 37424 4519 37426 4528
rect 37372 4490 37424 4496
rect 37094 4312 37150 4321
rect 37476 4282 37504 4626
rect 37832 4480 37884 4486
rect 37832 4422 37884 4428
rect 37094 4247 37150 4256
rect 37464 4276 37516 4282
rect 37464 4218 37516 4224
rect 37372 3936 37424 3942
rect 37372 3878 37424 3884
rect 37384 3602 37412 3878
rect 37476 3670 37504 4218
rect 37844 3738 37872 4422
rect 38120 4282 38148 4694
rect 38108 4276 38160 4282
rect 38108 4218 38160 4224
rect 38212 3913 38240 4966
rect 39132 4826 39160 4966
rect 39120 4820 39172 4826
rect 39120 4762 39172 4768
rect 38292 4752 38344 4758
rect 38290 4720 38292 4729
rect 38344 4720 38346 4729
rect 38290 4655 38346 4664
rect 38304 4146 38332 4655
rect 39868 4146 39896 6054
rect 40696 5778 40724 7278
rect 41144 7268 41196 7274
rect 41144 7210 41196 7216
rect 41156 7002 41184 7210
rect 41144 6996 41196 7002
rect 41144 6938 41196 6944
rect 42076 6089 42104 9522
rect 42444 9178 42472 10066
rect 42800 9648 42852 9654
rect 42800 9590 42852 9596
rect 42616 9444 42668 9450
rect 42616 9386 42668 9392
rect 42524 9376 42576 9382
rect 42524 9318 42576 9324
rect 42432 9172 42484 9178
rect 42432 9114 42484 9120
rect 42432 9036 42484 9042
rect 42432 8978 42484 8984
rect 42444 8634 42472 8978
rect 42432 8628 42484 8634
rect 42432 8570 42484 8576
rect 42536 8090 42564 9318
rect 42524 8084 42576 8090
rect 42524 8026 42576 8032
rect 42536 7546 42564 8026
rect 42524 7540 42576 7546
rect 42524 7482 42576 7488
rect 42628 6866 42656 9386
rect 42812 8566 42840 9590
rect 43180 9518 43208 11018
rect 43444 11008 43496 11014
rect 43444 10950 43496 10956
rect 43456 10198 43484 10950
rect 43640 10538 43668 11222
rect 43628 10532 43680 10538
rect 43628 10474 43680 10480
rect 43640 10441 43668 10474
rect 44088 10464 44140 10470
rect 43626 10432 43682 10441
rect 44192 10418 44220 11494
rect 44140 10412 44220 10418
rect 44088 10406 44220 10412
rect 44100 10390 44220 10406
rect 43626 10367 43682 10376
rect 43444 10192 43496 10198
rect 43444 10134 43496 10140
rect 43904 10192 43956 10198
rect 43904 10134 43956 10140
rect 43456 9722 43484 10134
rect 43628 10056 43680 10062
rect 43628 9998 43680 10004
rect 43444 9716 43496 9722
rect 43444 9658 43496 9664
rect 43168 9512 43220 9518
rect 43168 9454 43220 9460
rect 43640 8838 43668 9998
rect 43916 9654 43944 10134
rect 43904 9648 43956 9654
rect 43904 9590 43956 9596
rect 44192 8974 44220 10390
rect 46938 10432 46994 10441
rect 46938 10367 46994 10376
rect 46952 10266 46980 10367
rect 46940 10260 46992 10266
rect 46940 10202 46992 10208
rect 46938 10160 46994 10169
rect 45836 10124 45888 10130
rect 46938 10095 46994 10104
rect 47398 10160 47454 10169
rect 47398 10095 47454 10104
rect 45836 10066 45888 10072
rect 45560 10056 45612 10062
rect 45560 9998 45612 10004
rect 44272 9920 44324 9926
rect 44272 9862 44324 9868
rect 45100 9920 45152 9926
rect 45100 9862 45152 9868
rect 44284 9518 44312 9862
rect 44272 9512 44324 9518
rect 44272 9454 44324 9460
rect 45112 9450 45140 9862
rect 44824 9444 44876 9450
rect 44824 9386 44876 9392
rect 45100 9444 45152 9450
rect 45100 9386 45152 9392
rect 44836 9178 44864 9386
rect 45008 9376 45060 9382
rect 45008 9318 45060 9324
rect 44824 9172 44876 9178
rect 44824 9114 44876 9120
rect 45020 9110 45048 9318
rect 45008 9104 45060 9110
rect 45008 9046 45060 9052
rect 44180 8968 44232 8974
rect 44180 8910 44232 8916
rect 44824 8968 44876 8974
rect 44824 8910 44876 8916
rect 43628 8832 43680 8838
rect 43628 8774 43680 8780
rect 42800 8560 42852 8566
rect 43640 8537 43668 8774
rect 42800 8502 42852 8508
rect 43626 8528 43682 8537
rect 43626 8463 43628 8472
rect 43680 8463 43682 8472
rect 43628 8434 43680 8440
rect 43076 8356 43128 8362
rect 43076 8298 43128 8304
rect 43088 7750 43116 8298
rect 44836 8294 44864 8910
rect 44824 8288 44876 8294
rect 44824 8230 44876 8236
rect 43628 8084 43680 8090
rect 43628 8026 43680 8032
rect 43076 7744 43128 7750
rect 43076 7686 43128 7692
rect 42616 6860 42668 6866
rect 42616 6802 42668 6808
rect 42628 6458 42656 6802
rect 43088 6458 43116 7686
rect 43640 7342 43668 8026
rect 44836 7886 44864 8230
rect 44824 7880 44876 7886
rect 44824 7822 44876 7828
rect 43628 7336 43680 7342
rect 43628 7278 43680 7284
rect 44836 7274 44864 7822
rect 43444 7268 43496 7274
rect 43444 7210 43496 7216
rect 44824 7268 44876 7274
rect 44824 7210 44876 7216
rect 43352 6792 43404 6798
rect 43456 6746 43484 7210
rect 44180 7200 44232 7206
rect 44180 7142 44232 7148
rect 44192 6866 44220 7142
rect 45112 7041 45140 9386
rect 45572 9382 45600 9998
rect 45848 9518 45876 10066
rect 46952 9654 46980 10095
rect 47412 9654 47440 10095
rect 46940 9648 46992 9654
rect 46940 9590 46992 9596
rect 47400 9648 47452 9654
rect 47400 9590 47452 9596
rect 45836 9512 45888 9518
rect 45836 9454 45888 9460
rect 46480 9512 46532 9518
rect 46480 9454 46532 9460
rect 45192 9376 45244 9382
rect 45192 9318 45244 9324
rect 45560 9376 45612 9382
rect 45560 9318 45612 9324
rect 45204 9042 45232 9318
rect 46492 9178 46520 9454
rect 46480 9172 46532 9178
rect 46480 9114 46532 9120
rect 45560 9104 45612 9110
rect 45560 9046 45612 9052
rect 45192 9036 45244 9042
rect 45192 8978 45244 8984
rect 45572 8294 45600 9046
rect 46940 8560 46992 8566
rect 46938 8528 46940 8537
rect 46992 8528 46994 8537
rect 46938 8463 46994 8472
rect 47398 8528 47454 8537
rect 47398 8463 47400 8472
rect 47452 8463 47454 8472
rect 47400 8434 47452 8440
rect 45560 8288 45612 8294
rect 45560 8230 45612 8236
rect 45572 8090 45600 8230
rect 45560 8084 45612 8090
rect 45560 8026 45612 8032
rect 45376 7948 45428 7954
rect 45376 7890 45428 7896
rect 44362 7032 44418 7041
rect 44362 6967 44418 6976
rect 45098 7032 45154 7041
rect 45098 6967 45154 6976
rect 44180 6860 44232 6866
rect 44180 6802 44232 6808
rect 43404 6740 43484 6746
rect 43352 6734 43484 6740
rect 43364 6718 43484 6734
rect 42616 6452 42668 6458
rect 42616 6394 42668 6400
rect 43076 6452 43128 6458
rect 43076 6394 43128 6400
rect 43456 6390 43484 6718
rect 43444 6384 43496 6390
rect 43444 6326 43496 6332
rect 44376 6254 44404 6967
rect 44732 6860 44784 6866
rect 44732 6802 44784 6808
rect 44744 6662 44772 6802
rect 45388 6662 45416 7890
rect 45836 7200 45888 7206
rect 45836 7142 45888 7148
rect 46940 7200 46992 7206
rect 46940 7142 46992 7148
rect 47400 7200 47452 7206
rect 47400 7142 47452 7148
rect 45848 6798 45876 7142
rect 46952 7041 46980 7142
rect 47412 7041 47440 7142
rect 46938 7032 46994 7041
rect 46938 6967 46994 6976
rect 47398 7032 47454 7041
rect 47398 6967 47454 6976
rect 46112 6860 46164 6866
rect 46112 6802 46164 6808
rect 45836 6792 45888 6798
rect 45888 6740 45968 6746
rect 45836 6734 45968 6740
rect 45848 6718 45968 6734
rect 44732 6656 44784 6662
rect 44732 6598 44784 6604
rect 45376 6656 45428 6662
rect 45376 6598 45428 6604
rect 44364 6248 44416 6254
rect 44364 6190 44416 6196
rect 43812 6112 43864 6118
rect 42062 6080 42118 6089
rect 43812 6054 43864 6060
rect 42062 6015 42118 6024
rect 42076 5914 42104 6015
rect 43824 5914 43852 6054
rect 44376 5914 44404 6190
rect 44744 6118 44772 6598
rect 45388 6322 45416 6598
rect 45376 6316 45428 6322
rect 45376 6258 45428 6264
rect 45940 6118 45968 6718
rect 46124 6458 46152 6802
rect 46112 6452 46164 6458
rect 46112 6394 46164 6400
rect 44732 6112 44784 6118
rect 45928 6112 45980 6118
rect 44732 6054 44784 6060
rect 45926 6080 45928 6089
rect 45980 6080 45982 6089
rect 45926 6015 45982 6024
rect 49238 6080 49294 6089
rect 49238 6015 49294 6024
rect 42064 5908 42116 5914
rect 42064 5850 42116 5856
rect 43812 5908 43864 5914
rect 43812 5850 43864 5856
rect 44364 5908 44416 5914
rect 44364 5850 44416 5856
rect 40684 5772 40736 5778
rect 40604 5732 40684 5760
rect 39948 5568 40000 5574
rect 40000 5516 40080 5522
rect 39948 5510 40080 5516
rect 39960 5494 40080 5510
rect 40052 4729 40080 5494
rect 40604 5166 40632 5732
rect 40684 5714 40736 5720
rect 40960 5772 41012 5778
rect 40960 5714 41012 5720
rect 40684 5568 40736 5574
rect 40684 5510 40736 5516
rect 40592 5160 40644 5166
rect 40592 5102 40644 5108
rect 40604 4826 40632 5102
rect 40696 5098 40724 5510
rect 40684 5092 40736 5098
rect 40684 5034 40736 5040
rect 40592 4820 40644 4826
rect 40592 4762 40644 4768
rect 40038 4720 40094 4729
rect 40038 4655 40094 4664
rect 38292 4140 38344 4146
rect 38292 4082 38344 4088
rect 39856 4140 39908 4146
rect 39856 4082 39908 4088
rect 40052 4010 40080 4655
rect 40500 4480 40552 4486
rect 40500 4422 40552 4428
rect 40512 4321 40540 4422
rect 40498 4312 40554 4321
rect 40498 4247 40554 4256
rect 40408 4140 40460 4146
rect 40408 4082 40460 4088
rect 40040 4004 40092 4010
rect 40040 3946 40092 3952
rect 39396 3936 39448 3942
rect 38198 3904 38254 3913
rect 39396 3878 39448 3884
rect 38198 3839 38254 3848
rect 37832 3732 37884 3738
rect 37832 3674 37884 3680
rect 39408 3670 39436 3878
rect 37464 3664 37516 3670
rect 37464 3606 37516 3612
rect 39396 3664 39448 3670
rect 39396 3606 39448 3612
rect 40224 3664 40276 3670
rect 40224 3606 40276 3612
rect 37372 3596 37424 3602
rect 37372 3538 37424 3544
rect 37384 3194 37412 3538
rect 37372 3188 37424 3194
rect 37372 3130 37424 3136
rect 36268 3120 36320 3126
rect 36266 3088 36268 3097
rect 36320 3088 36322 3097
rect 36266 3023 36322 3032
rect 37476 2990 37504 3606
rect 38568 3528 38620 3534
rect 38568 3470 38620 3476
rect 37832 3392 37884 3398
rect 37832 3334 37884 3340
rect 37464 2984 37516 2990
rect 36634 2952 36690 2961
rect 37464 2926 37516 2932
rect 36634 2887 36690 2896
rect 37280 2916 37332 2922
rect 36648 2514 36676 2887
rect 37280 2858 37332 2864
rect 37292 2650 37320 2858
rect 37844 2825 37872 3334
rect 38580 2854 38608 3470
rect 39408 3194 39436 3606
rect 39764 3392 39816 3398
rect 39764 3334 39816 3340
rect 39396 3188 39448 3194
rect 39396 3130 39448 3136
rect 38568 2848 38620 2854
rect 37830 2816 37886 2825
rect 38568 2790 38620 2796
rect 37830 2751 37886 2760
rect 37280 2644 37332 2650
rect 37280 2586 37332 2592
rect 38580 2582 38608 2790
rect 38568 2576 38620 2582
rect 38568 2518 38620 2524
rect 36636 2508 36688 2514
rect 36636 2450 36688 2456
rect 37096 2508 37148 2514
rect 37096 2450 37148 2456
rect 36174 1456 36230 1465
rect 36174 1391 36230 1400
rect 37108 480 37136 2450
rect 38200 2372 38252 2378
rect 38200 2314 38252 2320
rect 38212 1170 38240 2314
rect 38212 1142 38424 1170
rect 38396 480 38424 1142
rect 39776 480 39804 3334
rect 40040 2916 40092 2922
rect 40040 2858 40092 2864
rect 40052 2650 40080 2858
rect 40040 2644 40092 2650
rect 40040 2586 40092 2592
rect 40236 2378 40264 3606
rect 40420 2650 40448 4082
rect 40512 4078 40540 4247
rect 40500 4072 40552 4078
rect 40500 4014 40552 4020
rect 40604 3210 40632 4762
rect 40696 3534 40724 5034
rect 40972 5030 41000 5714
rect 40960 5024 41012 5030
rect 40960 4966 41012 4972
rect 40972 4826 41000 4966
rect 40960 4820 41012 4826
rect 40960 4762 41012 4768
rect 40776 4072 40828 4078
rect 40776 4014 40828 4020
rect 40788 3738 40816 4014
rect 41052 3936 41104 3942
rect 41050 3904 41052 3913
rect 42340 3936 42392 3942
rect 41104 3904 41106 3913
rect 41050 3839 41106 3848
rect 41418 3904 41474 3913
rect 42340 3878 42392 3884
rect 41418 3839 41474 3848
rect 40776 3732 40828 3738
rect 40776 3674 40828 3680
rect 41432 3641 41460 3839
rect 41418 3632 41474 3641
rect 41418 3567 41474 3576
rect 40684 3528 40736 3534
rect 40684 3470 40736 3476
rect 40512 3194 40632 3210
rect 40696 3194 40724 3470
rect 41052 3392 41104 3398
rect 41052 3334 41104 3340
rect 41144 3392 41196 3398
rect 41144 3334 41196 3340
rect 40500 3188 40632 3194
rect 40552 3182 40632 3188
rect 40684 3188 40736 3194
rect 40500 3130 40552 3136
rect 40684 3130 40736 3136
rect 41064 2922 41092 3334
rect 41052 2916 41104 2922
rect 41052 2858 41104 2864
rect 40408 2644 40460 2650
rect 40408 2586 40460 2592
rect 40224 2372 40276 2378
rect 40224 2314 40276 2320
rect 41156 480 41184 3334
rect 41328 2916 41380 2922
rect 41328 2858 41380 2864
rect 41340 2530 41368 2858
rect 42352 2582 42380 3878
rect 47858 3632 47914 3641
rect 47858 3567 47914 3576
rect 42706 2816 42762 2825
rect 42706 2751 42762 2760
rect 42340 2576 42392 2582
rect 41340 2514 41460 2530
rect 42340 2518 42392 2524
rect 42720 2514 42748 2751
rect 41340 2508 41472 2514
rect 41340 2502 41420 2508
rect 41420 2450 41472 2456
rect 42432 2508 42484 2514
rect 42432 2450 42484 2456
rect 42708 2508 42760 2514
rect 42708 2450 42760 2456
rect 45192 2508 45244 2514
rect 45192 2450 45244 2456
rect 42444 480 42472 2450
rect 43812 2372 43864 2378
rect 43812 2314 43864 2320
rect 43824 480 43852 2314
rect 45204 2310 45232 2450
rect 46480 2372 46532 2378
rect 46480 2314 46532 2320
rect 45192 2304 45244 2310
rect 45192 2246 45244 2252
rect 45204 480 45232 2246
rect 46492 480 46520 2314
rect 47872 480 47900 3567
rect 49252 480 49280 6015
rect 36082 96 36138 105
rect 36082 31 36138 40
rect 37094 0 37150 480
rect 38382 0 38438 480
rect 39762 0 39818 480
rect 41142 0 41198 480
rect 42430 0 42486 480
rect 43810 0 43866 480
rect 45190 0 45246 480
rect 46478 0 46534 480
rect 47858 0 47914 480
rect 49238 0 49294 480
<< via2 >>
rect 4220 46810 4276 46812
rect 4300 46810 4356 46812
rect 4380 46810 4436 46812
rect 4460 46810 4516 46812
rect 4220 46758 4246 46810
rect 4246 46758 4276 46810
rect 4300 46758 4310 46810
rect 4310 46758 4356 46810
rect 4380 46758 4426 46810
rect 4426 46758 4436 46810
rect 4460 46758 4490 46810
rect 4490 46758 4516 46810
rect 4220 46756 4276 46758
rect 4300 46756 4356 46758
rect 4380 46756 4436 46758
rect 4460 46756 4516 46758
rect 4220 45722 4276 45724
rect 4300 45722 4356 45724
rect 4380 45722 4436 45724
rect 4460 45722 4516 45724
rect 4220 45670 4246 45722
rect 4246 45670 4276 45722
rect 4300 45670 4310 45722
rect 4310 45670 4356 45722
rect 4380 45670 4426 45722
rect 4426 45670 4436 45722
rect 4460 45670 4490 45722
rect 4490 45670 4516 45722
rect 4220 45668 4276 45670
rect 4300 45668 4356 45670
rect 4380 45668 4436 45670
rect 4460 45668 4516 45670
rect 4220 44634 4276 44636
rect 4300 44634 4356 44636
rect 4380 44634 4436 44636
rect 4460 44634 4516 44636
rect 4220 44582 4246 44634
rect 4246 44582 4276 44634
rect 4300 44582 4310 44634
rect 4310 44582 4356 44634
rect 4380 44582 4426 44634
rect 4426 44582 4436 44634
rect 4460 44582 4490 44634
rect 4490 44582 4516 44634
rect 4220 44580 4276 44582
rect 4300 44580 4356 44582
rect 4380 44580 4436 44582
rect 4460 44580 4516 44582
rect 4220 43546 4276 43548
rect 4300 43546 4356 43548
rect 4380 43546 4436 43548
rect 4460 43546 4516 43548
rect 4220 43494 4246 43546
rect 4246 43494 4276 43546
rect 4300 43494 4310 43546
rect 4310 43494 4356 43546
rect 4380 43494 4426 43546
rect 4426 43494 4436 43546
rect 4460 43494 4490 43546
rect 4490 43494 4516 43546
rect 4220 43492 4276 43494
rect 4300 43492 4356 43494
rect 4380 43492 4436 43494
rect 4460 43492 4516 43494
rect 4220 42458 4276 42460
rect 4300 42458 4356 42460
rect 4380 42458 4436 42460
rect 4460 42458 4516 42460
rect 4220 42406 4246 42458
rect 4246 42406 4276 42458
rect 4300 42406 4310 42458
rect 4310 42406 4356 42458
rect 4380 42406 4426 42458
rect 4426 42406 4436 42458
rect 4460 42406 4490 42458
rect 4490 42406 4516 42458
rect 4220 42404 4276 42406
rect 4300 42404 4356 42406
rect 4380 42404 4436 42406
rect 4460 42404 4516 42406
rect 4220 41370 4276 41372
rect 4300 41370 4356 41372
rect 4380 41370 4436 41372
rect 4460 41370 4516 41372
rect 4220 41318 4246 41370
rect 4246 41318 4276 41370
rect 4300 41318 4310 41370
rect 4310 41318 4356 41370
rect 4380 41318 4426 41370
rect 4426 41318 4436 41370
rect 4460 41318 4490 41370
rect 4490 41318 4516 41370
rect 4220 41316 4276 41318
rect 4300 41316 4356 41318
rect 4380 41316 4436 41318
rect 4460 41316 4516 41318
rect 4220 40282 4276 40284
rect 4300 40282 4356 40284
rect 4380 40282 4436 40284
rect 4460 40282 4516 40284
rect 4220 40230 4246 40282
rect 4246 40230 4276 40282
rect 4300 40230 4310 40282
rect 4310 40230 4356 40282
rect 4380 40230 4426 40282
rect 4426 40230 4436 40282
rect 4460 40230 4490 40282
rect 4490 40230 4516 40282
rect 4220 40228 4276 40230
rect 4300 40228 4356 40230
rect 4380 40228 4436 40230
rect 4460 40228 4516 40230
rect 4220 39194 4276 39196
rect 4300 39194 4356 39196
rect 4380 39194 4436 39196
rect 4460 39194 4516 39196
rect 4220 39142 4246 39194
rect 4246 39142 4276 39194
rect 4300 39142 4310 39194
rect 4310 39142 4356 39194
rect 4380 39142 4426 39194
rect 4426 39142 4436 39194
rect 4460 39142 4490 39194
rect 4490 39142 4516 39194
rect 4220 39140 4276 39142
rect 4300 39140 4356 39142
rect 4380 39140 4436 39142
rect 4460 39140 4516 39142
rect 4220 38106 4276 38108
rect 4300 38106 4356 38108
rect 4380 38106 4436 38108
rect 4460 38106 4516 38108
rect 4220 38054 4246 38106
rect 4246 38054 4276 38106
rect 4300 38054 4310 38106
rect 4310 38054 4356 38106
rect 4380 38054 4426 38106
rect 4426 38054 4436 38106
rect 4460 38054 4490 38106
rect 4490 38054 4516 38106
rect 4220 38052 4276 38054
rect 4300 38052 4356 38054
rect 4380 38052 4436 38054
rect 4460 38052 4516 38054
rect 3422 37576 3478 37632
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4246 37018
rect 4246 36966 4276 37018
rect 4300 36966 4310 37018
rect 4310 36966 4356 37018
rect 4380 36966 4426 37018
rect 4426 36966 4436 37018
rect 4460 36966 4490 37018
rect 4490 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4246 35930
rect 4246 35878 4276 35930
rect 4300 35878 4310 35930
rect 4310 35878 4356 35930
rect 4380 35878 4426 35930
rect 4426 35878 4436 35930
rect 4460 35878 4490 35930
rect 4490 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4246 34842
rect 4246 34790 4276 34842
rect 4300 34790 4310 34842
rect 4310 34790 4356 34842
rect 4380 34790 4426 34842
rect 4426 34790 4436 34842
rect 4460 34790 4490 34842
rect 4490 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4246 33754
rect 4246 33702 4276 33754
rect 4300 33702 4310 33754
rect 4310 33702 4356 33754
rect 4380 33702 4426 33754
rect 4426 33702 4436 33754
rect 4460 33702 4490 33754
rect 4490 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4246 32666
rect 4246 32614 4276 32666
rect 4300 32614 4310 32666
rect 4310 32614 4356 32666
rect 4380 32614 4426 32666
rect 4426 32614 4436 32666
rect 4460 32614 4490 32666
rect 4490 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4246 31578
rect 4246 31526 4276 31578
rect 4300 31526 4310 31578
rect 4310 31526 4356 31578
rect 4380 31526 4426 31578
rect 4426 31526 4436 31578
rect 4460 31526 4490 31578
rect 4490 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4246 30490
rect 4246 30438 4276 30490
rect 4300 30438 4310 30490
rect 4310 30438 4356 30490
rect 4380 30438 4426 30490
rect 4426 30438 4436 30490
rect 4460 30438 4490 30490
rect 4490 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4246 29402
rect 4246 29350 4276 29402
rect 4300 29350 4310 29402
rect 4310 29350 4356 29402
rect 4380 29350 4426 29402
rect 4426 29350 4436 29402
rect 4460 29350 4490 29402
rect 4490 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4246 28314
rect 4246 28262 4276 28314
rect 4300 28262 4310 28314
rect 4310 28262 4356 28314
rect 4380 28262 4426 28314
rect 4426 28262 4436 28314
rect 4460 28262 4490 28314
rect 4490 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4246 27226
rect 4246 27174 4276 27226
rect 4300 27174 4310 27226
rect 4310 27174 4356 27226
rect 4380 27174 4426 27226
rect 4426 27174 4436 27226
rect 4460 27174 4490 27226
rect 4490 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4246 26138
rect 4246 26086 4276 26138
rect 4300 26086 4310 26138
rect 4310 26086 4356 26138
rect 4380 26086 4426 26138
rect 4426 26086 4436 26138
rect 4460 26086 4490 26138
rect 4490 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 19580 47354 19636 47356
rect 19660 47354 19716 47356
rect 19740 47354 19796 47356
rect 19820 47354 19876 47356
rect 19580 47302 19606 47354
rect 19606 47302 19636 47354
rect 19660 47302 19670 47354
rect 19670 47302 19716 47354
rect 19740 47302 19786 47354
rect 19786 47302 19796 47354
rect 19820 47302 19850 47354
rect 19850 47302 19876 47354
rect 19580 47300 19636 47302
rect 19660 47300 19716 47302
rect 19740 47300 19796 47302
rect 19820 47300 19876 47302
rect 19580 46266 19636 46268
rect 19660 46266 19716 46268
rect 19740 46266 19796 46268
rect 19820 46266 19876 46268
rect 19580 46214 19606 46266
rect 19606 46214 19636 46266
rect 19660 46214 19670 46266
rect 19670 46214 19716 46266
rect 19740 46214 19786 46266
rect 19786 46214 19796 46266
rect 19820 46214 19850 46266
rect 19850 46214 19876 46266
rect 19580 46212 19636 46214
rect 19660 46212 19716 46214
rect 19740 46212 19796 46214
rect 19820 46212 19876 46214
rect 34940 46810 34996 46812
rect 35020 46810 35076 46812
rect 35100 46810 35156 46812
rect 35180 46810 35236 46812
rect 34940 46758 34966 46810
rect 34966 46758 34996 46810
rect 35020 46758 35030 46810
rect 35030 46758 35076 46810
rect 35100 46758 35146 46810
rect 35146 46758 35156 46810
rect 35180 46758 35210 46810
rect 35210 46758 35236 46810
rect 34940 46756 34996 46758
rect 35020 46756 35076 46758
rect 35100 46756 35156 46758
rect 35180 46756 35236 46758
rect 34940 45722 34996 45724
rect 35020 45722 35076 45724
rect 35100 45722 35156 45724
rect 35180 45722 35236 45724
rect 34940 45670 34966 45722
rect 34966 45670 34996 45722
rect 35020 45670 35030 45722
rect 35030 45670 35076 45722
rect 35100 45670 35146 45722
rect 35146 45670 35156 45722
rect 35180 45670 35210 45722
rect 35210 45670 35236 45722
rect 34940 45668 34996 45670
rect 35020 45668 35076 45670
rect 35100 45668 35156 45670
rect 35180 45668 35236 45670
rect 24950 45600 25006 45656
rect 28078 45600 28134 45656
rect 19580 45178 19636 45180
rect 19660 45178 19716 45180
rect 19740 45178 19796 45180
rect 19820 45178 19876 45180
rect 19580 45126 19606 45178
rect 19606 45126 19636 45178
rect 19660 45126 19670 45178
rect 19670 45126 19716 45178
rect 19740 45126 19786 45178
rect 19786 45126 19796 45178
rect 19820 45126 19850 45178
rect 19850 45126 19876 45178
rect 19580 45124 19636 45126
rect 19660 45124 19716 45126
rect 19740 45124 19796 45126
rect 19820 45124 19876 45126
rect 19580 44090 19636 44092
rect 19660 44090 19716 44092
rect 19740 44090 19796 44092
rect 19820 44090 19876 44092
rect 19580 44038 19606 44090
rect 19606 44038 19636 44090
rect 19660 44038 19670 44090
rect 19670 44038 19716 44090
rect 19740 44038 19786 44090
rect 19786 44038 19796 44090
rect 19820 44038 19850 44090
rect 19850 44038 19876 44090
rect 19580 44036 19636 44038
rect 19660 44036 19716 44038
rect 19740 44036 19796 44038
rect 19820 44036 19876 44038
rect 19580 43002 19636 43004
rect 19660 43002 19716 43004
rect 19740 43002 19796 43004
rect 19820 43002 19876 43004
rect 19580 42950 19606 43002
rect 19606 42950 19636 43002
rect 19660 42950 19670 43002
rect 19670 42950 19716 43002
rect 19740 42950 19786 43002
rect 19786 42950 19796 43002
rect 19820 42950 19850 43002
rect 19850 42950 19876 43002
rect 19580 42948 19636 42950
rect 19660 42948 19716 42950
rect 19740 42948 19796 42950
rect 19820 42948 19876 42950
rect 19580 41914 19636 41916
rect 19660 41914 19716 41916
rect 19740 41914 19796 41916
rect 19820 41914 19876 41916
rect 19580 41862 19606 41914
rect 19606 41862 19636 41914
rect 19660 41862 19670 41914
rect 19670 41862 19716 41914
rect 19740 41862 19786 41914
rect 19786 41862 19796 41914
rect 19820 41862 19850 41914
rect 19850 41862 19876 41914
rect 19580 41860 19636 41862
rect 19660 41860 19716 41862
rect 19740 41860 19796 41862
rect 19820 41860 19876 41862
rect 19580 40826 19636 40828
rect 19660 40826 19716 40828
rect 19740 40826 19796 40828
rect 19820 40826 19876 40828
rect 19580 40774 19606 40826
rect 19606 40774 19636 40826
rect 19660 40774 19670 40826
rect 19670 40774 19716 40826
rect 19740 40774 19786 40826
rect 19786 40774 19796 40826
rect 19820 40774 19850 40826
rect 19850 40774 19876 40826
rect 19580 40772 19636 40774
rect 19660 40772 19716 40774
rect 19740 40772 19796 40774
rect 19820 40772 19876 40774
rect 19580 39738 19636 39740
rect 19660 39738 19716 39740
rect 19740 39738 19796 39740
rect 19820 39738 19876 39740
rect 19580 39686 19606 39738
rect 19606 39686 19636 39738
rect 19660 39686 19670 39738
rect 19670 39686 19716 39738
rect 19740 39686 19786 39738
rect 19786 39686 19796 39738
rect 19820 39686 19850 39738
rect 19850 39686 19876 39738
rect 19580 39684 19636 39686
rect 19660 39684 19716 39686
rect 19740 39684 19796 39686
rect 19820 39684 19876 39686
rect 19580 38650 19636 38652
rect 19660 38650 19716 38652
rect 19740 38650 19796 38652
rect 19820 38650 19876 38652
rect 19580 38598 19606 38650
rect 19606 38598 19636 38650
rect 19660 38598 19670 38650
rect 19670 38598 19716 38650
rect 19740 38598 19786 38650
rect 19786 38598 19796 38650
rect 19820 38598 19850 38650
rect 19850 38598 19876 38650
rect 19580 38596 19636 38598
rect 19660 38596 19716 38598
rect 19740 38596 19796 38598
rect 19820 38596 19876 38598
rect 19580 37562 19636 37564
rect 19660 37562 19716 37564
rect 19740 37562 19796 37564
rect 19820 37562 19876 37564
rect 19580 37510 19606 37562
rect 19606 37510 19636 37562
rect 19660 37510 19670 37562
rect 19670 37510 19716 37562
rect 19740 37510 19786 37562
rect 19786 37510 19796 37562
rect 19820 37510 19850 37562
rect 19850 37510 19876 37562
rect 19580 37508 19636 37510
rect 19660 37508 19716 37510
rect 19740 37508 19796 37510
rect 19820 37508 19876 37510
rect 19580 36474 19636 36476
rect 19660 36474 19716 36476
rect 19740 36474 19796 36476
rect 19820 36474 19876 36476
rect 19580 36422 19606 36474
rect 19606 36422 19636 36474
rect 19660 36422 19670 36474
rect 19670 36422 19716 36474
rect 19740 36422 19786 36474
rect 19786 36422 19796 36474
rect 19820 36422 19850 36474
rect 19850 36422 19876 36474
rect 19580 36420 19636 36422
rect 19660 36420 19716 36422
rect 19740 36420 19796 36422
rect 19820 36420 19876 36422
rect 19580 35386 19636 35388
rect 19660 35386 19716 35388
rect 19740 35386 19796 35388
rect 19820 35386 19876 35388
rect 19580 35334 19606 35386
rect 19606 35334 19636 35386
rect 19660 35334 19670 35386
rect 19670 35334 19716 35386
rect 19740 35334 19786 35386
rect 19786 35334 19796 35386
rect 19820 35334 19850 35386
rect 19850 35334 19876 35386
rect 19580 35332 19636 35334
rect 19660 35332 19716 35334
rect 19740 35332 19796 35334
rect 19820 35332 19876 35334
rect 19580 34298 19636 34300
rect 19660 34298 19716 34300
rect 19740 34298 19796 34300
rect 19820 34298 19876 34300
rect 19580 34246 19606 34298
rect 19606 34246 19636 34298
rect 19660 34246 19670 34298
rect 19670 34246 19716 34298
rect 19740 34246 19786 34298
rect 19786 34246 19796 34298
rect 19820 34246 19850 34298
rect 19850 34246 19876 34298
rect 19580 34244 19636 34246
rect 19660 34244 19716 34246
rect 19740 34244 19796 34246
rect 19820 34244 19876 34246
rect 19580 33210 19636 33212
rect 19660 33210 19716 33212
rect 19740 33210 19796 33212
rect 19820 33210 19876 33212
rect 19580 33158 19606 33210
rect 19606 33158 19636 33210
rect 19660 33158 19670 33210
rect 19670 33158 19716 33210
rect 19740 33158 19786 33210
rect 19786 33158 19796 33210
rect 19820 33158 19850 33210
rect 19850 33158 19876 33210
rect 19580 33156 19636 33158
rect 19660 33156 19716 33158
rect 19740 33156 19796 33158
rect 19820 33156 19876 33158
rect 19580 32122 19636 32124
rect 19660 32122 19716 32124
rect 19740 32122 19796 32124
rect 19820 32122 19876 32124
rect 19580 32070 19606 32122
rect 19606 32070 19636 32122
rect 19660 32070 19670 32122
rect 19670 32070 19716 32122
rect 19740 32070 19786 32122
rect 19786 32070 19796 32122
rect 19820 32070 19850 32122
rect 19850 32070 19876 32122
rect 19580 32068 19636 32070
rect 19660 32068 19716 32070
rect 19740 32068 19796 32070
rect 19820 32068 19876 32070
rect 19580 31034 19636 31036
rect 19660 31034 19716 31036
rect 19740 31034 19796 31036
rect 19820 31034 19876 31036
rect 19580 30982 19606 31034
rect 19606 30982 19636 31034
rect 19660 30982 19670 31034
rect 19670 30982 19716 31034
rect 19740 30982 19786 31034
rect 19786 30982 19796 31034
rect 19820 30982 19850 31034
rect 19850 30982 19876 31034
rect 19580 30980 19636 30982
rect 19660 30980 19716 30982
rect 19740 30980 19796 30982
rect 19820 30980 19876 30982
rect 19580 29946 19636 29948
rect 19660 29946 19716 29948
rect 19740 29946 19796 29948
rect 19820 29946 19876 29948
rect 19580 29894 19606 29946
rect 19606 29894 19636 29946
rect 19660 29894 19670 29946
rect 19670 29894 19716 29946
rect 19740 29894 19786 29946
rect 19786 29894 19796 29946
rect 19820 29894 19850 29946
rect 19850 29894 19876 29946
rect 19580 29892 19636 29894
rect 19660 29892 19716 29894
rect 19740 29892 19796 29894
rect 19820 29892 19876 29894
rect 19580 28858 19636 28860
rect 19660 28858 19716 28860
rect 19740 28858 19796 28860
rect 19820 28858 19876 28860
rect 19580 28806 19606 28858
rect 19606 28806 19636 28858
rect 19660 28806 19670 28858
rect 19670 28806 19716 28858
rect 19740 28806 19786 28858
rect 19786 28806 19796 28858
rect 19820 28806 19850 28858
rect 19850 28806 19876 28858
rect 19580 28804 19636 28806
rect 19660 28804 19716 28806
rect 19740 28804 19796 28806
rect 19820 28804 19876 28806
rect 19580 27770 19636 27772
rect 19660 27770 19716 27772
rect 19740 27770 19796 27772
rect 19820 27770 19876 27772
rect 19580 27718 19606 27770
rect 19606 27718 19636 27770
rect 19660 27718 19670 27770
rect 19670 27718 19716 27770
rect 19740 27718 19786 27770
rect 19786 27718 19796 27770
rect 19820 27718 19850 27770
rect 19850 27718 19876 27770
rect 19580 27716 19636 27718
rect 19660 27716 19716 27718
rect 19740 27716 19796 27718
rect 19820 27716 19876 27718
rect 19580 26682 19636 26684
rect 19660 26682 19716 26684
rect 19740 26682 19796 26684
rect 19820 26682 19876 26684
rect 19580 26630 19606 26682
rect 19606 26630 19636 26682
rect 19660 26630 19670 26682
rect 19670 26630 19716 26682
rect 19740 26630 19786 26682
rect 19786 26630 19796 26682
rect 19820 26630 19850 26682
rect 19850 26630 19876 26682
rect 19580 26628 19636 26630
rect 19660 26628 19716 26630
rect 19740 26628 19796 26630
rect 19820 26628 19876 26630
rect 19580 25594 19636 25596
rect 19660 25594 19716 25596
rect 19740 25594 19796 25596
rect 19820 25594 19876 25596
rect 19580 25542 19606 25594
rect 19606 25542 19636 25594
rect 19660 25542 19670 25594
rect 19670 25542 19716 25594
rect 19740 25542 19786 25594
rect 19786 25542 19796 25594
rect 19820 25542 19850 25594
rect 19850 25542 19876 25594
rect 19580 25540 19636 25542
rect 19660 25540 19716 25542
rect 19740 25540 19796 25542
rect 19820 25540 19876 25542
rect 19580 24506 19636 24508
rect 19660 24506 19716 24508
rect 19740 24506 19796 24508
rect 19820 24506 19876 24508
rect 19580 24454 19606 24506
rect 19606 24454 19636 24506
rect 19660 24454 19670 24506
rect 19670 24454 19716 24506
rect 19740 24454 19786 24506
rect 19786 24454 19796 24506
rect 19820 24454 19850 24506
rect 19850 24454 19876 24506
rect 19580 24452 19636 24454
rect 19660 24452 19716 24454
rect 19740 24452 19796 24454
rect 19820 24452 19876 24454
rect 19580 23418 19636 23420
rect 19660 23418 19716 23420
rect 19740 23418 19796 23420
rect 19820 23418 19876 23420
rect 19580 23366 19606 23418
rect 19606 23366 19636 23418
rect 19660 23366 19670 23418
rect 19670 23366 19716 23418
rect 19740 23366 19786 23418
rect 19786 23366 19796 23418
rect 19820 23366 19850 23418
rect 19850 23366 19876 23418
rect 19580 23364 19636 23366
rect 19660 23364 19716 23366
rect 19740 23364 19796 23366
rect 19820 23364 19876 23366
rect 19580 22330 19636 22332
rect 19660 22330 19716 22332
rect 19740 22330 19796 22332
rect 19820 22330 19876 22332
rect 19580 22278 19606 22330
rect 19606 22278 19636 22330
rect 19660 22278 19670 22330
rect 19670 22278 19716 22330
rect 19740 22278 19786 22330
rect 19786 22278 19796 22330
rect 19820 22278 19850 22330
rect 19850 22278 19876 22330
rect 19580 22276 19636 22278
rect 19660 22276 19716 22278
rect 19740 22276 19796 22278
rect 19820 22276 19876 22278
rect 8298 21392 8354 21448
rect 19580 21242 19636 21244
rect 19660 21242 19716 21244
rect 19740 21242 19796 21244
rect 19820 21242 19876 21244
rect 19580 21190 19606 21242
rect 19606 21190 19636 21242
rect 19660 21190 19670 21242
rect 19670 21190 19716 21242
rect 19740 21190 19786 21242
rect 19786 21190 19796 21242
rect 19820 21190 19850 21242
rect 19850 21190 19876 21242
rect 19580 21188 19636 21190
rect 19660 21188 19716 21190
rect 19740 21188 19796 21190
rect 19820 21188 19876 21190
rect 34940 44634 34996 44636
rect 35020 44634 35076 44636
rect 35100 44634 35156 44636
rect 35180 44634 35236 44636
rect 34940 44582 34966 44634
rect 34966 44582 34996 44634
rect 35020 44582 35030 44634
rect 35030 44582 35076 44634
rect 35100 44582 35146 44634
rect 35146 44582 35156 44634
rect 35180 44582 35210 44634
rect 35210 44582 35236 44634
rect 34940 44580 34996 44582
rect 35020 44580 35076 44582
rect 35100 44580 35156 44582
rect 35180 44580 35236 44582
rect 34940 43546 34996 43548
rect 35020 43546 35076 43548
rect 35100 43546 35156 43548
rect 35180 43546 35236 43548
rect 34940 43494 34966 43546
rect 34966 43494 34996 43546
rect 35020 43494 35030 43546
rect 35030 43494 35076 43546
rect 35100 43494 35146 43546
rect 35146 43494 35156 43546
rect 35180 43494 35210 43546
rect 35210 43494 35236 43546
rect 34940 43492 34996 43494
rect 35020 43492 35076 43494
rect 35100 43492 35156 43494
rect 35180 43492 35236 43494
rect 34940 42458 34996 42460
rect 35020 42458 35076 42460
rect 35100 42458 35156 42460
rect 35180 42458 35236 42460
rect 34940 42406 34966 42458
rect 34966 42406 34996 42458
rect 35020 42406 35030 42458
rect 35030 42406 35076 42458
rect 35100 42406 35146 42458
rect 35146 42406 35156 42458
rect 35180 42406 35210 42458
rect 35210 42406 35236 42458
rect 34940 42404 34996 42406
rect 35020 42404 35076 42406
rect 35100 42404 35156 42406
rect 35180 42404 35236 42406
rect 34940 41370 34996 41372
rect 35020 41370 35076 41372
rect 35100 41370 35156 41372
rect 35180 41370 35236 41372
rect 34940 41318 34966 41370
rect 34966 41318 34996 41370
rect 35020 41318 35030 41370
rect 35030 41318 35076 41370
rect 35100 41318 35146 41370
rect 35146 41318 35156 41370
rect 35180 41318 35210 41370
rect 35210 41318 35236 41370
rect 34940 41316 34996 41318
rect 35020 41316 35076 41318
rect 35100 41316 35156 41318
rect 35180 41316 35236 41318
rect 46938 49136 46994 49192
rect 46754 47640 46810 47696
rect 46846 46008 46902 46064
rect 34940 40282 34996 40284
rect 35020 40282 35076 40284
rect 35100 40282 35156 40284
rect 35180 40282 35236 40284
rect 34940 40230 34966 40282
rect 34966 40230 34996 40282
rect 35020 40230 35030 40282
rect 35030 40230 35076 40282
rect 35100 40230 35146 40282
rect 35146 40230 35156 40282
rect 35180 40230 35210 40282
rect 35210 40230 35236 40282
rect 34940 40228 34996 40230
rect 35020 40228 35076 40230
rect 35100 40228 35156 40230
rect 35180 40228 35236 40230
rect 34940 39194 34996 39196
rect 35020 39194 35076 39196
rect 35100 39194 35156 39196
rect 35180 39194 35236 39196
rect 34940 39142 34966 39194
rect 34966 39142 34996 39194
rect 35020 39142 35030 39194
rect 35030 39142 35076 39194
rect 35100 39142 35146 39194
rect 35146 39142 35156 39194
rect 35180 39142 35210 39194
rect 35210 39142 35236 39194
rect 34940 39140 34996 39142
rect 35020 39140 35076 39142
rect 35100 39140 35156 39142
rect 35180 39140 35236 39142
rect 34940 38106 34996 38108
rect 35020 38106 35076 38108
rect 35100 38106 35156 38108
rect 35180 38106 35236 38108
rect 34940 38054 34966 38106
rect 34966 38054 34996 38106
rect 35020 38054 35030 38106
rect 35030 38054 35076 38106
rect 35100 38054 35146 38106
rect 35146 38054 35156 38106
rect 35180 38054 35210 38106
rect 35210 38054 35236 38106
rect 34940 38052 34996 38054
rect 35020 38052 35076 38054
rect 35100 38052 35156 38054
rect 35180 38052 35236 38054
rect 34940 37018 34996 37020
rect 35020 37018 35076 37020
rect 35100 37018 35156 37020
rect 35180 37018 35236 37020
rect 34940 36966 34966 37018
rect 34966 36966 34996 37018
rect 35020 36966 35030 37018
rect 35030 36966 35076 37018
rect 35100 36966 35146 37018
rect 35146 36966 35156 37018
rect 35180 36966 35210 37018
rect 35210 36966 35236 37018
rect 34940 36964 34996 36966
rect 35020 36964 35076 36966
rect 35100 36964 35156 36966
rect 35180 36964 35236 36966
rect 34940 35930 34996 35932
rect 35020 35930 35076 35932
rect 35100 35930 35156 35932
rect 35180 35930 35236 35932
rect 34940 35878 34966 35930
rect 34966 35878 34996 35930
rect 35020 35878 35030 35930
rect 35030 35878 35076 35930
rect 35100 35878 35146 35930
rect 35146 35878 35156 35930
rect 35180 35878 35210 35930
rect 35210 35878 35236 35930
rect 34940 35876 34996 35878
rect 35020 35876 35076 35878
rect 35100 35876 35156 35878
rect 35180 35876 35236 35878
rect 34940 34842 34996 34844
rect 35020 34842 35076 34844
rect 35100 34842 35156 34844
rect 35180 34842 35236 34844
rect 34940 34790 34966 34842
rect 34966 34790 34996 34842
rect 35020 34790 35030 34842
rect 35030 34790 35076 34842
rect 35100 34790 35146 34842
rect 35146 34790 35156 34842
rect 35180 34790 35210 34842
rect 35210 34790 35236 34842
rect 34940 34788 34996 34790
rect 35020 34788 35076 34790
rect 35100 34788 35156 34790
rect 35180 34788 35236 34790
rect 34940 33754 34996 33756
rect 35020 33754 35076 33756
rect 35100 33754 35156 33756
rect 35180 33754 35236 33756
rect 34940 33702 34966 33754
rect 34966 33702 34996 33754
rect 35020 33702 35030 33754
rect 35030 33702 35076 33754
rect 35100 33702 35146 33754
rect 35146 33702 35156 33754
rect 35180 33702 35210 33754
rect 35210 33702 35236 33754
rect 34940 33700 34996 33702
rect 35020 33700 35076 33702
rect 35100 33700 35156 33702
rect 35180 33700 35236 33702
rect 34940 32666 34996 32668
rect 35020 32666 35076 32668
rect 35100 32666 35156 32668
rect 35180 32666 35236 32668
rect 34940 32614 34966 32666
rect 34966 32614 34996 32666
rect 35020 32614 35030 32666
rect 35030 32614 35076 32666
rect 35100 32614 35146 32666
rect 35146 32614 35156 32666
rect 35180 32614 35210 32666
rect 35210 32614 35236 32666
rect 34940 32612 34996 32614
rect 35020 32612 35076 32614
rect 35100 32612 35156 32614
rect 35180 32612 35236 32614
rect 34940 31578 34996 31580
rect 35020 31578 35076 31580
rect 35100 31578 35156 31580
rect 35180 31578 35236 31580
rect 34940 31526 34966 31578
rect 34966 31526 34996 31578
rect 35020 31526 35030 31578
rect 35030 31526 35076 31578
rect 35100 31526 35146 31578
rect 35146 31526 35156 31578
rect 35180 31526 35210 31578
rect 35210 31526 35236 31578
rect 34940 31524 34996 31526
rect 35020 31524 35076 31526
rect 35100 31524 35156 31526
rect 35180 31524 35236 31526
rect 34940 30490 34996 30492
rect 35020 30490 35076 30492
rect 35100 30490 35156 30492
rect 35180 30490 35236 30492
rect 34940 30438 34966 30490
rect 34966 30438 34996 30490
rect 35020 30438 35030 30490
rect 35030 30438 35076 30490
rect 35100 30438 35146 30490
rect 35146 30438 35156 30490
rect 35180 30438 35210 30490
rect 35210 30438 35236 30490
rect 34940 30436 34996 30438
rect 35020 30436 35076 30438
rect 35100 30436 35156 30438
rect 35180 30436 35236 30438
rect 34940 29402 34996 29404
rect 35020 29402 35076 29404
rect 35100 29402 35156 29404
rect 35180 29402 35236 29404
rect 34940 29350 34966 29402
rect 34966 29350 34996 29402
rect 35020 29350 35030 29402
rect 35030 29350 35076 29402
rect 35100 29350 35146 29402
rect 35146 29350 35156 29402
rect 35180 29350 35210 29402
rect 35210 29350 35236 29402
rect 34940 29348 34996 29350
rect 35020 29348 35076 29350
rect 35100 29348 35156 29350
rect 35180 29348 35236 29350
rect 39578 29300 39634 29336
rect 39578 29280 39580 29300
rect 39580 29280 39632 29300
rect 39632 29280 39634 29300
rect 34940 28314 34996 28316
rect 35020 28314 35076 28316
rect 35100 28314 35156 28316
rect 35180 28314 35236 28316
rect 34940 28262 34966 28314
rect 34966 28262 34996 28314
rect 35020 28262 35030 28314
rect 35030 28262 35076 28314
rect 35100 28262 35146 28314
rect 35146 28262 35156 28314
rect 35180 28262 35210 28314
rect 35210 28262 35236 28314
rect 34940 28260 34996 28262
rect 35020 28260 35076 28262
rect 35100 28260 35156 28262
rect 35180 28260 35236 28262
rect 34940 27226 34996 27228
rect 35020 27226 35076 27228
rect 35100 27226 35156 27228
rect 35180 27226 35236 27228
rect 34940 27174 34966 27226
rect 34966 27174 34996 27226
rect 35020 27174 35030 27226
rect 35030 27174 35076 27226
rect 35100 27174 35146 27226
rect 35146 27174 35156 27226
rect 35180 27174 35210 27226
rect 35210 27174 35236 27226
rect 34940 27172 34996 27174
rect 35020 27172 35076 27174
rect 35100 27172 35156 27174
rect 35180 27172 35236 27174
rect 38382 27124 38438 27160
rect 38382 27104 38384 27124
rect 38384 27104 38436 27124
rect 38436 27104 38438 27124
rect 34940 26138 34996 26140
rect 35020 26138 35076 26140
rect 35100 26138 35156 26140
rect 35180 26138 35236 26140
rect 34940 26086 34966 26138
rect 34966 26086 34996 26138
rect 35020 26086 35030 26138
rect 35030 26086 35076 26138
rect 35100 26086 35146 26138
rect 35146 26086 35156 26138
rect 35180 26086 35210 26138
rect 35210 26086 35236 26138
rect 34940 26084 34996 26086
rect 35020 26084 35076 26086
rect 35100 26084 35156 26086
rect 35180 26084 35236 26086
rect 35990 25220 36046 25256
rect 35990 25200 35992 25220
rect 35992 25200 36044 25220
rect 36044 25200 36046 25220
rect 34940 25050 34996 25052
rect 35020 25050 35076 25052
rect 35100 25050 35156 25052
rect 35180 25050 35236 25052
rect 34940 24998 34966 25050
rect 34966 24998 34996 25050
rect 35020 24998 35030 25050
rect 35030 24998 35076 25050
rect 35100 24998 35146 25050
rect 35146 24998 35156 25050
rect 35180 24998 35210 25050
rect 35210 24998 35236 25050
rect 34940 24996 34996 24998
rect 35020 24996 35076 24998
rect 35100 24996 35156 24998
rect 35180 24996 35236 24998
rect 31298 24112 31354 24168
rect 34940 23962 34996 23964
rect 35020 23962 35076 23964
rect 35100 23962 35156 23964
rect 35180 23962 35236 23964
rect 34940 23910 34966 23962
rect 34966 23910 34996 23962
rect 35020 23910 35030 23962
rect 35030 23910 35076 23962
rect 35100 23910 35146 23962
rect 35146 23910 35156 23962
rect 35180 23910 35210 23962
rect 35210 23910 35236 23962
rect 34940 23908 34996 23910
rect 35020 23908 35076 23910
rect 35100 23908 35156 23910
rect 35180 23908 35236 23910
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 27618 20576 27674 20632
rect 29642 21412 29698 21448
rect 30286 21936 30342 21992
rect 29642 21392 29644 21412
rect 29644 21392 29696 21412
rect 29696 21392 29698 21412
rect 28262 20712 28318 20768
rect 33598 23044 33654 23080
rect 33598 23024 33600 23044
rect 33600 23024 33652 23044
rect 33652 23024 33654 23044
rect 34940 22874 34996 22876
rect 35020 22874 35076 22876
rect 35100 22874 35156 22876
rect 35180 22874 35236 22876
rect 34940 22822 34966 22874
rect 34966 22822 34996 22874
rect 35020 22822 35030 22874
rect 35030 22822 35076 22874
rect 35100 22822 35146 22874
rect 35146 22822 35156 22874
rect 35180 22822 35210 22874
rect 35210 22822 35236 22874
rect 34940 22820 34996 22822
rect 35020 22820 35076 22822
rect 35100 22820 35156 22822
rect 35180 22820 35236 22822
rect 38198 25608 38254 25664
rect 36174 22924 36176 22944
rect 36176 22924 36228 22944
rect 36228 22924 36230 22944
rect 36174 22888 36230 22924
rect 36634 22888 36690 22944
rect 19580 20154 19636 20156
rect 19660 20154 19716 20156
rect 19740 20154 19796 20156
rect 19820 20154 19876 20156
rect 19580 20102 19606 20154
rect 19606 20102 19636 20154
rect 19660 20102 19670 20154
rect 19670 20102 19716 20154
rect 19740 20102 19786 20154
rect 19786 20102 19796 20154
rect 19820 20102 19850 20154
rect 19850 20102 19876 20154
rect 19580 20100 19636 20102
rect 19660 20100 19716 20102
rect 19740 20100 19796 20102
rect 19820 20100 19876 20102
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 19580 19066 19636 19068
rect 19660 19066 19716 19068
rect 19740 19066 19796 19068
rect 19820 19066 19876 19068
rect 19580 19014 19606 19066
rect 19606 19014 19636 19066
rect 19660 19014 19670 19066
rect 19670 19014 19716 19066
rect 19740 19014 19786 19066
rect 19786 19014 19796 19066
rect 19820 19014 19850 19066
rect 19850 19014 19876 19066
rect 19580 19012 19636 19014
rect 19660 19012 19716 19014
rect 19740 19012 19796 19014
rect 19820 19012 19876 19014
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 19580 17978 19636 17980
rect 19660 17978 19716 17980
rect 19740 17978 19796 17980
rect 19820 17978 19876 17980
rect 19580 17926 19606 17978
rect 19606 17926 19636 17978
rect 19660 17926 19670 17978
rect 19670 17926 19716 17978
rect 19740 17926 19786 17978
rect 19786 17926 19796 17978
rect 19820 17926 19850 17978
rect 19850 17926 19876 17978
rect 19580 17924 19636 17926
rect 19660 17924 19716 17926
rect 19740 17924 19796 17926
rect 19820 17924 19876 17926
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 3422 17040 3478 17096
rect 23478 17060 23534 17096
rect 23478 17040 23480 17060
rect 23480 17040 23532 17060
rect 23532 17040 23534 17060
rect 19580 16890 19636 16892
rect 19660 16890 19716 16892
rect 19740 16890 19796 16892
rect 19820 16890 19876 16892
rect 19580 16838 19606 16890
rect 19606 16838 19636 16890
rect 19660 16838 19670 16890
rect 19670 16838 19716 16890
rect 19740 16838 19786 16890
rect 19786 16838 19796 16890
rect 19820 16838 19850 16890
rect 19850 16838 19876 16890
rect 19580 16836 19636 16838
rect 19660 16836 19716 16838
rect 19740 16836 19796 16838
rect 19820 16836 19876 16838
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 26514 16768 26570 16824
rect 19580 15802 19636 15804
rect 19660 15802 19716 15804
rect 19740 15802 19796 15804
rect 19820 15802 19876 15804
rect 19580 15750 19606 15802
rect 19606 15750 19636 15802
rect 19660 15750 19670 15802
rect 19670 15750 19716 15802
rect 19740 15750 19786 15802
rect 19786 15750 19796 15802
rect 19820 15750 19850 15802
rect 19850 15750 19876 15802
rect 19580 15748 19636 15750
rect 19660 15748 19716 15750
rect 19740 15748 19796 15750
rect 19820 15748 19876 15750
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 19580 14714 19636 14716
rect 19660 14714 19716 14716
rect 19740 14714 19796 14716
rect 19820 14714 19876 14716
rect 19580 14662 19606 14714
rect 19606 14662 19636 14714
rect 19660 14662 19670 14714
rect 19670 14662 19716 14714
rect 19740 14662 19786 14714
rect 19786 14662 19796 14714
rect 19820 14662 19850 14714
rect 19850 14662 19876 14714
rect 19580 14660 19636 14662
rect 19660 14660 19716 14662
rect 19740 14660 19796 14662
rect 19820 14660 19876 14662
rect 20258 14456 20314 14512
rect 8390 14340 8446 14376
rect 8390 14320 8392 14340
rect 8392 14320 8444 14340
rect 8444 14320 8446 14340
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 7010 12724 7012 12744
rect 7012 12724 7064 12744
rect 7064 12724 7066 12744
rect 7010 12688 7066 12724
rect 5446 11600 5502 11656
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 5262 10804 5318 10840
rect 5262 10784 5264 10804
rect 5264 10784 5316 10804
rect 5316 10784 5318 10804
rect 5354 10124 5410 10160
rect 5354 10104 5356 10124
rect 5356 10104 5408 10124
rect 5408 10104 5410 10124
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 8298 12724 8300 12744
rect 8300 12724 8352 12744
rect 8352 12724 8354 12744
rect 8298 12688 8354 12724
rect 19580 13626 19636 13628
rect 19660 13626 19716 13628
rect 19740 13626 19796 13628
rect 19820 13626 19876 13628
rect 19580 13574 19606 13626
rect 19606 13574 19636 13626
rect 19660 13574 19670 13626
rect 19670 13574 19716 13626
rect 19740 13574 19786 13626
rect 19786 13574 19796 13626
rect 19820 13574 19850 13626
rect 19850 13574 19876 13626
rect 19580 13572 19636 13574
rect 19660 13572 19716 13574
rect 19740 13572 19796 13574
rect 19820 13572 19876 13574
rect 9954 12300 10010 12336
rect 19580 12538 19636 12540
rect 19660 12538 19716 12540
rect 19740 12538 19796 12540
rect 19820 12538 19876 12540
rect 19580 12486 19606 12538
rect 19606 12486 19636 12538
rect 19660 12486 19670 12538
rect 19670 12486 19716 12538
rect 19740 12486 19786 12538
rect 19786 12486 19796 12538
rect 19820 12486 19850 12538
rect 19850 12486 19876 12538
rect 19580 12484 19636 12486
rect 19660 12484 19716 12486
rect 19740 12484 19796 12486
rect 19820 12484 19876 12486
rect 9954 12280 9956 12300
rect 9956 12280 10008 12300
rect 10008 12280 10010 12300
rect 6918 10104 6974 10160
rect 662 3032 718 3088
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 2502 3460 2558 3496
rect 2502 3440 2504 3460
rect 2504 3440 2556 3460
rect 2556 3440 2558 3460
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 4710 3440 4766 3496
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 11150 11636 11152 11656
rect 11152 11636 11204 11656
rect 11204 11636 11206 11656
rect 11150 11600 11206 11636
rect 10414 11076 10470 11112
rect 10414 11056 10416 11076
rect 10416 11056 10468 11076
rect 10468 11056 10470 11076
rect 11058 10804 11114 10840
rect 11058 10784 11060 10804
rect 11060 10784 11112 10804
rect 11112 10784 11114 10804
rect 6274 6704 6330 6760
rect 9586 7268 9642 7304
rect 9586 7248 9588 7268
rect 9588 7248 9640 7268
rect 9640 7248 9642 7268
rect 5998 3848 6054 3904
rect 8666 6180 8722 6216
rect 8666 6160 8668 6180
rect 8668 6160 8720 6180
rect 8720 6160 8722 6180
rect 9586 4800 9642 4856
rect 8206 4548 8262 4584
rect 8206 4528 8208 4548
rect 8208 4528 8260 4548
rect 8260 4528 8262 4548
rect 7838 3984 7894 4040
rect 8758 4004 8814 4040
rect 7562 2760 7618 2816
rect 8758 3984 8760 4004
rect 8760 3984 8812 4004
rect 8812 3984 8814 4004
rect 11426 10684 11428 10704
rect 11428 10684 11480 10704
rect 11480 10684 11482 10704
rect 11426 10648 11482 10684
rect 12530 11464 12586 11520
rect 12990 11056 13046 11112
rect 18878 12280 18934 12336
rect 20442 12824 20498 12880
rect 15474 11500 15476 11520
rect 15476 11500 15528 11520
rect 15528 11500 15530 11520
rect 15474 11464 15530 11500
rect 20994 12824 21050 12880
rect 12254 9560 12310 9616
rect 11794 7248 11850 7304
rect 10046 6704 10102 6760
rect 11334 6160 11390 6216
rect 11058 5636 11114 5672
rect 11058 5616 11060 5636
rect 11060 5616 11112 5636
rect 11112 5616 11114 5636
rect 15106 8336 15162 8392
rect 10230 4256 10286 4312
rect 11518 4528 11574 4584
rect 11702 4820 11758 4856
rect 11702 4800 11704 4820
rect 11704 4800 11756 4820
rect 11756 4800 11758 4820
rect 11610 4392 11666 4448
rect 11978 4156 11980 4176
rect 11980 4156 12032 4176
rect 12032 4156 12034 4176
rect 11978 4120 12034 4156
rect 13358 4256 13414 4312
rect 9954 3848 10010 3904
rect 10322 3884 10324 3904
rect 10324 3884 10376 3904
rect 10376 3884 10378 3904
rect 10322 3848 10378 3884
rect 10046 2760 10102 2816
rect 12806 3848 12862 3904
rect 15658 9560 15714 9616
rect 19580 11450 19636 11452
rect 19660 11450 19716 11452
rect 19740 11450 19796 11452
rect 19820 11450 19876 11452
rect 19580 11398 19606 11450
rect 19606 11398 19636 11450
rect 19660 11398 19670 11450
rect 19670 11398 19716 11450
rect 19740 11398 19786 11450
rect 19786 11398 19796 11450
rect 19820 11398 19850 11450
rect 19850 11398 19876 11450
rect 19580 11396 19636 11398
rect 19660 11396 19716 11398
rect 19740 11396 19796 11398
rect 19820 11396 19876 11398
rect 16946 8356 17002 8392
rect 16946 8336 16948 8356
rect 16948 8336 17000 8356
rect 17000 8336 17002 8356
rect 13910 4392 13966 4448
rect 13818 4256 13874 4312
rect 16118 4392 16174 4448
rect 17406 5616 17462 5672
rect 16486 3848 16542 3904
rect 15474 3460 15530 3496
rect 15474 3440 15476 3460
rect 15476 3440 15528 3460
rect 15528 3440 15530 3460
rect 16486 3340 16488 3360
rect 16488 3340 16540 3360
rect 16540 3340 16542 3360
rect 16486 3304 16542 3340
rect 16854 2896 16910 2952
rect 18142 3984 18198 4040
rect 18694 3304 18750 3360
rect 20258 10668 20314 10704
rect 20258 10648 20260 10668
rect 20260 10648 20312 10668
rect 20312 10648 20314 10668
rect 20442 10648 20498 10704
rect 19580 10362 19636 10364
rect 19660 10362 19716 10364
rect 19740 10362 19796 10364
rect 19820 10362 19876 10364
rect 19580 10310 19606 10362
rect 19606 10310 19636 10362
rect 19660 10310 19670 10362
rect 19670 10310 19716 10362
rect 19740 10310 19786 10362
rect 19786 10310 19796 10362
rect 19820 10310 19850 10362
rect 19850 10310 19876 10362
rect 19580 10308 19636 10310
rect 19660 10308 19716 10310
rect 19740 10308 19796 10310
rect 19820 10308 19876 10310
rect 22282 12280 22338 12336
rect 21362 11892 21418 11928
rect 21362 11872 21364 11892
rect 21364 11872 21416 11892
rect 21416 11872 21418 11892
rect 25042 11892 25098 11928
rect 25042 11872 25044 11892
rect 25044 11872 25096 11892
rect 25096 11872 25098 11892
rect 23662 11192 23718 11248
rect 22098 10648 22154 10704
rect 19580 9274 19636 9276
rect 19660 9274 19716 9276
rect 19740 9274 19796 9276
rect 19820 9274 19876 9276
rect 19580 9222 19606 9274
rect 19606 9222 19636 9274
rect 19660 9222 19670 9274
rect 19670 9222 19716 9274
rect 19740 9222 19786 9274
rect 19786 9222 19796 9274
rect 19820 9222 19850 9274
rect 19850 9222 19876 9274
rect 19580 9220 19636 9222
rect 19660 9220 19716 9222
rect 19740 9220 19796 9222
rect 19820 9220 19876 9222
rect 19580 8186 19636 8188
rect 19660 8186 19716 8188
rect 19740 8186 19796 8188
rect 19820 8186 19876 8188
rect 19580 8134 19606 8186
rect 19606 8134 19636 8186
rect 19660 8134 19670 8186
rect 19670 8134 19716 8186
rect 19740 8134 19786 8186
rect 19786 8134 19796 8186
rect 19820 8134 19850 8186
rect 19850 8134 19876 8186
rect 19580 8132 19636 8134
rect 19660 8132 19716 8134
rect 19740 8132 19796 8134
rect 19820 8132 19876 8134
rect 26606 11212 26662 11248
rect 26606 11192 26608 11212
rect 26608 11192 26660 11212
rect 26660 11192 26662 11212
rect 25410 10260 25466 10296
rect 25410 10240 25412 10260
rect 25412 10240 25464 10260
rect 25464 10240 25466 10260
rect 19580 7098 19636 7100
rect 19660 7098 19716 7100
rect 19740 7098 19796 7100
rect 19820 7098 19876 7100
rect 19580 7046 19606 7098
rect 19606 7046 19636 7098
rect 19660 7046 19670 7098
rect 19670 7046 19716 7098
rect 19740 7046 19786 7098
rect 19786 7046 19796 7098
rect 19820 7046 19850 7098
rect 19850 7046 19876 7098
rect 19580 7044 19636 7046
rect 19660 7044 19716 7046
rect 19740 7044 19796 7046
rect 19820 7044 19876 7046
rect 19580 6010 19636 6012
rect 19660 6010 19716 6012
rect 19740 6010 19796 6012
rect 19820 6010 19876 6012
rect 19580 5958 19606 6010
rect 19606 5958 19636 6010
rect 19660 5958 19670 6010
rect 19670 5958 19716 6010
rect 19740 5958 19786 6010
rect 19786 5958 19796 6010
rect 19820 5958 19850 6010
rect 19850 5958 19876 6010
rect 19580 5956 19636 5958
rect 19660 5956 19716 5958
rect 19740 5956 19796 5958
rect 19820 5956 19876 5958
rect 20994 5888 21050 5944
rect 19580 4922 19636 4924
rect 19660 4922 19716 4924
rect 19740 4922 19796 4924
rect 19820 4922 19876 4924
rect 19580 4870 19606 4922
rect 19606 4870 19636 4922
rect 19660 4870 19670 4922
rect 19670 4870 19716 4922
rect 19740 4870 19786 4922
rect 19786 4870 19796 4922
rect 19820 4870 19850 4922
rect 19850 4870 19876 4922
rect 19580 4868 19636 4870
rect 19660 4868 19716 4870
rect 19740 4868 19796 4870
rect 19820 4868 19876 4870
rect 19982 4800 20038 4856
rect 19338 4120 19394 4176
rect 19338 3848 19394 3904
rect 19580 3834 19636 3836
rect 19660 3834 19716 3836
rect 19740 3834 19796 3836
rect 19820 3834 19876 3836
rect 19580 3782 19606 3834
rect 19606 3782 19636 3834
rect 19660 3782 19670 3834
rect 19670 3782 19716 3834
rect 19740 3782 19786 3834
rect 19786 3782 19796 3834
rect 19820 3782 19850 3834
rect 19850 3782 19876 3834
rect 19580 3780 19636 3782
rect 19660 3780 19716 3782
rect 19740 3780 19796 3782
rect 19820 3780 19876 3782
rect 19430 3576 19486 3632
rect 19246 3168 19302 3224
rect 21086 5480 21142 5536
rect 22558 5652 22560 5672
rect 22560 5652 22612 5672
rect 22612 5652 22614 5672
rect 22558 5616 22614 5652
rect 22558 4820 22614 4856
rect 22558 4800 22560 4820
rect 22560 4800 22612 4820
rect 22612 4800 22614 4820
rect 20718 3460 20774 3496
rect 31022 20712 31078 20768
rect 32402 20576 32458 20632
rect 34610 21936 34666 21992
rect 34940 21786 34996 21788
rect 35020 21786 35076 21788
rect 35100 21786 35156 21788
rect 35180 21786 35236 21788
rect 34940 21734 34966 21786
rect 34966 21734 34996 21786
rect 35020 21734 35030 21786
rect 35030 21734 35076 21786
rect 35100 21734 35146 21786
rect 35146 21734 35156 21786
rect 35180 21734 35210 21786
rect 35210 21734 35236 21786
rect 34940 21732 34996 21734
rect 35020 21732 35076 21734
rect 35100 21732 35156 21734
rect 35180 21732 35236 21734
rect 32770 20032 32826 20088
rect 34940 20698 34996 20700
rect 35020 20698 35076 20700
rect 35100 20698 35156 20700
rect 35180 20698 35236 20700
rect 34940 20646 34966 20698
rect 34966 20646 34996 20698
rect 35020 20646 35030 20698
rect 35030 20646 35076 20698
rect 35100 20646 35146 20698
rect 35146 20646 35156 20698
rect 35180 20646 35210 20698
rect 35210 20646 35236 20698
rect 34940 20644 34996 20646
rect 35020 20644 35076 20646
rect 35100 20644 35156 20646
rect 35180 20644 35236 20646
rect 35622 20576 35678 20632
rect 32402 19352 32458 19408
rect 29918 16768 29974 16824
rect 30378 16768 30434 16824
rect 30286 13776 30342 13832
rect 31758 13776 31814 13832
rect 27526 12824 27582 12880
rect 31022 12588 31024 12608
rect 31024 12588 31076 12608
rect 31076 12588 31078 12608
rect 31022 12552 31078 12588
rect 29642 11872 29698 11928
rect 27250 10648 27306 10704
rect 27986 10240 28042 10296
rect 28814 10240 28870 10296
rect 26054 10140 26056 10160
rect 26056 10140 26108 10160
rect 26108 10140 26110 10160
rect 26054 10104 26110 10140
rect 25502 10004 25504 10024
rect 25504 10004 25556 10024
rect 25556 10004 25558 10024
rect 25502 9968 25558 10004
rect 27158 9968 27214 10024
rect 23846 5480 23902 5536
rect 23754 5364 23810 5400
rect 23754 5344 23756 5364
rect 23756 5344 23808 5364
rect 23808 5344 23810 5364
rect 23110 4120 23166 4176
rect 23110 3884 23112 3904
rect 23112 3884 23164 3904
rect 23164 3884 23166 3904
rect 23110 3848 23166 3884
rect 20718 3440 20720 3460
rect 20720 3440 20772 3460
rect 20772 3440 20774 3460
rect 22190 3304 22246 3360
rect 19580 2746 19636 2748
rect 19660 2746 19716 2748
rect 19740 2746 19796 2748
rect 19820 2746 19876 2748
rect 19580 2694 19606 2746
rect 19606 2694 19636 2746
rect 19660 2694 19670 2746
rect 19670 2694 19716 2746
rect 19740 2694 19786 2746
rect 19786 2694 19796 2746
rect 19820 2694 19850 2746
rect 19850 2694 19876 2746
rect 19580 2692 19636 2694
rect 19660 2692 19716 2694
rect 19740 2692 19796 2694
rect 19820 2692 19876 2694
rect 20902 2760 20958 2816
rect 22282 2916 22338 2952
rect 22282 2896 22284 2916
rect 22284 2896 22336 2916
rect 22336 2896 22338 2916
rect 23754 3848 23810 3904
rect 26238 6332 26240 6352
rect 26240 6332 26292 6352
rect 26292 6332 26294 6352
rect 26238 6296 26294 6332
rect 25594 5616 25650 5672
rect 25594 4564 25596 4584
rect 25596 4564 25648 4584
rect 25648 4564 25650 4584
rect 25594 4528 25650 4564
rect 26054 4120 26110 4176
rect 24766 4020 24768 4040
rect 24768 4020 24820 4040
rect 24820 4020 24822 4040
rect 24766 3984 24822 4020
rect 25686 3984 25742 4040
rect 24582 3576 24638 3632
rect 23846 3460 23902 3496
rect 23846 3440 23848 3460
rect 23848 3440 23900 3460
rect 23900 3440 23902 3460
rect 25594 2796 25596 2816
rect 25596 2796 25648 2816
rect 25648 2796 25650 2816
rect 25594 2760 25650 2796
rect 27710 7420 27712 7440
rect 27712 7420 27764 7440
rect 27764 7420 27766 7440
rect 27710 7384 27766 7420
rect 30470 10240 30526 10296
rect 28170 7248 28226 7304
rect 26514 4528 26570 4584
rect 30746 7248 30802 7304
rect 29274 5344 29330 5400
rect 26422 3848 26478 3904
rect 26238 3168 26294 3224
rect 27710 3984 27766 4040
rect 26790 3032 26846 3088
rect 28078 3884 28080 3904
rect 28080 3884 28132 3904
rect 28132 3884 28134 3904
rect 28078 3848 28134 3884
rect 28170 3576 28226 3632
rect 27618 3460 27674 3496
rect 27618 3440 27620 3460
rect 27620 3440 27672 3460
rect 27672 3440 27674 3460
rect 30930 5888 30986 5944
rect 28446 3168 28502 3224
rect 29090 3068 29092 3088
rect 29092 3068 29144 3088
rect 29144 3068 29146 3088
rect 29090 3032 29146 3068
rect 30194 2896 30250 2952
rect 30470 3848 30526 3904
rect 30378 3712 30434 3768
rect 31850 4548 31906 4584
rect 31850 4528 31852 4548
rect 31852 4528 31904 4548
rect 31904 4528 31906 4548
rect 32126 11892 32182 11928
rect 32126 11872 32128 11892
rect 32128 11872 32180 11892
rect 32180 11872 32182 11892
rect 32402 6316 32458 6352
rect 32402 6296 32404 6316
rect 32404 6296 32456 6316
rect 32456 6296 32458 6316
rect 34794 20032 34850 20088
rect 34978 19916 35034 19952
rect 34978 19896 34980 19916
rect 34980 19896 35032 19916
rect 35032 19896 35034 19916
rect 34702 19352 34758 19408
rect 34940 19610 34996 19612
rect 35020 19610 35076 19612
rect 35100 19610 35156 19612
rect 35180 19610 35236 19612
rect 34940 19558 34966 19610
rect 34966 19558 34996 19610
rect 35020 19558 35030 19610
rect 35030 19558 35076 19610
rect 35100 19558 35146 19610
rect 35146 19558 35156 19610
rect 35180 19558 35210 19610
rect 35210 19558 35236 19610
rect 34940 19556 34996 19558
rect 35020 19556 35076 19558
rect 35100 19556 35156 19558
rect 35180 19556 35236 19558
rect 34940 18522 34996 18524
rect 35020 18522 35076 18524
rect 35100 18522 35156 18524
rect 35180 18522 35236 18524
rect 34940 18470 34966 18522
rect 34966 18470 34996 18522
rect 35020 18470 35030 18522
rect 35030 18470 35076 18522
rect 35100 18470 35146 18522
rect 35146 18470 35156 18522
rect 35180 18470 35210 18522
rect 35210 18470 35236 18522
rect 34940 18468 34996 18470
rect 35020 18468 35076 18470
rect 35100 18468 35156 18470
rect 35180 18468 35236 18470
rect 34940 17434 34996 17436
rect 35020 17434 35076 17436
rect 35100 17434 35156 17436
rect 35180 17434 35236 17436
rect 34940 17382 34966 17434
rect 34966 17382 34996 17434
rect 35020 17382 35030 17434
rect 35030 17382 35076 17434
rect 35100 17382 35146 17434
rect 35146 17382 35156 17434
rect 35180 17382 35210 17434
rect 35210 17382 35236 17434
rect 34940 17380 34996 17382
rect 35020 17380 35076 17382
rect 35100 17380 35156 17382
rect 35180 17380 35236 17382
rect 34940 16346 34996 16348
rect 35020 16346 35076 16348
rect 35100 16346 35156 16348
rect 35180 16346 35236 16348
rect 34940 16294 34966 16346
rect 34966 16294 34996 16346
rect 35020 16294 35030 16346
rect 35030 16294 35076 16346
rect 35100 16294 35146 16346
rect 35146 16294 35156 16346
rect 35180 16294 35210 16346
rect 35210 16294 35236 16346
rect 34940 16292 34996 16294
rect 35020 16292 35076 16294
rect 35100 16292 35156 16294
rect 35180 16292 35236 16294
rect 34940 15258 34996 15260
rect 35020 15258 35076 15260
rect 35100 15258 35156 15260
rect 35180 15258 35236 15260
rect 34940 15206 34966 15258
rect 34966 15206 34996 15258
rect 35020 15206 35030 15258
rect 35030 15206 35076 15258
rect 35100 15206 35146 15258
rect 35146 15206 35156 15258
rect 35180 15206 35210 15258
rect 35210 15206 35236 15258
rect 34940 15204 34996 15206
rect 35020 15204 35076 15206
rect 35100 15204 35156 15206
rect 35180 15204 35236 15206
rect 34940 14170 34996 14172
rect 35020 14170 35076 14172
rect 35100 14170 35156 14172
rect 35180 14170 35236 14172
rect 34940 14118 34966 14170
rect 34966 14118 34996 14170
rect 35020 14118 35030 14170
rect 35030 14118 35076 14170
rect 35100 14118 35146 14170
rect 35146 14118 35156 14170
rect 35180 14118 35210 14170
rect 35210 14118 35236 14170
rect 34940 14116 34996 14118
rect 35020 14116 35076 14118
rect 35100 14116 35156 14118
rect 35180 14116 35236 14118
rect 35162 13812 35164 13832
rect 35164 13812 35216 13832
rect 35216 13812 35218 13832
rect 35162 13776 35218 13812
rect 35622 18844 35624 18864
rect 35624 18844 35676 18864
rect 35676 18844 35678 18864
rect 35622 18808 35678 18844
rect 35530 17212 35532 17232
rect 35532 17212 35584 17232
rect 35584 17212 35586 17232
rect 35530 17176 35586 17212
rect 39578 25472 39634 25528
rect 38658 24692 38660 24712
rect 38660 24692 38712 24712
rect 38712 24692 38714 24712
rect 38658 24656 38714 24692
rect 41234 28872 41290 28928
rect 42062 28872 42118 28928
rect 41694 27920 41750 27976
rect 40590 25608 40646 25664
rect 41970 25472 42026 25528
rect 41050 24792 41106 24848
rect 40314 24112 40370 24168
rect 43626 30640 43682 30696
rect 42430 29280 42486 29336
rect 42246 27412 42248 27432
rect 42248 27412 42300 27432
rect 42300 27412 42302 27432
rect 42246 27376 42302 27412
rect 42338 24656 42394 24712
rect 44546 27956 44548 27976
rect 44548 27956 44600 27976
rect 44600 27956 44602 27976
rect 44546 27920 44602 27956
rect 45190 27376 45246 27432
rect 45282 26732 45284 26752
rect 45284 26732 45336 26752
rect 45336 26732 45338 26752
rect 45282 26696 45338 26732
rect 45190 26324 45192 26344
rect 45192 26324 45244 26344
rect 45244 26324 45246 26344
rect 45190 26288 45246 26324
rect 45650 24792 45706 24848
rect 43442 24112 43498 24168
rect 40498 22924 40500 22944
rect 40500 22924 40552 22944
rect 40552 22924 40554 22944
rect 40498 22888 40554 22924
rect 36174 14456 36230 14512
rect 38198 20712 38254 20768
rect 38290 20032 38346 20088
rect 37278 17176 37334 17232
rect 38106 18828 38162 18864
rect 38106 18808 38108 18828
rect 38108 18808 38160 18828
rect 38160 18808 38162 18828
rect 39854 19896 39910 19952
rect 41602 21972 41604 21992
rect 41604 21972 41656 21992
rect 41656 21972 41658 21992
rect 41602 21936 41658 21972
rect 40590 20596 40646 20632
rect 40590 20576 40592 20596
rect 40592 20576 40644 20596
rect 40644 20576 40646 20596
rect 40774 20748 40776 20768
rect 40776 20748 40828 20768
rect 40828 20748 40830 20768
rect 40774 20712 40830 20748
rect 38566 19252 38568 19272
rect 38568 19252 38620 19272
rect 38620 19252 38622 19272
rect 38566 19216 38622 19252
rect 36634 14320 36690 14376
rect 35714 13812 35716 13832
rect 35716 13812 35768 13832
rect 35768 13812 35770 13832
rect 35714 13776 35770 13812
rect 34940 13082 34996 13084
rect 35020 13082 35076 13084
rect 35100 13082 35156 13084
rect 35180 13082 35236 13084
rect 34940 13030 34966 13082
rect 34966 13030 34996 13082
rect 35020 13030 35030 13082
rect 35030 13030 35076 13082
rect 35100 13030 35146 13082
rect 35146 13030 35156 13082
rect 35180 13030 35210 13082
rect 35210 13030 35236 13082
rect 34940 13028 34996 13030
rect 35020 13028 35076 13030
rect 35100 13028 35156 13030
rect 35180 13028 35236 13030
rect 34940 11994 34996 11996
rect 35020 11994 35076 11996
rect 35100 11994 35156 11996
rect 35180 11994 35236 11996
rect 34940 11942 34966 11994
rect 34966 11942 34996 11994
rect 35020 11942 35030 11994
rect 35030 11942 35076 11994
rect 35100 11942 35146 11994
rect 35146 11942 35156 11994
rect 35180 11942 35210 11994
rect 35210 11942 35236 11994
rect 34940 11940 34996 11942
rect 35020 11940 35076 11942
rect 35100 11940 35156 11942
rect 35180 11940 35236 11942
rect 34940 10906 34996 10908
rect 35020 10906 35076 10908
rect 35100 10906 35156 10908
rect 35180 10906 35236 10908
rect 34940 10854 34966 10906
rect 34966 10854 34996 10906
rect 35020 10854 35030 10906
rect 35030 10854 35076 10906
rect 35100 10854 35146 10906
rect 35146 10854 35156 10906
rect 35180 10854 35210 10906
rect 35210 10854 35236 10906
rect 34940 10852 34996 10854
rect 35020 10852 35076 10854
rect 35100 10852 35156 10854
rect 35180 10852 35236 10854
rect 33230 10104 33286 10160
rect 34940 9818 34996 9820
rect 35020 9818 35076 9820
rect 35100 9818 35156 9820
rect 35180 9818 35236 9820
rect 34940 9766 34966 9818
rect 34966 9766 34996 9818
rect 35020 9766 35030 9818
rect 35030 9766 35076 9818
rect 35100 9766 35146 9818
rect 35146 9766 35156 9818
rect 35180 9766 35210 9818
rect 35210 9766 35236 9818
rect 34940 9764 34996 9766
rect 35020 9764 35076 9766
rect 35100 9764 35156 9766
rect 35180 9764 35236 9766
rect 35438 9696 35494 9752
rect 34940 8730 34996 8732
rect 35020 8730 35076 8732
rect 35100 8730 35156 8732
rect 35180 8730 35236 8732
rect 34940 8678 34966 8730
rect 34966 8678 34996 8730
rect 35020 8678 35030 8730
rect 35030 8678 35076 8730
rect 35100 8678 35146 8730
rect 35146 8678 35156 8730
rect 35180 8678 35210 8730
rect 35210 8678 35236 8730
rect 34940 8676 34996 8678
rect 35020 8676 35076 8678
rect 35100 8676 35156 8678
rect 35180 8676 35236 8678
rect 34940 7642 34996 7644
rect 35020 7642 35076 7644
rect 35100 7642 35156 7644
rect 35180 7642 35236 7644
rect 34940 7590 34966 7642
rect 34966 7590 34996 7642
rect 35020 7590 35030 7642
rect 35030 7590 35076 7642
rect 35100 7590 35146 7642
rect 35146 7590 35156 7642
rect 35180 7590 35210 7642
rect 35210 7590 35236 7642
rect 34940 7588 34996 7590
rect 35020 7588 35076 7590
rect 35100 7588 35156 7590
rect 35180 7588 35236 7590
rect 33598 7384 33654 7440
rect 33322 6180 33378 6216
rect 33322 6160 33324 6180
rect 33324 6160 33376 6180
rect 33376 6160 33378 6180
rect 34940 6554 34996 6556
rect 35020 6554 35076 6556
rect 35100 6554 35156 6556
rect 35180 6554 35236 6556
rect 34940 6502 34966 6554
rect 34966 6502 34996 6554
rect 35020 6502 35030 6554
rect 35030 6502 35076 6554
rect 35100 6502 35146 6554
rect 35146 6502 35156 6554
rect 35180 6502 35210 6554
rect 35210 6502 35236 6554
rect 34940 6500 34996 6502
rect 35020 6500 35076 6502
rect 35100 6500 35156 6502
rect 35180 6500 35236 6502
rect 34940 5466 34996 5468
rect 35020 5466 35076 5468
rect 35100 5466 35156 5468
rect 35180 5466 35236 5468
rect 34940 5414 34966 5466
rect 34966 5414 34996 5466
rect 35020 5414 35030 5466
rect 35030 5414 35076 5466
rect 35100 5414 35146 5466
rect 35146 5414 35156 5466
rect 35180 5414 35210 5466
rect 35210 5414 35236 5466
rect 34940 5412 34996 5414
rect 35020 5412 35076 5414
rect 35100 5412 35156 5414
rect 35180 5412 35236 5414
rect 35530 5616 35586 5672
rect 32954 4120 33010 4176
rect 33966 4528 34022 4584
rect 32678 3984 32734 4040
rect 32034 3848 32090 3904
rect 31942 3596 31998 3632
rect 31942 3576 31944 3596
rect 31944 3576 31996 3596
rect 31996 3576 31998 3596
rect 33046 3712 33102 3768
rect 32126 3304 32182 3360
rect 32678 3168 32734 3224
rect 31114 2760 31170 2816
rect 33046 2760 33102 2816
rect 34518 3732 34574 3768
rect 34518 3712 34520 3732
rect 34520 3712 34572 3732
rect 34572 3712 34574 3732
rect 34940 4378 34996 4380
rect 35020 4378 35076 4380
rect 35100 4378 35156 4380
rect 35180 4378 35236 4380
rect 34940 4326 34966 4378
rect 34966 4326 34996 4378
rect 35020 4326 35030 4378
rect 35030 4326 35076 4378
rect 35100 4326 35146 4378
rect 35146 4326 35156 4378
rect 35180 4326 35210 4378
rect 35210 4326 35236 4378
rect 34940 4324 34996 4326
rect 35020 4324 35076 4326
rect 35100 4324 35156 4326
rect 35180 4324 35236 4326
rect 34940 3290 34996 3292
rect 35020 3290 35076 3292
rect 35100 3290 35156 3292
rect 35180 3290 35236 3292
rect 34940 3238 34966 3290
rect 34966 3238 34996 3290
rect 35020 3238 35030 3290
rect 35030 3238 35076 3290
rect 35100 3238 35146 3290
rect 35146 3238 35156 3290
rect 35180 3238 35210 3290
rect 35210 3238 35236 3290
rect 34940 3236 34996 3238
rect 35020 3236 35076 3238
rect 35100 3236 35156 3238
rect 35180 3236 35236 3238
rect 34940 2202 34996 2204
rect 35020 2202 35076 2204
rect 35100 2202 35156 2204
rect 35180 2202 35236 2204
rect 34940 2150 34966 2202
rect 34966 2150 34996 2202
rect 35020 2150 35030 2202
rect 35030 2150 35076 2202
rect 35100 2150 35146 2202
rect 35146 2150 35156 2202
rect 35180 2150 35210 2202
rect 35210 2150 35236 2202
rect 34940 2148 34996 2150
rect 35020 2148 35076 2150
rect 35100 2148 35156 2150
rect 35180 2148 35236 2150
rect 41142 18536 41198 18592
rect 46110 25200 46166 25256
rect 47398 44532 47454 44568
rect 47398 44512 47400 44532
rect 47400 44512 47452 44532
rect 47452 44512 47454 44532
rect 46938 42880 46994 42936
rect 46754 41384 46810 41440
rect 46938 39752 46994 39808
rect 46754 38256 46810 38312
rect 46938 36624 46994 36680
rect 46754 35148 46810 35184
rect 46754 35128 46756 35148
rect 46756 35128 46808 35148
rect 46808 35128 46810 35148
rect 46754 32000 46810 32056
rect 46662 27104 46718 27160
rect 46938 33496 46994 33552
rect 47214 30660 47270 30696
rect 47214 30640 47216 30660
rect 47216 30640 47268 30660
rect 47268 30640 47270 30660
rect 46938 30368 46994 30424
rect 47306 28872 47362 28928
rect 46938 27240 46994 27296
rect 45926 20576 45982 20632
rect 42890 18572 42892 18592
rect 42892 18572 42944 18592
rect 42944 18572 42946 18592
rect 42890 18536 42946 18572
rect 42614 17332 42670 17368
rect 42614 17312 42616 17332
rect 42616 17312 42668 17332
rect 42668 17312 42670 17332
rect 42246 15816 42302 15872
rect 40958 10240 41014 10296
rect 37738 9716 37794 9752
rect 37738 9696 37740 9716
rect 37740 9696 37792 9716
rect 37792 9696 37794 9716
rect 42338 15308 42340 15328
rect 42340 15308 42392 15328
rect 42392 15308 42394 15328
rect 42338 15272 42394 15308
rect 47030 26696 47086 26752
rect 47214 26288 47270 26344
rect 46754 23024 46810 23080
rect 47306 25744 47362 25800
rect 47306 22652 47308 22672
rect 47308 22652 47360 22672
rect 47360 22652 47362 22672
rect 47306 22616 47362 22652
rect 46754 21004 46810 21040
rect 46754 20984 46756 21004
rect 46756 20984 46808 21004
rect 46808 20984 46810 21004
rect 47490 21956 47546 21992
rect 47490 21936 47492 21956
rect 47492 21936 47544 21956
rect 47544 21936 47546 21956
rect 47306 19508 47362 19544
rect 47306 19488 47308 19508
rect 47308 19488 47360 19508
rect 47360 19488 47362 19508
rect 46478 19216 46534 19272
rect 44362 18420 44418 18456
rect 44362 18400 44364 18420
rect 44364 18400 44416 18420
rect 44416 18400 44418 18420
rect 43718 15816 43774 15872
rect 47490 18400 47546 18456
rect 46754 17856 46810 17912
rect 47122 17312 47178 17368
rect 44270 15852 44272 15872
rect 44272 15852 44324 15872
rect 44324 15852 44326 15872
rect 44270 15816 44326 15852
rect 43994 15136 44050 15192
rect 46846 16360 46902 16416
rect 46570 15272 46626 15328
rect 46938 15136 46994 15192
rect 42706 11636 42708 11656
rect 42708 11636 42760 11656
rect 42760 11636 42762 11656
rect 42706 11600 42762 11636
rect 47214 14728 47270 14784
rect 47490 13232 47546 13288
rect 43074 10260 43130 10296
rect 43074 10240 43076 10260
rect 43076 10240 43128 10260
rect 43128 10240 43130 10260
rect 42062 10140 42064 10160
rect 42064 10140 42116 10160
rect 42116 10140 42118 10160
rect 42062 10104 42118 10140
rect 39210 8472 39266 8528
rect 39302 6196 39304 6216
rect 39304 6196 39356 6216
rect 39356 6196 39358 6216
rect 39302 6160 39358 6196
rect 38290 6024 38346 6080
rect 38106 5616 38162 5672
rect 37370 4548 37426 4584
rect 37370 4528 37372 4548
rect 37372 4528 37424 4548
rect 37424 4528 37426 4548
rect 37094 4256 37150 4312
rect 38290 4700 38292 4720
rect 38292 4700 38344 4720
rect 38344 4700 38346 4720
rect 38290 4664 38346 4700
rect 43626 10376 43682 10432
rect 46938 10376 46994 10432
rect 46938 10104 46994 10160
rect 47398 10104 47454 10160
rect 43626 8492 43682 8528
rect 43626 8472 43628 8492
rect 43628 8472 43680 8492
rect 43680 8472 43682 8492
rect 46938 8508 46940 8528
rect 46940 8508 46992 8528
rect 46992 8508 46994 8528
rect 46938 8472 46994 8508
rect 47398 8492 47454 8528
rect 47398 8472 47400 8492
rect 47400 8472 47452 8492
rect 47452 8472 47454 8492
rect 44362 6976 44418 7032
rect 45098 6976 45154 7032
rect 46938 6976 46994 7032
rect 47398 6976 47454 7032
rect 42062 6024 42118 6080
rect 45926 6060 45928 6080
rect 45928 6060 45980 6080
rect 45980 6060 45982 6080
rect 45926 6024 45982 6060
rect 49238 6024 49294 6080
rect 40038 4664 40094 4720
rect 40498 4256 40554 4312
rect 38198 3848 38254 3904
rect 36266 3068 36268 3088
rect 36268 3068 36320 3088
rect 36320 3068 36322 3088
rect 36266 3032 36322 3068
rect 36634 2896 36690 2952
rect 37830 2760 37886 2816
rect 36174 1400 36230 1456
rect 41050 3884 41052 3904
rect 41052 3884 41104 3904
rect 41104 3884 41106 3904
rect 41050 3848 41106 3884
rect 41418 3848 41474 3904
rect 41418 3576 41474 3632
rect 47858 3576 47914 3632
rect 42706 2760 42762 2816
rect 36082 40 36138 96
<< metal3 >>
rect 46933 49194 46999 49197
rect 49520 49194 50000 49224
rect 46933 49192 50000 49194
rect 46933 49136 46938 49192
rect 46994 49136 50000 49192
rect 46933 49134 50000 49136
rect 46933 49131 46999 49134
rect 49520 49104 50000 49134
rect 46749 47698 46815 47701
rect 49520 47698 50000 47728
rect 46749 47696 50000 47698
rect 46749 47640 46754 47696
rect 46810 47640 50000 47696
rect 46749 47638 50000 47640
rect 46749 47635 46815 47638
rect 49520 47608 50000 47638
rect 19568 47360 19888 47361
rect 19568 47296 19576 47360
rect 19640 47296 19656 47360
rect 19720 47296 19736 47360
rect 19800 47296 19816 47360
rect 19880 47296 19888 47360
rect 19568 47295 19888 47296
rect 4208 46816 4528 46817
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 46751 4528 46752
rect 34928 46816 35248 46817
rect 34928 46752 34936 46816
rect 35000 46752 35016 46816
rect 35080 46752 35096 46816
rect 35160 46752 35176 46816
rect 35240 46752 35248 46816
rect 34928 46751 35248 46752
rect 19568 46272 19888 46273
rect 19568 46208 19576 46272
rect 19640 46208 19656 46272
rect 19720 46208 19736 46272
rect 19800 46208 19816 46272
rect 19880 46208 19888 46272
rect 19568 46207 19888 46208
rect 46841 46066 46907 46069
rect 49520 46066 50000 46096
rect 46841 46064 50000 46066
rect 46841 46008 46846 46064
rect 46902 46008 50000 46064
rect 46841 46006 50000 46008
rect 46841 46003 46907 46006
rect 49520 45976 50000 46006
rect 4208 45728 4528 45729
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 45663 4528 45664
rect 34928 45728 35248 45729
rect 34928 45664 34936 45728
rect 35000 45664 35016 45728
rect 35080 45664 35096 45728
rect 35160 45664 35176 45728
rect 35240 45664 35248 45728
rect 34928 45663 35248 45664
rect 24945 45658 25011 45661
rect 28073 45658 28139 45661
rect 24945 45656 28139 45658
rect 24945 45600 24950 45656
rect 25006 45600 28078 45656
rect 28134 45600 28139 45656
rect 24945 45598 28139 45600
rect 24945 45595 25011 45598
rect 28073 45595 28139 45598
rect 19568 45184 19888 45185
rect 19568 45120 19576 45184
rect 19640 45120 19656 45184
rect 19720 45120 19736 45184
rect 19800 45120 19816 45184
rect 19880 45120 19888 45184
rect 19568 45119 19888 45120
rect 4208 44640 4528 44641
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 44575 4528 44576
rect 34928 44640 35248 44641
rect 34928 44576 34936 44640
rect 35000 44576 35016 44640
rect 35080 44576 35096 44640
rect 35160 44576 35176 44640
rect 35240 44576 35248 44640
rect 34928 44575 35248 44576
rect 47393 44570 47459 44573
rect 49520 44570 50000 44600
rect 47393 44568 50000 44570
rect 47393 44512 47398 44568
rect 47454 44512 50000 44568
rect 47393 44510 50000 44512
rect 47393 44507 47459 44510
rect 49520 44480 50000 44510
rect 19568 44096 19888 44097
rect 19568 44032 19576 44096
rect 19640 44032 19656 44096
rect 19720 44032 19736 44096
rect 19800 44032 19816 44096
rect 19880 44032 19888 44096
rect 19568 44031 19888 44032
rect 4208 43552 4528 43553
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 43487 4528 43488
rect 34928 43552 35248 43553
rect 34928 43488 34936 43552
rect 35000 43488 35016 43552
rect 35080 43488 35096 43552
rect 35160 43488 35176 43552
rect 35240 43488 35248 43552
rect 34928 43487 35248 43488
rect 19568 43008 19888 43009
rect 19568 42944 19576 43008
rect 19640 42944 19656 43008
rect 19720 42944 19736 43008
rect 19800 42944 19816 43008
rect 19880 42944 19888 43008
rect 19568 42943 19888 42944
rect 46933 42938 46999 42941
rect 49520 42938 50000 42968
rect 46933 42936 50000 42938
rect 46933 42880 46938 42936
rect 46994 42880 50000 42936
rect 46933 42878 50000 42880
rect 46933 42875 46999 42878
rect 49520 42848 50000 42878
rect 4208 42464 4528 42465
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 42399 4528 42400
rect 34928 42464 35248 42465
rect 34928 42400 34936 42464
rect 35000 42400 35016 42464
rect 35080 42400 35096 42464
rect 35160 42400 35176 42464
rect 35240 42400 35248 42464
rect 34928 42399 35248 42400
rect 19568 41920 19888 41921
rect 19568 41856 19576 41920
rect 19640 41856 19656 41920
rect 19720 41856 19736 41920
rect 19800 41856 19816 41920
rect 19880 41856 19888 41920
rect 19568 41855 19888 41856
rect 46749 41442 46815 41445
rect 49520 41442 50000 41472
rect 46749 41440 50000 41442
rect 46749 41384 46754 41440
rect 46810 41384 50000 41440
rect 46749 41382 50000 41384
rect 46749 41379 46815 41382
rect 4208 41376 4528 41377
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 41311 4528 41312
rect 34928 41376 35248 41377
rect 34928 41312 34936 41376
rect 35000 41312 35016 41376
rect 35080 41312 35096 41376
rect 35160 41312 35176 41376
rect 35240 41312 35248 41376
rect 49520 41352 50000 41382
rect 34928 41311 35248 41312
rect 19568 40832 19888 40833
rect 19568 40768 19576 40832
rect 19640 40768 19656 40832
rect 19720 40768 19736 40832
rect 19800 40768 19816 40832
rect 19880 40768 19888 40832
rect 19568 40767 19888 40768
rect 4208 40288 4528 40289
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 40223 4528 40224
rect 34928 40288 35248 40289
rect 34928 40224 34936 40288
rect 35000 40224 35016 40288
rect 35080 40224 35096 40288
rect 35160 40224 35176 40288
rect 35240 40224 35248 40288
rect 34928 40223 35248 40224
rect 46933 39810 46999 39813
rect 49520 39810 50000 39840
rect 46933 39808 50000 39810
rect 46933 39752 46938 39808
rect 46994 39752 50000 39808
rect 46933 39750 50000 39752
rect 46933 39747 46999 39750
rect 19568 39744 19888 39745
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 49520 39720 50000 39750
rect 19568 39679 19888 39680
rect 4208 39200 4528 39201
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 39135 4528 39136
rect 34928 39200 35248 39201
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 39135 35248 39136
rect 19568 38656 19888 38657
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 38591 19888 38592
rect 46749 38314 46815 38317
rect 49520 38314 50000 38344
rect 46749 38312 50000 38314
rect 46749 38256 46754 38312
rect 46810 38256 50000 38312
rect 46749 38254 50000 38256
rect 46749 38251 46815 38254
rect 49520 38224 50000 38254
rect 4208 38112 4528 38113
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 38047 4528 38048
rect 34928 38112 35248 38113
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 38047 35248 38048
rect 0 37634 480 37664
rect 3417 37634 3483 37637
rect 0 37632 3483 37634
rect 0 37576 3422 37632
rect 3478 37576 3483 37632
rect 0 37574 3483 37576
rect 0 37544 480 37574
rect 3417 37571 3483 37574
rect 19568 37568 19888 37569
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 37503 19888 37504
rect 4208 37024 4528 37025
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 34928 37024 35248 37025
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 36959 35248 36960
rect 46933 36682 46999 36685
rect 49520 36682 50000 36712
rect 46933 36680 50000 36682
rect 46933 36624 46938 36680
rect 46994 36624 50000 36680
rect 46933 36622 50000 36624
rect 46933 36619 46999 36622
rect 49520 36592 50000 36622
rect 19568 36480 19888 36481
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 36415 19888 36416
rect 4208 35936 4528 35937
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 34928 35936 35248 35937
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 35871 35248 35872
rect 19568 35392 19888 35393
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 35327 19888 35328
rect 46749 35186 46815 35189
rect 49520 35186 50000 35216
rect 46749 35184 50000 35186
rect 46749 35128 46754 35184
rect 46810 35128 50000 35184
rect 46749 35126 50000 35128
rect 46749 35123 46815 35126
rect 49520 35096 50000 35126
rect 4208 34848 4528 34849
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 34928 34848 35248 34849
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 34783 35248 34784
rect 19568 34304 19888 34305
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 34239 19888 34240
rect 4208 33760 4528 33761
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 34928 33760 35248 33761
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 33695 35248 33696
rect 46933 33554 46999 33557
rect 49520 33554 50000 33584
rect 46933 33552 50000 33554
rect 46933 33496 46938 33552
rect 46994 33496 50000 33552
rect 46933 33494 50000 33496
rect 46933 33491 46999 33494
rect 49520 33464 50000 33494
rect 19568 33216 19888 33217
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 33151 19888 33152
rect 4208 32672 4528 32673
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 34928 32672 35248 32673
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 32607 35248 32608
rect 19568 32128 19888 32129
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 32063 19888 32064
rect 46749 32058 46815 32061
rect 49520 32058 50000 32088
rect 46749 32056 50000 32058
rect 46749 32000 46754 32056
rect 46810 32000 50000 32056
rect 46749 31998 50000 32000
rect 46749 31995 46815 31998
rect 49520 31968 50000 31998
rect 4208 31584 4528 31585
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 34928 31584 35248 31585
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 31519 35248 31520
rect 19568 31040 19888 31041
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 30975 19888 30976
rect 43621 30698 43687 30701
rect 47209 30698 47275 30701
rect 43621 30696 47275 30698
rect 43621 30640 43626 30696
rect 43682 30640 47214 30696
rect 47270 30640 47275 30696
rect 43621 30638 47275 30640
rect 43621 30635 43687 30638
rect 47209 30635 47275 30638
rect 4208 30496 4528 30497
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 34928 30496 35248 30497
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 30431 35248 30432
rect 46933 30426 46999 30429
rect 49520 30426 50000 30456
rect 46933 30424 50000 30426
rect 46933 30368 46938 30424
rect 46994 30368 50000 30424
rect 46933 30366 50000 30368
rect 46933 30363 46999 30366
rect 49520 30336 50000 30366
rect 19568 29952 19888 29953
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 29887 19888 29888
rect 4208 29408 4528 29409
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 34928 29408 35248 29409
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 29343 35248 29344
rect 39573 29338 39639 29341
rect 42425 29338 42491 29341
rect 39573 29336 42491 29338
rect 39573 29280 39578 29336
rect 39634 29280 42430 29336
rect 42486 29280 42491 29336
rect 39573 29278 42491 29280
rect 39573 29275 39639 29278
rect 42425 29275 42491 29278
rect 41229 28930 41295 28933
rect 42057 28930 42123 28933
rect 41229 28928 42123 28930
rect 41229 28872 41234 28928
rect 41290 28872 42062 28928
rect 42118 28872 42123 28928
rect 41229 28870 42123 28872
rect 41229 28867 41295 28870
rect 42057 28867 42123 28870
rect 47301 28930 47367 28933
rect 49520 28930 50000 28960
rect 47301 28928 50000 28930
rect 47301 28872 47306 28928
rect 47362 28872 50000 28928
rect 47301 28870 50000 28872
rect 47301 28867 47367 28870
rect 19568 28864 19888 28865
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 49520 28840 50000 28870
rect 19568 28799 19888 28800
rect 4208 28320 4528 28321
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 34928 28320 35248 28321
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 28255 35248 28256
rect 41689 27978 41755 27981
rect 44541 27978 44607 27981
rect 41689 27976 44607 27978
rect 41689 27920 41694 27976
rect 41750 27920 44546 27976
rect 44602 27920 44607 27976
rect 41689 27918 44607 27920
rect 41689 27915 41755 27918
rect 44541 27915 44607 27918
rect 19568 27776 19888 27777
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 27711 19888 27712
rect 42241 27434 42307 27437
rect 45185 27434 45251 27437
rect 42241 27432 45251 27434
rect 42241 27376 42246 27432
rect 42302 27376 45190 27432
rect 45246 27376 45251 27432
rect 42241 27374 45251 27376
rect 42241 27371 42307 27374
rect 45185 27371 45251 27374
rect 46933 27298 46999 27301
rect 49520 27298 50000 27328
rect 46933 27296 50000 27298
rect 46933 27240 46938 27296
rect 46994 27240 50000 27296
rect 46933 27238 50000 27240
rect 46933 27235 46999 27238
rect 4208 27232 4528 27233
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 34928 27232 35248 27233
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 49520 27208 50000 27238
rect 34928 27167 35248 27168
rect 38377 27162 38443 27165
rect 46657 27162 46723 27165
rect 38377 27160 46723 27162
rect 38377 27104 38382 27160
rect 38438 27104 46662 27160
rect 46718 27104 46723 27160
rect 38377 27102 46723 27104
rect 38377 27099 38443 27102
rect 46657 27099 46723 27102
rect 45277 26754 45343 26757
rect 47025 26754 47091 26757
rect 45277 26752 47091 26754
rect 45277 26696 45282 26752
rect 45338 26696 47030 26752
rect 47086 26696 47091 26752
rect 45277 26694 47091 26696
rect 45277 26691 45343 26694
rect 47025 26691 47091 26694
rect 19568 26688 19888 26689
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 26623 19888 26624
rect 45185 26346 45251 26349
rect 47209 26346 47275 26349
rect 45185 26344 47275 26346
rect 45185 26288 45190 26344
rect 45246 26288 47214 26344
rect 47270 26288 47275 26344
rect 45185 26286 47275 26288
rect 45185 26283 45251 26286
rect 47209 26283 47275 26286
rect 4208 26144 4528 26145
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect 34928 26144 35248 26145
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 26079 35248 26080
rect 47301 25802 47367 25805
rect 49520 25802 50000 25832
rect 47301 25800 50000 25802
rect 47301 25744 47306 25800
rect 47362 25744 50000 25800
rect 47301 25742 50000 25744
rect 47301 25739 47367 25742
rect 49520 25712 50000 25742
rect 38193 25666 38259 25669
rect 40585 25666 40651 25669
rect 38193 25664 40651 25666
rect 38193 25608 38198 25664
rect 38254 25608 40590 25664
rect 40646 25608 40651 25664
rect 38193 25606 40651 25608
rect 38193 25603 38259 25606
rect 40585 25603 40651 25606
rect 19568 25600 19888 25601
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 25535 19888 25536
rect 39573 25530 39639 25533
rect 41965 25530 42031 25533
rect 39573 25528 42031 25530
rect 39573 25472 39578 25528
rect 39634 25472 41970 25528
rect 42026 25472 42031 25528
rect 39573 25470 42031 25472
rect 39573 25467 39639 25470
rect 41965 25467 42031 25470
rect 35985 25258 36051 25261
rect 46105 25258 46171 25261
rect 35985 25256 46171 25258
rect 35985 25200 35990 25256
rect 36046 25200 46110 25256
rect 46166 25200 46171 25256
rect 35985 25198 46171 25200
rect 35985 25195 36051 25198
rect 46105 25195 46171 25198
rect 4208 25056 4528 25057
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 34928 25056 35248 25057
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 24991 35248 24992
rect 41045 24850 41111 24853
rect 45645 24850 45711 24853
rect 41045 24848 45711 24850
rect 41045 24792 41050 24848
rect 41106 24792 45650 24848
rect 45706 24792 45711 24848
rect 41045 24790 45711 24792
rect 41045 24787 41111 24790
rect 45645 24787 45711 24790
rect 38653 24714 38719 24717
rect 42333 24714 42399 24717
rect 38653 24712 42399 24714
rect 38653 24656 38658 24712
rect 38714 24656 42338 24712
rect 42394 24656 42399 24712
rect 38653 24654 42399 24656
rect 38653 24651 38719 24654
rect 42333 24651 42399 24654
rect 19568 24512 19888 24513
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 24447 19888 24448
rect 31293 24170 31359 24173
rect 40309 24170 40375 24173
rect 31293 24168 40375 24170
rect 31293 24112 31298 24168
rect 31354 24112 40314 24168
rect 40370 24112 40375 24168
rect 31293 24110 40375 24112
rect 31293 24107 31359 24110
rect 40309 24107 40375 24110
rect 43437 24170 43503 24173
rect 49520 24170 50000 24200
rect 43437 24168 50000 24170
rect 43437 24112 43442 24168
rect 43498 24112 50000 24168
rect 43437 24110 50000 24112
rect 43437 24107 43503 24110
rect 49520 24080 50000 24110
rect 4208 23968 4528 23969
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 34928 23968 35248 23969
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 23903 35248 23904
rect 19568 23424 19888 23425
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 23359 19888 23360
rect 33593 23082 33659 23085
rect 46749 23082 46815 23085
rect 33593 23080 46815 23082
rect 33593 23024 33598 23080
rect 33654 23024 46754 23080
rect 46810 23024 46815 23080
rect 33593 23022 46815 23024
rect 33593 23019 33659 23022
rect 46749 23019 46815 23022
rect 36169 22946 36235 22949
rect 36629 22946 36695 22949
rect 40493 22946 40559 22949
rect 36169 22944 40559 22946
rect 36169 22888 36174 22944
rect 36230 22888 36634 22944
rect 36690 22888 40498 22944
rect 40554 22888 40559 22944
rect 36169 22886 40559 22888
rect 36169 22883 36235 22886
rect 36629 22883 36695 22886
rect 40493 22883 40559 22886
rect 4208 22880 4528 22881
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect 34928 22880 35248 22881
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 22815 35248 22816
rect 47301 22674 47367 22677
rect 49520 22674 50000 22704
rect 47301 22672 50000 22674
rect 47301 22616 47306 22672
rect 47362 22616 50000 22672
rect 47301 22614 50000 22616
rect 47301 22611 47367 22614
rect 49520 22584 50000 22614
rect 19568 22336 19888 22337
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 22271 19888 22272
rect 30281 21994 30347 21997
rect 34605 21994 34671 21997
rect 30281 21992 34671 21994
rect 30281 21936 30286 21992
rect 30342 21936 34610 21992
rect 34666 21936 34671 21992
rect 30281 21934 34671 21936
rect 30281 21931 30347 21934
rect 34605 21931 34671 21934
rect 41597 21994 41663 21997
rect 47485 21994 47551 21997
rect 41597 21992 47551 21994
rect 41597 21936 41602 21992
rect 41658 21936 47490 21992
rect 47546 21936 47551 21992
rect 41597 21934 47551 21936
rect 41597 21931 41663 21934
rect 47485 21931 47551 21934
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 34928 21792 35248 21793
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 21727 35248 21728
rect 8293 21450 8359 21453
rect 29637 21450 29703 21453
rect 8293 21448 29703 21450
rect 8293 21392 8298 21448
rect 8354 21392 29642 21448
rect 29698 21392 29703 21448
rect 8293 21390 29703 21392
rect 8293 21387 8359 21390
rect 29637 21387 29703 21390
rect 19568 21248 19888 21249
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 21183 19888 21184
rect 46749 21042 46815 21045
rect 49520 21042 50000 21072
rect 46749 21040 50000 21042
rect 46749 20984 46754 21040
rect 46810 20984 50000 21040
rect 46749 20982 50000 20984
rect 46749 20979 46815 20982
rect 49520 20952 50000 20982
rect 28257 20770 28323 20773
rect 31017 20770 31083 20773
rect 38193 20770 38259 20773
rect 40769 20770 40835 20773
rect 28257 20768 31083 20770
rect 28257 20712 28262 20768
rect 28318 20712 31022 20768
rect 31078 20712 31083 20768
rect 28257 20710 31083 20712
rect 28257 20707 28323 20710
rect 31017 20707 31083 20710
rect 38150 20768 40835 20770
rect 38150 20712 38198 20768
rect 38254 20712 40774 20768
rect 40830 20712 40835 20768
rect 38150 20710 40835 20712
rect 38150 20707 38259 20710
rect 40769 20707 40835 20710
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 34928 20704 35248 20705
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 20639 35248 20640
rect 27613 20634 27679 20637
rect 32397 20634 32463 20637
rect 27613 20632 32463 20634
rect 27613 20576 27618 20632
rect 27674 20576 32402 20632
rect 32458 20576 32463 20632
rect 27613 20574 32463 20576
rect 27613 20571 27679 20574
rect 32397 20571 32463 20574
rect 35617 20634 35683 20637
rect 38150 20634 38210 20707
rect 35617 20632 38210 20634
rect 35617 20576 35622 20632
rect 35678 20576 38210 20632
rect 35617 20574 38210 20576
rect 40585 20634 40651 20637
rect 45921 20634 45987 20637
rect 40585 20632 45987 20634
rect 40585 20576 40590 20632
rect 40646 20576 45926 20632
rect 45982 20576 45987 20632
rect 40585 20574 45987 20576
rect 35617 20571 35683 20574
rect 40585 20571 40651 20574
rect 45921 20571 45987 20574
rect 19568 20160 19888 20161
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 20095 19888 20096
rect 32765 20090 32831 20093
rect 34789 20090 34855 20093
rect 38285 20090 38351 20093
rect 32765 20088 38351 20090
rect 32765 20032 32770 20088
rect 32826 20032 34794 20088
rect 34850 20032 38290 20088
rect 38346 20032 38351 20088
rect 32765 20030 38351 20032
rect 32765 20027 32831 20030
rect 34789 20027 34855 20030
rect 38285 20027 38351 20030
rect 34973 19954 35039 19957
rect 39849 19954 39915 19957
rect 34973 19952 39915 19954
rect 34973 19896 34978 19952
rect 35034 19896 39854 19952
rect 39910 19896 39915 19952
rect 34973 19894 39915 19896
rect 34973 19891 35039 19894
rect 39849 19891 39915 19894
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 34928 19616 35248 19617
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 19551 35248 19552
rect 47301 19546 47367 19549
rect 49520 19546 50000 19576
rect 47301 19544 50000 19546
rect 47301 19488 47306 19544
rect 47362 19488 50000 19544
rect 47301 19486 50000 19488
rect 47301 19483 47367 19486
rect 49520 19456 50000 19486
rect 32397 19410 32463 19413
rect 34697 19410 34763 19413
rect 32397 19408 34763 19410
rect 32397 19352 32402 19408
rect 32458 19352 34702 19408
rect 34758 19352 34763 19408
rect 32397 19350 34763 19352
rect 32397 19347 32463 19350
rect 34697 19347 34763 19350
rect 38561 19274 38627 19277
rect 46473 19274 46539 19277
rect 38561 19272 46539 19274
rect 38561 19216 38566 19272
rect 38622 19216 46478 19272
rect 46534 19216 46539 19272
rect 38561 19214 46539 19216
rect 38561 19211 38627 19214
rect 46473 19211 46539 19214
rect 19568 19072 19888 19073
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 19007 19888 19008
rect 35617 18866 35683 18869
rect 38101 18866 38167 18869
rect 35617 18864 38167 18866
rect 35617 18808 35622 18864
rect 35678 18808 38106 18864
rect 38162 18808 38167 18864
rect 35617 18806 38167 18808
rect 35617 18803 35683 18806
rect 38101 18803 38167 18806
rect 41137 18594 41203 18597
rect 42885 18594 42951 18597
rect 41137 18592 42951 18594
rect 41137 18536 41142 18592
rect 41198 18536 42890 18592
rect 42946 18536 42951 18592
rect 41137 18534 42951 18536
rect 41137 18531 41203 18534
rect 42885 18531 42951 18534
rect 4208 18528 4528 18529
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 34928 18528 35248 18529
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 18463 35248 18464
rect 44357 18458 44423 18461
rect 47485 18458 47551 18461
rect 44357 18456 47551 18458
rect 44357 18400 44362 18456
rect 44418 18400 47490 18456
rect 47546 18400 47551 18456
rect 44357 18398 47551 18400
rect 44357 18395 44423 18398
rect 47485 18395 47551 18398
rect 19568 17984 19888 17985
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 17919 19888 17920
rect 46749 17914 46815 17917
rect 49520 17914 50000 17944
rect 46749 17912 50000 17914
rect 46749 17856 46754 17912
rect 46810 17856 50000 17912
rect 46749 17854 50000 17856
rect 46749 17851 46815 17854
rect 49520 17824 50000 17854
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 34928 17440 35248 17441
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 17375 35248 17376
rect 42609 17370 42675 17373
rect 47117 17370 47183 17373
rect 42609 17368 47183 17370
rect 42609 17312 42614 17368
rect 42670 17312 47122 17368
rect 47178 17312 47183 17368
rect 42609 17310 47183 17312
rect 42609 17307 42675 17310
rect 47117 17307 47183 17310
rect 35525 17234 35591 17237
rect 37273 17234 37339 17237
rect 35525 17232 37339 17234
rect 35525 17176 35530 17232
rect 35586 17176 37278 17232
rect 37334 17176 37339 17232
rect 35525 17174 37339 17176
rect 35525 17171 35591 17174
rect 37273 17171 37339 17174
rect 3417 17098 3483 17101
rect 23473 17098 23539 17101
rect 3417 17096 23539 17098
rect 3417 17040 3422 17096
rect 3478 17040 23478 17096
rect 23534 17040 23539 17096
rect 3417 17038 23539 17040
rect 3417 17035 3483 17038
rect 23473 17035 23539 17038
rect 19568 16896 19888 16897
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 16831 19888 16832
rect 26509 16826 26575 16829
rect 29913 16826 29979 16829
rect 30373 16826 30439 16829
rect 26509 16824 30439 16826
rect 26509 16768 26514 16824
rect 26570 16768 29918 16824
rect 29974 16768 30378 16824
rect 30434 16768 30439 16824
rect 26509 16766 30439 16768
rect 26509 16763 26575 16766
rect 29913 16763 29979 16766
rect 30373 16763 30439 16766
rect 46841 16418 46907 16421
rect 49520 16418 50000 16448
rect 46841 16416 50000 16418
rect 46841 16360 46846 16416
rect 46902 16360 50000 16416
rect 46841 16358 50000 16360
rect 46841 16355 46907 16358
rect 4208 16352 4528 16353
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 34928 16352 35248 16353
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 49520 16328 50000 16358
rect 34928 16287 35248 16288
rect 42241 15874 42307 15877
rect 43713 15874 43779 15877
rect 44265 15874 44331 15877
rect 42241 15872 44331 15874
rect 42241 15816 42246 15872
rect 42302 15816 43718 15872
rect 43774 15816 44270 15872
rect 44326 15816 44331 15872
rect 42241 15814 44331 15816
rect 42241 15811 42307 15814
rect 43713 15811 43779 15814
rect 44265 15811 44331 15814
rect 19568 15808 19888 15809
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 15743 19888 15744
rect 42333 15330 42399 15333
rect 46565 15330 46631 15333
rect 42333 15328 46631 15330
rect 42333 15272 42338 15328
rect 42394 15272 46570 15328
rect 46626 15272 46631 15328
rect 42333 15270 46631 15272
rect 42333 15267 42399 15270
rect 46565 15267 46631 15270
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 34928 15264 35248 15265
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 15199 35248 15200
rect 43989 15194 44055 15197
rect 46933 15194 46999 15197
rect 43989 15192 46999 15194
rect 43989 15136 43994 15192
rect 44050 15136 46938 15192
rect 46994 15136 46999 15192
rect 43989 15134 46999 15136
rect 43989 15131 44055 15134
rect 46933 15131 46999 15134
rect 47209 14786 47275 14789
rect 49520 14786 50000 14816
rect 47209 14784 50000 14786
rect 47209 14728 47214 14784
rect 47270 14728 50000 14784
rect 47209 14726 50000 14728
rect 47209 14723 47275 14726
rect 19568 14720 19888 14721
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 49520 14696 50000 14726
rect 19568 14655 19888 14656
rect 20253 14514 20319 14517
rect 36169 14514 36235 14517
rect 20253 14512 36235 14514
rect 20253 14456 20258 14512
rect 20314 14456 36174 14512
rect 36230 14456 36235 14512
rect 20253 14454 36235 14456
rect 20253 14451 20319 14454
rect 36169 14451 36235 14454
rect 8385 14378 8451 14381
rect 36629 14378 36695 14381
rect 8385 14376 36695 14378
rect 8385 14320 8390 14376
rect 8446 14320 36634 14376
rect 36690 14320 36695 14376
rect 8385 14318 36695 14320
rect 8385 14315 8451 14318
rect 36629 14315 36695 14318
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 34928 14176 35248 14177
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 14111 35248 14112
rect 30281 13834 30347 13837
rect 31753 13834 31819 13837
rect 30281 13832 31819 13834
rect 30281 13776 30286 13832
rect 30342 13776 31758 13832
rect 31814 13776 31819 13832
rect 30281 13774 31819 13776
rect 30281 13771 30347 13774
rect 31753 13771 31819 13774
rect 35157 13834 35223 13837
rect 35709 13834 35775 13837
rect 35157 13832 35775 13834
rect 35157 13776 35162 13832
rect 35218 13776 35714 13832
rect 35770 13776 35775 13832
rect 35157 13774 35775 13776
rect 35157 13771 35223 13774
rect 35709 13771 35775 13774
rect 19568 13632 19888 13633
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 13567 19888 13568
rect 47485 13290 47551 13293
rect 49520 13290 50000 13320
rect 47485 13288 50000 13290
rect 47485 13232 47490 13288
rect 47546 13232 50000 13288
rect 47485 13230 50000 13232
rect 47485 13227 47551 13230
rect 49520 13200 50000 13230
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 34928 13088 35248 13089
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 13023 35248 13024
rect 20437 12882 20503 12885
rect 20989 12882 21055 12885
rect 27521 12882 27587 12885
rect 20437 12880 27587 12882
rect 20437 12824 20442 12880
rect 20498 12824 20994 12880
rect 21050 12824 27526 12880
rect 27582 12824 27587 12880
rect 20437 12822 27587 12824
rect 20437 12819 20503 12822
rect 20989 12819 21055 12822
rect 27521 12819 27587 12822
rect 7005 12746 7071 12749
rect 8293 12746 8359 12749
rect 7005 12744 8359 12746
rect 7005 12688 7010 12744
rect 7066 12688 8298 12744
rect 8354 12688 8359 12744
rect 7005 12686 8359 12688
rect 7005 12683 7071 12686
rect 8293 12683 8359 12686
rect 0 12520 480 12640
rect 31017 12612 31083 12613
rect 30966 12548 30972 12612
rect 31036 12610 31083 12612
rect 31036 12608 31128 12610
rect 31078 12552 31128 12608
rect 31036 12550 31128 12552
rect 31036 12548 31083 12550
rect 31017 12547 31083 12548
rect 19568 12544 19888 12545
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 12479 19888 12480
rect 9949 12338 10015 12341
rect 18873 12338 18939 12341
rect 22277 12338 22343 12341
rect 9949 12336 22343 12338
rect 9949 12280 9954 12336
rect 10010 12280 18878 12336
rect 18934 12280 22282 12336
rect 22338 12280 22343 12336
rect 9949 12278 22343 12280
rect 9949 12275 10015 12278
rect 18873 12275 18939 12278
rect 22277 12275 22343 12278
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 34928 12000 35248 12001
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 11935 35248 11936
rect 21357 11930 21423 11933
rect 25037 11930 25103 11933
rect 21357 11928 25103 11930
rect 21357 11872 21362 11928
rect 21418 11872 25042 11928
rect 25098 11872 25103 11928
rect 21357 11870 25103 11872
rect 21357 11867 21423 11870
rect 25037 11867 25103 11870
rect 29637 11930 29703 11933
rect 32121 11930 32187 11933
rect 29637 11928 32187 11930
rect 29637 11872 29642 11928
rect 29698 11872 32126 11928
rect 32182 11872 32187 11928
rect 29637 11870 32187 11872
rect 29637 11867 29703 11870
rect 32121 11867 32187 11870
rect 5441 11658 5507 11661
rect 11145 11658 11211 11661
rect 5441 11656 11211 11658
rect 5441 11600 5446 11656
rect 5502 11600 11150 11656
rect 11206 11600 11211 11656
rect 5441 11598 11211 11600
rect 5441 11595 5507 11598
rect 11145 11595 11211 11598
rect 42701 11658 42767 11661
rect 49520 11658 50000 11688
rect 42701 11656 50000 11658
rect 42701 11600 42706 11656
rect 42762 11600 50000 11656
rect 42701 11598 50000 11600
rect 42701 11595 42767 11598
rect 49520 11568 50000 11598
rect 12525 11522 12591 11525
rect 15469 11522 15535 11525
rect 12525 11520 15535 11522
rect 12525 11464 12530 11520
rect 12586 11464 15474 11520
rect 15530 11464 15535 11520
rect 12525 11462 15535 11464
rect 12525 11459 12591 11462
rect 15469 11459 15535 11462
rect 19568 11456 19888 11457
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 11391 19888 11392
rect 23657 11250 23723 11253
rect 26601 11250 26667 11253
rect 23657 11248 26667 11250
rect 23657 11192 23662 11248
rect 23718 11192 26606 11248
rect 26662 11192 26667 11248
rect 23657 11190 26667 11192
rect 23657 11187 23723 11190
rect 26601 11187 26667 11190
rect 10409 11114 10475 11117
rect 12985 11114 13051 11117
rect 10409 11112 13051 11114
rect 10409 11056 10414 11112
rect 10470 11056 12990 11112
rect 13046 11056 13051 11112
rect 10409 11054 13051 11056
rect 10409 11051 10475 11054
rect 12985 11051 13051 11054
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 34928 10912 35248 10913
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 10847 35248 10848
rect 5257 10842 5323 10845
rect 11053 10842 11119 10845
rect 5257 10840 11119 10842
rect 5257 10784 5262 10840
rect 5318 10784 11058 10840
rect 11114 10784 11119 10840
rect 5257 10782 11119 10784
rect 5257 10779 5323 10782
rect 11053 10779 11119 10782
rect 11421 10706 11487 10709
rect 20253 10706 20319 10709
rect 11421 10704 20319 10706
rect 11421 10648 11426 10704
rect 11482 10648 20258 10704
rect 20314 10648 20319 10704
rect 11421 10646 20319 10648
rect 11421 10643 11487 10646
rect 20253 10643 20319 10646
rect 20437 10706 20503 10709
rect 22093 10706 22159 10709
rect 27245 10706 27311 10709
rect 20437 10704 27311 10706
rect 20437 10648 20442 10704
rect 20498 10648 22098 10704
rect 22154 10648 27250 10704
rect 27306 10648 27311 10704
rect 20437 10646 27311 10648
rect 20437 10643 20503 10646
rect 22093 10643 22159 10646
rect 27245 10643 27311 10646
rect 43621 10434 43687 10437
rect 46933 10434 46999 10437
rect 43621 10432 46999 10434
rect 43621 10376 43626 10432
rect 43682 10376 46938 10432
rect 46994 10376 46999 10432
rect 43621 10374 46999 10376
rect 43621 10371 43687 10374
rect 46933 10371 46999 10374
rect 19568 10368 19888 10369
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 10303 19888 10304
rect 25405 10298 25471 10301
rect 27981 10298 28047 10301
rect 25405 10296 28047 10298
rect 25405 10240 25410 10296
rect 25466 10240 27986 10296
rect 28042 10240 28047 10296
rect 25405 10238 28047 10240
rect 25405 10235 25471 10238
rect 27981 10235 28047 10238
rect 28809 10298 28875 10301
rect 30465 10298 30531 10301
rect 28809 10296 30531 10298
rect 28809 10240 28814 10296
rect 28870 10240 30470 10296
rect 30526 10240 30531 10296
rect 28809 10238 30531 10240
rect 28809 10235 28875 10238
rect 30465 10235 30531 10238
rect 40953 10298 41019 10301
rect 43069 10298 43135 10301
rect 40953 10296 43135 10298
rect 40953 10240 40958 10296
rect 41014 10240 43074 10296
rect 43130 10240 43135 10296
rect 40953 10238 43135 10240
rect 40953 10235 41019 10238
rect 43069 10235 43135 10238
rect 5349 10162 5415 10165
rect 6913 10162 6979 10165
rect 5349 10160 6979 10162
rect 5349 10104 5354 10160
rect 5410 10104 6918 10160
rect 6974 10104 6979 10160
rect 5349 10102 6979 10104
rect 5349 10099 5415 10102
rect 6913 10099 6979 10102
rect 26049 10162 26115 10165
rect 33225 10162 33291 10165
rect 26049 10160 33291 10162
rect 26049 10104 26054 10160
rect 26110 10104 33230 10160
rect 33286 10104 33291 10160
rect 26049 10102 33291 10104
rect 26049 10099 26115 10102
rect 33225 10099 33291 10102
rect 42057 10162 42123 10165
rect 46933 10162 46999 10165
rect 42057 10160 46999 10162
rect 42057 10104 42062 10160
rect 42118 10104 46938 10160
rect 46994 10104 46999 10160
rect 42057 10102 46999 10104
rect 42057 10099 42123 10102
rect 46933 10099 46999 10102
rect 47393 10162 47459 10165
rect 49520 10162 50000 10192
rect 47393 10160 50000 10162
rect 47393 10104 47398 10160
rect 47454 10104 50000 10160
rect 47393 10102 50000 10104
rect 47393 10099 47459 10102
rect 49520 10072 50000 10102
rect 25497 10026 25563 10029
rect 27153 10026 27219 10029
rect 25497 10024 27219 10026
rect 25497 9968 25502 10024
rect 25558 9968 27158 10024
rect 27214 9968 27219 10024
rect 25497 9966 27219 9968
rect 25497 9963 25563 9966
rect 27153 9963 27219 9966
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 34928 9824 35248 9825
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 9759 35248 9760
rect 35433 9754 35499 9757
rect 37733 9754 37799 9757
rect 35433 9752 37799 9754
rect 35433 9696 35438 9752
rect 35494 9696 37738 9752
rect 37794 9696 37799 9752
rect 35433 9694 37799 9696
rect 35433 9691 35499 9694
rect 37733 9691 37799 9694
rect 12249 9618 12315 9621
rect 15653 9618 15719 9621
rect 12249 9616 15719 9618
rect 12249 9560 12254 9616
rect 12310 9560 15658 9616
rect 15714 9560 15719 9616
rect 12249 9558 15719 9560
rect 12249 9555 12315 9558
rect 15653 9555 15719 9558
rect 19568 9280 19888 9281
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 9215 19888 9216
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 34928 8736 35248 8737
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 8671 35248 8672
rect 39205 8530 39271 8533
rect 43621 8530 43687 8533
rect 46933 8530 46999 8533
rect 39205 8528 46999 8530
rect 39205 8472 39210 8528
rect 39266 8472 43626 8528
rect 43682 8472 46938 8528
rect 46994 8472 46999 8528
rect 39205 8470 46999 8472
rect 39205 8467 39271 8470
rect 43621 8467 43687 8470
rect 46933 8467 46999 8470
rect 47393 8530 47459 8533
rect 49520 8530 50000 8560
rect 47393 8528 50000 8530
rect 47393 8472 47398 8528
rect 47454 8472 50000 8528
rect 47393 8470 50000 8472
rect 47393 8467 47459 8470
rect 49520 8440 50000 8470
rect 15101 8394 15167 8397
rect 16941 8394 17007 8397
rect 15101 8392 17007 8394
rect 15101 8336 15106 8392
rect 15162 8336 16946 8392
rect 17002 8336 17007 8392
rect 15101 8334 17007 8336
rect 15101 8331 15167 8334
rect 16941 8331 17007 8334
rect 19568 8192 19888 8193
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 8127 19888 8128
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 34928 7648 35248 7649
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 7583 35248 7584
rect 27705 7442 27771 7445
rect 33593 7442 33659 7445
rect 27705 7440 33659 7442
rect 27705 7384 27710 7440
rect 27766 7384 33598 7440
rect 33654 7384 33659 7440
rect 27705 7382 33659 7384
rect 27705 7379 27771 7382
rect 33593 7379 33659 7382
rect 9581 7306 9647 7309
rect 11789 7306 11855 7309
rect 9581 7304 11855 7306
rect 9581 7248 9586 7304
rect 9642 7248 11794 7304
rect 11850 7248 11855 7304
rect 9581 7246 11855 7248
rect 9581 7243 9647 7246
rect 11789 7243 11855 7246
rect 28165 7306 28231 7309
rect 30741 7306 30807 7309
rect 28165 7304 30807 7306
rect 28165 7248 28170 7304
rect 28226 7248 30746 7304
rect 30802 7248 30807 7304
rect 28165 7246 30807 7248
rect 28165 7243 28231 7246
rect 30741 7243 30807 7246
rect 19568 7104 19888 7105
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 7039 19888 7040
rect 44357 7034 44423 7037
rect 45093 7034 45159 7037
rect 46933 7034 46999 7037
rect 44357 7032 46999 7034
rect 44357 6976 44362 7032
rect 44418 6976 45098 7032
rect 45154 6976 46938 7032
rect 46994 6976 46999 7032
rect 44357 6974 46999 6976
rect 44357 6971 44423 6974
rect 45093 6971 45159 6974
rect 46933 6971 46999 6974
rect 47393 7034 47459 7037
rect 49520 7034 50000 7064
rect 47393 7032 50000 7034
rect 47393 6976 47398 7032
rect 47454 6976 50000 7032
rect 47393 6974 50000 6976
rect 47393 6971 47459 6974
rect 49520 6944 50000 6974
rect 6269 6762 6335 6765
rect 10041 6762 10107 6765
rect 6269 6760 10107 6762
rect 6269 6704 6274 6760
rect 6330 6704 10046 6760
rect 10102 6704 10107 6760
rect 6269 6702 10107 6704
rect 6269 6699 6335 6702
rect 10041 6699 10107 6702
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 34928 6560 35248 6561
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 6495 35248 6496
rect 26233 6354 26299 6357
rect 32397 6354 32463 6357
rect 26233 6352 32463 6354
rect 26233 6296 26238 6352
rect 26294 6296 32402 6352
rect 32458 6296 32463 6352
rect 26233 6294 32463 6296
rect 26233 6291 26299 6294
rect 32397 6291 32463 6294
rect 8661 6218 8727 6221
rect 11329 6218 11395 6221
rect 8661 6216 11395 6218
rect 8661 6160 8666 6216
rect 8722 6160 11334 6216
rect 11390 6160 11395 6216
rect 8661 6158 11395 6160
rect 8661 6155 8727 6158
rect 11329 6155 11395 6158
rect 33317 6218 33383 6221
rect 39297 6218 39363 6221
rect 33317 6216 39363 6218
rect 33317 6160 33322 6216
rect 33378 6160 39302 6216
rect 39358 6160 39363 6216
rect 33317 6158 39363 6160
rect 33317 6155 33383 6158
rect 39297 6155 39363 6158
rect 38285 6082 38351 6085
rect 42057 6082 42123 6085
rect 38285 6080 42123 6082
rect 38285 6024 38290 6080
rect 38346 6024 42062 6080
rect 42118 6024 42123 6080
rect 38285 6022 42123 6024
rect 38285 6019 38351 6022
rect 42057 6019 42123 6022
rect 45921 6082 45987 6085
rect 49233 6082 49299 6085
rect 45921 6080 49299 6082
rect 45921 6024 45926 6080
rect 45982 6024 49238 6080
rect 49294 6024 49299 6080
rect 45921 6022 49299 6024
rect 45921 6019 45987 6022
rect 49233 6019 49299 6022
rect 19568 6016 19888 6017
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 5951 19888 5952
rect 20989 5946 21055 5949
rect 30925 5946 30991 5949
rect 20989 5944 30991 5946
rect 20989 5888 20994 5944
rect 21050 5888 30930 5944
rect 30986 5888 30991 5944
rect 20989 5886 30991 5888
rect 20989 5883 21055 5886
rect 30925 5883 30991 5886
rect 11053 5674 11119 5677
rect 17401 5674 17467 5677
rect 11053 5672 17467 5674
rect 11053 5616 11058 5672
rect 11114 5616 17406 5672
rect 17462 5616 17467 5672
rect 11053 5614 17467 5616
rect 11053 5611 11119 5614
rect 17401 5611 17467 5614
rect 22553 5674 22619 5677
rect 25589 5674 25655 5677
rect 22553 5672 25655 5674
rect 22553 5616 22558 5672
rect 22614 5616 25594 5672
rect 25650 5616 25655 5672
rect 22553 5614 25655 5616
rect 22553 5611 22619 5614
rect 25589 5611 25655 5614
rect 35525 5674 35591 5677
rect 38101 5674 38167 5677
rect 35525 5672 38167 5674
rect 35525 5616 35530 5672
rect 35586 5616 38106 5672
rect 38162 5616 38167 5672
rect 35525 5614 38167 5616
rect 35525 5611 35591 5614
rect 38101 5611 38167 5614
rect 21081 5538 21147 5541
rect 23841 5538 23907 5541
rect 21081 5536 23907 5538
rect 21081 5480 21086 5536
rect 21142 5480 23846 5536
rect 23902 5480 23907 5536
rect 21081 5478 23907 5480
rect 21081 5475 21147 5478
rect 23841 5475 23907 5478
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 34928 5472 35248 5473
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 5407 35248 5408
rect 23749 5402 23815 5405
rect 29269 5402 29335 5405
rect 49520 5402 50000 5432
rect 23749 5400 29335 5402
rect 23749 5344 23754 5400
rect 23810 5344 29274 5400
rect 29330 5344 29335 5400
rect 23749 5342 29335 5344
rect 23749 5339 23815 5342
rect 29269 5339 29335 5342
rect 49374 5342 50000 5402
rect 19568 4928 19888 4929
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 4863 19888 4864
rect 9581 4858 9647 4861
rect 11697 4858 11763 4861
rect 9581 4856 11763 4858
rect 9581 4800 9586 4856
rect 9642 4800 11702 4856
rect 11758 4800 11763 4856
rect 9581 4798 11763 4800
rect 9581 4795 9647 4798
rect 11697 4795 11763 4798
rect 19977 4858 20043 4861
rect 22553 4858 22619 4861
rect 19977 4856 22619 4858
rect 19977 4800 19982 4856
rect 20038 4800 22558 4856
rect 22614 4800 22619 4856
rect 19977 4798 22619 4800
rect 19977 4795 20043 4798
rect 22553 4795 22619 4798
rect 38285 4722 38351 4725
rect 40033 4722 40099 4725
rect 38285 4720 40099 4722
rect 38285 4664 38290 4720
rect 38346 4664 40038 4720
rect 40094 4664 40099 4720
rect 38285 4662 40099 4664
rect 38285 4659 38351 4662
rect 40033 4659 40099 4662
rect 8201 4586 8267 4589
rect 11513 4586 11579 4589
rect 8201 4584 11579 4586
rect 8201 4528 8206 4584
rect 8262 4528 11518 4584
rect 11574 4528 11579 4584
rect 8201 4526 11579 4528
rect 8201 4523 8267 4526
rect 11513 4523 11579 4526
rect 25589 4586 25655 4589
rect 26509 4586 26575 4589
rect 31845 4586 31911 4589
rect 25589 4584 31911 4586
rect 25589 4528 25594 4584
rect 25650 4528 26514 4584
rect 26570 4528 31850 4584
rect 31906 4528 31911 4584
rect 25589 4526 31911 4528
rect 25589 4523 25655 4526
rect 26509 4523 26575 4526
rect 31845 4523 31911 4526
rect 33961 4586 34027 4589
rect 37365 4586 37431 4589
rect 33961 4584 37431 4586
rect 33961 4528 33966 4584
rect 34022 4528 37370 4584
rect 37426 4528 37431 4584
rect 33961 4526 37431 4528
rect 33961 4523 34027 4526
rect 37365 4523 37431 4526
rect 11605 4450 11671 4453
rect 13905 4450 13971 4453
rect 16113 4450 16179 4453
rect 11605 4448 16179 4450
rect 11605 4392 11610 4448
rect 11666 4392 13910 4448
rect 13966 4392 16118 4448
rect 16174 4392 16179 4448
rect 11605 4390 16179 4392
rect 11605 4387 11671 4390
rect 13905 4387 13971 4390
rect 16113 4387 16179 4390
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 34928 4384 35248 4385
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 4319 35248 4320
rect 10225 4314 10291 4317
rect 13353 4314 13419 4317
rect 13813 4314 13879 4317
rect 10225 4312 13879 4314
rect 10225 4256 10230 4312
rect 10286 4256 13358 4312
rect 13414 4256 13818 4312
rect 13874 4256 13879 4312
rect 10225 4254 13879 4256
rect 10225 4251 10291 4254
rect 13353 4251 13419 4254
rect 13813 4251 13879 4254
rect 37089 4314 37155 4317
rect 40493 4314 40559 4317
rect 37089 4312 40559 4314
rect 37089 4256 37094 4312
rect 37150 4256 40498 4312
rect 40554 4256 40559 4312
rect 37089 4254 40559 4256
rect 37089 4251 37155 4254
rect 40493 4251 40559 4254
rect 11973 4178 12039 4181
rect 19333 4178 19399 4181
rect 11973 4176 19399 4178
rect 11973 4120 11978 4176
rect 12034 4120 19338 4176
rect 19394 4120 19399 4176
rect 11973 4118 19399 4120
rect 11973 4115 12039 4118
rect 19333 4115 19399 4118
rect 23105 4178 23171 4181
rect 26049 4178 26115 4181
rect 23105 4176 26115 4178
rect 23105 4120 23110 4176
rect 23166 4120 26054 4176
rect 26110 4120 26115 4176
rect 23105 4118 26115 4120
rect 23105 4115 23171 4118
rect 26049 4115 26115 4118
rect 32949 4178 33015 4181
rect 49374 4178 49434 5342
rect 49520 5312 50000 5342
rect 32949 4176 49434 4178
rect 32949 4120 32954 4176
rect 33010 4120 49434 4176
rect 32949 4118 49434 4120
rect 32949 4115 33015 4118
rect 7833 4042 7899 4045
rect 8753 4042 8819 4045
rect 7833 4040 8819 4042
rect 7833 3984 7838 4040
rect 7894 3984 8758 4040
rect 8814 3984 8819 4040
rect 7833 3982 8819 3984
rect 7833 3979 7899 3982
rect 8753 3979 8819 3982
rect 18137 4042 18203 4045
rect 24761 4042 24827 4045
rect 18137 4040 24827 4042
rect 18137 3984 18142 4040
rect 18198 3984 24766 4040
rect 24822 3984 24827 4040
rect 18137 3982 24827 3984
rect 18137 3979 18203 3982
rect 24761 3979 24827 3982
rect 25681 4042 25747 4045
rect 27705 4042 27771 4045
rect 25681 4040 27771 4042
rect 25681 3984 25686 4040
rect 25742 3984 27710 4040
rect 27766 3984 27771 4040
rect 25681 3982 27771 3984
rect 25681 3979 25747 3982
rect 27705 3979 27771 3982
rect 32673 4042 32739 4045
rect 32673 4040 38210 4042
rect 32673 3984 32678 4040
rect 32734 3984 38210 4040
rect 32673 3982 38210 3984
rect 32673 3979 32739 3982
rect 38150 3909 38210 3982
rect 5993 3906 6059 3909
rect 9949 3906 10015 3909
rect 5993 3904 10015 3906
rect 5993 3848 5998 3904
rect 6054 3848 9954 3904
rect 10010 3848 10015 3904
rect 5993 3846 10015 3848
rect 5993 3843 6059 3846
rect 9949 3843 10015 3846
rect 10317 3906 10383 3909
rect 12801 3906 12867 3909
rect 10317 3904 12867 3906
rect 10317 3848 10322 3904
rect 10378 3848 12806 3904
rect 12862 3848 12867 3904
rect 10317 3846 12867 3848
rect 10317 3843 10383 3846
rect 12801 3843 12867 3846
rect 16481 3906 16547 3909
rect 19333 3906 19399 3909
rect 16481 3904 19399 3906
rect 16481 3848 16486 3904
rect 16542 3848 19338 3904
rect 19394 3848 19399 3904
rect 16481 3846 19399 3848
rect 16481 3843 16547 3846
rect 19333 3843 19399 3846
rect 23105 3906 23171 3909
rect 23749 3906 23815 3909
rect 26417 3906 26483 3909
rect 23105 3904 26483 3906
rect 23105 3848 23110 3904
rect 23166 3848 23754 3904
rect 23810 3848 26422 3904
rect 26478 3848 26483 3904
rect 23105 3846 26483 3848
rect 23105 3843 23171 3846
rect 23749 3843 23815 3846
rect 26417 3843 26483 3846
rect 28073 3906 28139 3909
rect 30465 3906 30531 3909
rect 28073 3904 30531 3906
rect 28073 3848 28078 3904
rect 28134 3848 30470 3904
rect 30526 3848 30531 3904
rect 28073 3846 30531 3848
rect 28073 3843 28139 3846
rect 30465 3843 30531 3846
rect 32029 3906 32095 3909
rect 38150 3906 38259 3909
rect 41045 3906 41111 3909
rect 41413 3906 41479 3909
rect 49520 3906 50000 3936
rect 32029 3904 34714 3906
rect 32029 3848 32034 3904
rect 32090 3848 34714 3904
rect 32029 3846 34714 3848
rect 38150 3904 41479 3906
rect 38150 3848 38198 3904
rect 38254 3848 41050 3904
rect 41106 3848 41418 3904
rect 41474 3848 41479 3904
rect 38150 3846 41479 3848
rect 32029 3843 32095 3846
rect 19568 3840 19888 3841
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 3775 19888 3776
rect 30373 3772 30439 3773
rect 30373 3770 30420 3772
rect 30328 3768 30420 3770
rect 30328 3712 30378 3768
rect 30328 3710 30420 3712
rect 30373 3708 30420 3710
rect 30484 3708 30490 3772
rect 33041 3770 33107 3773
rect 34513 3770 34579 3773
rect 33041 3768 34579 3770
rect 33041 3712 33046 3768
rect 33102 3712 34518 3768
rect 34574 3712 34579 3768
rect 33041 3710 34579 3712
rect 34654 3770 34714 3846
rect 38193 3843 38259 3846
rect 41045 3843 41111 3846
rect 41413 3843 41479 3846
rect 45510 3846 50000 3906
rect 45510 3770 45570 3846
rect 49520 3816 50000 3846
rect 34654 3710 45570 3770
rect 30373 3707 30439 3708
rect 33041 3707 33107 3710
rect 34513 3707 34579 3710
rect 19425 3634 19491 3637
rect 24577 3634 24643 3637
rect 19425 3632 24643 3634
rect 19425 3576 19430 3632
rect 19486 3576 24582 3632
rect 24638 3576 24643 3632
rect 19425 3574 24643 3576
rect 19425 3571 19491 3574
rect 24577 3571 24643 3574
rect 28165 3634 28231 3637
rect 31937 3634 32003 3637
rect 28165 3632 32003 3634
rect 28165 3576 28170 3632
rect 28226 3576 31942 3632
rect 31998 3576 32003 3632
rect 28165 3574 32003 3576
rect 28165 3571 28231 3574
rect 31937 3571 32003 3574
rect 41413 3634 41479 3637
rect 47853 3634 47919 3637
rect 41413 3632 47919 3634
rect 41413 3576 41418 3632
rect 41474 3576 47858 3632
rect 47914 3576 47919 3632
rect 41413 3574 47919 3576
rect 41413 3571 41479 3574
rect 47853 3571 47919 3574
rect 2497 3498 2563 3501
rect 4705 3498 4771 3501
rect 2497 3496 4771 3498
rect 2497 3440 2502 3496
rect 2558 3440 4710 3496
rect 4766 3440 4771 3496
rect 2497 3438 4771 3440
rect 2497 3435 2563 3438
rect 4705 3435 4771 3438
rect 15469 3498 15535 3501
rect 20713 3498 20779 3501
rect 20846 3498 20852 3500
rect 15469 3496 20852 3498
rect 15469 3440 15474 3496
rect 15530 3440 20718 3496
rect 20774 3440 20852 3496
rect 15469 3438 20852 3440
rect 15469 3435 15535 3438
rect 20713 3435 20779 3438
rect 20846 3436 20852 3438
rect 20916 3436 20922 3500
rect 23841 3498 23907 3501
rect 27613 3498 27679 3501
rect 23841 3496 27679 3498
rect 23841 3440 23846 3496
rect 23902 3440 27618 3496
rect 27674 3440 27679 3496
rect 23841 3438 27679 3440
rect 23841 3435 23907 3438
rect 27613 3435 27679 3438
rect 16481 3362 16547 3365
rect 18689 3362 18755 3365
rect 16481 3360 18755 3362
rect 16481 3304 16486 3360
rect 16542 3304 18694 3360
rect 18750 3304 18755 3360
rect 16481 3302 18755 3304
rect 16481 3299 16547 3302
rect 18689 3299 18755 3302
rect 22185 3362 22251 3365
rect 32121 3362 32187 3365
rect 22185 3360 32187 3362
rect 22185 3304 22190 3360
rect 22246 3304 32126 3360
rect 32182 3304 32187 3360
rect 22185 3302 32187 3304
rect 22185 3299 22251 3302
rect 32121 3299 32187 3302
rect 4208 3296 4528 3297
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 34928 3296 35248 3297
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 3231 35248 3232
rect 19241 3226 19307 3229
rect 26233 3226 26299 3229
rect 28441 3226 28507 3229
rect 32673 3226 32739 3229
rect 19241 3224 28507 3226
rect 19241 3168 19246 3224
rect 19302 3168 26238 3224
rect 26294 3168 28446 3224
rect 28502 3168 28507 3224
rect 19241 3166 28507 3168
rect 19241 3163 19307 3166
rect 26233 3163 26299 3166
rect 28441 3163 28507 3166
rect 28582 3224 32739 3226
rect 28582 3168 32678 3224
rect 32734 3168 32739 3224
rect 28582 3166 32739 3168
rect 657 3090 723 3093
rect 790 3090 796 3092
rect 657 3088 796 3090
rect 657 3032 662 3088
rect 718 3032 796 3088
rect 657 3030 796 3032
rect 657 3027 723 3030
rect 790 3028 796 3030
rect 860 3028 866 3092
rect 26785 3090 26851 3093
rect 28582 3090 28642 3166
rect 32673 3163 32739 3166
rect 26785 3088 28642 3090
rect 26785 3032 26790 3088
rect 26846 3032 28642 3088
rect 26785 3030 28642 3032
rect 29085 3090 29151 3093
rect 36261 3090 36327 3093
rect 29085 3088 36327 3090
rect 29085 3032 29090 3088
rect 29146 3032 36266 3088
rect 36322 3032 36327 3088
rect 29085 3030 36327 3032
rect 26785 3027 26851 3030
rect 29085 3027 29151 3030
rect 36261 3027 36327 3030
rect 16849 2954 16915 2957
rect 22277 2954 22343 2957
rect 16849 2952 22343 2954
rect 16849 2896 16854 2952
rect 16910 2896 22282 2952
rect 22338 2896 22343 2952
rect 16849 2894 22343 2896
rect 16849 2891 16915 2894
rect 22277 2891 22343 2894
rect 30189 2954 30255 2957
rect 36629 2954 36695 2957
rect 30189 2952 36695 2954
rect 30189 2896 30194 2952
rect 30250 2896 36634 2952
rect 36690 2896 36695 2952
rect 30189 2894 36695 2896
rect 30189 2891 30255 2894
rect 36629 2891 36695 2894
rect 7557 2818 7623 2821
rect 10041 2818 10107 2821
rect 7557 2816 10107 2818
rect 7557 2760 7562 2816
rect 7618 2760 10046 2816
rect 10102 2760 10107 2816
rect 7557 2758 10107 2760
rect 7557 2755 7623 2758
rect 10041 2755 10107 2758
rect 20897 2818 20963 2821
rect 25589 2818 25655 2821
rect 20897 2816 25655 2818
rect 20897 2760 20902 2816
rect 20958 2760 25594 2816
rect 25650 2760 25655 2816
rect 20897 2758 25655 2760
rect 20897 2755 20963 2758
rect 25589 2755 25655 2758
rect 31109 2818 31175 2821
rect 33041 2818 33107 2821
rect 31109 2816 33107 2818
rect 31109 2760 31114 2816
rect 31170 2760 33046 2816
rect 33102 2760 33107 2816
rect 31109 2758 33107 2760
rect 31109 2755 31175 2758
rect 33041 2755 33107 2758
rect 37825 2818 37891 2821
rect 42701 2818 42767 2821
rect 37825 2816 42767 2818
rect 37825 2760 37830 2816
rect 37886 2760 42706 2816
rect 42762 2760 42767 2816
rect 37825 2758 42767 2760
rect 37825 2755 37891 2758
rect 42701 2755 42767 2758
rect 19568 2752 19888 2753
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2687 19888 2688
rect 49520 2274 50000 2304
rect 47534 2214 50000 2274
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 34928 2208 35248 2209
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2143 35248 2144
rect 36169 1458 36235 1461
rect 47534 1458 47594 2214
rect 49520 2184 50000 2214
rect 36169 1456 47594 1458
rect 36169 1400 36174 1456
rect 36230 1400 47594 1456
rect 36169 1398 47594 1400
rect 36169 1395 36235 1398
rect 49520 778 50000 808
rect 47534 718 50000 778
rect 36077 98 36143 101
rect 47534 98 47594 718
rect 49520 688 50000 718
rect 36077 96 47594 98
rect 36077 40 36082 96
rect 36138 40 47594 96
rect 36077 38 47594 40
rect 36077 35 36143 38
<< via3 >>
rect 19576 47356 19640 47360
rect 19576 47300 19580 47356
rect 19580 47300 19636 47356
rect 19636 47300 19640 47356
rect 19576 47296 19640 47300
rect 19656 47356 19720 47360
rect 19656 47300 19660 47356
rect 19660 47300 19716 47356
rect 19716 47300 19720 47356
rect 19656 47296 19720 47300
rect 19736 47356 19800 47360
rect 19736 47300 19740 47356
rect 19740 47300 19796 47356
rect 19796 47300 19800 47356
rect 19736 47296 19800 47300
rect 19816 47356 19880 47360
rect 19816 47300 19820 47356
rect 19820 47300 19876 47356
rect 19876 47300 19880 47356
rect 19816 47296 19880 47300
rect 4216 46812 4280 46816
rect 4216 46756 4220 46812
rect 4220 46756 4276 46812
rect 4276 46756 4280 46812
rect 4216 46752 4280 46756
rect 4296 46812 4360 46816
rect 4296 46756 4300 46812
rect 4300 46756 4356 46812
rect 4356 46756 4360 46812
rect 4296 46752 4360 46756
rect 4376 46812 4440 46816
rect 4376 46756 4380 46812
rect 4380 46756 4436 46812
rect 4436 46756 4440 46812
rect 4376 46752 4440 46756
rect 4456 46812 4520 46816
rect 4456 46756 4460 46812
rect 4460 46756 4516 46812
rect 4516 46756 4520 46812
rect 4456 46752 4520 46756
rect 34936 46812 35000 46816
rect 34936 46756 34940 46812
rect 34940 46756 34996 46812
rect 34996 46756 35000 46812
rect 34936 46752 35000 46756
rect 35016 46812 35080 46816
rect 35016 46756 35020 46812
rect 35020 46756 35076 46812
rect 35076 46756 35080 46812
rect 35016 46752 35080 46756
rect 35096 46812 35160 46816
rect 35096 46756 35100 46812
rect 35100 46756 35156 46812
rect 35156 46756 35160 46812
rect 35096 46752 35160 46756
rect 35176 46812 35240 46816
rect 35176 46756 35180 46812
rect 35180 46756 35236 46812
rect 35236 46756 35240 46812
rect 35176 46752 35240 46756
rect 19576 46268 19640 46272
rect 19576 46212 19580 46268
rect 19580 46212 19636 46268
rect 19636 46212 19640 46268
rect 19576 46208 19640 46212
rect 19656 46268 19720 46272
rect 19656 46212 19660 46268
rect 19660 46212 19716 46268
rect 19716 46212 19720 46268
rect 19656 46208 19720 46212
rect 19736 46268 19800 46272
rect 19736 46212 19740 46268
rect 19740 46212 19796 46268
rect 19796 46212 19800 46268
rect 19736 46208 19800 46212
rect 19816 46268 19880 46272
rect 19816 46212 19820 46268
rect 19820 46212 19876 46268
rect 19876 46212 19880 46268
rect 19816 46208 19880 46212
rect 4216 45724 4280 45728
rect 4216 45668 4220 45724
rect 4220 45668 4276 45724
rect 4276 45668 4280 45724
rect 4216 45664 4280 45668
rect 4296 45724 4360 45728
rect 4296 45668 4300 45724
rect 4300 45668 4356 45724
rect 4356 45668 4360 45724
rect 4296 45664 4360 45668
rect 4376 45724 4440 45728
rect 4376 45668 4380 45724
rect 4380 45668 4436 45724
rect 4436 45668 4440 45724
rect 4376 45664 4440 45668
rect 4456 45724 4520 45728
rect 4456 45668 4460 45724
rect 4460 45668 4516 45724
rect 4516 45668 4520 45724
rect 4456 45664 4520 45668
rect 34936 45724 35000 45728
rect 34936 45668 34940 45724
rect 34940 45668 34996 45724
rect 34996 45668 35000 45724
rect 34936 45664 35000 45668
rect 35016 45724 35080 45728
rect 35016 45668 35020 45724
rect 35020 45668 35076 45724
rect 35076 45668 35080 45724
rect 35016 45664 35080 45668
rect 35096 45724 35160 45728
rect 35096 45668 35100 45724
rect 35100 45668 35156 45724
rect 35156 45668 35160 45724
rect 35096 45664 35160 45668
rect 35176 45724 35240 45728
rect 35176 45668 35180 45724
rect 35180 45668 35236 45724
rect 35236 45668 35240 45724
rect 35176 45664 35240 45668
rect 19576 45180 19640 45184
rect 19576 45124 19580 45180
rect 19580 45124 19636 45180
rect 19636 45124 19640 45180
rect 19576 45120 19640 45124
rect 19656 45180 19720 45184
rect 19656 45124 19660 45180
rect 19660 45124 19716 45180
rect 19716 45124 19720 45180
rect 19656 45120 19720 45124
rect 19736 45180 19800 45184
rect 19736 45124 19740 45180
rect 19740 45124 19796 45180
rect 19796 45124 19800 45180
rect 19736 45120 19800 45124
rect 19816 45180 19880 45184
rect 19816 45124 19820 45180
rect 19820 45124 19876 45180
rect 19876 45124 19880 45180
rect 19816 45120 19880 45124
rect 4216 44636 4280 44640
rect 4216 44580 4220 44636
rect 4220 44580 4276 44636
rect 4276 44580 4280 44636
rect 4216 44576 4280 44580
rect 4296 44636 4360 44640
rect 4296 44580 4300 44636
rect 4300 44580 4356 44636
rect 4356 44580 4360 44636
rect 4296 44576 4360 44580
rect 4376 44636 4440 44640
rect 4376 44580 4380 44636
rect 4380 44580 4436 44636
rect 4436 44580 4440 44636
rect 4376 44576 4440 44580
rect 4456 44636 4520 44640
rect 4456 44580 4460 44636
rect 4460 44580 4516 44636
rect 4516 44580 4520 44636
rect 4456 44576 4520 44580
rect 34936 44636 35000 44640
rect 34936 44580 34940 44636
rect 34940 44580 34996 44636
rect 34996 44580 35000 44636
rect 34936 44576 35000 44580
rect 35016 44636 35080 44640
rect 35016 44580 35020 44636
rect 35020 44580 35076 44636
rect 35076 44580 35080 44636
rect 35016 44576 35080 44580
rect 35096 44636 35160 44640
rect 35096 44580 35100 44636
rect 35100 44580 35156 44636
rect 35156 44580 35160 44636
rect 35096 44576 35160 44580
rect 35176 44636 35240 44640
rect 35176 44580 35180 44636
rect 35180 44580 35236 44636
rect 35236 44580 35240 44636
rect 35176 44576 35240 44580
rect 19576 44092 19640 44096
rect 19576 44036 19580 44092
rect 19580 44036 19636 44092
rect 19636 44036 19640 44092
rect 19576 44032 19640 44036
rect 19656 44092 19720 44096
rect 19656 44036 19660 44092
rect 19660 44036 19716 44092
rect 19716 44036 19720 44092
rect 19656 44032 19720 44036
rect 19736 44092 19800 44096
rect 19736 44036 19740 44092
rect 19740 44036 19796 44092
rect 19796 44036 19800 44092
rect 19736 44032 19800 44036
rect 19816 44092 19880 44096
rect 19816 44036 19820 44092
rect 19820 44036 19876 44092
rect 19876 44036 19880 44092
rect 19816 44032 19880 44036
rect 4216 43548 4280 43552
rect 4216 43492 4220 43548
rect 4220 43492 4276 43548
rect 4276 43492 4280 43548
rect 4216 43488 4280 43492
rect 4296 43548 4360 43552
rect 4296 43492 4300 43548
rect 4300 43492 4356 43548
rect 4356 43492 4360 43548
rect 4296 43488 4360 43492
rect 4376 43548 4440 43552
rect 4376 43492 4380 43548
rect 4380 43492 4436 43548
rect 4436 43492 4440 43548
rect 4376 43488 4440 43492
rect 4456 43548 4520 43552
rect 4456 43492 4460 43548
rect 4460 43492 4516 43548
rect 4516 43492 4520 43548
rect 4456 43488 4520 43492
rect 34936 43548 35000 43552
rect 34936 43492 34940 43548
rect 34940 43492 34996 43548
rect 34996 43492 35000 43548
rect 34936 43488 35000 43492
rect 35016 43548 35080 43552
rect 35016 43492 35020 43548
rect 35020 43492 35076 43548
rect 35076 43492 35080 43548
rect 35016 43488 35080 43492
rect 35096 43548 35160 43552
rect 35096 43492 35100 43548
rect 35100 43492 35156 43548
rect 35156 43492 35160 43548
rect 35096 43488 35160 43492
rect 35176 43548 35240 43552
rect 35176 43492 35180 43548
rect 35180 43492 35236 43548
rect 35236 43492 35240 43548
rect 35176 43488 35240 43492
rect 19576 43004 19640 43008
rect 19576 42948 19580 43004
rect 19580 42948 19636 43004
rect 19636 42948 19640 43004
rect 19576 42944 19640 42948
rect 19656 43004 19720 43008
rect 19656 42948 19660 43004
rect 19660 42948 19716 43004
rect 19716 42948 19720 43004
rect 19656 42944 19720 42948
rect 19736 43004 19800 43008
rect 19736 42948 19740 43004
rect 19740 42948 19796 43004
rect 19796 42948 19800 43004
rect 19736 42944 19800 42948
rect 19816 43004 19880 43008
rect 19816 42948 19820 43004
rect 19820 42948 19876 43004
rect 19876 42948 19880 43004
rect 19816 42944 19880 42948
rect 4216 42460 4280 42464
rect 4216 42404 4220 42460
rect 4220 42404 4276 42460
rect 4276 42404 4280 42460
rect 4216 42400 4280 42404
rect 4296 42460 4360 42464
rect 4296 42404 4300 42460
rect 4300 42404 4356 42460
rect 4356 42404 4360 42460
rect 4296 42400 4360 42404
rect 4376 42460 4440 42464
rect 4376 42404 4380 42460
rect 4380 42404 4436 42460
rect 4436 42404 4440 42460
rect 4376 42400 4440 42404
rect 4456 42460 4520 42464
rect 4456 42404 4460 42460
rect 4460 42404 4516 42460
rect 4516 42404 4520 42460
rect 4456 42400 4520 42404
rect 34936 42460 35000 42464
rect 34936 42404 34940 42460
rect 34940 42404 34996 42460
rect 34996 42404 35000 42460
rect 34936 42400 35000 42404
rect 35016 42460 35080 42464
rect 35016 42404 35020 42460
rect 35020 42404 35076 42460
rect 35076 42404 35080 42460
rect 35016 42400 35080 42404
rect 35096 42460 35160 42464
rect 35096 42404 35100 42460
rect 35100 42404 35156 42460
rect 35156 42404 35160 42460
rect 35096 42400 35160 42404
rect 35176 42460 35240 42464
rect 35176 42404 35180 42460
rect 35180 42404 35236 42460
rect 35236 42404 35240 42460
rect 35176 42400 35240 42404
rect 19576 41916 19640 41920
rect 19576 41860 19580 41916
rect 19580 41860 19636 41916
rect 19636 41860 19640 41916
rect 19576 41856 19640 41860
rect 19656 41916 19720 41920
rect 19656 41860 19660 41916
rect 19660 41860 19716 41916
rect 19716 41860 19720 41916
rect 19656 41856 19720 41860
rect 19736 41916 19800 41920
rect 19736 41860 19740 41916
rect 19740 41860 19796 41916
rect 19796 41860 19800 41916
rect 19736 41856 19800 41860
rect 19816 41916 19880 41920
rect 19816 41860 19820 41916
rect 19820 41860 19876 41916
rect 19876 41860 19880 41916
rect 19816 41856 19880 41860
rect 4216 41372 4280 41376
rect 4216 41316 4220 41372
rect 4220 41316 4276 41372
rect 4276 41316 4280 41372
rect 4216 41312 4280 41316
rect 4296 41372 4360 41376
rect 4296 41316 4300 41372
rect 4300 41316 4356 41372
rect 4356 41316 4360 41372
rect 4296 41312 4360 41316
rect 4376 41372 4440 41376
rect 4376 41316 4380 41372
rect 4380 41316 4436 41372
rect 4436 41316 4440 41372
rect 4376 41312 4440 41316
rect 4456 41372 4520 41376
rect 4456 41316 4460 41372
rect 4460 41316 4516 41372
rect 4516 41316 4520 41372
rect 4456 41312 4520 41316
rect 34936 41372 35000 41376
rect 34936 41316 34940 41372
rect 34940 41316 34996 41372
rect 34996 41316 35000 41372
rect 34936 41312 35000 41316
rect 35016 41372 35080 41376
rect 35016 41316 35020 41372
rect 35020 41316 35076 41372
rect 35076 41316 35080 41372
rect 35016 41312 35080 41316
rect 35096 41372 35160 41376
rect 35096 41316 35100 41372
rect 35100 41316 35156 41372
rect 35156 41316 35160 41372
rect 35096 41312 35160 41316
rect 35176 41372 35240 41376
rect 35176 41316 35180 41372
rect 35180 41316 35236 41372
rect 35236 41316 35240 41372
rect 35176 41312 35240 41316
rect 19576 40828 19640 40832
rect 19576 40772 19580 40828
rect 19580 40772 19636 40828
rect 19636 40772 19640 40828
rect 19576 40768 19640 40772
rect 19656 40828 19720 40832
rect 19656 40772 19660 40828
rect 19660 40772 19716 40828
rect 19716 40772 19720 40828
rect 19656 40768 19720 40772
rect 19736 40828 19800 40832
rect 19736 40772 19740 40828
rect 19740 40772 19796 40828
rect 19796 40772 19800 40828
rect 19736 40768 19800 40772
rect 19816 40828 19880 40832
rect 19816 40772 19820 40828
rect 19820 40772 19876 40828
rect 19876 40772 19880 40828
rect 19816 40768 19880 40772
rect 4216 40284 4280 40288
rect 4216 40228 4220 40284
rect 4220 40228 4276 40284
rect 4276 40228 4280 40284
rect 4216 40224 4280 40228
rect 4296 40284 4360 40288
rect 4296 40228 4300 40284
rect 4300 40228 4356 40284
rect 4356 40228 4360 40284
rect 4296 40224 4360 40228
rect 4376 40284 4440 40288
rect 4376 40228 4380 40284
rect 4380 40228 4436 40284
rect 4436 40228 4440 40284
rect 4376 40224 4440 40228
rect 4456 40284 4520 40288
rect 4456 40228 4460 40284
rect 4460 40228 4516 40284
rect 4516 40228 4520 40284
rect 4456 40224 4520 40228
rect 34936 40284 35000 40288
rect 34936 40228 34940 40284
rect 34940 40228 34996 40284
rect 34996 40228 35000 40284
rect 34936 40224 35000 40228
rect 35016 40284 35080 40288
rect 35016 40228 35020 40284
rect 35020 40228 35076 40284
rect 35076 40228 35080 40284
rect 35016 40224 35080 40228
rect 35096 40284 35160 40288
rect 35096 40228 35100 40284
rect 35100 40228 35156 40284
rect 35156 40228 35160 40284
rect 35096 40224 35160 40228
rect 35176 40284 35240 40288
rect 35176 40228 35180 40284
rect 35180 40228 35236 40284
rect 35236 40228 35240 40284
rect 35176 40224 35240 40228
rect 19576 39740 19640 39744
rect 19576 39684 19580 39740
rect 19580 39684 19636 39740
rect 19636 39684 19640 39740
rect 19576 39680 19640 39684
rect 19656 39740 19720 39744
rect 19656 39684 19660 39740
rect 19660 39684 19716 39740
rect 19716 39684 19720 39740
rect 19656 39680 19720 39684
rect 19736 39740 19800 39744
rect 19736 39684 19740 39740
rect 19740 39684 19796 39740
rect 19796 39684 19800 39740
rect 19736 39680 19800 39684
rect 19816 39740 19880 39744
rect 19816 39684 19820 39740
rect 19820 39684 19876 39740
rect 19876 39684 19880 39740
rect 19816 39680 19880 39684
rect 4216 39196 4280 39200
rect 4216 39140 4220 39196
rect 4220 39140 4276 39196
rect 4276 39140 4280 39196
rect 4216 39136 4280 39140
rect 4296 39196 4360 39200
rect 4296 39140 4300 39196
rect 4300 39140 4356 39196
rect 4356 39140 4360 39196
rect 4296 39136 4360 39140
rect 4376 39196 4440 39200
rect 4376 39140 4380 39196
rect 4380 39140 4436 39196
rect 4436 39140 4440 39196
rect 4376 39136 4440 39140
rect 4456 39196 4520 39200
rect 4456 39140 4460 39196
rect 4460 39140 4516 39196
rect 4516 39140 4520 39196
rect 4456 39136 4520 39140
rect 34936 39196 35000 39200
rect 34936 39140 34940 39196
rect 34940 39140 34996 39196
rect 34996 39140 35000 39196
rect 34936 39136 35000 39140
rect 35016 39196 35080 39200
rect 35016 39140 35020 39196
rect 35020 39140 35076 39196
rect 35076 39140 35080 39196
rect 35016 39136 35080 39140
rect 35096 39196 35160 39200
rect 35096 39140 35100 39196
rect 35100 39140 35156 39196
rect 35156 39140 35160 39196
rect 35096 39136 35160 39140
rect 35176 39196 35240 39200
rect 35176 39140 35180 39196
rect 35180 39140 35236 39196
rect 35236 39140 35240 39196
rect 35176 39136 35240 39140
rect 19576 38652 19640 38656
rect 19576 38596 19580 38652
rect 19580 38596 19636 38652
rect 19636 38596 19640 38652
rect 19576 38592 19640 38596
rect 19656 38652 19720 38656
rect 19656 38596 19660 38652
rect 19660 38596 19716 38652
rect 19716 38596 19720 38652
rect 19656 38592 19720 38596
rect 19736 38652 19800 38656
rect 19736 38596 19740 38652
rect 19740 38596 19796 38652
rect 19796 38596 19800 38652
rect 19736 38592 19800 38596
rect 19816 38652 19880 38656
rect 19816 38596 19820 38652
rect 19820 38596 19876 38652
rect 19876 38596 19880 38652
rect 19816 38592 19880 38596
rect 4216 38108 4280 38112
rect 4216 38052 4220 38108
rect 4220 38052 4276 38108
rect 4276 38052 4280 38108
rect 4216 38048 4280 38052
rect 4296 38108 4360 38112
rect 4296 38052 4300 38108
rect 4300 38052 4356 38108
rect 4356 38052 4360 38108
rect 4296 38048 4360 38052
rect 4376 38108 4440 38112
rect 4376 38052 4380 38108
rect 4380 38052 4436 38108
rect 4436 38052 4440 38108
rect 4376 38048 4440 38052
rect 4456 38108 4520 38112
rect 4456 38052 4460 38108
rect 4460 38052 4516 38108
rect 4516 38052 4520 38108
rect 4456 38048 4520 38052
rect 34936 38108 35000 38112
rect 34936 38052 34940 38108
rect 34940 38052 34996 38108
rect 34996 38052 35000 38108
rect 34936 38048 35000 38052
rect 35016 38108 35080 38112
rect 35016 38052 35020 38108
rect 35020 38052 35076 38108
rect 35076 38052 35080 38108
rect 35016 38048 35080 38052
rect 35096 38108 35160 38112
rect 35096 38052 35100 38108
rect 35100 38052 35156 38108
rect 35156 38052 35160 38108
rect 35096 38048 35160 38052
rect 35176 38108 35240 38112
rect 35176 38052 35180 38108
rect 35180 38052 35236 38108
rect 35236 38052 35240 38108
rect 35176 38048 35240 38052
rect 19576 37564 19640 37568
rect 19576 37508 19580 37564
rect 19580 37508 19636 37564
rect 19636 37508 19640 37564
rect 19576 37504 19640 37508
rect 19656 37564 19720 37568
rect 19656 37508 19660 37564
rect 19660 37508 19716 37564
rect 19716 37508 19720 37564
rect 19656 37504 19720 37508
rect 19736 37564 19800 37568
rect 19736 37508 19740 37564
rect 19740 37508 19796 37564
rect 19796 37508 19800 37564
rect 19736 37504 19800 37508
rect 19816 37564 19880 37568
rect 19816 37508 19820 37564
rect 19820 37508 19876 37564
rect 19876 37508 19880 37564
rect 19816 37504 19880 37508
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 34936 37020 35000 37024
rect 34936 36964 34940 37020
rect 34940 36964 34996 37020
rect 34996 36964 35000 37020
rect 34936 36960 35000 36964
rect 35016 37020 35080 37024
rect 35016 36964 35020 37020
rect 35020 36964 35076 37020
rect 35076 36964 35080 37020
rect 35016 36960 35080 36964
rect 35096 37020 35160 37024
rect 35096 36964 35100 37020
rect 35100 36964 35156 37020
rect 35156 36964 35160 37020
rect 35096 36960 35160 36964
rect 35176 37020 35240 37024
rect 35176 36964 35180 37020
rect 35180 36964 35236 37020
rect 35236 36964 35240 37020
rect 35176 36960 35240 36964
rect 19576 36476 19640 36480
rect 19576 36420 19580 36476
rect 19580 36420 19636 36476
rect 19636 36420 19640 36476
rect 19576 36416 19640 36420
rect 19656 36476 19720 36480
rect 19656 36420 19660 36476
rect 19660 36420 19716 36476
rect 19716 36420 19720 36476
rect 19656 36416 19720 36420
rect 19736 36476 19800 36480
rect 19736 36420 19740 36476
rect 19740 36420 19796 36476
rect 19796 36420 19800 36476
rect 19736 36416 19800 36420
rect 19816 36476 19880 36480
rect 19816 36420 19820 36476
rect 19820 36420 19876 36476
rect 19876 36420 19880 36476
rect 19816 36416 19880 36420
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 34936 35932 35000 35936
rect 34936 35876 34940 35932
rect 34940 35876 34996 35932
rect 34996 35876 35000 35932
rect 34936 35872 35000 35876
rect 35016 35932 35080 35936
rect 35016 35876 35020 35932
rect 35020 35876 35076 35932
rect 35076 35876 35080 35932
rect 35016 35872 35080 35876
rect 35096 35932 35160 35936
rect 35096 35876 35100 35932
rect 35100 35876 35156 35932
rect 35156 35876 35160 35932
rect 35096 35872 35160 35876
rect 35176 35932 35240 35936
rect 35176 35876 35180 35932
rect 35180 35876 35236 35932
rect 35236 35876 35240 35932
rect 35176 35872 35240 35876
rect 19576 35388 19640 35392
rect 19576 35332 19580 35388
rect 19580 35332 19636 35388
rect 19636 35332 19640 35388
rect 19576 35328 19640 35332
rect 19656 35388 19720 35392
rect 19656 35332 19660 35388
rect 19660 35332 19716 35388
rect 19716 35332 19720 35388
rect 19656 35328 19720 35332
rect 19736 35388 19800 35392
rect 19736 35332 19740 35388
rect 19740 35332 19796 35388
rect 19796 35332 19800 35388
rect 19736 35328 19800 35332
rect 19816 35388 19880 35392
rect 19816 35332 19820 35388
rect 19820 35332 19876 35388
rect 19876 35332 19880 35388
rect 19816 35328 19880 35332
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 34936 34844 35000 34848
rect 34936 34788 34940 34844
rect 34940 34788 34996 34844
rect 34996 34788 35000 34844
rect 34936 34784 35000 34788
rect 35016 34844 35080 34848
rect 35016 34788 35020 34844
rect 35020 34788 35076 34844
rect 35076 34788 35080 34844
rect 35016 34784 35080 34788
rect 35096 34844 35160 34848
rect 35096 34788 35100 34844
rect 35100 34788 35156 34844
rect 35156 34788 35160 34844
rect 35096 34784 35160 34788
rect 35176 34844 35240 34848
rect 35176 34788 35180 34844
rect 35180 34788 35236 34844
rect 35236 34788 35240 34844
rect 35176 34784 35240 34788
rect 19576 34300 19640 34304
rect 19576 34244 19580 34300
rect 19580 34244 19636 34300
rect 19636 34244 19640 34300
rect 19576 34240 19640 34244
rect 19656 34300 19720 34304
rect 19656 34244 19660 34300
rect 19660 34244 19716 34300
rect 19716 34244 19720 34300
rect 19656 34240 19720 34244
rect 19736 34300 19800 34304
rect 19736 34244 19740 34300
rect 19740 34244 19796 34300
rect 19796 34244 19800 34300
rect 19736 34240 19800 34244
rect 19816 34300 19880 34304
rect 19816 34244 19820 34300
rect 19820 34244 19876 34300
rect 19876 34244 19880 34300
rect 19816 34240 19880 34244
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 34936 33756 35000 33760
rect 34936 33700 34940 33756
rect 34940 33700 34996 33756
rect 34996 33700 35000 33756
rect 34936 33696 35000 33700
rect 35016 33756 35080 33760
rect 35016 33700 35020 33756
rect 35020 33700 35076 33756
rect 35076 33700 35080 33756
rect 35016 33696 35080 33700
rect 35096 33756 35160 33760
rect 35096 33700 35100 33756
rect 35100 33700 35156 33756
rect 35156 33700 35160 33756
rect 35096 33696 35160 33700
rect 35176 33756 35240 33760
rect 35176 33700 35180 33756
rect 35180 33700 35236 33756
rect 35236 33700 35240 33756
rect 35176 33696 35240 33700
rect 19576 33212 19640 33216
rect 19576 33156 19580 33212
rect 19580 33156 19636 33212
rect 19636 33156 19640 33212
rect 19576 33152 19640 33156
rect 19656 33212 19720 33216
rect 19656 33156 19660 33212
rect 19660 33156 19716 33212
rect 19716 33156 19720 33212
rect 19656 33152 19720 33156
rect 19736 33212 19800 33216
rect 19736 33156 19740 33212
rect 19740 33156 19796 33212
rect 19796 33156 19800 33212
rect 19736 33152 19800 33156
rect 19816 33212 19880 33216
rect 19816 33156 19820 33212
rect 19820 33156 19876 33212
rect 19876 33156 19880 33212
rect 19816 33152 19880 33156
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 34936 32668 35000 32672
rect 34936 32612 34940 32668
rect 34940 32612 34996 32668
rect 34996 32612 35000 32668
rect 34936 32608 35000 32612
rect 35016 32668 35080 32672
rect 35016 32612 35020 32668
rect 35020 32612 35076 32668
rect 35076 32612 35080 32668
rect 35016 32608 35080 32612
rect 35096 32668 35160 32672
rect 35096 32612 35100 32668
rect 35100 32612 35156 32668
rect 35156 32612 35160 32668
rect 35096 32608 35160 32612
rect 35176 32668 35240 32672
rect 35176 32612 35180 32668
rect 35180 32612 35236 32668
rect 35236 32612 35240 32668
rect 35176 32608 35240 32612
rect 19576 32124 19640 32128
rect 19576 32068 19580 32124
rect 19580 32068 19636 32124
rect 19636 32068 19640 32124
rect 19576 32064 19640 32068
rect 19656 32124 19720 32128
rect 19656 32068 19660 32124
rect 19660 32068 19716 32124
rect 19716 32068 19720 32124
rect 19656 32064 19720 32068
rect 19736 32124 19800 32128
rect 19736 32068 19740 32124
rect 19740 32068 19796 32124
rect 19796 32068 19800 32124
rect 19736 32064 19800 32068
rect 19816 32124 19880 32128
rect 19816 32068 19820 32124
rect 19820 32068 19876 32124
rect 19876 32068 19880 32124
rect 19816 32064 19880 32068
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 34936 31580 35000 31584
rect 34936 31524 34940 31580
rect 34940 31524 34996 31580
rect 34996 31524 35000 31580
rect 34936 31520 35000 31524
rect 35016 31580 35080 31584
rect 35016 31524 35020 31580
rect 35020 31524 35076 31580
rect 35076 31524 35080 31580
rect 35016 31520 35080 31524
rect 35096 31580 35160 31584
rect 35096 31524 35100 31580
rect 35100 31524 35156 31580
rect 35156 31524 35160 31580
rect 35096 31520 35160 31524
rect 35176 31580 35240 31584
rect 35176 31524 35180 31580
rect 35180 31524 35236 31580
rect 35236 31524 35240 31580
rect 35176 31520 35240 31524
rect 19576 31036 19640 31040
rect 19576 30980 19580 31036
rect 19580 30980 19636 31036
rect 19636 30980 19640 31036
rect 19576 30976 19640 30980
rect 19656 31036 19720 31040
rect 19656 30980 19660 31036
rect 19660 30980 19716 31036
rect 19716 30980 19720 31036
rect 19656 30976 19720 30980
rect 19736 31036 19800 31040
rect 19736 30980 19740 31036
rect 19740 30980 19796 31036
rect 19796 30980 19800 31036
rect 19736 30976 19800 30980
rect 19816 31036 19880 31040
rect 19816 30980 19820 31036
rect 19820 30980 19876 31036
rect 19876 30980 19880 31036
rect 19816 30976 19880 30980
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 34936 30492 35000 30496
rect 34936 30436 34940 30492
rect 34940 30436 34996 30492
rect 34996 30436 35000 30492
rect 34936 30432 35000 30436
rect 35016 30492 35080 30496
rect 35016 30436 35020 30492
rect 35020 30436 35076 30492
rect 35076 30436 35080 30492
rect 35016 30432 35080 30436
rect 35096 30492 35160 30496
rect 35096 30436 35100 30492
rect 35100 30436 35156 30492
rect 35156 30436 35160 30492
rect 35096 30432 35160 30436
rect 35176 30492 35240 30496
rect 35176 30436 35180 30492
rect 35180 30436 35236 30492
rect 35236 30436 35240 30492
rect 35176 30432 35240 30436
rect 19576 29948 19640 29952
rect 19576 29892 19580 29948
rect 19580 29892 19636 29948
rect 19636 29892 19640 29948
rect 19576 29888 19640 29892
rect 19656 29948 19720 29952
rect 19656 29892 19660 29948
rect 19660 29892 19716 29948
rect 19716 29892 19720 29948
rect 19656 29888 19720 29892
rect 19736 29948 19800 29952
rect 19736 29892 19740 29948
rect 19740 29892 19796 29948
rect 19796 29892 19800 29948
rect 19736 29888 19800 29892
rect 19816 29948 19880 29952
rect 19816 29892 19820 29948
rect 19820 29892 19876 29948
rect 19876 29892 19880 29948
rect 19816 29888 19880 29892
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 34936 29404 35000 29408
rect 34936 29348 34940 29404
rect 34940 29348 34996 29404
rect 34996 29348 35000 29404
rect 34936 29344 35000 29348
rect 35016 29404 35080 29408
rect 35016 29348 35020 29404
rect 35020 29348 35076 29404
rect 35076 29348 35080 29404
rect 35016 29344 35080 29348
rect 35096 29404 35160 29408
rect 35096 29348 35100 29404
rect 35100 29348 35156 29404
rect 35156 29348 35160 29404
rect 35096 29344 35160 29348
rect 35176 29404 35240 29408
rect 35176 29348 35180 29404
rect 35180 29348 35236 29404
rect 35236 29348 35240 29404
rect 35176 29344 35240 29348
rect 19576 28860 19640 28864
rect 19576 28804 19580 28860
rect 19580 28804 19636 28860
rect 19636 28804 19640 28860
rect 19576 28800 19640 28804
rect 19656 28860 19720 28864
rect 19656 28804 19660 28860
rect 19660 28804 19716 28860
rect 19716 28804 19720 28860
rect 19656 28800 19720 28804
rect 19736 28860 19800 28864
rect 19736 28804 19740 28860
rect 19740 28804 19796 28860
rect 19796 28804 19800 28860
rect 19736 28800 19800 28804
rect 19816 28860 19880 28864
rect 19816 28804 19820 28860
rect 19820 28804 19876 28860
rect 19876 28804 19880 28860
rect 19816 28800 19880 28804
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 34936 28316 35000 28320
rect 34936 28260 34940 28316
rect 34940 28260 34996 28316
rect 34996 28260 35000 28316
rect 34936 28256 35000 28260
rect 35016 28316 35080 28320
rect 35016 28260 35020 28316
rect 35020 28260 35076 28316
rect 35076 28260 35080 28316
rect 35016 28256 35080 28260
rect 35096 28316 35160 28320
rect 35096 28260 35100 28316
rect 35100 28260 35156 28316
rect 35156 28260 35160 28316
rect 35096 28256 35160 28260
rect 35176 28316 35240 28320
rect 35176 28260 35180 28316
rect 35180 28260 35236 28316
rect 35236 28260 35240 28316
rect 35176 28256 35240 28260
rect 19576 27772 19640 27776
rect 19576 27716 19580 27772
rect 19580 27716 19636 27772
rect 19636 27716 19640 27772
rect 19576 27712 19640 27716
rect 19656 27772 19720 27776
rect 19656 27716 19660 27772
rect 19660 27716 19716 27772
rect 19716 27716 19720 27772
rect 19656 27712 19720 27716
rect 19736 27772 19800 27776
rect 19736 27716 19740 27772
rect 19740 27716 19796 27772
rect 19796 27716 19800 27772
rect 19736 27712 19800 27716
rect 19816 27772 19880 27776
rect 19816 27716 19820 27772
rect 19820 27716 19876 27772
rect 19876 27716 19880 27772
rect 19816 27712 19880 27716
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 34936 27228 35000 27232
rect 34936 27172 34940 27228
rect 34940 27172 34996 27228
rect 34996 27172 35000 27228
rect 34936 27168 35000 27172
rect 35016 27228 35080 27232
rect 35016 27172 35020 27228
rect 35020 27172 35076 27228
rect 35076 27172 35080 27228
rect 35016 27168 35080 27172
rect 35096 27228 35160 27232
rect 35096 27172 35100 27228
rect 35100 27172 35156 27228
rect 35156 27172 35160 27228
rect 35096 27168 35160 27172
rect 35176 27228 35240 27232
rect 35176 27172 35180 27228
rect 35180 27172 35236 27228
rect 35236 27172 35240 27228
rect 35176 27168 35240 27172
rect 19576 26684 19640 26688
rect 19576 26628 19580 26684
rect 19580 26628 19636 26684
rect 19636 26628 19640 26684
rect 19576 26624 19640 26628
rect 19656 26684 19720 26688
rect 19656 26628 19660 26684
rect 19660 26628 19716 26684
rect 19716 26628 19720 26684
rect 19656 26624 19720 26628
rect 19736 26684 19800 26688
rect 19736 26628 19740 26684
rect 19740 26628 19796 26684
rect 19796 26628 19800 26684
rect 19736 26624 19800 26628
rect 19816 26684 19880 26688
rect 19816 26628 19820 26684
rect 19820 26628 19876 26684
rect 19876 26628 19880 26684
rect 19816 26624 19880 26628
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 34936 26140 35000 26144
rect 34936 26084 34940 26140
rect 34940 26084 34996 26140
rect 34996 26084 35000 26140
rect 34936 26080 35000 26084
rect 35016 26140 35080 26144
rect 35016 26084 35020 26140
rect 35020 26084 35076 26140
rect 35076 26084 35080 26140
rect 35016 26080 35080 26084
rect 35096 26140 35160 26144
rect 35096 26084 35100 26140
rect 35100 26084 35156 26140
rect 35156 26084 35160 26140
rect 35096 26080 35160 26084
rect 35176 26140 35240 26144
rect 35176 26084 35180 26140
rect 35180 26084 35236 26140
rect 35236 26084 35240 26140
rect 35176 26080 35240 26084
rect 19576 25596 19640 25600
rect 19576 25540 19580 25596
rect 19580 25540 19636 25596
rect 19636 25540 19640 25596
rect 19576 25536 19640 25540
rect 19656 25596 19720 25600
rect 19656 25540 19660 25596
rect 19660 25540 19716 25596
rect 19716 25540 19720 25596
rect 19656 25536 19720 25540
rect 19736 25596 19800 25600
rect 19736 25540 19740 25596
rect 19740 25540 19796 25596
rect 19796 25540 19800 25596
rect 19736 25536 19800 25540
rect 19816 25596 19880 25600
rect 19816 25540 19820 25596
rect 19820 25540 19876 25596
rect 19876 25540 19880 25596
rect 19816 25536 19880 25540
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 34936 25052 35000 25056
rect 34936 24996 34940 25052
rect 34940 24996 34996 25052
rect 34996 24996 35000 25052
rect 34936 24992 35000 24996
rect 35016 25052 35080 25056
rect 35016 24996 35020 25052
rect 35020 24996 35076 25052
rect 35076 24996 35080 25052
rect 35016 24992 35080 24996
rect 35096 25052 35160 25056
rect 35096 24996 35100 25052
rect 35100 24996 35156 25052
rect 35156 24996 35160 25052
rect 35096 24992 35160 24996
rect 35176 25052 35240 25056
rect 35176 24996 35180 25052
rect 35180 24996 35236 25052
rect 35236 24996 35240 25052
rect 35176 24992 35240 24996
rect 19576 24508 19640 24512
rect 19576 24452 19580 24508
rect 19580 24452 19636 24508
rect 19636 24452 19640 24508
rect 19576 24448 19640 24452
rect 19656 24508 19720 24512
rect 19656 24452 19660 24508
rect 19660 24452 19716 24508
rect 19716 24452 19720 24508
rect 19656 24448 19720 24452
rect 19736 24508 19800 24512
rect 19736 24452 19740 24508
rect 19740 24452 19796 24508
rect 19796 24452 19800 24508
rect 19736 24448 19800 24452
rect 19816 24508 19880 24512
rect 19816 24452 19820 24508
rect 19820 24452 19876 24508
rect 19876 24452 19880 24508
rect 19816 24448 19880 24452
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 34936 23964 35000 23968
rect 34936 23908 34940 23964
rect 34940 23908 34996 23964
rect 34996 23908 35000 23964
rect 34936 23904 35000 23908
rect 35016 23964 35080 23968
rect 35016 23908 35020 23964
rect 35020 23908 35076 23964
rect 35076 23908 35080 23964
rect 35016 23904 35080 23908
rect 35096 23964 35160 23968
rect 35096 23908 35100 23964
rect 35100 23908 35156 23964
rect 35156 23908 35160 23964
rect 35096 23904 35160 23908
rect 35176 23964 35240 23968
rect 35176 23908 35180 23964
rect 35180 23908 35236 23964
rect 35236 23908 35240 23964
rect 35176 23904 35240 23908
rect 19576 23420 19640 23424
rect 19576 23364 19580 23420
rect 19580 23364 19636 23420
rect 19636 23364 19640 23420
rect 19576 23360 19640 23364
rect 19656 23420 19720 23424
rect 19656 23364 19660 23420
rect 19660 23364 19716 23420
rect 19716 23364 19720 23420
rect 19656 23360 19720 23364
rect 19736 23420 19800 23424
rect 19736 23364 19740 23420
rect 19740 23364 19796 23420
rect 19796 23364 19800 23420
rect 19736 23360 19800 23364
rect 19816 23420 19880 23424
rect 19816 23364 19820 23420
rect 19820 23364 19876 23420
rect 19876 23364 19880 23420
rect 19816 23360 19880 23364
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 34936 22876 35000 22880
rect 34936 22820 34940 22876
rect 34940 22820 34996 22876
rect 34996 22820 35000 22876
rect 34936 22816 35000 22820
rect 35016 22876 35080 22880
rect 35016 22820 35020 22876
rect 35020 22820 35076 22876
rect 35076 22820 35080 22876
rect 35016 22816 35080 22820
rect 35096 22876 35160 22880
rect 35096 22820 35100 22876
rect 35100 22820 35156 22876
rect 35156 22820 35160 22876
rect 35096 22816 35160 22820
rect 35176 22876 35240 22880
rect 35176 22820 35180 22876
rect 35180 22820 35236 22876
rect 35236 22820 35240 22876
rect 35176 22816 35240 22820
rect 19576 22332 19640 22336
rect 19576 22276 19580 22332
rect 19580 22276 19636 22332
rect 19636 22276 19640 22332
rect 19576 22272 19640 22276
rect 19656 22332 19720 22336
rect 19656 22276 19660 22332
rect 19660 22276 19716 22332
rect 19716 22276 19720 22332
rect 19656 22272 19720 22276
rect 19736 22332 19800 22336
rect 19736 22276 19740 22332
rect 19740 22276 19796 22332
rect 19796 22276 19800 22332
rect 19736 22272 19800 22276
rect 19816 22332 19880 22336
rect 19816 22276 19820 22332
rect 19820 22276 19876 22332
rect 19876 22276 19880 22332
rect 19816 22272 19880 22276
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 34936 21788 35000 21792
rect 34936 21732 34940 21788
rect 34940 21732 34996 21788
rect 34996 21732 35000 21788
rect 34936 21728 35000 21732
rect 35016 21788 35080 21792
rect 35016 21732 35020 21788
rect 35020 21732 35076 21788
rect 35076 21732 35080 21788
rect 35016 21728 35080 21732
rect 35096 21788 35160 21792
rect 35096 21732 35100 21788
rect 35100 21732 35156 21788
rect 35156 21732 35160 21788
rect 35096 21728 35160 21732
rect 35176 21788 35240 21792
rect 35176 21732 35180 21788
rect 35180 21732 35236 21788
rect 35236 21732 35240 21788
rect 35176 21728 35240 21732
rect 19576 21244 19640 21248
rect 19576 21188 19580 21244
rect 19580 21188 19636 21244
rect 19636 21188 19640 21244
rect 19576 21184 19640 21188
rect 19656 21244 19720 21248
rect 19656 21188 19660 21244
rect 19660 21188 19716 21244
rect 19716 21188 19720 21244
rect 19656 21184 19720 21188
rect 19736 21244 19800 21248
rect 19736 21188 19740 21244
rect 19740 21188 19796 21244
rect 19796 21188 19800 21244
rect 19736 21184 19800 21188
rect 19816 21244 19880 21248
rect 19816 21188 19820 21244
rect 19820 21188 19876 21244
rect 19876 21188 19880 21244
rect 19816 21184 19880 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 34936 20700 35000 20704
rect 34936 20644 34940 20700
rect 34940 20644 34996 20700
rect 34996 20644 35000 20700
rect 34936 20640 35000 20644
rect 35016 20700 35080 20704
rect 35016 20644 35020 20700
rect 35020 20644 35076 20700
rect 35076 20644 35080 20700
rect 35016 20640 35080 20644
rect 35096 20700 35160 20704
rect 35096 20644 35100 20700
rect 35100 20644 35156 20700
rect 35156 20644 35160 20700
rect 35096 20640 35160 20644
rect 35176 20700 35240 20704
rect 35176 20644 35180 20700
rect 35180 20644 35236 20700
rect 35236 20644 35240 20700
rect 35176 20640 35240 20644
rect 19576 20156 19640 20160
rect 19576 20100 19580 20156
rect 19580 20100 19636 20156
rect 19636 20100 19640 20156
rect 19576 20096 19640 20100
rect 19656 20156 19720 20160
rect 19656 20100 19660 20156
rect 19660 20100 19716 20156
rect 19716 20100 19720 20156
rect 19656 20096 19720 20100
rect 19736 20156 19800 20160
rect 19736 20100 19740 20156
rect 19740 20100 19796 20156
rect 19796 20100 19800 20156
rect 19736 20096 19800 20100
rect 19816 20156 19880 20160
rect 19816 20100 19820 20156
rect 19820 20100 19876 20156
rect 19876 20100 19880 20156
rect 19816 20096 19880 20100
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 34936 19612 35000 19616
rect 34936 19556 34940 19612
rect 34940 19556 34996 19612
rect 34996 19556 35000 19612
rect 34936 19552 35000 19556
rect 35016 19612 35080 19616
rect 35016 19556 35020 19612
rect 35020 19556 35076 19612
rect 35076 19556 35080 19612
rect 35016 19552 35080 19556
rect 35096 19612 35160 19616
rect 35096 19556 35100 19612
rect 35100 19556 35156 19612
rect 35156 19556 35160 19612
rect 35096 19552 35160 19556
rect 35176 19612 35240 19616
rect 35176 19556 35180 19612
rect 35180 19556 35236 19612
rect 35236 19556 35240 19612
rect 35176 19552 35240 19556
rect 19576 19068 19640 19072
rect 19576 19012 19580 19068
rect 19580 19012 19636 19068
rect 19636 19012 19640 19068
rect 19576 19008 19640 19012
rect 19656 19068 19720 19072
rect 19656 19012 19660 19068
rect 19660 19012 19716 19068
rect 19716 19012 19720 19068
rect 19656 19008 19720 19012
rect 19736 19068 19800 19072
rect 19736 19012 19740 19068
rect 19740 19012 19796 19068
rect 19796 19012 19800 19068
rect 19736 19008 19800 19012
rect 19816 19068 19880 19072
rect 19816 19012 19820 19068
rect 19820 19012 19876 19068
rect 19876 19012 19880 19068
rect 19816 19008 19880 19012
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 34936 18524 35000 18528
rect 34936 18468 34940 18524
rect 34940 18468 34996 18524
rect 34996 18468 35000 18524
rect 34936 18464 35000 18468
rect 35016 18524 35080 18528
rect 35016 18468 35020 18524
rect 35020 18468 35076 18524
rect 35076 18468 35080 18524
rect 35016 18464 35080 18468
rect 35096 18524 35160 18528
rect 35096 18468 35100 18524
rect 35100 18468 35156 18524
rect 35156 18468 35160 18524
rect 35096 18464 35160 18468
rect 35176 18524 35240 18528
rect 35176 18468 35180 18524
rect 35180 18468 35236 18524
rect 35236 18468 35240 18524
rect 35176 18464 35240 18468
rect 19576 17980 19640 17984
rect 19576 17924 19580 17980
rect 19580 17924 19636 17980
rect 19636 17924 19640 17980
rect 19576 17920 19640 17924
rect 19656 17980 19720 17984
rect 19656 17924 19660 17980
rect 19660 17924 19716 17980
rect 19716 17924 19720 17980
rect 19656 17920 19720 17924
rect 19736 17980 19800 17984
rect 19736 17924 19740 17980
rect 19740 17924 19796 17980
rect 19796 17924 19800 17980
rect 19736 17920 19800 17924
rect 19816 17980 19880 17984
rect 19816 17924 19820 17980
rect 19820 17924 19876 17980
rect 19876 17924 19880 17980
rect 19816 17920 19880 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 34936 17436 35000 17440
rect 34936 17380 34940 17436
rect 34940 17380 34996 17436
rect 34996 17380 35000 17436
rect 34936 17376 35000 17380
rect 35016 17436 35080 17440
rect 35016 17380 35020 17436
rect 35020 17380 35076 17436
rect 35076 17380 35080 17436
rect 35016 17376 35080 17380
rect 35096 17436 35160 17440
rect 35096 17380 35100 17436
rect 35100 17380 35156 17436
rect 35156 17380 35160 17436
rect 35096 17376 35160 17380
rect 35176 17436 35240 17440
rect 35176 17380 35180 17436
rect 35180 17380 35236 17436
rect 35236 17380 35240 17436
rect 35176 17376 35240 17380
rect 19576 16892 19640 16896
rect 19576 16836 19580 16892
rect 19580 16836 19636 16892
rect 19636 16836 19640 16892
rect 19576 16832 19640 16836
rect 19656 16892 19720 16896
rect 19656 16836 19660 16892
rect 19660 16836 19716 16892
rect 19716 16836 19720 16892
rect 19656 16832 19720 16836
rect 19736 16892 19800 16896
rect 19736 16836 19740 16892
rect 19740 16836 19796 16892
rect 19796 16836 19800 16892
rect 19736 16832 19800 16836
rect 19816 16892 19880 16896
rect 19816 16836 19820 16892
rect 19820 16836 19876 16892
rect 19876 16836 19880 16892
rect 19816 16832 19880 16836
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 34936 16348 35000 16352
rect 34936 16292 34940 16348
rect 34940 16292 34996 16348
rect 34996 16292 35000 16348
rect 34936 16288 35000 16292
rect 35016 16348 35080 16352
rect 35016 16292 35020 16348
rect 35020 16292 35076 16348
rect 35076 16292 35080 16348
rect 35016 16288 35080 16292
rect 35096 16348 35160 16352
rect 35096 16292 35100 16348
rect 35100 16292 35156 16348
rect 35156 16292 35160 16348
rect 35096 16288 35160 16292
rect 35176 16348 35240 16352
rect 35176 16292 35180 16348
rect 35180 16292 35236 16348
rect 35236 16292 35240 16348
rect 35176 16288 35240 16292
rect 19576 15804 19640 15808
rect 19576 15748 19580 15804
rect 19580 15748 19636 15804
rect 19636 15748 19640 15804
rect 19576 15744 19640 15748
rect 19656 15804 19720 15808
rect 19656 15748 19660 15804
rect 19660 15748 19716 15804
rect 19716 15748 19720 15804
rect 19656 15744 19720 15748
rect 19736 15804 19800 15808
rect 19736 15748 19740 15804
rect 19740 15748 19796 15804
rect 19796 15748 19800 15804
rect 19736 15744 19800 15748
rect 19816 15804 19880 15808
rect 19816 15748 19820 15804
rect 19820 15748 19876 15804
rect 19876 15748 19880 15804
rect 19816 15744 19880 15748
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 34936 15260 35000 15264
rect 34936 15204 34940 15260
rect 34940 15204 34996 15260
rect 34996 15204 35000 15260
rect 34936 15200 35000 15204
rect 35016 15260 35080 15264
rect 35016 15204 35020 15260
rect 35020 15204 35076 15260
rect 35076 15204 35080 15260
rect 35016 15200 35080 15204
rect 35096 15260 35160 15264
rect 35096 15204 35100 15260
rect 35100 15204 35156 15260
rect 35156 15204 35160 15260
rect 35096 15200 35160 15204
rect 35176 15260 35240 15264
rect 35176 15204 35180 15260
rect 35180 15204 35236 15260
rect 35236 15204 35240 15260
rect 35176 15200 35240 15204
rect 19576 14716 19640 14720
rect 19576 14660 19580 14716
rect 19580 14660 19636 14716
rect 19636 14660 19640 14716
rect 19576 14656 19640 14660
rect 19656 14716 19720 14720
rect 19656 14660 19660 14716
rect 19660 14660 19716 14716
rect 19716 14660 19720 14716
rect 19656 14656 19720 14660
rect 19736 14716 19800 14720
rect 19736 14660 19740 14716
rect 19740 14660 19796 14716
rect 19796 14660 19800 14716
rect 19736 14656 19800 14660
rect 19816 14716 19880 14720
rect 19816 14660 19820 14716
rect 19820 14660 19876 14716
rect 19876 14660 19880 14716
rect 19816 14656 19880 14660
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 34936 14172 35000 14176
rect 34936 14116 34940 14172
rect 34940 14116 34996 14172
rect 34996 14116 35000 14172
rect 34936 14112 35000 14116
rect 35016 14172 35080 14176
rect 35016 14116 35020 14172
rect 35020 14116 35076 14172
rect 35076 14116 35080 14172
rect 35016 14112 35080 14116
rect 35096 14172 35160 14176
rect 35096 14116 35100 14172
rect 35100 14116 35156 14172
rect 35156 14116 35160 14172
rect 35096 14112 35160 14116
rect 35176 14172 35240 14176
rect 35176 14116 35180 14172
rect 35180 14116 35236 14172
rect 35236 14116 35240 14172
rect 35176 14112 35240 14116
rect 19576 13628 19640 13632
rect 19576 13572 19580 13628
rect 19580 13572 19636 13628
rect 19636 13572 19640 13628
rect 19576 13568 19640 13572
rect 19656 13628 19720 13632
rect 19656 13572 19660 13628
rect 19660 13572 19716 13628
rect 19716 13572 19720 13628
rect 19656 13568 19720 13572
rect 19736 13628 19800 13632
rect 19736 13572 19740 13628
rect 19740 13572 19796 13628
rect 19796 13572 19800 13628
rect 19736 13568 19800 13572
rect 19816 13628 19880 13632
rect 19816 13572 19820 13628
rect 19820 13572 19876 13628
rect 19876 13572 19880 13628
rect 19816 13568 19880 13572
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 34936 13084 35000 13088
rect 34936 13028 34940 13084
rect 34940 13028 34996 13084
rect 34996 13028 35000 13084
rect 34936 13024 35000 13028
rect 35016 13084 35080 13088
rect 35016 13028 35020 13084
rect 35020 13028 35076 13084
rect 35076 13028 35080 13084
rect 35016 13024 35080 13028
rect 35096 13084 35160 13088
rect 35096 13028 35100 13084
rect 35100 13028 35156 13084
rect 35156 13028 35160 13084
rect 35096 13024 35160 13028
rect 35176 13084 35240 13088
rect 35176 13028 35180 13084
rect 35180 13028 35236 13084
rect 35236 13028 35240 13084
rect 35176 13024 35240 13028
rect 30972 12608 31036 12612
rect 30972 12552 31022 12608
rect 31022 12552 31036 12608
rect 30972 12548 31036 12552
rect 19576 12540 19640 12544
rect 19576 12484 19580 12540
rect 19580 12484 19636 12540
rect 19636 12484 19640 12540
rect 19576 12480 19640 12484
rect 19656 12540 19720 12544
rect 19656 12484 19660 12540
rect 19660 12484 19716 12540
rect 19716 12484 19720 12540
rect 19656 12480 19720 12484
rect 19736 12540 19800 12544
rect 19736 12484 19740 12540
rect 19740 12484 19796 12540
rect 19796 12484 19800 12540
rect 19736 12480 19800 12484
rect 19816 12540 19880 12544
rect 19816 12484 19820 12540
rect 19820 12484 19876 12540
rect 19876 12484 19880 12540
rect 19816 12480 19880 12484
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 34936 11996 35000 12000
rect 34936 11940 34940 11996
rect 34940 11940 34996 11996
rect 34996 11940 35000 11996
rect 34936 11936 35000 11940
rect 35016 11996 35080 12000
rect 35016 11940 35020 11996
rect 35020 11940 35076 11996
rect 35076 11940 35080 11996
rect 35016 11936 35080 11940
rect 35096 11996 35160 12000
rect 35096 11940 35100 11996
rect 35100 11940 35156 11996
rect 35156 11940 35160 11996
rect 35096 11936 35160 11940
rect 35176 11996 35240 12000
rect 35176 11940 35180 11996
rect 35180 11940 35236 11996
rect 35236 11940 35240 11996
rect 35176 11936 35240 11940
rect 19576 11452 19640 11456
rect 19576 11396 19580 11452
rect 19580 11396 19636 11452
rect 19636 11396 19640 11452
rect 19576 11392 19640 11396
rect 19656 11452 19720 11456
rect 19656 11396 19660 11452
rect 19660 11396 19716 11452
rect 19716 11396 19720 11452
rect 19656 11392 19720 11396
rect 19736 11452 19800 11456
rect 19736 11396 19740 11452
rect 19740 11396 19796 11452
rect 19796 11396 19800 11452
rect 19736 11392 19800 11396
rect 19816 11452 19880 11456
rect 19816 11396 19820 11452
rect 19820 11396 19876 11452
rect 19876 11396 19880 11452
rect 19816 11392 19880 11396
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 34936 10908 35000 10912
rect 34936 10852 34940 10908
rect 34940 10852 34996 10908
rect 34996 10852 35000 10908
rect 34936 10848 35000 10852
rect 35016 10908 35080 10912
rect 35016 10852 35020 10908
rect 35020 10852 35076 10908
rect 35076 10852 35080 10908
rect 35016 10848 35080 10852
rect 35096 10908 35160 10912
rect 35096 10852 35100 10908
rect 35100 10852 35156 10908
rect 35156 10852 35160 10908
rect 35096 10848 35160 10852
rect 35176 10908 35240 10912
rect 35176 10852 35180 10908
rect 35180 10852 35236 10908
rect 35236 10852 35240 10908
rect 35176 10848 35240 10852
rect 19576 10364 19640 10368
rect 19576 10308 19580 10364
rect 19580 10308 19636 10364
rect 19636 10308 19640 10364
rect 19576 10304 19640 10308
rect 19656 10364 19720 10368
rect 19656 10308 19660 10364
rect 19660 10308 19716 10364
rect 19716 10308 19720 10364
rect 19656 10304 19720 10308
rect 19736 10364 19800 10368
rect 19736 10308 19740 10364
rect 19740 10308 19796 10364
rect 19796 10308 19800 10364
rect 19736 10304 19800 10308
rect 19816 10364 19880 10368
rect 19816 10308 19820 10364
rect 19820 10308 19876 10364
rect 19876 10308 19880 10364
rect 19816 10304 19880 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 34936 9820 35000 9824
rect 34936 9764 34940 9820
rect 34940 9764 34996 9820
rect 34996 9764 35000 9820
rect 34936 9760 35000 9764
rect 35016 9820 35080 9824
rect 35016 9764 35020 9820
rect 35020 9764 35076 9820
rect 35076 9764 35080 9820
rect 35016 9760 35080 9764
rect 35096 9820 35160 9824
rect 35096 9764 35100 9820
rect 35100 9764 35156 9820
rect 35156 9764 35160 9820
rect 35096 9760 35160 9764
rect 35176 9820 35240 9824
rect 35176 9764 35180 9820
rect 35180 9764 35236 9820
rect 35236 9764 35240 9820
rect 35176 9760 35240 9764
rect 19576 9276 19640 9280
rect 19576 9220 19580 9276
rect 19580 9220 19636 9276
rect 19636 9220 19640 9276
rect 19576 9216 19640 9220
rect 19656 9276 19720 9280
rect 19656 9220 19660 9276
rect 19660 9220 19716 9276
rect 19716 9220 19720 9276
rect 19656 9216 19720 9220
rect 19736 9276 19800 9280
rect 19736 9220 19740 9276
rect 19740 9220 19796 9276
rect 19796 9220 19800 9276
rect 19736 9216 19800 9220
rect 19816 9276 19880 9280
rect 19816 9220 19820 9276
rect 19820 9220 19876 9276
rect 19876 9220 19880 9276
rect 19816 9216 19880 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 34936 8732 35000 8736
rect 34936 8676 34940 8732
rect 34940 8676 34996 8732
rect 34996 8676 35000 8732
rect 34936 8672 35000 8676
rect 35016 8732 35080 8736
rect 35016 8676 35020 8732
rect 35020 8676 35076 8732
rect 35076 8676 35080 8732
rect 35016 8672 35080 8676
rect 35096 8732 35160 8736
rect 35096 8676 35100 8732
rect 35100 8676 35156 8732
rect 35156 8676 35160 8732
rect 35096 8672 35160 8676
rect 35176 8732 35240 8736
rect 35176 8676 35180 8732
rect 35180 8676 35236 8732
rect 35236 8676 35240 8732
rect 35176 8672 35240 8676
rect 19576 8188 19640 8192
rect 19576 8132 19580 8188
rect 19580 8132 19636 8188
rect 19636 8132 19640 8188
rect 19576 8128 19640 8132
rect 19656 8188 19720 8192
rect 19656 8132 19660 8188
rect 19660 8132 19716 8188
rect 19716 8132 19720 8188
rect 19656 8128 19720 8132
rect 19736 8188 19800 8192
rect 19736 8132 19740 8188
rect 19740 8132 19796 8188
rect 19796 8132 19800 8188
rect 19736 8128 19800 8132
rect 19816 8188 19880 8192
rect 19816 8132 19820 8188
rect 19820 8132 19876 8188
rect 19876 8132 19880 8188
rect 19816 8128 19880 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 34936 7644 35000 7648
rect 34936 7588 34940 7644
rect 34940 7588 34996 7644
rect 34996 7588 35000 7644
rect 34936 7584 35000 7588
rect 35016 7644 35080 7648
rect 35016 7588 35020 7644
rect 35020 7588 35076 7644
rect 35076 7588 35080 7644
rect 35016 7584 35080 7588
rect 35096 7644 35160 7648
rect 35096 7588 35100 7644
rect 35100 7588 35156 7644
rect 35156 7588 35160 7644
rect 35096 7584 35160 7588
rect 35176 7644 35240 7648
rect 35176 7588 35180 7644
rect 35180 7588 35236 7644
rect 35236 7588 35240 7644
rect 35176 7584 35240 7588
rect 19576 7100 19640 7104
rect 19576 7044 19580 7100
rect 19580 7044 19636 7100
rect 19636 7044 19640 7100
rect 19576 7040 19640 7044
rect 19656 7100 19720 7104
rect 19656 7044 19660 7100
rect 19660 7044 19716 7100
rect 19716 7044 19720 7100
rect 19656 7040 19720 7044
rect 19736 7100 19800 7104
rect 19736 7044 19740 7100
rect 19740 7044 19796 7100
rect 19796 7044 19800 7100
rect 19736 7040 19800 7044
rect 19816 7100 19880 7104
rect 19816 7044 19820 7100
rect 19820 7044 19876 7100
rect 19876 7044 19880 7100
rect 19816 7040 19880 7044
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 34936 6556 35000 6560
rect 34936 6500 34940 6556
rect 34940 6500 34996 6556
rect 34996 6500 35000 6556
rect 34936 6496 35000 6500
rect 35016 6556 35080 6560
rect 35016 6500 35020 6556
rect 35020 6500 35076 6556
rect 35076 6500 35080 6556
rect 35016 6496 35080 6500
rect 35096 6556 35160 6560
rect 35096 6500 35100 6556
rect 35100 6500 35156 6556
rect 35156 6500 35160 6556
rect 35096 6496 35160 6500
rect 35176 6556 35240 6560
rect 35176 6500 35180 6556
rect 35180 6500 35236 6556
rect 35236 6500 35240 6556
rect 35176 6496 35240 6500
rect 19576 6012 19640 6016
rect 19576 5956 19580 6012
rect 19580 5956 19636 6012
rect 19636 5956 19640 6012
rect 19576 5952 19640 5956
rect 19656 6012 19720 6016
rect 19656 5956 19660 6012
rect 19660 5956 19716 6012
rect 19716 5956 19720 6012
rect 19656 5952 19720 5956
rect 19736 6012 19800 6016
rect 19736 5956 19740 6012
rect 19740 5956 19796 6012
rect 19796 5956 19800 6012
rect 19736 5952 19800 5956
rect 19816 6012 19880 6016
rect 19816 5956 19820 6012
rect 19820 5956 19876 6012
rect 19876 5956 19880 6012
rect 19816 5952 19880 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 34936 5468 35000 5472
rect 34936 5412 34940 5468
rect 34940 5412 34996 5468
rect 34996 5412 35000 5468
rect 34936 5408 35000 5412
rect 35016 5468 35080 5472
rect 35016 5412 35020 5468
rect 35020 5412 35076 5468
rect 35076 5412 35080 5468
rect 35016 5408 35080 5412
rect 35096 5468 35160 5472
rect 35096 5412 35100 5468
rect 35100 5412 35156 5468
rect 35156 5412 35160 5468
rect 35096 5408 35160 5412
rect 35176 5468 35240 5472
rect 35176 5412 35180 5468
rect 35180 5412 35236 5468
rect 35236 5412 35240 5468
rect 35176 5408 35240 5412
rect 19576 4924 19640 4928
rect 19576 4868 19580 4924
rect 19580 4868 19636 4924
rect 19636 4868 19640 4924
rect 19576 4864 19640 4868
rect 19656 4924 19720 4928
rect 19656 4868 19660 4924
rect 19660 4868 19716 4924
rect 19716 4868 19720 4924
rect 19656 4864 19720 4868
rect 19736 4924 19800 4928
rect 19736 4868 19740 4924
rect 19740 4868 19796 4924
rect 19796 4868 19800 4924
rect 19736 4864 19800 4868
rect 19816 4924 19880 4928
rect 19816 4868 19820 4924
rect 19820 4868 19876 4924
rect 19876 4868 19880 4924
rect 19816 4864 19880 4868
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 34936 4380 35000 4384
rect 34936 4324 34940 4380
rect 34940 4324 34996 4380
rect 34996 4324 35000 4380
rect 34936 4320 35000 4324
rect 35016 4380 35080 4384
rect 35016 4324 35020 4380
rect 35020 4324 35076 4380
rect 35076 4324 35080 4380
rect 35016 4320 35080 4324
rect 35096 4380 35160 4384
rect 35096 4324 35100 4380
rect 35100 4324 35156 4380
rect 35156 4324 35160 4380
rect 35096 4320 35160 4324
rect 35176 4380 35240 4384
rect 35176 4324 35180 4380
rect 35180 4324 35236 4380
rect 35236 4324 35240 4380
rect 35176 4320 35240 4324
rect 19576 3836 19640 3840
rect 19576 3780 19580 3836
rect 19580 3780 19636 3836
rect 19636 3780 19640 3836
rect 19576 3776 19640 3780
rect 19656 3836 19720 3840
rect 19656 3780 19660 3836
rect 19660 3780 19716 3836
rect 19716 3780 19720 3836
rect 19656 3776 19720 3780
rect 19736 3836 19800 3840
rect 19736 3780 19740 3836
rect 19740 3780 19796 3836
rect 19796 3780 19800 3836
rect 19736 3776 19800 3780
rect 19816 3836 19880 3840
rect 19816 3780 19820 3836
rect 19820 3780 19876 3836
rect 19876 3780 19880 3836
rect 19816 3776 19880 3780
rect 30420 3768 30484 3772
rect 30420 3712 30434 3768
rect 30434 3712 30484 3768
rect 30420 3708 30484 3712
rect 20852 3436 20916 3500
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 34936 3292 35000 3296
rect 34936 3236 34940 3292
rect 34940 3236 34996 3292
rect 34996 3236 35000 3292
rect 34936 3232 35000 3236
rect 35016 3292 35080 3296
rect 35016 3236 35020 3292
rect 35020 3236 35076 3292
rect 35076 3236 35080 3292
rect 35016 3232 35080 3236
rect 35096 3292 35160 3296
rect 35096 3236 35100 3292
rect 35100 3236 35156 3292
rect 35156 3236 35160 3292
rect 35096 3232 35160 3236
rect 35176 3292 35240 3296
rect 35176 3236 35180 3292
rect 35180 3236 35236 3292
rect 35236 3236 35240 3292
rect 35176 3232 35240 3236
rect 796 3028 860 3092
rect 19576 2748 19640 2752
rect 19576 2692 19580 2748
rect 19580 2692 19636 2748
rect 19636 2692 19640 2748
rect 19576 2688 19640 2692
rect 19656 2748 19720 2752
rect 19656 2692 19660 2748
rect 19660 2692 19716 2748
rect 19716 2692 19720 2748
rect 19656 2688 19720 2692
rect 19736 2748 19800 2752
rect 19736 2692 19740 2748
rect 19740 2692 19796 2748
rect 19796 2692 19800 2748
rect 19736 2688 19800 2692
rect 19816 2748 19880 2752
rect 19816 2692 19820 2748
rect 19820 2692 19876 2748
rect 19876 2692 19880 2748
rect 19816 2688 19880 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
rect 34936 2204 35000 2208
rect 34936 2148 34940 2204
rect 34940 2148 34996 2204
rect 34996 2148 35000 2204
rect 34936 2144 35000 2148
rect 35016 2204 35080 2208
rect 35016 2148 35020 2204
rect 35020 2148 35076 2204
rect 35076 2148 35080 2204
rect 35016 2144 35080 2148
rect 35096 2204 35160 2208
rect 35096 2148 35100 2204
rect 35100 2148 35156 2204
rect 35156 2148 35160 2204
rect 35096 2144 35160 2148
rect 35176 2204 35240 2208
rect 35176 2148 35180 2204
rect 35180 2148 35236 2204
rect 35236 2148 35240 2204
rect 35176 2144 35240 2148
<< metal4 >>
rect 4208 46816 4528 47376
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 45728 4528 46752
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 44640 4528 45664
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 43552 4528 44576
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 42464 4528 43488
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 41376 4528 42400
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 40288 4528 41312
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 39200 4528 40224
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 38112 4528 39136
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 37024 4528 38048
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 35936 4528 36960
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5472 4528 6496
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 4384 4528 5408
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2128 4528 2144
rect 19568 47360 19888 47376
rect 19568 47296 19576 47360
rect 19640 47296 19656 47360
rect 19720 47296 19736 47360
rect 19800 47296 19816 47360
rect 19880 47296 19888 47360
rect 19568 46272 19888 47296
rect 19568 46208 19576 46272
rect 19640 46208 19656 46272
rect 19720 46208 19736 46272
rect 19800 46208 19816 46272
rect 19880 46208 19888 46272
rect 19568 45184 19888 46208
rect 19568 45120 19576 45184
rect 19640 45120 19656 45184
rect 19720 45120 19736 45184
rect 19800 45120 19816 45184
rect 19880 45120 19888 45184
rect 19568 44096 19888 45120
rect 19568 44032 19576 44096
rect 19640 44032 19656 44096
rect 19720 44032 19736 44096
rect 19800 44032 19816 44096
rect 19880 44032 19888 44096
rect 19568 43008 19888 44032
rect 19568 42944 19576 43008
rect 19640 42944 19656 43008
rect 19720 42944 19736 43008
rect 19800 42944 19816 43008
rect 19880 42944 19888 43008
rect 19568 41920 19888 42944
rect 19568 41856 19576 41920
rect 19640 41856 19656 41920
rect 19720 41856 19736 41920
rect 19800 41856 19816 41920
rect 19880 41856 19888 41920
rect 19568 40832 19888 41856
rect 19568 40768 19576 40832
rect 19640 40768 19656 40832
rect 19720 40768 19736 40832
rect 19800 40768 19816 40832
rect 19880 40768 19888 40832
rect 19568 39744 19888 40768
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 19568 38656 19888 39680
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 37568 19888 38592
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 36480 19888 37504
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 35392 19888 36416
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 34304 19888 35328
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 33216 19888 34240
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 32128 19888 33152
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 31040 19888 32064
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 29952 19888 30976
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 28864 19888 29888
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 27776 19888 28800
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 26688 19888 27712
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 25600 19888 26624
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 24512 19888 25536
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 23424 19888 24448
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 22336 19888 23360
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 21248 19888 22272
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 20160 19888 21184
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 19072 19888 20096
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 17984 19888 19008
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 16896 19888 17920
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 15808 19888 16832
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 14720 19888 15744
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 13632 19888 14656
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 12544 19888 13568
rect 34928 46816 35248 47376
rect 34928 46752 34936 46816
rect 35000 46752 35016 46816
rect 35080 46752 35096 46816
rect 35160 46752 35176 46816
rect 35240 46752 35248 46816
rect 34928 45728 35248 46752
rect 34928 45664 34936 45728
rect 35000 45664 35016 45728
rect 35080 45664 35096 45728
rect 35160 45664 35176 45728
rect 35240 45664 35248 45728
rect 34928 44640 35248 45664
rect 34928 44576 34936 44640
rect 35000 44576 35016 44640
rect 35080 44576 35096 44640
rect 35160 44576 35176 44640
rect 35240 44576 35248 44640
rect 34928 43552 35248 44576
rect 34928 43488 34936 43552
rect 35000 43488 35016 43552
rect 35080 43488 35096 43552
rect 35160 43488 35176 43552
rect 35240 43488 35248 43552
rect 34928 42464 35248 43488
rect 34928 42400 34936 42464
rect 35000 42400 35016 42464
rect 35080 42400 35096 42464
rect 35160 42400 35176 42464
rect 35240 42400 35248 42464
rect 34928 41376 35248 42400
rect 34928 41312 34936 41376
rect 35000 41312 35016 41376
rect 35080 41312 35096 41376
rect 35160 41312 35176 41376
rect 35240 41312 35248 41376
rect 34928 40288 35248 41312
rect 34928 40224 34936 40288
rect 35000 40224 35016 40288
rect 35080 40224 35096 40288
rect 35160 40224 35176 40288
rect 35240 40224 35248 40288
rect 34928 39200 35248 40224
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 38112 35248 39136
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 37024 35248 38048
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 35936 35248 36960
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 34848 35248 35872
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 33760 35248 34784
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 32672 35248 33696
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 31584 35248 32608
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 30496 35248 31520
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 29408 35248 30432
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 28320 35248 29344
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 27232 35248 28256
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 26144 35248 27168
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 25056 35248 26080
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 23968 35248 24992
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 22880 35248 23904
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 21792 35248 22816
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 20704 35248 21728
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 19616 35248 20640
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 18528 35248 19552
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 17440 35248 18464
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 16352 35248 17376
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 15264 35248 16288
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 14176 35248 15200
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 13088 35248 14112
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 30971 12612 31037 12613
rect 30971 12548 30972 12612
rect 31036 12548 31037 12612
rect 30971 12547 31037 12548
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 11456 19888 12480
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 10368 19888 11392
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 9280 19888 10304
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 8192 19888 9216
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 7104 19888 8128
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 6016 19888 7040
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 4928 19888 5952
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 3840 19888 4864
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 2752 19888 3776
rect 20854 3501 20914 3622
rect 20851 3500 20917 3501
rect 20851 3436 20852 3500
rect 20916 3436 20917 3500
rect 20851 3435 20917 3436
rect 30974 3178 31034 12547
rect 34928 12000 35248 13024
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 10912 35248 11936
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 9824 35248 10848
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 8736 35248 9760
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 7648 35248 8672
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 6560 35248 7584
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 5472 35248 6496
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 4384 35248 5408
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 3296 35248 4320
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2128 19888 2688
rect 34928 2208 35248 3232
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2128 35248 2144
<< via4 >>
rect 710 3092 946 3178
rect 710 3028 796 3092
rect 796 3028 860 3092
rect 860 3028 946 3092
rect 710 2942 946 3028
rect 20766 3622 21002 3858
rect 30334 3772 30570 3858
rect 30334 3708 30420 3772
rect 30420 3708 30484 3772
rect 30484 3708 30570 3772
rect 30334 3622 30570 3708
rect 30886 2942 31122 3178
<< metal5 >>
rect 20724 3858 30612 3900
rect 20724 3622 20766 3858
rect 21002 3622 30334 3858
rect 30570 3622 30612 3858
rect 20724 3580 30612 3622
rect 668 3178 31164 3220
rect 668 2942 710 3178
rect 946 2942 30886 3178
rect 31122 2942 31164 3178
rect 668 2900 31164 2942
use scs8hd_fill_1  FILLER_1_11 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2116 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_7 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_3
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2208 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
timestamp 1586364061
transform 1 0 1564 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_14
timestamp 1586364061
transform 1 0 2392 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
timestamp 1586364061
transform 1 0 2576 0 1 2720
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2760 0 1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
timestamp 1586364061
transform 1 0 1472 0 -1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_1_37
timestamp 1586364061
transform 1 0 4508 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_166 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_45
timestamp 1586364061
transform 1 0 5244 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_41
timestamp 1586364061
transform 1 0 4876 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1586364061
transform 1 0 5428 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 5060 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5612 0 1 2720
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
timestamp 1586364061
transform 1 0 4324 0 -1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_71
timestamp 1586364061
transform 1 0 7636 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_67
timestamp 1586364061
transform 1 0 7268 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
timestamp 1586364061
transform 1 0 7820 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
timestamp 1586364061
transform 1 0 7176 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 7452 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
timestamp 1586364061
transform 1 0 7360 0 1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_0_84
timestamp 1586364061
transform 1 0 8832 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1586364061
transform 1 0 9016 0 -1 2720
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_91
timestamp 1586364061
transform 1 0 9476 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_87
timestamp 1586364061
transform 1 0 9108 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_88
timestamp 1586364061
transform 1 0 9200 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
timestamp 1586364061
transform 1 0 9292 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
timestamp 1586364061
transform 1 0 9660 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
timestamp 1586364061
transform 1 0 9844 0 1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
timestamp 1586364061
transform 1 0 11684 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_113
timestamp 1586364061
transform 1 0 11500 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_117
timestamp 1586364061
transform 1 0 11868 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_121
timestamp 1586364061
transform 1 0 12236 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_0_130
timestamp 1586364061
transform 1 0 13064 0 -1 2720
box -38 -48 222 592
use scs8hd_or2_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 498 592
use scs8hd_decap_6  FILLER_0_134 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
timestamp 1586364061
transform 1 0 13248 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_142
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_140
timestamp 1586364061
transform 1 0 13984 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
timestamp 1586364061
transform 1 0 14076 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 14260 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_1_146
timestamp 1586364061
transform 1 0 14536 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
timestamp 1586364061
transform 1 0 14812 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
timestamp 1586364061
transform 1 0 14996 0 1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
timestamp 1586364061
transform 1 0 15732 0 -1 2720
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 16928 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_170
timestamp 1586364061
transform 1 0 16744 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_178
timestamp 1586364061
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_174
timestamp 1586364061
transform 1 0 17112 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use scs8hd_decap_4  FILLER_1_197
timestamp 1586364061
transform 1 0 19228 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_193
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
timestamp 1586364061
transform 1 0 18584 0 -1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_0_209
timestamp 1586364061
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_222
timestamp 1586364061
transform 1 0 21528 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 21436 0 -1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
timestamp 1586364061
transform 1 0 19780 0 1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_1_235
timestamp 1586364061
transform 1 0 22724 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_226
timestamp 1586364061
transform 1 0 21896 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 21712 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
timestamp 1586364061
transform 1 0 22080 0 1 2720
box -38 -48 222 592
use scs8hd_or2_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
timestamp 1586364061
transform 1 0 22264 0 1 2720
box -38 -48 498 592
use scs8hd_decap_3  FILLER_1_239
timestamp 1586364061
transform 1 0 23092 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_244
timestamp 1586364061
transform 1 0 23552 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_240
timestamp 1586364061
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
timestamp 1586364061
transform 1 0 22908 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1786 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 26220 0 1 2720
box -38 -48 2246 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 24288 0 -1 2720
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 26036 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 25576 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_0_271
timestamp 1586364061
transform 1 0 26036 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_264
timestamp 1586364061
transform 1 0 25392 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_268
timestamp 1586364061
transform 1 0 25760 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_278
timestamp 1586364061
transform 1 0 26680 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_275
timestamp 1586364061
transform 1 0 26404 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 26496 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 26864 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_0_289
timestamp 1586364061
transform 1 0 27692 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 27876 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_297
timestamp 1586364061
transform 1 0 28428 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_293
timestamp 1586364061
transform 1 0 28060 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 28244 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _65_
timestamp 1586364061
transform 1 0 28428 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 28612 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_301
timestamp 1586364061
transform 1 0 28796 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_301
timestamp 1586364061
transform 1 0 28796 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__65__A
timestamp 1586364061
transform 1 0 28980 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 28980 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_305
timestamp 1586364061
transform 1 0 29164 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 29440 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 29532 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_306
timestamp 1586364061
transform 1 0 29256 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_311
timestamp 1586364061
transform 1 0 29716 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 29900 0 1 2720
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 30084 0 1 2720
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 29716 0 -1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_1_328
timestamp 1586364061
transform 1 0 31280 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_324
timestamp 1586364061
transform 1 0 30912 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_335
timestamp 1586364061
transform 1 0 31924 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_330
timestamp 1586364061
transform 1 0 31464 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 31464 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 31740 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__67__A
timestamp 1586364061
transform 1 0 31096 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_342
timestamp 1586364061
transform 1 0 32568 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_339
timestamp 1586364061
transform 1 0 32292 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 32108 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 32844 0 -1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 31648 0 1 2720
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_1_359
timestamp 1586364061
transform 1 0 34132 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_355
timestamp 1586364061
transform 1 0 33764 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_351
timestamp 1586364061
transform 1 0 33396 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 34224 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 33580 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_362
timestamp 1586364061
transform 1 0 34408 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_371
timestamp 1586364061
transform 1 0 35236 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_368
timestamp 1586364061
transform 1 0 34960 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_364
timestamp 1586364061
transform 1 0 34592 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 35052 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 34592 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 34868 0 1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_0_381
timestamp 1586364061
transform 1 0 36156 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_377
timestamp 1586364061
transform 1 0 35788 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 36340 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__68__A
timestamp 1586364061
transform 1 0 35972 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _68_
timestamp 1586364061
transform 1 0 35420 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_2  _69_
timestamp 1586364061
transform 1 0 36616 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 36800 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_385
timestamp 1586364061
transform 1 0 36524 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_386
timestamp 1586364061
transform 1 0 36616 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__69__A
timestamp 1586364061
transform 1 0 37168 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 37168 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_390
timestamp 1586364061
transform 1 0 36984 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_394
timestamp 1586364061
transform 1 0 37352 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_390
timestamp 1586364061
transform 1 0 36984 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 37628 0 -1 2720
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 37352 0 1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 38272 0 -1 2720
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 37996 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 39652 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 39284 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_399
timestamp 1586364061
transform 1 0 37812 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_413
timestamp 1586364061
transform 1 0 39100 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_417
timestamp 1586364061
transform 1 0 39468 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_421
timestamp 1586364061
transform 1 0 39836 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_430
timestamp 1586364061
transform 1 0 40664 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_427
timestamp 1586364061
transform 1 0 40388 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_423
timestamp 1586364061
transform 1 0 40020 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 40480 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 40204 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 40848 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 40388 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 41032 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_444
timestamp 1586364061
transform 1 0 41952 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 42136 0 -1 2720
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 41124 0 -1 2720
box -38 -48 866 592
use scs8hd_decap_12  FILLER_1_447 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 42228 0 1 2720
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 40480 0 1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_0_456
timestamp 1586364061
transform 1 0 43056 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_448
timestamp 1586364061
transform 1 0 42320 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__71__A
timestamp 1586364061
transform 1 0 43240 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _71_
timestamp 1586364061
transform 1 0 42688 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_0_466 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 43976 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_1  FILLER_0_464
timestamp 1586364061
transform 1 0 43792 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_460
timestamp 1586364061
transform 1 0 43424 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 43884 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_471
timestamp 1586364061
transform 1 0 44436 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_459
timestamp 1586364061
transform 1 0 43332 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_483
timestamp 1586364061
transform 1 0 45540 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_479
timestamp 1586364061
transform 1 0 45172 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_474
timestamp 1586364061
transform 1 0 44712 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__72__A
timestamp 1586364061
transform 1 0 45356 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _72_
timestamp 1586364061
transform 1 0 44804 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_487
timestamp 1586364061
transform 1 0 45908 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_495
timestamp 1586364061
transform 1 0 46644 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 46000 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 46736 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_489
timestamp 1586364061
transform 1 0 46092 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_483
timestamp 1586364061
transform 1 0 45540 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 48852 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 48852 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_497
timestamp 1586364061
transform 1 0 46828 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_509
timestamp 1586364061
transform 1 0 47932 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_0_515
timestamp 1586364061
transform 1 0 48484 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_501
timestamp 1586364061
transform 1 0 47196 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_1_513
timestamp 1586364061
transform 1 0 48300 0 1 2720
box -38 -48 314 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1586364061
transform 1 0 2392 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
timestamp 1586364061
transform 1 0 1564 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_7
timestamp 1586364061
transform 1 0 1748 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_11
timestamp 1586364061
transform 1 0 2116 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1586364061
transform 1 0 4600 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 5612 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 4416 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_47
timestamp 1586364061
transform 1 0 5428 0 -1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
timestamp 1586364061
transform 1 0 6164 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 5980 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_51
timestamp 1586364061
transform 1 0 5796 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_74
timestamp 1586364061
transform 1 0 7912 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 8096 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_78
timestamp 1586364061
transform 1 0 8280 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_82
timestamp 1586364061
transform 1 0 8648 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
timestamp 1586364061
transform 1 0 11316 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
timestamp 1586364061
transform 1 0 11132 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_102
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_106
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 314 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 13800 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 13248 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 13616 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_130
timestamp 1586364061
transform 1 0 13064 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_134
timestamp 1586364061
transform 1 0 13432 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_142
timestamp 1586364061
transform 1 0 14168 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_146
timestamp 1586364061
transform 1 0 14536 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_149
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1586364061
transform 1 0 15364 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
timestamp 1586364061
transform 1 0 16744 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_164
timestamp 1586364061
transform 1 0 16192 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_168
timestamp 1586364061
transform 1 0 16560 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_172
timestamp 1586364061
transform 1 0 16928 0 -1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
timestamp 1586364061
transform 1 0 17848 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 17664 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1586364061
transform 1 0 17112 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_176
timestamp 1586364061
transform 1 0 17296 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_201
timestamp 1586364061
transform 1 0 19596 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
timestamp 1586364061
transform 1 0 19780 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_205
timestamp 1586364061
transform 1 0 19964 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 20148 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_209
timestamp 1586364061
transform 1 0 20332 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_219
timestamp 1586364061
transform 1 0 21252 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 21436 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_223
timestamp 1586364061
transform 1 0 21620 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 866 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 23736 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 23552 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 23184 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 21804 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_236
timestamp 1586364061
transform 1 0 22816 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_242
timestamp 1586364061
transform 1 0 23368 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 26220 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 25852 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 24748 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 25116 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_255
timestamp 1586364061
transform 1 0 24564 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_259
timestamp 1586364061
transform 1 0 24932 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_267
timestamp 1586364061
transform 1 0 25668 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_271
timestamp 1586364061
transform 1 0 26036 0 -1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 28060 0 -1 3808
box -38 -48 1786 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 27600 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_285
timestamp 1586364061
transform 1 0 27324 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_2_290
timestamp 1586364061
transform 1 0 27784 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 30084 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 30452 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_312
timestamp 1586364061
transform 1 0 29808 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_317
timestamp 1586364061
transform 1 0 30268 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_321
timestamp 1586364061
transform 1 0 30636 0 -1 3808
box -38 -48 314 592
use scs8hd_buf_2  _67_
timestamp 1586364061
transform 1 0 30912 0 -1 3808
box -38 -48 406 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 32108 0 -1 3808
box -38 -48 2246 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 31832 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 31464 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_328
timestamp 1586364061
transform 1 0 31280 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_332
timestamp 1586364061
transform 1 0 31648 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 35052 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 34868 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 34500 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_361
timestamp 1586364061
transform 1 0 34316 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_365
timestamp 1586364061
transform 1 0 34684 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 37352 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 36984 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_378
timestamp 1586364061
transform 1 0 35880 0 -1 3808
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_2_392
timestamp 1586364061
transform 1 0 37168 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_396
timestamp 1586364061
transform 1 0 37536 0 -1 3808
box -38 -48 130 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 37720 0 -1 3808
box -38 -48 866 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 39652 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 39468 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 39100 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_407
timestamp 1586364061
transform 1 0 38548 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_2  FILLER_2_415
timestamp 1586364061
transform 1 0 39284 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _70_
timestamp 1586364061
transform 1 0 41216 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__70__A
timestamp 1586364061
transform 1 0 41768 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 40664 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 41032 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_428
timestamp 1586364061
transform 1 0 40480 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_432
timestamp 1586364061
transform 1 0 40848 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_440
timestamp 1586364061
transform 1 0 41584 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_444
timestamp 1586364061
transform 1 0 41952 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 43240 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_456
timestamp 1586364061
transform 1 0 43056 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_459
timestamp 1586364061
transform 1 0 43332 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_471
timestamp 1586364061
transform 1 0 44436 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_483
timestamp 1586364061
transform 1 0 45540 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_495
timestamp 1586364061
transform 1 0 46644 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 48852 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_507
timestamp 1586364061
transform 1 0 47748 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_515
timestamp 1586364061
transform 1 0 48484 0 -1 3808
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
timestamp 1586364061
transform 1 0 2576 0 1 3808
box -38 -48 1786 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
timestamp 1586364061
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_3_11
timestamp 1586364061
transform 1 0 2116 0 1 3808
box -38 -48 314 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_35
timestamp 1586364061
transform 1 0 4324 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_40
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 6992 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_68
timestamp 1586364061
transform 1 0 7360 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_72
timestamp 1586364061
transform 1 0 7728 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 7544 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1586364061
transform 1 0 8096 0 1 3808
box -38 -48 866 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 10212 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
timestamp 1586364061
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 9108 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_85
timestamp 1586364061
transform 1 0 8924 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_89
timestamp 1586364061
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_97
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_101
timestamp 1586364061
transform 1 0 10396 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_105
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 10856 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 11040 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_112
timestamp 1586364061
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_116
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_120
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1586364061
transform 1 0 12696 0 1 3808
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
timestamp 1586364061
transform 1 0 14260 0 1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
timestamp 1586364061
transform 1 0 14076 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
timestamp 1586364061
transform 1 0 13708 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_139
timestamp 1586364061
transform 1 0 13892 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
timestamp 1586364061
transform 1 0 16744 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1586364061
transform 1 0 16560 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
timestamp 1586364061
transform 1 0 16192 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_162
timestamp 1586364061
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_166
timestamp 1586364061
transform 1 0 16376 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1586364061
transform 1 0 17296 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_174
timestamp 1586364061
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_178
timestamp 1586364061
transform 1 0 17480 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_193
timestamp 1586364061
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_197
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 406 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1586364061
transform 1 0 21068 0 1 3808
box -38 -48 866 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 19964 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 20884 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 20516 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 19688 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_201
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_204
timestamp 1586364061
transform 1 0 19872 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_209
timestamp 1586364061
transform 1 0 20332 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_213
timestamp 1586364061
transform 1 0 20700 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_226
timestamp 1586364061
transform 1 0 21896 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 22080 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_230
timestamp 1586364061
transform 1 0 22264 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_236
timestamp 1586364061
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 22632 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 23000 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_240
timestamp 1586364061
transform 1 0 23184 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_buf_2  _64_
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_253
timestamp 1586364061
transform 1 0 24380 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_249
timestamp 1586364061
transform 1 0 24012 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__64__A
timestamp 1586364061
transform 1 0 24196 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 24564 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_261
timestamp 1586364061
transform 1 0 25116 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_265
timestamp 1586364061
transform 1 0 25484 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 25300 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_270
timestamp 1586364061
transform 1 0 25944 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1586364061
transform 1 0 25760 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 26128 0 1 3808
box -38 -48 222 592
use scs8hd_conb_1  _46_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 26312 0 1 3808
box -38 -48 314 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 27600 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 27416 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 26772 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_277
timestamp 1586364061
transform 1 0 26588 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_281
timestamp 1586364061
transform 1 0 26956 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_285
timestamp 1586364061
transform 1 0 27324 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_297
timestamp 1586364061
transform 1 0 28428 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_301
timestamp 1586364061
transform 1 0 28796 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 28612 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 28980 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use scs8hd_buf_2  _66_
timestamp 1586364061
transform 1 0 29256 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_310
timestamp 1586364061
transform 1 0 29624 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__66__A
timestamp 1586364061
transform 1 0 29808 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_314
timestamp 1586364061
transform 1 0 29992 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_322
timestamp 1586364061
transform 1 0 30728 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 30360 0 1 3808
box -38 -48 406 592
use scs8hd_conb_1  _44_
timestamp 1586364061
transform 1 0 31464 0 1 3808
box -38 -48 314 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 32568 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
timestamp 1586364061
transform 1 0 32108 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 30912 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
timestamp 1586364061
transform 1 0 31280 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_326
timestamp 1586364061
transform 1 0 31096 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_333
timestamp 1586364061
transform 1 0 31740 0 1 3808
box -38 -48 406 592
use scs8hd_decap_3  FILLER_3_339
timestamp 1586364061
transform 1 0 32292 0 1 3808
box -38 -48 314 592
use scs8hd_conb_1  _45_
timestamp 1586364061
transform 1 0 34868 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 33580 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 33948 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_351
timestamp 1586364061
transform 1 0 33396 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_355
timestamp 1586364061
transform 1 0 33764 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_359
timestamp 1586364061
transform 1 0 34132 0 1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_3_365
timestamp 1586364061
transform 1 0 34684 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_370
timestamp 1586364061
transform 1 0 35144 0 1 3808
box -38 -48 1142 592
use scs8hd_conb_1  _48_
timestamp 1586364061
transform 1 0 37444 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 37260 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_382
timestamp 1586364061
transform 1 0 36248 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_3_390
timestamp 1586364061
transform 1 0 36984 0 1 3808
box -38 -48 314 592
use scs8hd_conb_1  _49_
timestamp 1586364061
transform 1 0 39376 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 39836 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 37904 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 38272 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_398
timestamp 1586364061
transform 1 0 37720 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_402
timestamp 1586364061
transform 1 0 38088 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_406
timestamp 1586364061
transform 1 0 38456 0 1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_3_414
timestamp 1586364061
transform 1 0 39192 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_419
timestamp 1586364061
transform 1 0 39652 0 1 3808
box -38 -48 222 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 40480 0 1 3808
box -38 -48 2246 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 40388 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 40204 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_423
timestamp 1586364061
transform 1 0 40020 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_452
timestamp 1586364061
transform 1 0 42688 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_464
timestamp 1586364061
transform 1 0 43792 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 46000 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_476
timestamp 1586364061
transform 1 0 44896 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_489
timestamp 1586364061
transform 1 0 46092 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 48852 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_501
timestamp 1586364061
transform 1 0 47196 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_3_513
timestamp 1586364061
transform 1 0 48300 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
timestamp 1586364061
transform 1 0 3128 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
timestamp 1586364061
transform 1 0 2576 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_18
timestamp 1586364061
transform 1 0 2760 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_6  FILLER_4_24
timestamp 1586364061
transform 1 0 3312 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_2  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_30
timestamp 1586364061
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 4232 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_40
timestamp 1586364061
transform 1 0 4784 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_36
timestamp 1586364061
transform 1 0 4416 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 4600 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_46
timestamp 1586364061
transform 1 0 5336 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1586364061
transform 1 0 5520 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 7452 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_57
timestamp 1586364061
transform 1 0 6348 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_4_71
timestamp 1586364061
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1586364061
transform 1 0 8004 0 -1 4896
box -38 -48 866 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 10028 0 -1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_4  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 406 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1586364061
transform 1 0 11132 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 10948 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
timestamp 1586364061
transform 1 0 12328 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_101
timestamp 1586364061
transform 1 0 10396 0 -1 4896
box -38 -48 590 592
use scs8hd_decap_4  FILLER_4_118
timestamp 1586364061
transform 1 0 11960 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_124
timestamp 1586364061
transform 1 0 12512 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1586364061
transform 1 0 13616 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1586364061
transform 1 0 12696 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1586364061
transform 1 0 13064 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 13432 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_128
timestamp 1586364061
transform 1 0 12880 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_132
timestamp 1586364061
transform 1 0 13248 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_149
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1586364061
transform 1 0 16560 0 -1 4896
box -38 -48 866 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 15824 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_158
timestamp 1586364061
transform 1 0 15640 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_162
timestamp 1586364061
transform 1 0 16008 0 -1 4896
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_177
timestamp 1586364061
transform 1 0 17388 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_185
timestamp 1586364061
transform 1 0 18124 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_188
timestamp 1586364061
transform 1 0 18400 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_192
timestamp 1586364061
transform 1 0 18768 0 -1 4896
box -38 -48 774 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 866 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 20240 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 19504 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_206
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_210
timestamp 1586364061
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 23000 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 22540 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 21896 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_224
timestamp 1586364061
transform 1 0 21712 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_228
timestamp 1586364061
transform 1 0 22080 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_232
timestamp 1586364061
transform 1 0 22448 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_235
timestamp 1586364061
transform 1 0 22724 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_247
timestamp 1586364061
transform 1 0 23828 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 24380 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 24012 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_255
timestamp 1586364061
transform 1 0 24564 0 -1 4896
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 24748 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_4  FILLER_4_261
timestamp 1586364061
transform 1 0 25116 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_267
timestamp 1586364061
transform 1 0 25668 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 25484 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_271
timestamp 1586364061
transform 1 0 26036 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1586364061
transform 1 0 25852 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1586364061
transform 1 0 26220 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 27600 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 28060 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_285
timestamp 1586364061
transform 1 0 27324 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_290
timestamp 1586364061
transform 1 0 27784 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_295
timestamp 1586364061
transform 1 0 28244 0 -1 4896
box -38 -48 774 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 29164 0 -1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1586364061
transform 1 0 28980 0 -1 4896
box -38 -48 222 592
use scs8hd_or2_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
timestamp 1586364061
transform 1 0 32108 0 -1 4896
box -38 -48 498 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 32752 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
timestamp 1586364061
transform 1 0 31280 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 31832 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_324
timestamp 1586364061
transform 1 0 30912 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_4  FILLER_4_330
timestamp 1586364061
transform 1 0 31464 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_342
timestamp 1586364061
transform 1 0 32568 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_346
timestamp 1586364061
transform 1 0 32936 0 -1 4896
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 33396 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 33120 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_350
timestamp 1586364061
transform 1 0 33304 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_355
timestamp 1586364061
transform 1 0 33764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_367
timestamp 1586364061
transform 1 0 34868 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 37444 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 36064 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 37076 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_379
timestamp 1586364061
transform 1 0 35972 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_382
timestamp 1586364061
transform 1 0 36248 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_390
timestamp 1586364061
transform 1 0 36984 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_393
timestamp 1586364061
transform 1 0 37260 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 37720 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 38732 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_407
timestamp 1586364061
transform 1 0 38548 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_411
timestamp 1586364061
transform 1 0 38916 0 -1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 40480 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 40848 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 41216 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_423
timestamp 1586364061
transform 1 0 40020 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_427
timestamp 1586364061
transform 1 0 40388 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_430
timestamp 1586364061
transform 1 0 40664 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_434
timestamp 1586364061
transform 1 0 41032 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_438
timestamp 1586364061
transform 1 0 41400 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 43240 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_450
timestamp 1586364061
transform 1 0 42504 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_12  FILLER_4_459
timestamp 1586364061
transform 1 0 43332 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_471
timestamp 1586364061
transform 1 0 44436 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_483
timestamp 1586364061
transform 1 0 45540 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_495
timestamp 1586364061
transform 1 0 46644 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 48852 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_507
timestamp 1586364061
transform 1 0 47748 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_515
timestamp 1586364061
transform 1 0 48484 0 -1 4896
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
timestamp 1586364061
transform 1 0 3128 0 1 4896
box -38 -48 1786 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
timestamp 1586364061
transform 1 0 2944 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_19
timestamp 1586364061
transform 1 0 2852 0 1 4896
box -38 -48 130 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
timestamp 1586364061
transform 1 0 5612 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 5060 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
timestamp 1586364061
transform 1 0 5428 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_41
timestamp 1586364061
transform 1 0 4876 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_45
timestamp 1586364061
transform 1 0 5244 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_66
timestamp 1586364061
transform 1 0 7176 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
timestamp 1586364061
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_70
timestamp 1586364061
transform 1 0 7544 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 130 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_90
timestamp 1586364061
transform 1 0 9384 0 1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_101
timestamp 1586364061
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_109
timestamp 1586364061
transform 1 0 11132 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_105
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10948 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
timestamp 1586364061
transform 1 0 13708 0 1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
timestamp 1586364061
transform 1 0 12972 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_127
timestamp 1586364061
transform 1 0 12788 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_131
timestamp 1586364061
transform 1 0 13156 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 16100 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_156
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_161
timestamp 1586364061
transform 1 0 15916 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_165
timestamp 1586364061
transform 1 0 16284 0 1 4896
box -38 -48 1142 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_193
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_197
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 406 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 19780 0 1 4896
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 21068 0 1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 20884 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 20516 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 19596 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_207
timestamp 1586364061
transform 1 0 20148 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_213
timestamp 1586364061
transform 1 0 20700 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_236
timestamp 1586364061
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_240
timestamp 1586364061
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1586364061
transform 1 0 26128 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 24656 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
timestamp 1586364061
transform 1 0 25944 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 25576 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 25208 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_254
timestamp 1586364061
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_258
timestamp 1586364061
transform 1 0 24840 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_264
timestamp 1586364061
transform 1 0 25392 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_268
timestamp 1586364061
transform 1 0 25760 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
timestamp 1586364061
transform 1 0 27140 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 27508 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_281
timestamp 1586364061
transform 1 0 26956 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_285
timestamp 1586364061
transform 1 0 27324 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_289
timestamp 1586364061
transform 1 0 27692 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_297
timestamp 1586364061
transform 1 0 28428 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1586364061
transform 1 0 29256 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
timestamp 1586364061
transform 1 0 28980 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
timestamp 1586364061
transform 1 0 28612 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1586364061
transform 1 0 30268 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1586364061
transform 1 0 30636 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_301
timestamp 1586364061
transform 1 0 28796 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_315
timestamp 1586364061
transform 1 0 30084 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_319
timestamp 1586364061
transform 1 0 30452 0 1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
timestamp 1586364061
transform 1 0 31280 0 1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
timestamp 1586364061
transform 1 0 31096 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_323
timestamp 1586364061
transform 1 0 30820 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_347
timestamp 1586364061
transform 1 0 33028 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 35052 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 33212 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 33580 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_351
timestamp 1586364061
transform 1 0 33396 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_355
timestamp 1586364061
transform 1 0 33764 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_5_363
timestamp 1586364061
transform 1 0 34500 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_367
timestamp 1586364061
transform 1 0 34868 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_371
timestamp 1586364061
transform 1 0 35236 0 1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 36064 0 1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 35880 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 35420 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_375
timestamp 1586364061
transform 1 0 35604 0 1 4896
box -38 -48 314 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 38548 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 37996 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 38364 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 39560 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_399
timestamp 1586364061
transform 1 0 37812 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_403
timestamp 1586364061
transform 1 0 38180 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_416
timestamp 1586364061
transform 1 0 39376 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_420
timestamp 1586364061
transform 1 0 39744 0 1 4896
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 40480 0 1 4896
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 40388 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 40204 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_424
timestamp 1586364061
transform 1 0 40112 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_447
timestamp 1586364061
transform 1 0 42228 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_459
timestamp 1586364061
transform 1 0 43332 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_471
timestamp 1586364061
transform 1 0 44436 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 46000 0 1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_5_483
timestamp 1586364061
transform 1 0 45540 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_487
timestamp 1586364061
transform 1 0 45908 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_489
timestamp 1586364061
transform 1 0 46092 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 48852 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_501
timestamp 1586364061
transform 1 0 47196 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_5_513
timestamp 1586364061
transform 1 0 48300 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_7_21
timestamp 1586364061
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_17
timestamp 1586364061
transform 1 0 2668 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_24
timestamp 1586364061
transform 1 0 3312 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_21
timestamp 1586364061
transform 1 0 3036 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
timestamp 1586364061
transform 1 0 3128 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
timestamp 1586364061
transform 1 0 3128 0 1 5984
box -38 -48 1786 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_30
timestamp 1586364061
transform 1 0 3864 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_41
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_6_49
timestamp 1586364061
transform 1 0 5612 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_7_41
timestamp 1586364061
transform 1 0 4876 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_7_49
timestamp 1586364061
transform 1 0 5612 0 1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_7_58
timestamp 1586364061
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_54
timestamp 1586364061
transform 1 0 6072 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
timestamp 1586364061
transform 1 0 6256 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
timestamp 1586364061
transform 1 0 5888 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_72
timestamp 1586364061
transform 1 0 7728 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_71
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 7544 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
timestamp 1586364061
transform 1 0 5888 0 -1 5984
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_7_85
timestamp 1586364061
transform 1 0 8924 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_83
timestamp 1586364061
transform 1 0 8740 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 8924 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 8188 0 -1 5984
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 8372 0 -1 5984
box -38 -48 406 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1586364061
transform 1 0 8096 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 9108 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_87
timestamp 1586364061
transform 1 0 9108 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_89
timestamp 1586364061
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 9844 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_97
timestamp 1586364061
transform 1 0 10028 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 10212 0 -1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 1786 592
use scs8hd_decap_6  FILLER_6_101
timestamp 1586364061
transform 1 0 10396 0 -1 5984
box -38 -48 590 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10948 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_116
timestamp 1586364061
transform 1 0 11776 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_112
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_116
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11960 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_120
timestamp 1586364061
transform 1 0 12144 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_120
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
timestamp 1586364061
transform 1 0 12512 0 -1 5984
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 12788 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1586364061
transform 1 0 12972 0 1 5984
box -38 -48 866 592
use scs8hd_decap_3  FILLER_7_142
timestamp 1586364061
transform 1 0 14168 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_138
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_143
timestamp 1586364061
transform 1 0 14260 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_147
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 14444 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14812 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_151
timestamp 1586364061
transform 1 0 14996 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_158
timestamp 1586364061
transform 1 0 15640 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
timestamp 1586364061
transform 1 0 15456 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 15180 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1586364061
transform 1 0 15364 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_164
timestamp 1586364061
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_168
timestamp 1586364061
transform 1 0 16560 0 1 5984
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15732 0 -1 5984
box -38 -48 1786 592
use scs8hd_decap_3  FILLER_7_180
timestamp 1586364061
transform 1 0 17664 0 1 5984
box -38 -48 314 592
use scs8hd_decap_6  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 18032 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_conb_1  _39_
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_198
timestamp 1586364061
transform 1 0 19320 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_195
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_187
timestamp 1586364061
transform 1 0 18308 0 1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18216 0 -1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 19688 0 1 5984
box -38 -48 1786 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 19504 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 21620 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_205
timestamp 1586364061
transform 1 0 19964 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_211
timestamp 1586364061
transform 1 0 20516 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_221
timestamp 1586364061
transform 1 0 21436 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_7_233
timestamp 1586364061
transform 1 0 22540 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_229
timestamp 1586364061
transform 1 0 22172 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_225
timestamp 1586364061
transform 1 0 21804 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_229
timestamp 1586364061
transform 1 0 22172 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_224
timestamp 1586364061
transform 1 0 21712 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 22356 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 21988 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 22356 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_241
timestamp 1586364061
transform 1 0 23276 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1786 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 22540 0 -1 5984
box -38 -48 2246 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1586364061
transform 1 0 26128 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 25944 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 26128 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_257
timestamp 1586364061
transform 1 0 24748 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_6_269
timestamp 1586364061
transform 1 0 25852 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_6  FILLER_7_264
timestamp 1586364061
transform 1 0 25392 0 1 5984
box -38 -48 590 592
use scs8hd_decap_4  FILLER_7_285
timestamp 1586364061
transform 1 0 27324 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_281
timestamp 1586364061
transform 1 0 26956 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_274
timestamp 1586364061
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
timestamp 1586364061
transform 1 0 27140 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_295
timestamp 1586364061
transform 1 0 28244 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_291
timestamp 1586364061
transform 1 0 27876 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_295
timestamp 1586364061
transform 1 0 28244 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
timestamp 1586364061
transform 1 0 28060 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
timestamp 1586364061
transform 1 0 27692 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
timestamp 1586364061
transform 1 0 29164 0 -1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 30268 0 1 5984
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 30084 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 29532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 28980 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_303
timestamp 1586364061
transform 1 0 28980 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_306
timestamp 1586364061
transform 1 0 29256 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_311
timestamp 1586364061
transform 1 0 29716 0 1 5984
box -38 -48 406 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1586364061
transform 1 0 32936 0 1 5984
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 32384 0 -1 5984
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 32752 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 32384 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_324
timestamp 1586364061
transform 1 0 30912 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_6_337
timestamp 1586364061
transform 1 0 32108 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_336
timestamp 1586364061
transform 1 0 32016 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_342
timestamp 1586364061
transform 1 0 32568 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_359
timestamp 1586364061
transform 1 0 34132 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_355
timestamp 1586364061
transform 1 0 33764 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_359
timestamp 1586364061
transform 1 0 34132 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 33948 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_367
timestamp 1586364061
transform 1 0 34868 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_7_363
timestamp 1586364061
transform 1 0 34500 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_363
timestamp 1586364061
transform 1 0 34500 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 34316 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 34592 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 35144 0 1 5984
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 34868 0 -1 5984
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_7_379
timestamp 1586364061
transform 1 0 35972 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 36156 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_389
timestamp 1586364061
transform 1 0 36892 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_383
timestamp 1586364061
transform 1 0 36340 0 1 5984
box -38 -48 406 592
use scs8hd_decap_8  FILLER_6_386
timestamp 1586364061
transform 1 0 36616 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 36708 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 37076 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_393
timestamp 1586364061
transform 1 0 37260 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_394
timestamp 1586364061
transform 1 0 37352 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 37444 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 37444 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 37628 0 1 5984
box -38 -48 866 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 39284 0 1 5984
box -38 -48 406 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 37720 0 -1 5984
box -38 -48 2246 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 39836 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_422
timestamp 1586364061
transform 1 0 39928 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_8  FILLER_7_406
timestamp 1586364061
transform 1 0 38456 0 1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_7_414
timestamp 1586364061
transform 1 0 39192 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_419
timestamp 1586364061
transform 1 0 39652 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 40664 0 -1 5984
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 40388 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 40480 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_423
timestamp 1586364061
transform 1 0 40020 0 1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_7_428
timestamp 1586364061
transform 1 0 40480 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_440
timestamp 1586364061
transform 1 0 41584 0 1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
timestamp 1586364061
transform 1 0 42596 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_448
timestamp 1586364061
transform 1 0 42320 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_453
timestamp 1586364061
transform 1 0 42780 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 43240 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
timestamp 1586364061
transform 1 0 43332 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1586364061
transform 1 0 42964 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_457
timestamp 1586364061
transform 1 0 43148 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_459
timestamp 1586364061
transform 1 0 43332 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_457
timestamp 1586364061
transform 1 0 43148 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_449
timestamp 1586364061
transform 1 0 42412 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_461
timestamp 1586364061
transform 1 0 43516 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_465
timestamp 1586364061
transform 1 0 43884 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1586364061
transform 1 0 44068 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1586364061
transform 1 0 43700 0 -1 5984
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1586364061
transform 1 0 43700 0 1 5984
box -38 -48 866 592
use scs8hd_decap_12  FILLER_6_469
timestamp 1586364061
transform 1 0 44252 0 -1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 46000 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
timestamp 1586364061
transform 1 0 45816 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
timestamp 1586364061
transform 1 0 46276 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_481
timestamp 1586364061
transform 1 0 45356 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_493
timestamp 1586364061
transform 1 0 46460 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_472
timestamp 1586364061
transform 1 0 44528 0 1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_484
timestamp 1586364061
transform 1 0 45632 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_489
timestamp 1586364061
transform 1 0 46092 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_493
timestamp 1586364061
transform 1 0 46460 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 48852 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 48852 0 1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_6_505
timestamp 1586364061
transform 1 0 47564 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_6_513
timestamp 1586364061
transform 1 0 48300 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_7_505
timestamp 1586364061
transform 1 0 47564 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_7_513
timestamp 1586364061
transform 1 0 48300 0 1 5984
box -38 -48 314 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 2852 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_8  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 5520 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_8_46
timestamp 1586364061
transform 1 0 5336 0 -1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
timestamp 1586364061
transform 1 0 5888 0 -1 7072
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_8_50
timestamp 1586364061
transform 1 0 5704 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_71
timestamp 1586364061
transform 1 0 7636 0 -1 7072
box -38 -48 406 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 9292 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 8096 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_75
timestamp 1586364061
transform 1 0 8004 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_78
timestamp 1586364061
transform 1 0 8280 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_86
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_91
timestamp 1586364061
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_4  FILLER_8_119
timestamp 1586364061
transform 1 0 12052 0 -1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 12788 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 13156 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_125
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_133
timestamp 1586364061
transform 1 0 13340 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_149
timestamp 1586364061
transform 1 0 14812 0 -1 7072
box -38 -48 130 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 406 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 14904 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_152
timestamp 1586364061
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_158
timestamp 1586364061
transform 1 0 15640 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_12  FILLER_8_170
timestamp 1586364061
transform 1 0 16744 0 -1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 18400 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_182
timestamp 1586364061
transform 1 0 17848 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_186
timestamp 1586364061
transform 1 0 18216 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use scs8hd_conb_1  _40_
timestamp 1586364061
transform 1 0 19780 0 -1 7072
box -38 -48 314 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 21068 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_206
timestamp 1586364061
transform 1 0 20056 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 222 592
use scs8hd_conb_1  _43_
timestamp 1586364061
transform 1 0 23920 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 23644 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_226
timestamp 1586364061
transform 1 0 21896 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_8_238
timestamp 1586364061
transform 1 0 23000 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_244
timestamp 1586364061
transform 1 0 23552 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_247
timestamp 1586364061
transform 1 0 23828 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 24840 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 26128 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_257
timestamp 1586364061
transform 1 0 24748 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_260
timestamp 1586364061
transform 1 0 25024 0 -1 7072
box -38 -48 1142 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
timestamp 1586364061
transform 1 0 27692 0 -1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 27508 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_274
timestamp 1586364061
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_8_280
timestamp 1586364061
transform 1 0 26864 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_286
timestamp 1586364061
transform 1 0 27416 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 30268 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 29624 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 30636 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_308
timestamp 1586364061
transform 1 0 29440 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_312
timestamp 1586364061
transform 1 0 29808 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_316
timestamp 1586364061
transform 1 0 30176 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_319
timestamp 1586364061
transform 1 0 30452 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 32660 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 31096 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 32476 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_323
timestamp 1586364061
transform 1 0 30820 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_328
timestamp 1586364061
transform 1 0 31280 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_4  FILLER_8_337
timestamp 1586364061
transform 1 0 32108 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_347
timestamp 1586364061
transform 1 0 33028 0 -1 7072
box -38 -48 222 592
use scs8hd_conb_1  _47_
timestamp 1586364061
transform 1 0 35328 0 -1 7072
box -38 -48 314 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 33764 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 35144 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 33212 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 33580 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_351
timestamp 1586364061
transform 1 0 33396 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_364
timestamp 1586364061
transform 1 0 34592 0 -1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_375
timestamp 1586364061
transform 1 0 35604 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_8_387
timestamp 1586364061
transform 1 0 36708 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_395
timestamp 1586364061
transform 1 0 37444 0 -1 7072
box -38 -48 222 592
use scs8hd_conb_1  _50_
timestamp 1586364061
transform 1 0 37812 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 38272 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_398
timestamp 1586364061
transform 1 0 37720 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_402
timestamp 1586364061
transform 1 0 38088 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_406
timestamp 1586364061
transform 1 0 38456 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_418
timestamp 1586364061
transform 1 0 39560 0 -1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
timestamp 1586364061
transform 1 0 41032 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_430
timestamp 1586364061
transform 1 0 40664 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_436
timestamp 1586364061
transform 1 0 41216 0 -1 7072
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
timestamp 1586364061
transform 1 0 43332 0 -1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 43240 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_448
timestamp 1586364061
transform 1 0 42320 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_456
timestamp 1586364061
transform 1 0 43056 0 -1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
timestamp 1586364061
transform 1 0 45816 0 -1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
timestamp 1586364061
transform 1 0 45264 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_478
timestamp 1586364061
transform 1 0 45080 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_482
timestamp 1586364061
transform 1 0 45448 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 48852 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_505
timestamp 1586364061
transform 1 0 47564 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_513
timestamp 1586364061
transform 1 0 48300 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 1564 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_7
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_19
timestamp 1586364061
transform 1 0 2852 0 1 7072
box -38 -48 1142 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
timestamp 1586364061
transform 1 0 4048 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
timestamp 1586364061
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_31
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_34
timestamp 1586364061
transform 1 0 4232 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_38
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 774 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 774 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 9292 0 1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 9108 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 8740 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_82
timestamp 1586364061
transform 1 0 8648 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_85
timestamp 1586364061
transform 1 0 8924 0 1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_108
timestamp 1586364061
transform 1 0 11040 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_112
timestamp 1586364061
transform 1 0 11408 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 14720 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_142
timestamp 1586364061
transform 1 0 14168 0 1 7072
box -38 -48 590 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1586364061
transform 1 0 14904 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 15916 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16284 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 16652 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_159
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_163
timestamp 1586364061
transform 1 0 16100 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_167
timestamp 1586364061
transform 1 0 16468 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_171
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_182
timestamp 1586364061
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_178
timestamp 1586364061
transform 1 0 17480 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 17296 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 17664 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_193
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use scs8hd_decap_6  FILLER_9_197
timestamp 1586364061
transform 1 0 19228 0 1 7072
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 20700 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 20516 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 20148 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 19780 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_205
timestamp 1586364061
transform 1 0 19964 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_209
timestamp 1586364061
transform 1 0 20332 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_222
timestamp 1586364061
transform 1 0 21528 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_230
timestamp 1586364061
transform 1 0 22264 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_226
timestamp 1586364061
transform 1 0 21896 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 22080 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 21712 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_234
timestamp 1586364061
transform 1 0 22632 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 22816 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_238
timestamp 1586364061
transform 1 0 23000 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_248
timestamp 1586364061
transform 1 0 23920 0 1 7072
box -38 -48 590 592
use scs8hd_conb_1  _41_
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 314 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
timestamp 1586364061
transform 1 0 25300 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 24472 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_256
timestamp 1586364061
transform 1 0 24656 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_260
timestamp 1586364061
transform 1 0 25024 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_267
timestamp 1586364061
transform 1 0 25668 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_271
timestamp 1586364061
transform 1 0 26036 0 1 7072
box -38 -48 406 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1586364061
transform 1 0 27600 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
timestamp 1586364061
transform 1 0 26496 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
timestamp 1586364061
transform 1 0 26864 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 27416 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_275
timestamp 1586364061
transform 1 0 26404 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_278
timestamp 1586364061
transform 1 0 26680 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_282
timestamp 1586364061
transform 1 0 27048 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_297
timestamp 1586364061
transform 1 0 28428 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1586364061
transform 1 0 29532 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 28980 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 28612 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 30544 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_301
timestamp 1586364061
transform 1 0 28796 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_306
timestamp 1586364061
transform 1 0 29256 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_318
timestamp 1586364061
transform 1 0 30360 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_322
timestamp 1586364061
transform 1 0 30728 0 1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 31096 0 1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 30912 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_345
timestamp 1586364061
transform 1 0 32844 0 1 7072
box -38 -48 774 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 33580 0 1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 34132 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_357
timestamp 1586364061
transform 1 0 33948 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_361
timestamp 1586364061
transform 1 0 34316 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_365
timestamp 1586364061
transform 1 0 34684 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_367
timestamp 1586364061
transform 1 0 34868 0 1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
timestamp 1586364061
transform 1 0 37628 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
timestamp 1586364061
transform 1 0 37260 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 36892 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_379
timestamp 1586364061
transform 1 0 35972 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_387
timestamp 1586364061
transform 1 0 36708 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_391
timestamp 1586364061
transform 1 0 37076 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_395
timestamp 1586364061
transform 1 0 37444 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1586364061
transform 1 0 37812 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
timestamp 1586364061
transform 1 0 39836 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 38824 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_408
timestamp 1586364061
transform 1 0 38640 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_412
timestamp 1586364061
transform 1 0 39008 0 1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_9_420
timestamp 1586364061
transform 1 0 39744 0 1 7072
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
timestamp 1586364061
transform 1 0 41032 0 1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 40388 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
timestamp 1586364061
transform 1 0 40848 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
timestamp 1586364061
transform 1 0 40204 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_423
timestamp 1586364061
transform 1 0 40020 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_428
timestamp 1586364061
transform 1 0 40480 0 1 7072
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
timestamp 1586364061
transform 1 0 43516 0 1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
timestamp 1586364061
transform 1 0 43332 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_453
timestamp 1586364061
transform 1 0 42780 0 1 7072
box -38 -48 590 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 46736 0 1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 46000 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
timestamp 1586364061
transform 1 0 45448 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_480
timestamp 1586364061
transform 1 0 45264 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_484
timestamp 1586364061
transform 1 0 45632 0 1 7072
box -38 -48 406 592
use scs8hd_decap_6  FILLER_9_489
timestamp 1586364061
transform 1 0 46092 0 1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_9_495
timestamp 1586364061
transform 1 0 46644 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 48852 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 47288 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_500
timestamp 1586364061
transform 1 0 47104 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_504
timestamp 1586364061
transform 1 0 47472 0 1 7072
box -38 -48 1142 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 1472 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_6  FILLER_10_8
timestamp 1586364061
transform 1 0 1840 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_14
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_17
timestamp 1586364061
transform 1 0 2668 0 -1 8160
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_29
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
timestamp 1586364061
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
timestamp 1586364061
transform 1 0 6440 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_51
timestamp 1586364061
transform 1 0 5796 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_57
timestamp 1586364061
transform 1 0 6348 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_60
timestamp 1586364061
transform 1 0 6624 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_64
timestamp 1586364061
transform 1 0 6992 0 -1 8160
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_76
timestamp 1586364061
transform 1 0 8096 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_10_88
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 406 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1586364061
transform 1 0 12420 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
timestamp 1586364061
transform 1 0 11960 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 11592 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_112
timestamp 1586364061
transform 1 0 11408 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_116
timestamp 1586364061
transform 1 0 11776 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_120
timestamp 1586364061
transform 1 0 12144 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_132
timestamp 1586364061
transform 1 0 13248 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_10_144
timestamp 1586364061
transform 1 0 14352 0 -1 8160
box -38 -48 590 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15916 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 16928 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 14904 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_152
timestamp 1586364061
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_6  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_160
timestamp 1586364061
transform 1 0 15824 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_170
timestamp 1586364061
transform 1 0 16744 0 -1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 17664 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_174
timestamp 1586364061
transform 1 0 17112 0 -1 8160
box -38 -48 406 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 21160 0 -1 8160
box -38 -48 2246 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 20516 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_199
timestamp 1586364061
transform 1 0 19412 0 -1 8160
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_10_213
timestamp 1586364061
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 23644 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_242
timestamp 1586364061
transform 1 0 23368 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_247
timestamp 1586364061
transform 1 0 23828 0 -1 8160
box -38 -48 774 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1586364061
transform 1 0 24840 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
timestamp 1586364061
transform 1 0 24656 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
timestamp 1586364061
transform 1 0 26128 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_255
timestamp 1586364061
transform 1 0 24564 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_267
timestamp 1586364061
transform 1 0 25668 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_271
timestamp 1586364061
transform 1 0 26036 0 -1 8160
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 28428 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_274
timestamp 1586364061
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_295
timestamp 1586364061
transform 1 0 28244 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1586364061
transform 1 0 28980 0 -1 8160
box -38 -48 866 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 30544 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 30176 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 28796 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_299
timestamp 1586364061
transform 1 0 28612 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_312
timestamp 1586364061
transform 1 0 29808 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_318
timestamp 1586364061
transform 1 0 30360 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 31740 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
timestamp 1586364061
transform 1 0 32292 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_324
timestamp 1586364061
transform 1 0 30912 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_332
timestamp 1586364061
transform 1 0 31648 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_335
timestamp 1586364061
transform 1 0 31924 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_337
timestamp 1586364061
transform 1 0 32108 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_341
timestamp 1586364061
transform 1 0 32476 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_353
timestamp 1586364061
transform 1 0 33580 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_365
timestamp 1586364061
transform 1 0 34684 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
timestamp 1586364061
transform 1 0 36432 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 35880 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_377
timestamp 1586364061
transform 1 0 35788 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_380
timestamp 1586364061
transform 1 0 36064 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_8  FILLER_10_386
timestamp 1586364061
transform 1 0 36616 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_10_394
timestamp 1586364061
transform 1 0 37352 0 -1 8160
box -38 -48 314 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
timestamp 1586364061
transform 1 0 37720 0 -1 8160
box -38 -48 1786 592
use scs8hd_decap_6  FILLER_10_417
timestamp 1586364061
transform 1 0 39468 0 -1 8160
box -38 -48 590 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
timestamp 1586364061
transform 1 0 40204 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 40020 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_444
timestamp 1586364061
transform 1 0 41952 0 -1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 43240 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
timestamp 1586364061
transform 1 0 43516 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 42964 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_452
timestamp 1586364061
transform 1 0 42688 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_457
timestamp 1586364061
transform 1 0 43148 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_459
timestamp 1586364061
transform 1 0 43332 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_463
timestamp 1586364061
transform 1 0 43700 0 -1 8160
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
timestamp 1586364061
transform 1 0 44804 0 -1 8160
box -38 -48 1786 592
use scs8hd_decap_12  FILLER_10_494
timestamp 1586364061
transform 1 0 46552 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 48852 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_506
timestamp 1586364061
transform 1 0 47656 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_514
timestamp 1586364061
transform 1 0 48392 0 -1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 1786 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
timestamp 1586364061
transform 1 0 2300 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 590 592
use scs8hd_fill_2  FILLER_11_11
timestamp 1586364061
transform 1 0 2116 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_34
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_38
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_42
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_46
timestamp 1586364061
transform 1 0 5336 0 1 8160
box -38 -48 774 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
timestamp 1586364061
transform 1 0 6440 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
timestamp 1586364061
transform 1 0 6072 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_56
timestamp 1586364061
transform 1 0 6256 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_60
timestamp 1586364061
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_81
timestamp 1586364061
transform 1 0 8556 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_93
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
timestamp 1586364061
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_105
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_111
timestamp 1586364061
transform 1 0 11316 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_142
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 774 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1586364061
transform 1 0 16284 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
timestamp 1586364061
transform 1 0 15272 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 16100 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
timestamp 1586364061
transform 1 0 14904 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_152
timestamp 1586364061
transform 1 0 15088 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_156
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_161
timestamp 1586364061
transform 1 0 15916 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_174
timestamp 1586364061
transform 1 0 17112 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_179
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 20516 0 1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 20332 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_203
timestamp 1586364061
transform 1 0 19780 0 1 8160
box -38 -48 590 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_230
timestamp 1586364061
transform 1 0 22264 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_234
timestamp 1586364061
transform 1 0 22632 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_238
timestamp 1586364061
transform 1 0 23000 0 1 8160
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
timestamp 1586364061
transform 1 0 26128 0 1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
timestamp 1586364061
transform 1 0 25944 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1586364061
transform 1 0 25576 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_264
timestamp 1586364061
transform 1 0 25392 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_268
timestamp 1586364061
transform 1 0 25760 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1586364061
transform 1 0 28060 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 28428 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_291
timestamp 1586364061
transform 1 0 27876 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_295
timestamp 1586364061
transform 1 0 28244 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1586364061
transform 1 0 30176 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 29992 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 29440 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 28980 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_299
timestamp 1586364061
transform 1 0 28612 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_306
timestamp 1586364061
transform 1 0 29256 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_310
timestamp 1586364061
transform 1 0 29624 0 1 8160
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 31740 0 1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
timestamp 1586364061
transform 1 0 31556 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_325
timestamp 1586364061
transform 1 0 31004 0 1 8160
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_352
timestamp 1586364061
transform 1 0 33488 0 1 8160
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_11_364
timestamp 1586364061
transform 1 0 34592 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_367
timestamp 1586364061
transform 1 0 34868 0 1 8160
box -38 -48 590 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
timestamp 1586364061
transform 1 0 36432 0 1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
timestamp 1586364061
transform 1 0 36248 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 35880 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 35512 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_373
timestamp 1586364061
transform 1 0 35420 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_376
timestamp 1586364061
transform 1 0 35696 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_380
timestamp 1586364061
transform 1 0 36064 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
timestamp 1586364061
transform 1 0 39836 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 39468 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 38548 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 38916 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_403
timestamp 1586364061
transform 1 0 38180 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_409
timestamp 1586364061
transform 1 0 38732 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_413
timestamp 1586364061
transform 1 0 39100 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_419
timestamp 1586364061
transform 1 0 39652 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
timestamp 1586364061
transform 1 0 40480 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 40388 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
timestamp 1586364061
transform 1 0 40204 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_423
timestamp 1586364061
transform 1 0 40020 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_447
timestamp 1586364061
transform 1 0 42228 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1586364061
transform 1 0 42964 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
timestamp 1586364061
transform 1 0 42412 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 42780 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_451
timestamp 1586364061
transform 1 0 42596 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_464
timestamp 1586364061
transform 1 0 43792 0 1 8160
box -38 -48 1142 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 46736 0 1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 46000 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
timestamp 1586364061
transform 1 0 45080 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
timestamp 1586364061
transform 1 0 45448 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_476
timestamp 1586364061
transform 1 0 44896 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_480
timestamp 1586364061
transform 1 0 45264 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_484
timestamp 1586364061
transform 1 0 45632 0 1 8160
box -38 -48 406 592
use scs8hd_decap_6  FILLER_11_489
timestamp 1586364061
transform 1 0 46092 0 1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_495
timestamp 1586364061
transform 1 0 46644 0 1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 48852 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 47288 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_500
timestamp 1586364061
transform 1 0 47104 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_504
timestamp 1586364061
transform 1 0 47472 0 1 8160
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_12_11
timestamp 1586364061
transform 1 0 2116 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_7
timestamp 1586364061
transform 1 0 1748 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
timestamp 1586364061
transform 1 0 1932 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
timestamp 1586364061
transform 1 0 1564 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 2668 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 2300 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_19
timestamp 1586364061
transform 1 0 2852 0 -1 9248
box -38 -48 1142 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_41
timestamp 1586364061
transform 1 0 4876 0 -1 9248
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
timestamp 1586364061
transform 1 0 6440 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_53
timestamp 1586364061
transform 1 0 5980 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_81
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_77
timestamp 1586364061
transform 1 0 8188 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1586364061
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_85
timestamp 1586364061
transform 1 0 8924 0 -1 9248
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1586364061
transform 1 0 8740 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_91
timestamp 1586364061
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_99
timestamp 1586364061
transform 1 0 10212 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
timestamp 1586364061
transform 1 0 10028 0 -1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
timestamp 1586364061
transform 1 0 11960 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
timestamp 1586364061
transform 1 0 10396 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_103
timestamp 1586364061
transform 1 0 10580 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_12_115
timestamp 1586364061
transform 1 0 11684 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
timestamp 1586364061
transform 1 0 14536 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_137
timestamp 1586364061
transform 1 0 13708 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_148
timestamp 1586364061
transform 1 0 14720 0 -1 9248
box -38 -48 314 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_173
timestamp 1586364061
transform 1 0 17020 0 -1 9248
box -38 -48 590 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 17756 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17572 0 -1 9248
box -38 -48 222 592
use scs8hd_conb_1  _42_
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_200
timestamp 1586364061
transform 1 0 19504 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_12_212
timestamp 1586364061
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_218
timestamp 1586364061
transform 1 0 21160 0 -1 9248
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 22264 0 -1 9248
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
timestamp 1586364061
transform 1 0 24656 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
timestamp 1586364061
transform 1 0 24472 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_249
timestamp 1586364061
transform 1 0 24012 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_253
timestamp 1586364061
transform 1 0 24380 0 -1 9248
box -38 -48 130 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 866 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1586364061
transform 1 0 27508 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 28520 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_285
timestamp 1586364061
transform 1 0 27324 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_296
timestamp 1586364061
transform 1 0 28336 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1586364061
transform 1 0 29072 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
timestamp 1586364061
transform 1 0 30084 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 28888 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 30452 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_300
timestamp 1586364061
transform 1 0 28704 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_313
timestamp 1586364061
transform 1 0 29900 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_317
timestamp 1586364061
transform 1 0 30268 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_321
timestamp 1586364061
transform 1 0 30636 0 -1 9248
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
timestamp 1586364061
transform 1 0 32108 0 -1 9248
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 31740 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_335
timestamp 1586364061
transform 1 0 31924 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 34868 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_356
timestamp 1586364061
transform 1 0 33856 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_12_364
timestamp 1586364061
transform 1 0 34592 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_12_369
timestamp 1586364061
transform 1 0 35052 0 -1 9248
box -38 -48 406 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1586364061
transform 1 0 35880 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 35512 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_373
timestamp 1586364061
transform 1 0 35420 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_376
timestamp 1586364061
transform 1 0 35696 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_387
timestamp 1586364061
transform 1 0 36708 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_395
timestamp 1586364061
transform 1 0 37444 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1586364061
transform 1 0 38548 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 39928 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 38364 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_398
timestamp 1586364061
transform 1 0 37720 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_404
timestamp 1586364061
transform 1 0 38272 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_12_416
timestamp 1586364061
transform 1 0 39376 0 -1 9248
box -38 -48 590 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1586364061
transform 1 0 40112 0 -1 9248
box -38 -48 866 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
timestamp 1586364061
transform 1 0 41768 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_12_433
timestamp 1586364061
transform 1 0 40940 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_441
timestamp 1586364061
transform 1 0 41676 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_446
timestamp 1586364061
transform 1 0 42136 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_454
timestamp 1586364061
transform 1 0 42872 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_450
timestamp 1586364061
transform 1 0 42504 0 -1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 42964 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
timestamp 1586364061
transform 1 0 42320 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_463
timestamp 1586364061
transform 1 0 43700 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_459
timestamp 1586364061
transform 1 0 43332 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_457
timestamp 1586364061
transform 1 0 43148 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 43516 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 43240 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1586364061
transform 1 0 44436 0 -1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
timestamp 1586364061
transform 1 0 45080 0 -1 9248
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_12_473
timestamp 1586364061
transform 1 0 44620 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_477
timestamp 1586364061
transform 1 0 44988 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 48852 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_497
timestamp 1586364061
transform 1 0 46828 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_12_509
timestamp 1586364061
transform 1 0 47932 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_515
timestamp 1586364061
transform 1 0 48484 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_7
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
timestamp 1586364061
transform 1 0 1564 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1586364061
transform 1 0 1932 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_22
timestamp 1586364061
transform 1 0 3128 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 3312 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_18
timestamp 1586364061
transform 1 0 2760 0 -1 10336
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_30
timestamp 1586364061
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_26
timestamp 1586364061
transform 1 0 3496 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 3680 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_286
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
timestamp 1586364061
transform 1 0 4140 0 -1 10336
box -38 -48 406 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1586364061
transform 1 0 3864 0 1 9248
box -38 -48 866 592
use scs8hd_decap_3  FILLER_14_41
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_37
timestamp 1586364061
transform 1 0 4508 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_43
timestamp 1586364061
transform 1 0 5060 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 4692 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
timestamp 1586364061
transform 1 0 4876 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
timestamp 1586364061
transform 1 0 5244 0 1 9248
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 5428 0 1 9248
box -38 -48 406 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
timestamp 1586364061
transform 1 0 5336 0 -1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 5888 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_55
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_50
timestamp 1586364061
transform 1 0 5704 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_54
timestamp 1586364061
transform 1 0 6072 0 -1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1586364061
transform 1 0 6440 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_60
timestamp 1586364061
transform 1 0 6624 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1586364061
transform 1 0 6440 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_3  FILLER_14_72
timestamp 1586364061
transform 1 0 7728 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_67
timestamp 1586364061
transform 1 0 7268 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_66
timestamp 1586364061
transform 1 0 7176 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1586364061
transform 1 0 6992 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
timestamp 1586364061
transform 1 0 7544 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
timestamp 1586364061
transform 1 0 7360 0 1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
timestamp 1586364061
transform 1 0 7544 0 1 9248
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1586364061
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1586364061
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_4  FILLER_14_88
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_95
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_89
timestamp 1586364061
transform 1 0 9292 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_287
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_or2_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 498 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_13_106
timestamp 1586364061
transform 1 0 10856 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_102
timestamp 1586364061
transform 1 0 10488 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
timestamp 1586364061
transform 1 0 10672 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_112
timestamp 1586364061
transform 1 0 11408 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1586364061
transform 1 0 12144 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_129
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_127
timestamp 1586364061
transform 1 0 12788 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 12972 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 12604 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13156 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_13_143
timestamp 1586364061
transform 1 0 14260 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
timestamp 1586364061
transform 1 0 14352 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_133
timestamp 1586364061
transform 1 0 13340 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_131
timestamp 1586364061
transform 1 0 13156 0 1 9248
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
timestamp 1586364061
transform 1 0 14536 0 1 9248
box -38 -48 1786 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_288
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 16468 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_165
timestamp 1586364061
transform 1 0 16284 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_169
timestamp 1586364061
transform 1 0 16652 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_173
timestamp 1586364061
transform 1 0 17020 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_163
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_185
timestamp 1586364061
transform 1 0 18124 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_181
timestamp 1586364061
transform 1 0 17756 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_175
timestamp 1586364061
transform 1 0 17204 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_181
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_conb_1  _36_
timestamp 1586364061
transform 1 0 17848 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_189
timestamp 1586364061
transform 1 0 18492 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 18676 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 18308 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_193
timestamp 1586364061
transform 1 0 18860 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_196
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_205
timestamp 1586364061
transform 1 0 19964 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_6  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 590 592
use scs8hd_decap_3  FILLER_14_211
timestamp 1586364061
transform 1 0 20516 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_217
timestamp 1586364061
transform 1 0 21068 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_214
timestamp 1586364061
transform 1 0 20792 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 20332 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 20884 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_289
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_221
timestamp 1586364061
transform 1 0 21436 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 21620 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 21252 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_231
timestamp 1586364061
transform 1 0 22356 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_228
timestamp 1586364061
transform 1 0 22080 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_224
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_234
timestamp 1586364061
transform 1 0 22632 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_231
timestamp 1586364061
transform 1 0 22356 0 1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_13_225
timestamp 1586364061
transform 1 0 21804 0 1 9248
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 22172 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 22448 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_3  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_242
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_238
timestamp 1586364061
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 23920 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_241
timestamp 1586364061
transform 1 0 23276 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_14_253
timestamp 1586364061
transform 1 0 24380 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_258
timestamp 1586364061
transform 1 0 24840 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_254
timestamp 1586364061
transform 1 0 24472 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_250
timestamp 1586364061
transform 1 0 24104 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 24656 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
timestamp 1586364061
transform 1 0 24288 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 24656 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
timestamp 1586364061
transform 1 0 25024 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1586364061
transform 1 0 24840 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_3  FILLER_14_272
timestamp 1586364061
transform 1 0 26128 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_267
timestamp 1586364061
transform 1 0 25668 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_clkbuf_1_0__f_clk_A
timestamp 1586364061
transform 1 0 25944 0 -1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
timestamp 1586364061
transform 1 0 25208 0 1 9248
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_285
timestamp 1586364061
transform 1 0 27324 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_281
timestamp 1586364061
transform 1 0 26956 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1586364061
transform 1 0 27140 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
timestamp 1586364061
transform 1 0 26680 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_290
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_296
timestamp 1586364061
transform 1 0 28336 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_292
timestamp 1586364061
transform 1 0 27968 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_297
timestamp 1586364061
transform 1 0 28428 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_289
timestamp 1586364061
transform 1 0 27692 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
timestamp 1586364061
transform 1 0 27876 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 27508 0 1 9248
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
timestamp 1586364061
transform 1 0 28060 0 1 9248
box -38 -48 406 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1586364061
transform 1 0 28428 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_12  FILLER_14_280
timestamp 1586364061
transform 1 0 26864 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_306
timestamp 1586364061
transform 1 0 29256 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_306
timestamp 1586364061
transform 1 0 29256 0 1 9248
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_301
timestamp 1586364061
transform 1 0 28796 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 28980 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 28612 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
timestamp 1586364061
transform 1 0 29440 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_312
timestamp 1586364061
transform 1 0 29808 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
timestamp 1586364061
transform 1 0 29900 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_322
timestamp 1586364061
transform 1 0 30728 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_310
timestamp 1586364061
transform 1 0 29624 0 -1 10336
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
timestamp 1586364061
transform 1 0 30084 0 1 9248
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_291
timestamp 1586364061
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_334
timestamp 1586364061
transform 1 0 31832 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_346
timestamp 1586364061
transform 1 0 32936 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_334
timestamp 1586364061
transform 1 0 31832 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_337
timestamp 1586364061
transform 1 0 32108 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_13_358
timestamp 1586364061
transform 1 0 34040 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 34224 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_361
timestamp 1586364061
transform 1 0 34316 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_13_371
timestamp 1586364061
transform 1 0 35236 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_367
timestamp 1586364061
transform 1 0 34868 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_362
timestamp 1586364061
transform 1 0 34408 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 34592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 35328 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1586364061
transform 1 0 34868 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_12  FILLER_14_349
timestamp 1586364061
transform 1 0 33212 0 -1 10336
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 35512 0 1 9248
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_292
timestamp 1586364061
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_393
timestamp 1586364061
transform 1 0 37260 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_397
timestamp 1586364061
transform 1 0 37628 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_376
timestamp 1586364061
transform 1 0 35696 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_388
timestamp 1586364061
transform 1 0 36800 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_396
timestamp 1586364061
transform 1 0 37536 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_14_407
timestamp 1586364061
transform 1 0 38548 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_404
timestamp 1586364061
transform 1 0 38272 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_400
timestamp 1586364061
transform 1 0 37904 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 38456 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 38088 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 37720 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1586364061
transform 1 0 37720 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_3  FILLER_14_412
timestamp 1586364061
transform 1 0 39008 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_13_417
timestamp 1586364061
transform 1 0 39468 0 1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_13_414
timestamp 1586364061
transform 1 0 39192 0 1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_13_408
timestamp 1586364061
transform 1 0 38640 0 1 9248
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
timestamp 1586364061
transform 1 0 39284 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 38824 0 -1 10336
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
timestamp 1586364061
transform 1 0 39284 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_419
timestamp 1586364061
transform 1 0 39652 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_14_431
timestamp 1586364061
transform 1 0 40756 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_13_432
timestamp 1586364061
transform 1 0 40848 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_428
timestamp 1586364061
transform 1 0 40480 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_425
timestamp 1586364061
transform 1 0 40204 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 40664 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 40388 0 1 9248
box -38 -48 130 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 40388 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_440
timestamp 1586364061
transform 1 0 41584 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_436
timestamp 1586364061
transform 1 0 41216 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_439
timestamp 1586364061
transform 1 0 41492 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_436
timestamp 1586364061
transform 1 0 41216 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 41032 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 41308 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 41400 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 41676 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_444
timestamp 1586364061
transform 1 0 41952 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_443
timestamp 1586364061
transform 1 0 41860 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 41768 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 42044 0 1 9248
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
timestamp 1586364061
transform 1 0 42136 0 -1 10336
box -38 -48 406 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1586364061
transform 1 0 42228 0 1 9248
box -38 -48 866 592
use scs8hd_decap_6  FILLER_14_450
timestamp 1586364061
transform 1 0 42504 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_3  FILLER_13_456
timestamp 1586364061
transform 1 0 43056 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1586364061
transform 1 0 43056 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_465
timestamp 1586364061
transform 1 0 43884 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_461
timestamp 1586364061
transform 1 0 43516 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 43700 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 43332 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_293
timestamp 1586364061
transform 1 0 43240 0 -1 10336
box -38 -48 130 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1586364061
transform 1 0 43332 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_3  FILLER_14_468
timestamp 1586364061
transform 1 0 44160 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1586364061
transform 1 0 44436 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1586364061
transform 1 0 44252 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1586364061
transform 1 0 44436 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_481
timestamp 1586364061
transform 1 0 45356 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_473
timestamp 1586364061
transform 1 0 44620 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_13_480
timestamp 1586364061
transform 1 0 45264 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
timestamp 1586364061
transform 1 0 45540 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_493
timestamp 1586364061
transform 1 0 46460 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_489
timestamp 1586364061
transform 1 0 46092 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_485
timestamp 1586364061
transform 1 0 45724 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
timestamp 1586364061
transform 1 0 46276 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 46000 0 1 9248
box -38 -48 130 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 46736 0 1 9248
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
timestamp 1586364061
transform 1 0 45540 0 -1 10336
box -38 -48 1786 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 48852 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 48852 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 47288 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_500
timestamp 1586364061
transform 1 0 47104 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_504
timestamp 1586364061
transform 1 0 47472 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_502
timestamp 1586364061
transform 1 0 47288 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_514
timestamp 1586364061
transform 1 0 48392 0 -1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
timestamp 1586364061
transform 1 0 1564 0 1 10336
box -38 -48 1786 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_24
timestamp 1586364061
transform 1 0 3312 0 1 10336
box -38 -48 774 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
timestamp 1586364061
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_32
timestamp 1586364061
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_36
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_40
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_294
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_71
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_75
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_102
timestamp 1586364061
transform 1 0 10488 0 1 10336
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 11040 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_295
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_136
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_148
timestamp 1586364061
transform 1 0 14720 0 1 10336
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_156
timestamp 1586364061
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_160
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_164
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 1142 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_296
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_176
timestamp 1586364061
transform 1 0 17296 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_193
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_197
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 590 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 20332 0 1 10336
box -38 -48 2246 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 20148 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 19780 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_205
timestamp 1586364061
transform 1 0 19964 0 1 10336
box -38 -48 222 592
use scs8hd_conb_1  _37_
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_297
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 22724 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_233
timestamp 1586364061
transform 1 0 22540 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_237
timestamp 1586364061
transform 1 0 22908 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_243
timestamp 1586364061
transform 1 0 23460 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_248
timestamp 1586364061
transform 1 0 23920 0 1 10336
box -38 -48 1142 592
use scs8hd_clkbuf_16  clkbuf_1_0__f_clk tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 25944 0 1 10336
box -38 -48 1878 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
timestamp 1586364061
transform 1 0 25760 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_260
timestamp 1586364061
transform 1 0 25024 0 1 10336
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
timestamp 1586364061
transform 1 0 28244 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_290
timestamp 1586364061
transform 1 0 27784 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_294
timestamp 1586364061
transform 1 0 28152 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_297
timestamp 1586364061
transform 1 0 28428 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
timestamp 1586364061
transform 1 0 29256 0 1 10336
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_298
timestamp 1586364061
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
timestamp 1586364061
transform 1 0 28980 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
timestamp 1586364061
transform 1 0 28612 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_301
timestamp 1586364061
transform 1 0 28796 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_325
timestamp 1586364061
transform 1 0 31004 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_337
timestamp 1586364061
transform 1 0 32108 0 1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_15_358
timestamp 1586364061
transform 1 0 34040 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_355
timestamp 1586364061
transform 1 0 33764 0 1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_15_349
timestamp 1586364061
transform 1 0 33212 0 1 10336
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 34224 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 33856 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_367
timestamp 1586364061
transform 1 0 34868 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_362
timestamp 1586364061
transform 1 0 34408 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 34592 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_299
timestamp 1586364061
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 34960 0 1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 37536 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_387
timestamp 1586364061
transform 1 0 36708 0 1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_15_395
timestamp 1586364061
transform 1 0 37444 0 1 10336
box -38 -48 130 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1586364061
transform 1 0 38824 0 1 10336
box -38 -48 866 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 37720 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 38640 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 38272 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 39836 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_402
timestamp 1586364061
transform 1 0 38088 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_406
timestamp 1586364061
transform 1 0 38456 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_419
timestamp 1586364061
transform 1 0 39652 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1586364061
transform 1 0 41400 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_300
timestamp 1586364061
transform 1 0 40388 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
timestamp 1586364061
transform 1 0 40664 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
timestamp 1586364061
transform 1 0 41032 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_423
timestamp 1586364061
transform 1 0 40020 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_428
timestamp 1586364061
transform 1 0 40480 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_432
timestamp 1586364061
transform 1 0 40848 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_436
timestamp 1586364061
transform 1 0 41216 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_447
timestamp 1586364061
transform 1 0 42228 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
timestamp 1586364061
transform 1 0 43332 0 1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
timestamp 1586364061
transform 1 0 43148 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
timestamp 1586364061
transform 1 0 42780 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1586364061
transform 1 0 42412 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_451
timestamp 1586364061
transform 1 0 42596 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_455
timestamp 1586364061
transform 1 0 42964 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_301
timestamp 1586364061
transform 1 0 46000 0 1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_15_478
timestamp 1586364061
transform 1 0 45080 0 1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_15_486
timestamp 1586364061
transform 1 0 45816 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_489
timestamp 1586364061
transform 1 0 46092 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 48852 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_501
timestamp 1586364061
transform 1 0 47196 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_15_513
timestamp 1586364061
transform 1 0 48300 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_7
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 1932 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
timestamp 1586364061
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_11
timestamp 1586364061
transform 1 0 2116 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
timestamp 1586364061
transform 1 0 2300 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_19
timestamp 1586364061
transform 1 0 2852 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 2668 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 3312 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1586364061
transform 1 0 5336 0 -1 11424
box -38 -48 866 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
timestamp 1586364061
transform 1 0 4232 0 -1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_302
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_26
timestamp 1586364061
transform 1 0 3496 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_30
timestamp 1586364061
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_38
timestamp 1586364061
transform 1 0 4600 0 -1 11424
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7452 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 7820 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 6440 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_55
timestamp 1586364061
transform 1 0 6164 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_60
timestamp 1586364061
transform 1 0 6624 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_64
timestamp 1586364061
transform 1 0 6992 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_71
timestamp 1586364061
transform 1 0 7636 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 10212 0 -1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_303
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
timestamp 1586364061
transform 1 0 8372 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_75
timestamp 1586364061
transform 1 0 8004 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_16_81
timestamp 1586364061
transform 1 0 8556 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  FILLER_16_89
timestamp 1586364061
transform 1 0 9292 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_6  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 590 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 11316 0 -1 11424
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_16_103
timestamp 1586364061
transform 1 0 10580 0 -1 11424
box -38 -48 774 592
use scs8hd_conb_1  _35_
timestamp 1586364061
transform 1 0 14168 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 13248 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_130
timestamp 1586364061
transform 1 0 13064 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_134
timestamp 1586364061
transform 1 0 13432 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_8  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 774 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15640 0 -1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_304
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18124 0 -1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 17940 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_177
timestamp 1586364061
transform 1 0 17388 0 -1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_305
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 20332 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_204
timestamp 1586364061
transform 1 0 19872 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_208
timestamp 1586364061
transform 1 0 20240 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_211
timestamp 1586364061
transform 1 0 20516 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 22172 0 -1 11424
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_248
timestamp 1586364061
transform 1 0 23920 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_260
timestamp 1586364061
transform 1 0 25024 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_16_272
timestamp 1586364061
transform 1 0 26128 0 -1 11424
box -38 -48 314 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
timestamp 1586364061
transform 1 0 26588 0 -1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_306
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_296
timestamp 1586364061
transform 1 0 28336 0 -1 11424
box -38 -48 774 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
timestamp 1586364061
transform 1 0 29072 0 -1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_307
timestamp 1586364061
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_323
timestamp 1586364061
transform 1 0 30820 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_16_335
timestamp 1586364061
transform 1 0 31924 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_337
timestamp 1586364061
transform 1 0 32108 0 -1 11424
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 33856 0 -1 11424
box -38 -48 1786 592
use scs8hd_decap_6  FILLER_16_349
timestamp 1586364061
transform 1 0 33212 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_355
timestamp 1586364061
transform 1 0 33764 0 -1 11424
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_308
timestamp 1586364061
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 35788 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 37444 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_375
timestamp 1586364061
transform 1 0 35604 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_379
timestamp 1586364061
transform 1 0 35972 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_16_391
timestamp 1586364061
transform 1 0 37076 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_406
timestamp 1586364061
transform 1 0 38456 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_402
timestamp 1586364061
transform 1 0 38088 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 38272 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 37720 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_414
timestamp 1586364061
transform 1 0 39192 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 38640 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 38824 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_16_422
timestamp 1586364061
transform 1 0 39928 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_418
timestamp 1586364061
transform 1 0 39560 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 39744 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 39376 0 -1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
timestamp 1586364061
transform 1 0 40664 0 -1 11424
box -38 -48 1786 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1586364061
transform 1 0 43332 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_309
timestamp 1586364061
transform 1 0 43240 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1586364061
transform 1 0 43056 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_449
timestamp 1586364061
transform 1 0 42412 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_455
timestamp 1586364061
transform 1 0 42964 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_468
timestamp 1586364061
transform 1 0 44160 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_480
timestamp 1586364061
transform 1 0 45264 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_492
timestamp 1586364061
transform 1 0 46368 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 48852 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_504
timestamp 1586364061
transform 1 0 47472 0 -1 11424
box -38 -48 1142 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 866 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1586364061
transform 1 0 3312 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
timestamp 1586364061
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 3128 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_16
timestamp 1586364061
transform 1 0 2576 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_20
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 5612 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
timestamp 1586364061
transform 1 0 4324 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 5428 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_33
timestamp 1586364061
transform 1 0 4140 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_37
timestamp 1586364061
transform 1 0 4508 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_41
timestamp 1586364061
transform 1 0 4876 0 1 11424
box -38 -48 590 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7452 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_310
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7268 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_66
timestamp 1586364061
transform 1 0 7176 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_78
timestamp 1586364061
transform 1 0 8280 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_17_90
timestamp 1586364061
transform 1 0 9384 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_95
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_99
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 774 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_311
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_107
timestamp 1586364061
transform 1 0 10948 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 774 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13340 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_131
timestamp 1586364061
transform 1 0 13156 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 16008 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 15456 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_154
timestamp 1586364061
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_158
timestamp 1586364061
transform 1 0 15640 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_171
timestamp 1586364061
transform 1 0 16836 0 1 11424
box -38 -48 774 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18952 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_312
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 18768 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 18216 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_179
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_188
timestamp 1586364061
transform 1 0 18400 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 21252 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_213
timestamp 1586364061
transform 1 0 20700 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_217
timestamp 1586364061
transform 1 0 21068 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_221
timestamp 1586364061
transform 1 0 21436 0 1 11424
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_313
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_233
timestamp 1586364061
transform 1 0 22540 0 1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_17_241
timestamp 1586364061
transform 1 0 23276 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_264
timestamp 1586364061
transform 1 0 25392 0 1 11424
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
timestamp 1586364061
transform 1 0 28336 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_276
timestamp 1586364061
transform 1 0 26496 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_288
timestamp 1586364061
transform 1 0 27600 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_298
timestamp 1586364061
transform 1 0 28520 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_314
timestamp 1586364061
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
timestamp 1586364061
transform 1 0 28704 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_302
timestamp 1586364061
transform 1 0 28888 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_306
timestamp 1586364061
transform 1 0 29256 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_318
timestamp 1586364061
transform 1 0 30360 0 1 11424
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
timestamp 1586364061
transform 1 0 32108 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
timestamp 1586364061
transform 1 0 32476 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_330
timestamp 1586364061
transform 1 0 31464 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_336
timestamp 1586364061
transform 1 0 32016 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_339
timestamp 1586364061
transform 1 0 32292 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_343
timestamp 1586364061
transform 1 0 32660 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_315
timestamp 1586364061
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
timestamp 1586364061
transform 1 0 34592 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
timestamp 1586364061
transform 1 0 35052 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
timestamp 1586364061
transform 1 0 34224 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_355
timestamp 1586364061
transform 1 0 33764 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_359
timestamp 1586364061
transform 1 0 34132 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_362
timestamp 1586364061
transform 1 0 34408 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_367
timestamp 1586364061
transform 1 0 34868 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_371
timestamp 1586364061
transform 1 0 35236 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 35420 0 1 11424
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 37628 0 1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 37444 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 35972 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 37076 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_377
timestamp 1586364061
transform 1 0 35788 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_381
timestamp 1586364061
transform 1 0 36156 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_389
timestamp 1586364061
transform 1 0 36892 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_393
timestamp 1586364061
transform 1 0 37260 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 39560 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 39928 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_416
timestamp 1586364061
transform 1 0 39376 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_420
timestamp 1586364061
transform 1 0 39744 0 1 11424
box -38 -48 222 592
use scs8hd_or2_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
timestamp 1586364061
transform 1 0 40756 0 1 11424
box -38 -48 498 592
use scs8hd_tapvpwrvgnd_1  PHY_316
timestamp 1586364061
transform 1 0 40388 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
timestamp 1586364061
transform 1 0 41400 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 41768 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_424
timestamp 1586364061
transform 1 0 40112 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_17_428
timestamp 1586364061
transform 1 0 40480 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_436
timestamp 1586364061
transform 1 0 41216 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_440
timestamp 1586364061
transform 1 0 41584 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_444
timestamp 1586364061
transform 1 0 41952 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_456
timestamp 1586364061
transform 1 0 43056 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_468
timestamp 1586364061
transform 1 0 44160 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_317
timestamp 1586364061
transform 1 0 46000 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
timestamp 1586364061
transform 1 0 44988 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
timestamp 1586364061
transform 1 0 45356 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_476
timestamp 1586364061
transform 1 0 44896 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_479
timestamp 1586364061
transform 1 0 45172 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_483
timestamp 1586364061
transform 1 0 45540 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_487
timestamp 1586364061
transform 1 0 45908 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_489
timestamp 1586364061
transform 1 0 46092 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 48852 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 47472 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_501
timestamp 1586364061
transform 1 0 47196 0 1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_17_506
timestamp 1586364061
transform 1 0 47656 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_514
timestamp 1586364061
transform 1 0 48392 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
timestamp 1586364061
transform 1 0 1472 0 -1 12512
box -38 -48 1786 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_318
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1586364061
transform 1 0 6532 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 7544 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 6348 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_51
timestamp 1586364061
transform 1 0 5796 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_72
timestamp 1586364061
transform 1 0 7728 0 -1 12512
box -38 -48 774 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_319
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_82
timestamp 1586364061
transform 1 0 8648 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_90
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_112
timestamp 1586364061
transform 1 0 11408 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_124
timestamp 1586364061
transform 1 0 12512 0 -1 12512
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 13524 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_132
timestamp 1586364061
transform 1 0 13248 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_137
timestamp 1586364061
transform 1 0 13708 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_18_149
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_320
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 16008 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_18_164
timestamp 1586364061
transform 1 0 16192 0 -1 12512
box -38 -48 1142 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 17940 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 18952 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 19320 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_176
timestamp 1586364061
transform 1 0 17296 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_182
timestamp 1586364061
transform 1 0 17848 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_192
timestamp 1586364061
transform 1 0 18768 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_196
timestamp 1586364061
transform 1 0 19136 0 -1 12512
box -38 -48 222 592
use scs8hd_conb_1  _38_
timestamp 1586364061
transform 1 0 19504 0 -1 12512
box -38 -48 314 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_321
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 19964 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 20332 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_203
timestamp 1586364061
transform 1 0 19780 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_207
timestamp 1586364061
transform 1 0 20148 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_211
timestamp 1586364061
transform 1 0 20516 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 23644 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_234
timestamp 1586364061
transform 1 0 22632 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_18_242
timestamp 1586364061
transform 1 0 23368 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_247
timestamp 1586364061
transform 1 0 23828 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_259
timestamp 1586364061
transform 1 0 24932 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_18_271
timestamp 1586364061
transform 1 0 26036 0 -1 12512
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
timestamp 1586364061
transform 1 0 28336 0 -1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_322
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_288
timestamp 1586364061
transform 1 0 27600 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_18_315
timestamp 1586364061
transform 1 0 30084 0 -1 12512
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
timestamp 1586364061
transform 1 0 32108 0 -1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_323
timestamp 1586364061
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 31832 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 31464 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_327
timestamp 1586364061
transform 1 0 31188 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_332
timestamp 1586364061
transform 1 0 31648 0 -1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
timestamp 1586364061
transform 1 0 34592 0 -1 12512
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
timestamp 1586364061
transform 1 0 34408 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_clkbuf_1_1__f_clk_A
timestamp 1586364061
transform 1 0 34040 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_356
timestamp 1586364061
transform 1 0 33856 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_360
timestamp 1586364061
transform 1 0 34224 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_324
timestamp 1586364061
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 36800 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 37444 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_383
timestamp 1586364061
transform 1 0 36340 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_387
timestamp 1586364061
transform 1 0 36708 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_390
timestamp 1586364061
transform 1 0 36984 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_394
timestamp 1586364061
transform 1 0 37352 0 -1 12512
box -38 -48 130 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1586364061
transform 1 0 39560 0 -1 12512
box -38 -48 866 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 37996 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  FILLER_18_398
timestamp 1586364061
transform 1 0 37720 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_410
timestamp 1586364061
transform 1 0 38824 0 -1 12512
box -38 -48 774 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 41124 0 -1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
timestamp 1586364061
transform 1 0 40756 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_427
timestamp 1586364061
transform 1 0 40388 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_433
timestamp 1586364061
transform 1 0 40940 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_439
timestamp 1586364061
transform 1 0 41492 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_325
timestamp 1586364061
transform 1 0 43240 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 43976 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 44344 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_451
timestamp 1586364061
transform 1 0 42596 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_457
timestamp 1586364061
transform 1 0 43148 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_18_459
timestamp 1586364061
transform 1 0 43332 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_465
timestamp 1586364061
transform 1 0 43884 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_468
timestamp 1586364061
transform 1 0 44160 0 -1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
timestamp 1586364061
transform 1 0 44988 0 -1 12512
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_18_472
timestamp 1586364061
transform 1 0 44528 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_476
timestamp 1586364061
transform 1 0 44896 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_496
timestamp 1586364061
transform 1 0 46736 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 47472 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 48852 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
timestamp 1586364061
transform 1 0 46920 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_500
timestamp 1586364061
transform 1 0 47104 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_18_508
timestamp 1586364061
transform 1 0 47840 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
timestamp 1586364061
transform 1 0 1932 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
timestamp 1586364061
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_6  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_4  FILLER_19_23
timestamp 1586364061
transform 1 0 3220 0 1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_11
timestamp 1586364061
transform 1 0 2116 0 -1 13600
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
timestamp 1586364061
transform 1 0 1472 0 1 12512
box -38 -48 1786 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
timestamp 1586364061
transform 1 0 4232 0 1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_334
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
timestamp 1586364061
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
timestamp 1586364061
transform 1 0 3680 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_30
timestamp 1586364061
transform 1 0 3864 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_41
timestamp 1586364061
transform 1 0 4876 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_20_53
timestamp 1586364061
transform 1 0 5980 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_19_60
timestamp 1586364061
transform 1 0 6624 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 6440 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_326
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_71
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 6440 0 -1 13600
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 8464 0 1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_335
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 8280 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_75
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_99
timestamp 1586364061
transform 1 0 10212 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_77
timestamp 1586364061
transform 1 0 8188 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_20_89
timestamp 1586364061
transform 1 0 9292 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_327
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_111
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_19_119
timestamp 1586364061
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_105
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_117
timestamp 1586364061
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_129
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_141
timestamp 1586364061
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_336
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_159
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_171
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_166
timestamp 1586364061
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_328
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_196
timestamp 1586364061
transform 1 0 19136 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_20_190
timestamp 1586364061
transform 1 0 18584 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_195
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_192
timestamp 1586364061
transform 1 0 18768 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 19228 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_12  FILLER_20_178
timestamp 1586364061
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 19872 0 1 12512
box -38 -48 2246 592
use scs8hd_tapvpwrvgnd_1  PHY_337
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 19688 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 20240 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_199
timestamp 1586364061
transform 1 0 19412 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_206
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_210
timestamp 1586364061
transform 1 0 20424 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_329
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_228
timestamp 1586364061
transform 1 0 22080 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_19_240
timestamp 1586364061
transform 1 0 23184 0 1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_227
timestamp 1586364061
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_239
timestamp 1586364061
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_251
timestamp 1586364061
transform 1 0 24196 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_263
timestamp 1586364061
transform 1 0 25300 0 -1 13600
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
timestamp 1586364061
transform 1 0 27140 0 -1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_338
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
timestamp 1586364061
transform 1 0 27140 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
timestamp 1586364061
transform 1 0 27508 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_281
timestamp 1586364061
transform 1 0 26956 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_285
timestamp 1586364061
transform 1 0 27324 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_289
timestamp 1586364061
transform 1 0 27692 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_20_282
timestamp 1586364061
transform 1 0 27048 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_308
timestamp 1586364061
transform 1 0 29440 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_302
timestamp 1586364061
transform 1 0 28888 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_4  FILLER_19_306
timestamp 1586364061
transform 1 0 29256 0 1 12512
box -38 -48 406 592
use scs8hd_decap_4  FILLER_19_301
timestamp 1586364061
transform 1 0 28796 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 29256 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
timestamp 1586364061
transform 1 0 29624 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_330
timestamp 1586364061
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_316
timestamp 1586364061
transform 1 0 30176 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_312
timestamp 1586364061
transform 1 0 29808 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
timestamp 1586364061
transform 1 0 29992 0 1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
timestamp 1586364061
transform 1 0 29624 0 -1 13600
box -38 -48 1786 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1586364061
transform 1 0 32108 0 -1 13600
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
timestamp 1586364061
transform 1 0 32936 0 1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_339
timestamp 1586364061
transform 1 0 32016 0 -1 13600
box -38 -48 130 592
use scs8hd_clkbuf_16  clkbuf_0_clk
timestamp 1586364061
transform 1 0 31096 0 1 12512
box -38 -48 1878 592
use scs8hd_diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1586364061
transform 1 0 30912 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 31832 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_329
timestamp 1586364061
transform 1 0 31372 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_333
timestamp 1586364061
transform 1 0 31740 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_346
timestamp 1586364061
transform 1 0 32936 0 -1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
timestamp 1586364061
transform 1 0 34868 0 1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_331
timestamp 1586364061
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use scs8hd_clkbuf_16  clkbuf_1_1__f_clk
timestamp 1586364061
transform 1 0 33764 0 -1 13600
box -38 -48 1878 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
timestamp 1586364061
transform 1 0 33120 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
timestamp 1586364061
transform 1 0 33488 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_365
timestamp 1586364061
transform 1 0 34684 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_350
timestamp 1586364061
transform 1 0 33304 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_354
timestamp 1586364061
transform 1 0 33672 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_383
timestamp 1586364061
transform 1 0 36340 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_379
timestamp 1586364061
transform 1 0 35972 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 36156 0 -1 13600
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 35604 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_394
timestamp 1586364061
transform 1 0 37352 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_390
timestamp 1586364061
transform 1 0 36984 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_387
timestamp 1586364061
transform 1 0 36708 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_386
timestamp 1586364061
transform 1 0 36616 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 37444 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 36800 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_340
timestamp 1586364061
transform 1 0 37628 0 -1 13600
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 36800 0 1 12512
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_20_407
timestamp 1586364061
transform 1 0 38548 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_407
timestamp 1586364061
transform 1 0 38548 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 38732 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 37720 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_6  FILLER_19_421
timestamp 1586364061
transform 1 0 39836 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_417
timestamp 1586364061
transform 1 0 39468 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_411
timestamp 1586364061
transform 1 0 38916 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
timestamp 1586364061
transform 1 0 39652 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
timestamp 1586364061
transform 1 0 39284 0 1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
timestamp 1586364061
transform 1 0 39284 0 -1 13600
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_20_434
timestamp 1586364061
transform 1 0 41032 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_432
timestamp 1586364061
transform 1 0 40848 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_428
timestamp 1586364061
transform 1 0 40480 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
timestamp 1586364061
transform 1 0 40940 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_332
timestamp 1586364061
transform 1 0 40388 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_435
timestamp 1586364061
transform 1 0 41124 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
timestamp 1586364061
transform 1 0 41216 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
timestamp 1586364061
transform 1 0 41308 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_438
timestamp 1586364061
transform 1 0 41400 0 -1 13600
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
timestamp 1586364061
transform 1 0 41492 0 1 12512
box -38 -48 1786 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1586364061
transform 1 0 43976 0 1 12512
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
timestamp 1586364061
transform 1 0 43332 0 -1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_341
timestamp 1586364061
transform 1 0 43240 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
timestamp 1586364061
transform 1 0 43424 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
timestamp 1586364061
transform 1 0 43792 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 43056 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_458
timestamp 1586364061
transform 1 0 43240 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_462
timestamp 1586364061
transform 1 0 43608 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_450
timestamp 1586364061
transform 1 0 42504 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_8  FILLER_20_478
timestamp 1586364061
transform 1 0 45080 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_484
timestamp 1586364061
transform 1 0 45632 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_479
timestamp 1586364061
transform 1 0 45172 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_475
timestamp 1586364061
transform 1 0 44804 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 44988 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
timestamp 1586364061
transform 1 0 45448 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_486
timestamp 1586364061
transform 1 0 45816 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
timestamp 1586364061
transform 1 0 45908 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
timestamp 1586364061
transform 1 0 45816 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_333
timestamp 1586364061
transform 1 0 46000 0 1 12512
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
timestamp 1586364061
transform 1 0 46092 0 -1 13600
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
timestamp 1586364061
transform 1 0 46092 0 1 12512
box -38 -48 1786 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 48852 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 48852 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_19_508
timestamp 1586364061
transform 1 0 47840 0 1 12512
box -38 -48 774 592
use scs8hd_decap_8  FILLER_20_508
timestamp 1586364061
transform 1 0 47840 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_31
timestamp 1586364061
transform 1 0 3956 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_34
timestamp 1586364061
transform 1 0 4232 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_46
timestamp 1586364061
transform 1 0 5336 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_342
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_21_58
timestamp 1586364061
transform 1 0 6440 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_21_74
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 8280 0 1 13600
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 8096 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_97
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_343
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_109
timestamp 1586364061
transform 1 0 11132 0 1 13600
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_21_121
timestamp 1586364061
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_135
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_147
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_159
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_171
timestamp 1586364061
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_344
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 19136 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_21_198
timestamp 1586364061
transform 1 0 19320 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 19688 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 19504 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_211
timestamp 1586364061
transform 1 0 20516 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_223
timestamp 1586364061
transform 1 0 21620 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_345
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_21_235
timestamp 1586364061
transform 1 0 22724 0 1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_21_243
timestamp 1586364061
transform 1 0 23460 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_257
timestamp 1586364061
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1586364061
transform 1 0 27508 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
timestamp 1586364061
transform 1 0 26588 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
timestamp 1586364061
transform 1 0 26956 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 27324 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 28520 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_279
timestamp 1586364061
transform 1 0 26772 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_283
timestamp 1586364061
transform 1 0 27140 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_296
timestamp 1586364061
transform 1 0 28336 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1586364061
transform 1 0 29624 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_346
timestamp 1586364061
transform 1 0 29164 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 29440 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 28980 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_300
timestamp 1586364061
transform 1 0 28704 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_306
timestamp 1586364061
transform 1 0 29256 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_319
timestamp 1586364061
transform 1 0 30452 0 1 13600
box -38 -48 406 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1586364061
transform 1 0 31648 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 32660 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1586364061
transform 1 0 33028 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
timestamp 1586364061
transform 1 0 30912 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 31464 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_323
timestamp 1586364061
transform 1 0 30820 0 1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_21_326
timestamp 1586364061
transform 1 0 31096 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_341
timestamp 1586364061
transform 1 0 32476 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_345
timestamp 1586364061
transform 1 0 32844 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1586364061
transform 1 0 33212 0 1 13600
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
timestamp 1586364061
transform 1 0 34868 0 1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_347
timestamp 1586364061
transform 1 0 34776 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
timestamp 1586364061
transform 1 0 34592 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
timestamp 1586364061
transform 1 0 34224 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_358
timestamp 1586364061
transform 1 0 34040 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_362
timestamp 1586364061
transform 1 0 34408 0 1 13600
box -38 -48 222 592
use scs8hd_conb_1  _55_
timestamp 1586364061
transform 1 0 37352 0 1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_21_386
timestamp 1586364061
transform 1 0 36616 0 1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_21_397
timestamp 1586364061
transform 1 0 37628 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 37812 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 38180 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 39836 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 39468 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_401
timestamp 1586364061
transform 1 0 37996 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_405
timestamp 1586364061
transform 1 0 38364 0 1 13600
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_21_419
timestamp 1586364061
transform 1 0 39652 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
timestamp 1586364061
transform 1 0 40480 0 1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_348
timestamp 1586364061
transform 1 0 40388 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
timestamp 1586364061
transform 1 0 40204 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_423
timestamp 1586364061
transform 1 0 40020 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_447
timestamp 1586364061
transform 1 0 42228 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
timestamp 1586364061
transform 1 0 43516 0 1 13600
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
timestamp 1586364061
transform 1 0 43332 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 42964 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
timestamp 1586364061
transform 1 0 42412 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_451
timestamp 1586364061
transform 1 0 42596 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_457
timestamp 1586364061
transform 1 0 43148 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1586364061
transform 1 0 46092 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_349
timestamp 1586364061
transform 1 0 46000 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1586364061
transform 1 0 45816 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 45448 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_480
timestamp 1586364061
transform 1 0 45264 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_484
timestamp 1586364061
transform 1 0 45632 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 48852 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 47104 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_498
timestamp 1586364061
transform 1 0 46920 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_502
timestamp 1586364061
transform 1 0 47288 0 1 13600
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_21_514
timestamp 1586364061
transform 1 0 48392 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_350
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_44
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_56
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_22_68
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_351
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 8280 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_76
timestamp 1586364061
transform 1 0 8096 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_80
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_105
timestamp 1586364061
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_117
timestamp 1586364061
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_129
timestamp 1586364061
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_141
timestamp 1586364061
transform 1 0 14076 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_352
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_166
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_178
timestamp 1586364061
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_190
timestamp 1586364061
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_353
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 19688 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_204
timestamp 1586364061
transform 1 0 19872 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_212
timestamp 1586364061
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_239
timestamp 1586364061
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_251
timestamp 1586364061
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_263
timestamp 1586364061
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
timestamp 1586364061
transform 1 0 26588 0 -1 14688
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_354
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_296
timestamp 1586364061
transform 1 0 28336 0 -1 14688
box -38 -48 406 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1586364061
transform 1 0 29256 0 -1 14688
box -38 -48 866 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
timestamp 1586364061
transform 1 0 30084 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 29072 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
timestamp 1586364061
transform 1 0 30636 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 28704 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_302
timestamp 1586364061
transform 1 0 28888 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_319
timestamp 1586364061
transform 1 0 30452 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_323
timestamp 1586364061
transform 1 0 30820 0 -1 14688
box -38 -48 130 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
timestamp 1586364061
transform 1 0 30912 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_332
timestamp 1586364061
transform 1 0 31648 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_328
timestamp 1586364061
transform 1 0 31280 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 31464 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_337
timestamp 1586364061
transform 1 0 32108 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 31832 0 -1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_355
timestamp 1586364061
transform 1 0 32016 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_342
timestamp 1586364061
transform 1 0 32568 0 -1 14688
box -38 -48 314 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 32200 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_347
timestamp 1586364061
transform 1 0 33028 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 32844 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_359
timestamp 1586364061
transform 1 0 34132 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_355
timestamp 1586364061
transform 1 0 33764 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_351
timestamp 1586364061
transform 1 0 33396 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1586364061
transform 1 0 33948 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 33580 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1586364061
transform 1 0 33212 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_369
timestamp 1586364061
transform 1 0 35052 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_365
timestamp 1586364061
transform 1 0 34684 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1586364061
transform 1 0 34500 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
timestamp 1586364061
transform 1 0 35144 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_372
timestamp 1586364061
transform 1 0 35328 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_356
timestamp 1586364061
transform 1 0 37628 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_384
timestamp 1586364061
transform 1 0 36432 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_22_396
timestamp 1586364061
transform 1 0 37536 0 -1 14688
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 37720 0 -1 14688
box -38 -48 1786 592
use scs8hd_decap_6  FILLER_22_417
timestamp 1586364061
transform 1 0 39468 0 -1 14688
box -38 -48 590 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1586364061
transform 1 0 40204 0 -1 14688
box -38 -48 866 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
timestamp 1586364061
transform 1 0 42044 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 41584 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 40020 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_434
timestamp 1586364061
transform 1 0 41032 0 -1 14688
box -38 -48 590 592
use scs8hd_decap_3  FILLER_22_442
timestamp 1586364061
transform 1 0 41768 0 -1 14688
box -38 -48 314 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1586364061
transform 1 0 43792 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_357
timestamp 1586364061
transform 1 0 43240 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
timestamp 1586364061
transform 1 0 43516 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 43056 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_449
timestamp 1586364061
transform 1 0 42412 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_455
timestamp 1586364061
transform 1 0 42964 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_459
timestamp 1586364061
transform 1 0 43332 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_463
timestamp 1586364061
transform 1 0 43700 0 -1 14688
box -38 -48 130 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 46736 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1586364061
transform 1 0 46092 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1586364061
transform 1 0 46460 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_473
timestamp 1586364061
transform 1 0 44620 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_22_485
timestamp 1586364061
transform 1 0 45724 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_491
timestamp 1586364061
transform 1 0 46276 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_495
timestamp 1586364061
transform 1 0 46644 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 48852 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_500
timestamp 1586364061
transform 1 0 47104 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_22_512
timestamp 1586364061
transform 1 0 48208 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_358
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_59
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_74
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_86
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_98
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_359
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_110
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_147
timestamp 1586364061
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_159
timestamp 1586364061
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_171
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_360
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_196
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_208
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_220
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_361
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_232
timestamp 1586364061
transform 1 0 22448 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_257
timestamp 1586364061
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_269
timestamp 1586364061
transform 1 0 25852 0 1 14688
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 28152 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 28520 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 27508 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_281
timestamp 1586364061
transform 1 0 26956 0 1 14688
box -38 -48 590 592
use scs8hd_decap_4  FILLER_23_289
timestamp 1586364061
transform 1 0 27692 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_293
timestamp 1586364061
transform 1 0 28060 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_296
timestamp 1586364061
transform 1 0 28336 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1586364061
transform 1 0 30268 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_362
timestamp 1586364061
transform 1 0 29164 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 30084 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 29624 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 28980 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_300
timestamp 1586364061
transform 1 0 28704 0 1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_23_306
timestamp 1586364061
transform 1 0 29256 0 1 14688
box -38 -48 406 592
use scs8hd_decap_3  FILLER_23_312
timestamp 1586364061
transform 1 0 29808 0 1 14688
box -38 -48 314 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1586364061
transform 1 0 31832 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 31648 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 32844 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 31280 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_326
timestamp 1586364061
transform 1 0 31096 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_330
timestamp 1586364061
transform 1 0 31464 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_343
timestamp 1586364061
transform 1 0 32660 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_347
timestamp 1586364061
transform 1 0 33028 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_359
timestamp 1586364061
transform 1 0 34132 0 1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_23_355
timestamp 1586364061
transform 1 0 33764 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
timestamp 1586364061
transform 1 0 33212 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1586364061
transform 1 0 34224 0 1 14688
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
timestamp 1586364061
transform 1 0 33396 0 1 14688
box -38 -48 406 592
use scs8hd_decap_3  FILLER_23_367
timestamp 1586364061
transform 1 0 34868 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_362
timestamp 1586364061
transform 1 0 34408 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
timestamp 1586364061
transform 1 0 34592 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_363
timestamp 1586364061
transform 1 0 34776 0 1 14688
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
timestamp 1586364061
transform 1 0 35144 0 1 14688
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_23_389
timestamp 1586364061
transform 1 0 36892 0 1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_23_397
timestamp 1586364061
transform 1 0 37628 0 1 14688
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
timestamp 1586364061
transform 1 0 37904 0 1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
timestamp 1586364061
transform 1 0 37720 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_419
timestamp 1586364061
transform 1 0 39652 0 1 14688
box -38 -48 590 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1586364061
transform 1 0 41584 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_364
timestamp 1586364061
transform 1 0 40388 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 40664 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 41032 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 41400 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 40204 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_428
timestamp 1586364061
transform 1 0 40480 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_432
timestamp 1586364061
transform 1 0 40848 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_436
timestamp 1586364061
transform 1 0 41216 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1586364061
transform 1 0 43148 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 44160 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 42964 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 42596 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_449
timestamp 1586364061
transform 1 0 42412 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_453
timestamp 1586364061
transform 1 0 42780 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_466
timestamp 1586364061
transform 1 0 43976 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_470
timestamp 1586364061
transform 1 0 44344 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_478
timestamp 1586364061
transform 1 0 45080 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_474
timestamp 1586364061
transform 1 0 44712 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 44896 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 44528 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_489
timestamp 1586364061
transform 1 0 46092 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
timestamp 1586364061
transform 1 0 45816 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_365
timestamp 1586364061
transform 1 0 46000 0 1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_23_493
timestamp 1586364061
transform 1 0 46460 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
timestamp 1586364061
transform 1 0 46276 0 1 14688
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 46736 0 1 14688
box -38 -48 406 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 48852 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 47288 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_500
timestamp 1586364061
transform 1 0 47104 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_504
timestamp 1586364061
transform 1 0 47472 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_366
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_56
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_367
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_105
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_117
timestamp 1586364061
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_129
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_141
timestamp 1586364061
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_368
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_166
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_178
timestamp 1586364061
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_190
timestamp 1586364061
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_369
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_202
timestamp 1586364061
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_239
timestamp 1586364061
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 25484 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_251
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_24_263
timestamp 1586364061
transform 1 0 25300 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_267
timestamp 1586364061
transform 1 0 25668 0 -1 15776
box -38 -48 774 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 28152 0 -1 15776
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_370
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 26864 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_282
timestamp 1586364061
transform 1 0 27048 0 -1 15776
box -38 -48 1142 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 30636 0 -1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 30268 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_313
timestamp 1586364061
transform 1 0 29900 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_319
timestamp 1586364061
transform 1 0 30452 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_329
timestamp 1586364061
transform 1 0 31372 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_325
timestamp 1586364061
transform 1 0 31004 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 31648 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 31188 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_341
timestamp 1586364061
transform 1 0 32476 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_337
timestamp 1586364061
transform 1 0 32108 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_334
timestamp 1586364061
transform 1 0 31832 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 32292 0 -1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_371
timestamp 1586364061
transform 1 0 32016 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_345
timestamp 1586364061
transform 1 0 32844 0 -1 15776
box -38 -48 130 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1586364061
transform 1 0 32936 0 -1 15776
box -38 -48 866 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1586364061
transform 1 0 34500 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1586364061
transform 1 0 34316 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_355
timestamp 1586364061
transform 1 0 33764 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_2  FILLER_24_372
timestamp 1586364061
transform 1 0 35328 0 -1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_372
timestamp 1586364061
transform 1 0 37628 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
timestamp 1586364061
transform 1 0 35512 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_376
timestamp 1586364061
transform 1 0 35696 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_24_388
timestamp 1586364061
transform 1 0 36800 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_1  FILLER_24_396
timestamp 1586364061
transform 1 0 37536 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 38824 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 39192 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
timestamp 1586364061
transform 1 0 37904 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_398
timestamp 1586364061
transform 1 0 37720 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_402
timestamp 1586364061
transform 1 0 38088 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_412
timestamp 1586364061
transform 1 0 39008 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_416
timestamp 1586364061
transform 1 0 39376 0 -1 15776
box -38 -48 1142 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1586364061
transform 1 0 40664 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 40480 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 41676 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_439
timestamp 1586364061
transform 1 0 41492 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_443
timestamp 1586364061
transform 1 0 41860 0 -1 15776
box -38 -48 1142 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1586364061
transform 1 0 43332 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_373
timestamp 1586364061
transform 1 0 43240 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 44436 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_455
timestamp 1586364061
transform 1 0 42964 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_468
timestamp 1586364061
transform 1 0 44160 0 -1 15776
box -38 -48 314 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
timestamp 1586364061
transform 1 0 46092 0 -1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
timestamp 1586364061
transform 1 0 45172 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 44804 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_473
timestamp 1586364061
transform 1 0 44620 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_477
timestamp 1586364061
transform 1 0 44988 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_481
timestamp 1586364061
transform 1 0 45356 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 48852 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_508
timestamp 1586364061
transform 1 0 47840 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_374
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_74
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_86
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_98
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_375
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_110
timestamp 1586364061
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_147
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_159
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_171
timestamp 1586364061
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_376
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_196
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_208
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_220
timestamp 1586364061
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_377
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_232
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 25484 0 1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 25300 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_257
timestamp 1586364061
transform 1 0 24748 0 1 15776
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 27416 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 28244 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_284
timestamp 1586364061
transform 1 0 27232 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_288
timestamp 1586364061
transform 1 0 27600 0 1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_25_294
timestamp 1586364061
transform 1 0 28152 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_297
timestamp 1586364061
transform 1 0 28428 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1586364061
transform 1 0 29256 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_378
timestamp 1586364061
transform 1 0 29164 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 28980 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 28612 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 30268 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 30636 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_301
timestamp 1586364061
transform 1 0 28796 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_315
timestamp 1586364061
transform 1 0 30084 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_319
timestamp 1586364061
transform 1 0 30452 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1586364061
transform 1 0 30820 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
timestamp 1586364061
transform 1 0 32108 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
timestamp 1586364061
transform 1 0 32476 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1586364061
transform 1 0 33028 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_332
timestamp 1586364061
transform 1 0 31648 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_336
timestamp 1586364061
transform 1 0 32016 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_339
timestamp 1586364061
transform 1 0 32292 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_343
timestamp 1586364061
transform 1 0 32660 0 1 15776
box -38 -48 406 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1586364061
transform 1 0 33212 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_379
timestamp 1586364061
transform 1 0 34776 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
timestamp 1586364061
transform 1 0 34224 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
timestamp 1586364061
transform 1 0 35328 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
timestamp 1586364061
transform 1 0 34592 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_358
timestamp 1586364061
transform 1 0 34040 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_362
timestamp 1586364061
transform 1 0 34408 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_367
timestamp 1586364061
transform 1 0 34868 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_371
timestamp 1586364061
transform 1 0 35236 0 1 15776
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
timestamp 1586364061
transform 1 0 35512 0 1 15776
box -38 -48 1786 592
use scs8hd_decap_6  FILLER_25_393
timestamp 1586364061
transform 1 0 37260 0 1 15776
box -38 -48 590 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1586364061
transform 1 0 38824 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 39836 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 38272 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 38640 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 37904 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_399
timestamp 1586364061
transform 1 0 37812 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_402
timestamp 1586364061
transform 1 0 38088 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_406
timestamp 1586364061
transform 1 0 38456 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_419
timestamp 1586364061
transform 1 0 39652 0 1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 40664 0 1 15776
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_380
timestamp 1586364061
transform 1 0 40388 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 40204 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_423
timestamp 1586364061
transform 1 0 40020 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_428
timestamp 1586364061
transform 1 0 40480 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_454
timestamp 1586364061
transform 1 0 42872 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_449
timestamp 1586364061
transform 1 0 42412 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 42688 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
timestamp 1586364061
transform 1 0 43056 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_466
timestamp 1586364061
transform 1 0 43976 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_462
timestamp 1586364061
transform 1 0 43608 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 43792 0 1 15776
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
timestamp 1586364061
transform 1 0 43240 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_470
timestamp 1586364061
transform 1 0 44344 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 44160 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1586364061
transform 1 0 44436 0 1 15776
box -38 -48 866 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1586364061
transform 1 0 46092 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_381
timestamp 1586364061
transform 1 0 46000 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
timestamp 1586364061
transform 1 0 45448 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1586364061
transform 1 0 45816 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_480
timestamp 1586364061
transform 1 0 45264 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_484
timestamp 1586364061
transform 1 0 45632 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 48852 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1586364061
transform 1 0 47104 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1586364061
transform 1 0 47472 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_498
timestamp 1586364061
transform 1 0 46920 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_502
timestamp 1586364061
transform 1 0 47288 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_506
timestamp 1586364061
transform 1 0 47656 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_514
timestamp 1586364061
transform 1 0 48392 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_382
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_390
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_383
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_80
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_86
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_98
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_391
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_105
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_117
timestamp 1586364061
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_110
timestamp 1586364061
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_129
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_141
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_135
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_147
timestamp 1586364061
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_384
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_166
timestamp 1586364061
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_159
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_171
timestamp 1586364061
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_392
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_178
timestamp 1586364061
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_190
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_385
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_202
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_220
timestamp 1586364061
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_232
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_240
timestamp 1586364061
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_245
timestamp 1586364061
transform 1 0 23644 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_26_239
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23736 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_393
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_248
timestamp 1586364061
transform 1 0 23920 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 23736 0 1 16864
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 26220 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 25852 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_260
timestamp 1586364061
transform 1 0 25024 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_26_272
timestamp 1586364061
transform 1 0 26128 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_27_265
timestamp 1586364061
transform 1 0 25484 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_271
timestamp 1586364061
transform 1 0 26036 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1586364061
transform 1 0 26404 0 1 16864
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 26864 0 -1 16864
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_386
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 26680 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_284
timestamp 1586364061
transform 1 0 27232 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_296
timestamp 1586364061
transform 1 0 28336 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_306
timestamp 1586364061
transform 1 0 29256 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_304
timestamp 1586364061
transform 1 0 29072 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_303
timestamp 1586364061
transform 1 0 28980 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_299
timestamp 1586364061
transform 1 0 28612 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 28796 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 29164 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_394
timestamp 1586364061
transform 1 0 29164 0 1 16864
box -38 -48 130 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1586364061
transform 1 0 29348 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_3  FILLER_27_310
timestamp 1586364061
transform 1 0 29624 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_316
timestamp 1586364061
transform 1 0 30176 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 29440 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 29900 0 1 16864
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 30084 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_319
timestamp 1586364061
transform 1 0 30452 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_320
timestamp 1586364061
transform 1 0 30544 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 30728 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 30360 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 30636 0 1 16864
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 30912 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_27_323
timestamp 1586364061
transform 1 0 30820 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_327
timestamp 1586364061
transform 1 0 31188 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 31648 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 31280 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 31464 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_328
timestamp 1586364061
transform 1 0 31280 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_332
timestamp 1586364061
transform 1 0 31648 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_330
timestamp 1586364061
transform 1 0 31464 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
timestamp 1586364061
transform 1 0 31832 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_342
timestamp 1586364061
transform 1 0 32568 0 -1 16864
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_387
timestamp 1586364061
transform 1 0 32016 0 -1 16864
box -38 -48 130 592
use scs8hd_or2_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
timestamp 1586364061
transform 1 0 32108 0 -1 16864
box -38 -48 498 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
timestamp 1586364061
transform 1 0 31832 0 1 16864
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_27_353
timestamp 1586364061
transform 1 0 33580 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_351
timestamp 1586364061
transform 1 0 33396 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_348
timestamp 1586364061
transform 1 0 33120 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1586364061
transform 1 0 33580 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1586364061
transform 1 0 33212 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_371
timestamp 1586364061
transform 1 0 35236 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_367
timestamp 1586364061
transform 1 0 34868 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_361
timestamp 1586364061
transform 1 0 34316 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 34592 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 35052 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_395
timestamp 1586364061
transform 1 0 34776 0 1 16864
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
timestamp 1586364061
transform 1 0 33764 0 -1 16864
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 35420 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_387
timestamp 1586364061
transform 1 0 36708 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_394
timestamp 1586364061
transform 1 0 37352 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_6  FILLER_26_386
timestamp 1586364061
transform 1 0 36616 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 37168 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 36984 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_388
timestamp 1586364061
transform 1 0 37628 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_375
timestamp 1586364061
transform 1 0 35604 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_374
timestamp 1586364061
transform 1 0 35512 0 -1 16864
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 37168 0 1 16864
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 38272 0 -1 16864
box -38 -48 1786 592
use scs8hd_decap_6  FILLER_26_398
timestamp 1586364061
transform 1 0 37720 0 -1 16864
box -38 -48 590 592
use scs8hd_decap_12  FILLER_27_411
timestamp 1586364061
transform 1 0 38916 0 1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_27_432
timestamp 1586364061
transform 1 0 40848 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_428
timestamp 1586364061
transform 1 0 40480 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_423
timestamp 1586364061
transform 1 0 40020 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_423
timestamp 1586364061
transform 1 0 40020 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 40204 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 40940 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 40572 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_396
timestamp 1586364061
transform 1 0 40388 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_444
timestamp 1586364061
transform 1 0 41952 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 42136 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1586364061
transform 1 0 41124 0 1 16864
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 40756 0 -1 16864
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_27_452
timestamp 1586364061
transform 1 0 42688 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_448
timestamp 1586364061
transform 1 0 42320 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_450
timestamp 1586364061
transform 1 0 42504 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 43056 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 42504 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 42872 0 1 16864
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 43056 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_464
timestamp 1586364061
transform 1 0 43792 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_460
timestamp 1586364061
transform 1 0 43424 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 43976 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 43608 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_389
timestamp 1586364061
transform 1 0 43240 0 -1 16864
box -38 -48 130 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1586364061
transform 1 0 43332 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_26_468
timestamp 1586364061
transform 1 0 44160 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
timestamp 1586364061
transform 1 0 44344 0 -1 16864
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
timestamp 1586364061
transform 1 0 44160 0 1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1586364061
transform 1 0 44712 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 44712 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_472
timestamp 1586364061
transform 1 0 44528 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_472
timestamp 1586364061
transform 1 0 44528 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1586364061
transform 1 0 45080 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_476
timestamp 1586364061
transform 1 0 44896 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_476
timestamp 1586364061
transform 1 0 44896 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
timestamp 1586364061
transform 1 0 45448 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_480
timestamp 1586364061
transform 1 0 45264 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_484
timestamp 1586364061
transform 1 0 45632 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
timestamp 1586364061
transform 1 0 45816 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_397
timestamp 1586364061
transform 1 0 46000 0 1 16864
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
timestamp 1586364061
transform 1 0 46092 0 1 16864
box -38 -48 1786 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
timestamp 1586364061
transform 1 0 45172 0 -1 16864
box -38 -48 1786 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 48852 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 48852 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
timestamp 1586364061
transform 1 0 47104 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_498
timestamp 1586364061
transform 1 0 46920 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_502
timestamp 1586364061
transform 1 0 47288 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_26_514
timestamp 1586364061
transform 1 0 48392 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_27_508
timestamp 1586364061
transform 1 0 47840 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_398
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_399
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_105
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_117
timestamp 1586364061
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_129
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_141
timestamp 1586364061
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_400
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_166
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_178
timestamp 1586364061
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_190
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_401
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_202
timestamp 1586364061
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_239
timestamp 1586364061
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_263
timestamp 1586364061
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_402
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_288
timestamp 1586364061
transform 1 0 27600 0 -1 17952
box -38 -48 1142 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 29072 0 -1 17952
box -38 -48 406 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 30176 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 29624 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 29992 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_300
timestamp 1586364061
transform 1 0 28704 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_308
timestamp 1586364061
transform 1 0 29440 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_312
timestamp 1586364061
transform 1 0 29808 0 -1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 32200 0 -1 17952
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_403
timestamp 1586364061
transform 1 0 32016 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
timestamp 1586364061
transform 1 0 31832 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_325
timestamp 1586364061
transform 1 0 31004 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_28_333
timestamp 1586364061
transform 1 0 31740 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_337
timestamp 1586364061
transform 1 0 32108 0 -1 17952
box -38 -48 130 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 34868 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_8  FILLER_28_357
timestamp 1586364061
transform 1 0 33948 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_365
timestamp 1586364061
transform 1 0 34684 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_404
timestamp 1586364061
transform 1 0 37628 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 35880 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_376
timestamp 1586364061
transform 1 0 35696 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_380
timestamp 1586364061
transform 1 0 36064 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_28_392
timestamp 1586364061
transform 1 0 37168 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_396
timestamp 1586364061
transform 1 0 37536 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_398
timestamp 1586364061
transform 1 0 37720 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_410
timestamp 1586364061
transform 1 0 38824 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_28_422
timestamp 1586364061
transform 1 0 39928 0 -1 17952
box -38 -48 774 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 42044 0 -1 17952
box -38 -48 406 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 40940 0 -1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 41492 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_430
timestamp 1586364061
transform 1 0 40664 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_437
timestamp 1586364061
transform 1 0 41308 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_441
timestamp 1586364061
transform 1 0 41676 0 -1 17952
box -38 -48 406 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 43332 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_405
timestamp 1586364061
transform 1 0 43240 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 42872 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_449
timestamp 1586364061
transform 1 0 42412 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_453
timestamp 1586364061
transform 1 0 42780 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_456
timestamp 1586364061
transform 1 0 43056 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_468
timestamp 1586364061
transform 1 0 44160 0 -1 17952
box -38 -48 774 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1586364061
transform 1 0 45172 0 -1 17952
box -38 -48 866 592
use scs8hd_or2_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
timestamp 1586364061
transform 1 0 46736 0 -1 17952
box -38 -48 498 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
timestamp 1586364061
transform 1 0 46184 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
timestamp 1586364061
transform 1 0 46552 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1586364061
transform 1 0 44988 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_476
timestamp 1586364061
transform 1 0 44896 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_488
timestamp 1586364061
transform 1 0 46000 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_492
timestamp 1586364061
transform 1 0 46368 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 48852 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
timestamp 1586364061
transform 1 0 47380 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_501
timestamp 1586364061
transform 1 0 47196 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_505
timestamp 1586364061
transform 1 0 47564 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  FILLER_28_513
timestamp 1586364061
transform 1 0 48300 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_39
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_406
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_98
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_407
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_110
timestamp 1586364061
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_147
timestamp 1586364061
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_159
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_171
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_408
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_220
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_409
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_232
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_281
timestamp 1586364061
transform 1 0 26956 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_29_293
timestamp 1586364061
transform 1 0 28060 0 1 17952
box -38 -48 590 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 29624 0 1 17952
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_410
timestamp 1586364061
transform 1 0 29164 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 29440 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 28980 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 28612 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_301
timestamp 1586364061
transform 1 0 28796 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_306
timestamp 1586364061
transform 1 0 29256 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_329
timestamp 1586364061
transform 1 0 31372 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_341
timestamp 1586364061
transform 1 0 32476 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_411
timestamp 1586364061
transform 1 0 34776 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 35052 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 34592 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 34224 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_353
timestamp 1586364061
transform 1 0 33580 0 1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_29_359
timestamp 1586364061
transform 1 0 34132 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_362
timestamp 1586364061
transform 1 0 34408 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_367
timestamp 1586364061
transform 1 0 34868 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_371
timestamp 1586364061
transform 1 0 35236 0 1 17952
box -38 -48 314 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 35696 0 1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 35512 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_395
timestamp 1586364061
transform 1 0 37444 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 37720 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 38088 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 38456 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 39836 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_400
timestamp 1586364061
transform 1 0 37904 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_404
timestamp 1586364061
transform 1 0 38272 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_408
timestamp 1586364061
transform 1 0 38640 0 1 17952
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_29_420
timestamp 1586364061
transform 1 0 39744 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_428
timestamp 1586364061
transform 1 0 40480 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_423
timestamp 1586364061
transform 1 0 40020 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 40204 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_412
timestamp 1586364061
transform 1 0 40388 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_432
timestamp 1586364061
transform 1 0 40848 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 41032 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 40664 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_436
timestamp 1586364061
transform 1 0 41216 0 1 17952
box -38 -48 590 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 41768 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_446
timestamp 1586364061
transform 1 0 42136 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1586364061
transform 1 0 42872 0 1 17952
box -38 -48 866 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 44436 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 43884 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 42688 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 42320 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 44252 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_450
timestamp 1586364061
transform 1 0 42504 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_463
timestamp 1586364061
transform 1 0 43700 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_467
timestamp 1586364061
transform 1 0 44068 0 1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
timestamp 1586364061
transform 1 0 46092 0 1 17952
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_413
timestamp 1586364061
transform 1 0 46000 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 45816 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 45448 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 44988 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_475
timestamp 1586364061
transform 1 0 44804 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_479
timestamp 1586364061
transform 1 0 45172 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_484
timestamp 1586364061
transform 1 0 45632 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 48852 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_508
timestamp 1586364061
transform 1 0 47840 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_414
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_415
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_141
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_416
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_417
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_202
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_418
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_288
timestamp 1586364061
transform 1 0 27600 0 -1 19040
box -38 -48 1142 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 29532 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 29348 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_300
timestamp 1586364061
transform 1 0 28704 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_30_306
timestamp 1586364061
transform 1 0 29256 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_318
timestamp 1586364061
transform 1 0 30360 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_419
timestamp 1586364061
transform 1 0 32016 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 32292 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_330
timestamp 1586364061
transform 1 0 31464 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_2  FILLER_30_337
timestamp 1586364061
transform 1 0 32108 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_341
timestamp 1586364061
transform 1 0 32476 0 -1 19040
box -38 -48 1142 592
use scs8hd_conb_1  _58_
timestamp 1586364061
transform 1 0 34040 0 -1 19040
box -38 -48 314 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 35052 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 34868 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 34500 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_353
timestamp 1586364061
transform 1 0 33580 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_357
timestamp 1586364061
transform 1 0 33948 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_361
timestamp 1586364061
transform 1 0 34316 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_365
timestamp 1586364061
transform 1 0 34684 0 -1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_420
timestamp 1586364061
transform 1 0 37628 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 37444 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_378
timestamp 1586364061
transform 1 0 35880 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_30_390
timestamp 1586364061
transform 1 0 36984 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_394
timestamp 1586364061
transform 1 0 37352 0 -1 19040
box -38 -48 130 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 37720 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 38732 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_407
timestamp 1586364061
transform 1 0 38548 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_411
timestamp 1586364061
transform 1 0 38916 0 -1 19040
box -38 -48 1142 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 40296 0 -1 19040
box -38 -48 2246 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 40112 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_423
timestamp 1586364061
transform 1 0 40020 0 -1 19040
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 43608 0 -1 19040
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_421
timestamp 1586364061
transform 1 0 43240 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 42872 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_450
timestamp 1586364061
transform 1 0 42504 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_30_456
timestamp 1586364061
transform 1 0 43056 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_459
timestamp 1586364061
transform 1 0 43332 0 -1 19040
box -38 -48 314 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 46092 0 -1 19040
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_30_481
timestamp 1586364061
transform 1 0 45356 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 48852 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_508
timestamp 1586364061
transform 1 0 47840 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_422
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_86
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_423
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_110
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_147
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_159
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_171
timestamp 1586364061
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_424
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_425
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_281
timestamp 1586364061
transform 1 0 26956 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_293
timestamp 1586364061
transform 1 0 28060 0 1 19040
box -38 -48 774 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 29716 0 1 19040
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_426
timestamp 1586364061
transform 1 0 29164 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 29532 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 28980 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_301
timestamp 1586364061
transform 1 0 28796 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_306
timestamp 1586364061
transform 1 0 29256 0 1 19040
box -38 -48 314 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 32200 0 1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 32016 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 31648 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_330
timestamp 1586364061
transform 1 0 31464 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_334
timestamp 1586364061
transform 1 0 31832 0 1 19040
box -38 -48 222 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 35052 0 1 19040
box -38 -48 2246 592
use scs8hd_tapvpwrvgnd_1  PHY_427
timestamp 1586364061
transform 1 0 34776 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 34592 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 34224 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_357
timestamp 1586364061
transform 1 0 33948 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_362
timestamp 1586364061
transform 1 0 34408 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_367
timestamp 1586364061
transform 1 0 34868 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_393
timestamp 1586364061
transform 1 0 37260 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_397
timestamp 1586364061
transform 1 0 37628 0 1 19040
box -38 -48 130 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 37996 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 37720 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 39008 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 39836 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 39376 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_400
timestamp 1586364061
transform 1 0 37904 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_410
timestamp 1586364061
transform 1 0 38824 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_414
timestamp 1586364061
transform 1 0 39192 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_418
timestamp 1586364061
transform 1 0 39560 0 1 19040
box -38 -48 314 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 40480 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_428
timestamp 1586364061
transform 1 0 40388 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 40204 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 41492 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 41860 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_423
timestamp 1586364061
transform 1 0 40020 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_437
timestamp 1586364061
transform 1 0 41308 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_441
timestamp 1586364061
transform 1 0 41676 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_445
timestamp 1586364061
transform 1 0 42044 0 1 19040
box -38 -48 774 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 43516 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 43332 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 42964 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_453
timestamp 1586364061
transform 1 0 42780 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_457
timestamp 1586364061
transform 1 0 43148 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_470
timestamp 1586364061
transform 1 0 44344 0 1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_429
timestamp 1586364061
transform 1 0 46000 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 44712 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 45080 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_476
timestamp 1586364061
transform 1 0 44896 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_480
timestamp 1586364061
transform 1 0 45264 0 1 19040
box -38 -48 774 592
use scs8hd_decap_12  FILLER_31_489
timestamp 1586364061
transform 1 0 46092 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 48852 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 47196 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_503
timestamp 1586364061
transform 1 0 47380 0 1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_31_515
timestamp 1586364061
transform 1 0 48484 0 1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_430
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_431
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_117
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_129
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_141
timestamp 1586364061
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_432
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_433
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_434
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_288
timestamp 1586364061
transform 1 0 27600 0 -1 20128
box -38 -48 1142 592
use scs8hd_conb_1  _51_
timestamp 1586364061
transform 1 0 29808 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 30360 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 30728 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 29624 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_300
timestamp 1586364061
transform 1 0 28704 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_32_308
timestamp 1586364061
transform 1 0 29440 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_315
timestamp 1586364061
transform 1 0 30084 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_320
timestamp 1586364061
transform 1 0 30544 0 -1 20128
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 32108 0 -1 20128
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_435
timestamp 1586364061
transform 1 0 32016 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 31096 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 32660 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_324
timestamp 1586364061
transform 1 0 30912 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_328
timestamp 1586364061
transform 1 0 31280 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_32_341
timestamp 1586364061
transform 1 0 32476 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_345
timestamp 1586364061
transform 1 0 32844 0 -1 20128
box -38 -48 314 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 34684 0 -1 20128
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 33120 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 33488 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 34500 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_350
timestamp 1586364061
transform 1 0 33304 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_354
timestamp 1586364061
transform 1 0 33672 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_32_362
timestamp 1586364061
transform 1 0 34408 0 -1 20128
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_436
timestamp 1586364061
transform 1 0 37628 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_384
timestamp 1586364061
transform 1 0 36432 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_32_396
timestamp 1586364061
transform 1 0 37536 0 -1 20128
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 37720 0 -1 20128
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_32_417
timestamp 1586364061
transform 1 0 39468 0 -1 20128
box -38 -48 774 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 40204 0 -1 20128
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 42228 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_444
timestamp 1586364061
transform 1 0 41952 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_449
timestamp 1586364061
transform 1 0 42412 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 42596 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_453
timestamp 1586364061
transform 1 0 42780 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_459
timestamp 1586364061
transform 1 0 43332 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_457
timestamp 1586364061
transform 1 0 43148 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 43516 0 -1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_437
timestamp 1586364061
transform 1 0 43240 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_466
timestamp 1586364061
transform 1 0 43976 0 -1 20128
box -38 -48 406 592
use scs8hd_conb_1  _59_
timestamp 1586364061
transform 1 0 43700 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_32_470
timestamp 1586364061
transform 1 0 44344 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 44436 0 -1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 44712 0 -1 20128
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_32_473
timestamp 1586364061
transform 1 0 44620 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_493
timestamp 1586364061
transform 1 0 46460 0 -1 20128
box -38 -48 774 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 47196 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 48852 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_505
timestamp 1586364061
transform 1 0 47564 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_3  FILLER_32_513
timestamp 1586364061
transform 1 0 48300 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_446
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_438
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_447
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_439
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_147
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_448
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_159
timestamp 1586364061
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_171
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_440
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_449
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_441
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_34_284
timestamp 1586364061
transform 1 0 27232 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_284
timestamp 1586364061
transform 1 0 27232 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_281
timestamp 1586364061
transform 1 0 26956 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 27048 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_450
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_296
timestamp 1586364061
transform 1 0 28336 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_292
timestamp 1586364061
transform 1 0 27968 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_288
timestamp 1586364061
transform 1 0 27600 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 28152 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 27784 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 27416 0 1 20128
box -38 -48 222 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 27416 0 -1 21216
box -38 -48 2246 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 29624 0 1 20128
box -38 -48 1786 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 30360 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_442
timestamp 1586364061
transform 1 0 29164 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 29440 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 29808 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_304
timestamp 1586364061
transform 1 0 29072 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_306
timestamp 1586364061
transform 1 0 29256 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_310
timestamp 1586364061
transform 1 0 29624 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_314
timestamp 1586364061
transform 1 0 29992 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_335
timestamp 1586364061
transform 1 0 31924 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_34_327
timestamp 1586364061
transform 1 0 31188 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_334
timestamp 1586364061
transform 1 0 31832 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_329
timestamp 1586364061
transform 1 0 31372 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 31648 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_337
timestamp 1586364061
transform 1 0 32108 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_4  FILLER_33_342
timestamp 1586364061
transform 1 0 32568 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_338
timestamp 1586364061
transform 1 0 32200 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 32016 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 32936 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 32384 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_451
timestamp 1586364061
transform 1 0 32016 0 -1 21216
box -38 -48 130 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 32384 0 -1 21216
box -38 -48 2246 592
use scs8hd_decap_8  FILLER_33_357
timestamp 1586364061
transform 1 0 33948 0 1 20128
box -38 -48 774 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 33120 0 1 20128
box -38 -48 866 592
use scs8hd_fill_1  FILLER_34_370
timestamp 1586364061
transform 1 0 35144 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_34_364
timestamp 1586364061
transform 1 0 34592 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_2  FILLER_33_367
timestamp 1586364061
transform 1 0 34868 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_365
timestamp 1586364061
transform 1 0 34684 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 35236 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 35052 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_443
timestamp 1586364061
transform 1 0 34776 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_371
timestamp 1586364061
transform 1 0 35236 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_379
timestamp 1586364061
transform 1 0 35972 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_34_373
timestamp 1586364061
transform 1 0 35420 0 -1 21216
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 36064 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_386
timestamp 1586364061
transform 1 0 36616 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_34_382
timestamp 1586364061
transform 1 0 36248 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_383
timestamp 1586364061
transform 1 0 36340 0 1 20128
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 36432 0 -1 21216
box -38 -48 222 592
use scs8hd_conb_1  _56_
timestamp 1586364061
transform 1 0 36892 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  FILLER_34_394
timestamp 1586364061
transform 1 0 37352 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_6  FILLER_33_392
timestamp 1586364061
transform 1 0 37168 0 1 20128
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_452
timestamp 1586364061
transform 1 0 37628 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_402
timestamp 1586364061
transform 1 0 38088 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_398
timestamp 1586364061
transform 1 0 37720 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 38272 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 37904 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 37720 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_418
timestamp 1586364061
transform 1 0 39560 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_419
timestamp 1586364061
transform 1 0 39652 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 39836 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_406
timestamp 1586364061
transform 1 0 38456 0 -1 21216
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 37904 0 1 20128
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_34_433
timestamp 1586364061
transform 1 0 40940 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_429
timestamp 1586364061
transform 1 0 40572 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_423
timestamp 1586364061
transform 1 0 40020 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 40204 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 40756 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_444
timestamp 1586364061
transform 1 0 40388 0 1 20128
box -38 -48 130 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 40480 0 1 20128
box -38 -48 866 592
use scs8hd_conb_1  _57_
timestamp 1586364061
transform 1 0 40296 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_6  FILLER_34_441
timestamp 1586364061
transform 1 0 41676 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_2  FILLER_34_437
timestamp 1586364061
transform 1 0 41308 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_441
timestamp 1586364061
transform 1 0 41676 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_437
timestamp 1586364061
transform 1 0 41308 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 41492 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 42228 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 41492 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 41124 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 42044 0 1 20128
box -38 -48 222 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 42228 0 1 20128
box -38 -48 2246 592
use scs8hd_fill_1  FILLER_34_455
timestamp 1586364061
transform 1 0 42964 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_34_449
timestamp 1586364061
transform 1 0 42412 0 -1 21216
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 43056 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_463
timestamp 1586364061
transform 1 0 43700 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_459
timestamp 1586364061
transform 1 0 43332 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 43884 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_453
timestamp 1586364061
transform 1 0 43240 0 -1 21216
box -38 -48 130 592
use scs8hd_conb_1  _62_
timestamp 1586364061
transform 1 0 43424 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_467
timestamp 1586364061
transform 1 0 44068 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_471
timestamp 1586364061
transform 1 0 44436 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 44252 0 -1 21216
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 44436 0 -1 21216
box -38 -48 866 592
use scs8hd_decap_8  FILLER_34_480
timestamp 1586364061
transform 1 0 45264 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_8  FILLER_33_479
timestamp 1586364061
transform 1 0 45172 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_475
timestamp 1586364061
transform 1 0 44804 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 44988 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 44620 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_488
timestamp 1586364061
transform 1 0 46000 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_33_489
timestamp 1586364061
transform 1 0 46092 0 1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_33_487
timestamp 1586364061
transform 1 0 45908 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 46092 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_445
timestamp 1586364061
transform 1 0 46000 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_495
timestamp 1586364061
transform 1 0 46644 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_491
timestamp 1586364061
transform 1 0 46276 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_495
timestamp 1586364061
transform 1 0 46644 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 46460 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 46736 0 1 20128
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 46736 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 48852 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 48852 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_498
timestamp 1586364061
transform 1 0 46920 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_33_510
timestamp 1586364061
transform 1 0 48024 0 1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_34_500
timestamp 1586364061
transform 1 0 47104 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_512
timestamp 1586364061
transform 1 0 48208 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_454
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_455
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_147
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_159
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_171
timestamp 1586364061
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_456
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_457
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 1142 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 27600 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 27416 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 27048 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_281
timestamp 1586364061
transform 1 0 26956 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_284
timestamp 1586364061
transform 1 0 27232 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_297
timestamp 1586364061
transform 1 0 28428 0 1 21216
box -38 -48 406 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 29256 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_458
timestamp 1586364061
transform 1 0 29164 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 28888 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 30268 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_301
timestamp 1586364061
transform 1 0 28796 0 1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_35_304
timestamp 1586364061
transform 1 0 29072 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_315
timestamp 1586364061
transform 1 0 30084 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_319
timestamp 1586364061
transform 1 0 30452 0 1 21216
box -38 -48 406 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 31096 0 1 21216
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 30912 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_323
timestamp 1586364061
transform 1 0 30820 0 1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_35_345
timestamp 1586364061
transform 1 0 32844 0 1 21216
box -38 -48 774 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 35236 0 1 21216
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_459
timestamp 1586364061
transform 1 0 34776 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 35052 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 33580 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 33948 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_355
timestamp 1586364061
transform 1 0 33764 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_359
timestamp 1586364061
transform 1 0 34132 0 1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_35_365
timestamp 1586364061
transform 1 0 34684 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_367
timestamp 1586364061
transform 1 0 34868 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 37536 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 37168 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_390
timestamp 1586364061
transform 1 0 36984 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_394
timestamp 1586364061
transform 1 0 37352 0 1 21216
box -38 -48 222 592
use scs8hd_conb_1  _34_
timestamp 1586364061
transform 1 0 37720 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 38180 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 38548 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 39836 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_401
timestamp 1586364061
transform 1 0 37996 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_405
timestamp 1586364061
transform 1 0 38364 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_409
timestamp 1586364061
transform 1 0 38732 0 1 21216
box -38 -48 1142 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 40756 0 1 21216
box -38 -48 2246 592
use scs8hd_tapvpwrvgnd_1  PHY_460
timestamp 1586364061
transform 1 0 40388 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 40204 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_423
timestamp 1586364061
transform 1 0 40020 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_428
timestamp 1586364061
transform 1 0 40480 0 1 21216
box -38 -48 314 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 43700 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 43332 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_455
timestamp 1586364061
transform 1 0 42964 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_461
timestamp 1586364061
transform 1 0 43516 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_484
timestamp 1586364061
transform 1 0 45632 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_480
timestamp 1586364061
transform 1 0 45264 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_476
timestamp 1586364061
transform 1 0 44896 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_472
timestamp 1586364061
transform 1 0 44528 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 45080 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 45448 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 44712 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 45816 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_461
timestamp 1586364061
transform 1 0 46000 0 1 21216
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 46092 0 1 21216
box -38 -48 1786 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 48852 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_508
timestamp 1586364061
transform 1 0 47840 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_462
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_463
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_117
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_129
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_141
timestamp 1586364061
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_464
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_166
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_178
timestamp 1586364061
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_190
timestamp 1586364061
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_465
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_202
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_conb_1  _54_
timestamp 1586364061
transform 1 0 27876 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_466
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 27600 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_36_290
timestamp 1586364061
transform 1 0 27784 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_36_294
timestamp 1586364061
transform 1 0 28152 0 -1 22304
box -38 -48 590 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 28888 0 -1 22304
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 28704 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_321
timestamp 1586364061
transform 1 0 30636 0 -1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_467
timestamp 1586364061
transform 1 0 32016 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 32292 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 31096 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_325
timestamp 1586364061
transform 1 0 31004 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_328
timestamp 1586364061
transform 1 0 31280 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_36_337
timestamp 1586364061
transform 1 0 32108 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_341
timestamp 1586364061
transform 1 0 32476 0 -1 22304
box -38 -48 774 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 33580 0 -1 22304
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 33396 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_349
timestamp 1586364061
transform 1 0 33212 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_372
timestamp 1586364061
transform 1 0 35328 0 -1 22304
box -38 -48 774 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 36064 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_468
timestamp 1586364061
transform 1 0 37628 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_389
timestamp 1586364061
transform 1 0 36892 0 -1 22304
box -38 -48 774 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 37904 0 -1 22304
box -38 -48 2246 592
use scs8hd_fill_2  FILLER_36_398
timestamp 1586364061
transform 1 0 37720 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 40940 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 40756 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 40388 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_424
timestamp 1586364061
transform 1 0 40112 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_36_429
timestamp 1586364061
transform 1 0 40572 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_36_442
timestamp 1586364061
transform 1 0 41768 0 -1 22304
box -38 -48 1142 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 43332 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_469
timestamp 1586364061
transform 1 0 43240 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_454
timestamp 1586364061
transform 1 0 42872 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_4  FILLER_36_468
timestamp 1586364061
transform 1 0 44160 0 -1 22304
box -38 -48 406 592
use scs8hd_conb_1  _60_
timestamp 1586364061
transform 1 0 45080 0 -1 22304
box -38 -48 314 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 46092 0 -1 22304
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 44620 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_472
timestamp 1586364061
transform 1 0 44528 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_36_475
timestamp 1586364061
transform 1 0 44804 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_481
timestamp 1586364061
transform 1 0 45356 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 48852 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_508
timestamp 1586364061
transform 1 0 47840 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_470
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_471
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_110
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_147
timestamp 1586364061
transform 1 0 14628 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_159
timestamp 1586364061
transform 1 0 15732 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_171
timestamp 1586364061
transform 1 0 16836 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_472
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_196
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_208
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_220
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_473
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_232
timestamp 1586364061
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_281
timestamp 1586364061
transform 1 0 26956 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_293
timestamp 1586364061
transform 1 0 28060 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_474
timestamp 1586364061
transform 1 0 29164 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 29440 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_306
timestamp 1586364061
transform 1 0 29256 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_310
timestamp 1586364061
transform 1 0 29624 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_322
timestamp 1586364061
transform 1 0 30728 0 1 22304
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 32292 0 1 22304
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 32108 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_334
timestamp 1586364061
transform 1 0 31832 0 1 22304
box -38 -48 314 592
use scs8hd_conb_1  _53_
timestamp 1586364061
transform 1 0 34868 0 1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_475
timestamp 1586364061
transform 1 0 34776 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 34224 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 34592 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_358
timestamp 1586364061
transform 1 0 34040 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_362
timestamp 1586364061
transform 1 0 34408 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_370
timestamp 1586364061
transform 1 0 35144 0 1 22304
box -38 -48 314 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 35972 0 1 22304
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 35788 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 35420 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_375
timestamp 1586364061
transform 1 0 35604 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 38456 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCE
timestamp 1586364061
transform 1 0 39468 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 38272 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__D
timestamp 1586364061
transform 1 0 37904 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__SCD
timestamp 1586364061
transform 1 0 39836 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_398
timestamp 1586364061
transform 1 0 37720 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_402
timestamp 1586364061
transform 1 0 38088 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_415
timestamp 1586364061
transform 1 0 39284 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_419
timestamp 1586364061
transform 1 0 39652 0 1 22304
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 40940 0 1 22304
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_476
timestamp 1586364061
transform 1 0 40388 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 40756 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 40204 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_423
timestamp 1586364061
transform 1 0 40020 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_428
timestamp 1586364061
transform 1 0 40480 0 1 22304
box -38 -48 314 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 43516 0 1 22304
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 43332 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_452
timestamp 1586364061
transform 1 0 42688 0 1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_37_458
timestamp 1586364061
transform 1 0 43240 0 1 22304
box -38 -48 130 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 46184 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_477
timestamp 1586364061
transform 1 0 46000 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 45448 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 45816 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_480
timestamp 1586364061
transform 1 0 45264 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_484
timestamp 1586364061
transform 1 0 45632 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_489
timestamp 1586364061
transform 1 0 46092 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 48852 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 47196 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_499
timestamp 1586364061
transform 1 0 47012 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_503
timestamp 1586364061
transform 1 0 47380 0 1 22304
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_37_515
timestamp 1586364061
transform 1 0 48484 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_478
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_479
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_141
timestamp 1586364061
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_480
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_166
timestamp 1586364061
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_178
timestamp 1586364061
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_190
timestamp 1586364061
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_481
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_202
timestamp 1586364061
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_263
timestamp 1586364061
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_482
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_288
timestamp 1586364061
transform 1 0 27600 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_300
timestamp 1586364061
transform 1 0 28704 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_312
timestamp 1586364061
transform 1 0 29808 0 -1 23392
box -38 -48 1142 592
use scs8hd_conb_1  _52_
timestamp 1586364061
transform 1 0 32108 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_483
timestamp 1586364061
transform 1 0 32016 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 31188 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_38_324
timestamp 1586364061
transform 1 0 30912 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_6  FILLER_38_329
timestamp 1586364061
transform 1 0 31372 0 -1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_38_335
timestamp 1586364061
transform 1 0 31924 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_340
timestamp 1586364061
transform 1 0 32384 0 -1 23392
box -38 -48 1142 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 33488 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_12  FILLER_38_361
timestamp 1586364061
transform 1 0 34316 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_484
timestamp 1586364061
transform 1 0 37628 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 36064 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 36432 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_373
timestamp 1586364061
transform 1 0 35420 0 -1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_38_379
timestamp 1586364061
transform 1 0 35972 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_382
timestamp 1586364061
transform 1 0 36248 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_386
timestamp 1586364061
transform 1 0 36616 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_3  FILLER_38_394
timestamp 1586364061
transform 1 0 37352 0 -1 23392
box -38 -48 314 592
use scs8hd_sdfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0_
timestamp 1586364061
transform 1 0 38640 0 -1 23392
box -38 -48 2246 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 38456 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_398
timestamp 1586364061
transform 1 0 37720 0 -1 23392
box -38 -48 774 592
use scs8hd_conb_1  _61_
timestamp 1586364061
transform 1 0 41584 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 41032 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_432
timestamp 1586364061
transform 1 0 40848 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_436
timestamp 1586364061
transform 1 0 41216 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_6  FILLER_38_443
timestamp 1586364061
transform 1 0 41860 0 -1 23392
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_485
timestamp 1586364061
transform 1 0 43240 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 42504 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 43516 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_449
timestamp 1586364061
transform 1 0 42412 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_6  FILLER_38_452
timestamp 1586364061
transform 1 0 42688 0 -1 23392
box -38 -48 590 592
use scs8hd_fill_2  FILLER_38_459
timestamp 1586364061
transform 1 0 43332 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_463
timestamp 1586364061
transform 1 0 43700 0 -1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_38_471
timestamp 1586364061
transform 1 0 44436 0 -1 23392
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 44620 0 -1 23392
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 46552 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_492
timestamp 1586364061
transform 1 0 46368 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_496
timestamp 1586364061
transform 1 0 46736 0 -1 23392
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 47104 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 48852 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 46920 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_504
timestamp 1586364061
transform 1 0 47472 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_15
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_494
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_27
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_39
timestamp 1586364061
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_486
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_51
timestamp 1586364061
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_495
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_487
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_110
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_135
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_147
timestamp 1586364061
transform 1 0 14628 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_496
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_159
timestamp 1586364061
transform 1 0 15732 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_171
timestamp 1586364061
transform 1 0 16836 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_488
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_196
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_497
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_208
timestamp 1586364061
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_220
timestamp 1586364061
transform 1 0 21344 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_489
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_232
timestamp 1586364061
transform 1 0 22448 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_257
timestamp 1586364061
transform 1 0 24748 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_269
timestamp 1586364061
transform 1 0 25852 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_263
timestamp 1586364061
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_498
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_281
timestamp 1586364061
transform 1 0 26956 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_293
timestamp 1586364061
transform 1 0 28060 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_288
timestamp 1586364061
transform 1 0 27600 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_490
timestamp 1586364061
transform 1 0 29164 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_306
timestamp 1586364061
transform 1 0 29256 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_39_318
timestamp 1586364061
transform 1 0 30360 0 1 23392
box -38 -48 590 592
use scs8hd_decap_12  FILLER_40_300
timestamp 1586364061
transform 1 0 28704 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_312
timestamp 1586364061
transform 1 0 29808 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_335
timestamp 1586364061
transform 1 0 31924 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_6  FILLER_40_329
timestamp 1586364061
transform 1 0 31372 0 -1 24480
box -38 -48 590 592
use scs8hd_decap_3  FILLER_40_324
timestamp 1586364061
transform 1 0 30912 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_1  FILLER_39_324
timestamp 1586364061
transform 1 0 30912 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 31188 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 31004 0 1 23392
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 31188 0 1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_499
timestamp 1586364061
transform 1 0 32016 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_337
timestamp 1586364061
transform 1 0 32108 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_336
timestamp 1586364061
transform 1 0 32016 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_39_360
timestamp 1586364061
transform 1 0 34224 0 1 23392
box -38 -48 590 592
use scs8hd_fill_2  FILLER_40_372
timestamp 1586364061
transform 1 0 35328 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_361
timestamp 1586364061
transform 1 0 34316 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_372
timestamp 1586364061
transform 1 0 35328 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_367
timestamp 1586364061
transform 1 0 34868 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 35144 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_491
timestamp 1586364061
transform 1 0 34776 0 1 23392
box -38 -48 130 592
use scs8hd_conb_1  _33_
timestamp 1586364061
transform 1 0 35052 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_349
timestamp 1586364061
transform 1 0 33212 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_348
timestamp 1586364061
transform 1 0 33120 0 1 23392
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_40_376
timestamp 1586364061
transform 1 0 35696 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_376
timestamp 1586364061
transform 1 0 35696 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 35512 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 35512 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 35880 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 35880 0 1 23392
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 36064 0 -1 24480
box -38 -48 866 592
use scs8hd_decap_8  FILLER_40_389
timestamp 1586364061
transform 1 0 36892 0 -1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_500
timestamp 1586364061
transform 1 0 37628 0 -1 24480
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 36064 0 1 23392
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 37904 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.scs8hd_sdfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 38640 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_399
timestamp 1586364061
transform 1 0 37812 0 1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_39_407
timestamp 1586364061
transform 1 0 38548 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_410
timestamp 1586364061
transform 1 0 38824 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_39_422
timestamp 1586364061
transform 1 0 39928 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_40_398
timestamp 1586364061
transform 1 0 37720 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_402
timestamp 1586364061
transform 1 0 38088 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_414
timestamp 1586364061
transform 1 0 39192 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_432
timestamp 1586364061
transform 1 0 40848 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_6  FILLER_40_426
timestamp 1586364061
transform 1 0 40296 0 -1 24480
box -38 -48 590 592
use scs8hd_decap_3  FILLER_39_428
timestamp 1586364061
transform 1 0 40480 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 40204 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 40756 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_492
timestamp 1586364061
transform 1 0 40388 0 1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_40_439
timestamp 1586364061
transform 1 0 41492 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_40_435
timestamp 1586364061
transform 1 0 41124 0 -1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 40940 0 -1 24480
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2_
timestamp 1586364061
transform 1 0 41584 0 -1 24480
box -38 -48 406 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 40940 0 1 23392
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_444
timestamp 1586364061
transform 1 0 41952 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_446
timestamp 1586364061
transform 1 0 42136 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_442
timestamp 1586364061
transform 1 0 41768 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_2__A
timestamp 1586364061
transform 1 0 41952 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 42136 0 -1 24480
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 42504 0 1 23392
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_501
timestamp 1586364061
transform 1 0 43240 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 42320 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 42504 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_469
timestamp 1586364061
transform 1 0 44252 0 1 23392
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_40_448
timestamp 1586364061
transform 1 0 42320 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_40_452
timestamp 1586364061
transform 1 0 42688 0 -1 24480
box -38 -48 590 592
use scs8hd_decap_12  FILLER_40_459
timestamp 1586364061
transform 1 0 43332 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_471
timestamp 1586364061
transform 1 0 44436 0 -1 24480
box -38 -48 774 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 45448 0 -1 24480
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_493
timestamp 1586364061
transform 1 0 46000 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 45448 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 45816 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 45172 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_481
timestamp 1586364061
transform 1 0 45356 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_484
timestamp 1586364061
transform 1 0 45632 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_489
timestamp 1586364061
transform 1 0 46092 0 1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_481
timestamp 1586364061
transform 1 0 45356 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 48852 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 48852 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_501
timestamp 1586364061
transform 1 0 47196 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_39_513
timestamp 1586364061
transform 1 0 48300 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_501
timestamp 1586364061
transform 1 0 47196 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_40_513
timestamp 1586364061
transform 1 0 48300 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_502
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_503
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_504
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_505
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_281
timestamp 1586364061
transform 1 0 26956 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_293
timestamp 1586364061
transform 1 0 28060 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_506
timestamp 1586364061
transform 1 0 29164 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_306
timestamp 1586364061
transform 1 0 29256 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_318
timestamp 1586364061
transform 1 0 30360 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_330
timestamp 1586364061
transform 1 0 31464 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_342
timestamp 1586364061
transform 1 0 32568 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_507
timestamp 1586364061
transform 1 0 34776 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 35328 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_354
timestamp 1586364061
transform 1 0 33672 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_41_367
timestamp 1586364061
transform 1 0 34868 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_371
timestamp 1586364061
transform 1 0 35236 0 1 24480
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 35512 0 1 24480
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_41_393
timestamp 1586364061
transform 1 0 37260 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_397
timestamp 1586364061
transform 1 0 37628 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_404
timestamp 1586364061
transform 1 0 38272 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_400
timestamp 1586364061
transform 1 0 37904 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 38088 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 37720 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1__A
timestamp 1586364061
transform 1 0 38456 0 1 24480
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_1_
timestamp 1586364061
transform 1 0 38640 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_417
timestamp 1586364061
transform 1 0 39468 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_412
timestamp 1586364061
transform 1 0 39008 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 39284 0 1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_41_421
timestamp 1586364061
transform 1 0 39836 0 1 24480
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 39652 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1586364061
transform 1 0 42136 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_508
timestamp 1586364061
transform 1 0 40388 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 41952 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 41584 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_428
timestamp 1586364061
transform 1 0 40480 0 1 24480
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_41_442
timestamp 1586364061
transform 1 0 41768 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__B
timestamp 1586364061
transform 1 0 43332 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0__A
timestamp 1586364061
transform 1 0 43700 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_455
timestamp 1586364061
transform 1 0 42964 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_461
timestamp 1586364061
transform 1 0 43516 0 1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_41_465
timestamp 1586364061
transform 1 0 43884 0 1 24480
box -38 -48 774 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 46092 0 1 24480
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_509
timestamp 1586364061
transform 1 0 46000 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 45816 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 45172 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 44804 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_473
timestamp 1586364061
transform 1 0 44620 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_477
timestamp 1586364061
transform 1 0 44988 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_481
timestamp 1586364061
transform 1 0 45356 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_485
timestamp 1586364061
transform 1 0 45724 0 1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 48852 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_508
timestamp 1586364061
transform 1 0 47840 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_510
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_68
timestamp 1586364061
transform 1 0 7360 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_511
timestamp 1586364061
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_80
timestamp 1586364061
transform 1 0 8464 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_93
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_105
timestamp 1586364061
transform 1 0 10764 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_117
timestamp 1586364061
transform 1 0 11868 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_129
timestamp 1586364061
transform 1 0 12972 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_141
timestamp 1586364061
transform 1 0 14076 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_512
timestamp 1586364061
transform 1 0 15180 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_154
timestamp 1586364061
transform 1 0 15272 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_166
timestamp 1586364061
transform 1 0 16376 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_178
timestamp 1586364061
transform 1 0 17480 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_190
timestamp 1586364061
transform 1 0 18584 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_513
timestamp 1586364061
transform 1 0 20792 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_202
timestamp 1586364061
transform 1 0 19688 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_215
timestamp 1586364061
transform 1 0 20884 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_227
timestamp 1586364061
transform 1 0 21988 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_239
timestamp 1586364061
transform 1 0 23092 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_251
timestamp 1586364061
transform 1 0 24196 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_263
timestamp 1586364061
transform 1 0 25300 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_514
timestamp 1586364061
transform 1 0 26404 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_276
timestamp 1586364061
transform 1 0 26496 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_288
timestamp 1586364061
transform 1 0 27600 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_300
timestamp 1586364061
transform 1 0 28704 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_312
timestamp 1586364061
transform 1 0 29808 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_515
timestamp 1586364061
transform 1 0 32016 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_324
timestamp 1586364061
transform 1 0 30912 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_337
timestamp 1586364061
transform 1 0 32108 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_349
timestamp 1586364061
transform 1 0 33212 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_361
timestamp 1586364061
transform 1 0 34316 0 -1 25568
box -38 -48 1142 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 35880 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_516
timestamp 1586364061
transform 1 0 37628 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 35696 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_42_373
timestamp 1586364061
transform 1 0 35420 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_8  FILLER_42_387
timestamp 1586364061
transform 1 0 36708 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_2  FILLER_42_395
timestamp 1586364061
transform 1 0 37444 0 -1 25568
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 39284 0 -1 25568
box -38 -48 1786 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 37720 0 -1 25568
box -38 -48 866 592
use scs8hd_decap_8  FILLER_42_407
timestamp 1586364061
transform 1 0 38548 0 -1 25568
box -38 -48 774 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 42136 0 -1 25568
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 41308 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 41676 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_42_434
timestamp 1586364061
transform 1 0 41032 0 -1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_42_439
timestamp 1586364061
transform 1 0 41492 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_42_443
timestamp 1586364061
transform 1 0 41860 0 -1 25568
box -38 -48 314 592
use scs8hd_or2_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.scs8hd_or2_1_0_
timestamp 1586364061
transform 1 0 43332 0 -1 25568
box -38 -48 498 592
use scs8hd_tapvpwrvgnd_1  PHY_517
timestamp 1586364061
transform 1 0 43240 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_450
timestamp 1586364061
transform 1 0 42504 0 -1 25568
box -38 -48 774 592
use scs8hd_decap_8  FILLER_42_464
timestamp 1586364061
transform 1 0 43792 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_1  FILLER_42_478
timestamp 1586364061
transform 1 0 45080 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_42_474
timestamp 1586364061
transform 1 0 44712 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3__A
timestamp 1586364061
transform 1 0 44896 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 44528 0 -1 25568
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1586364061
transform 1 0 45172 0 -1 25568
box -38 -48 866 592
use scs8hd_fill_2  FILLER_42_488
timestamp 1586364061
transform 1 0 46000 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 46184 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_492
timestamp 1586364061
transform 1 0 46368 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 46552 0 -1 25568
box -38 -48 222 592
use scs8hd_buf_2  _73_
timestamp 1586364061
transform 1 0 46736 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 48852 0 -1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__73__A
timestamp 1586364061
transform 1 0 47288 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_500
timestamp 1586364061
transform 1 0 47104 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_42_504
timestamp 1586364061
transform 1 0 47472 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_86
timestamp 1586364061
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_43_3
timestamp 1586364061
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_15
timestamp 1586364061
transform 1 0 2484 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_27
timestamp 1586364061
transform 1 0 3588 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_39
timestamp 1586364061
transform 1 0 4692 0 1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_518
timestamp 1586364061
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_43_51
timestamp 1586364061
transform 1 0 5796 0 1 25568
box -38 -48 774 592
use scs8hd_fill_2  FILLER_43_59
timestamp 1586364061
transform 1 0 6532 0 1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_43_62
timestamp 1586364061
transform 1 0 6808 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_74
timestamp 1586364061
transform 1 0 7912 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_86
timestamp 1586364061
transform 1 0 9016 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_98
timestamp 1586364061
transform 1 0 10120 0 1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_519
timestamp 1586364061
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_43_110
timestamp 1586364061
transform 1 0 11224 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_123
timestamp 1586364061
transform 1 0 12420 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_135
timestamp 1586364061
transform 1 0 13524 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_147
timestamp 1586364061
transform 1 0 14628 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_159
timestamp 1586364061
transform 1 0 15732 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_171
timestamp 1586364061
transform 1 0 16836 0 1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_520
timestamp 1586364061
transform 1 0 17940 0 1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_43_184
timestamp 1586364061
transform 1 0 18032 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_196
timestamp 1586364061
transform 1 0 19136 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_208
timestamp 1586364061
transform 1 0 20240 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_220
timestamp 1586364061
transform 1 0 21344 0 1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_521
timestamp 1586364061
transform 1 0 23552 0 1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_43_232
timestamp 1586364061
transform 1 0 22448 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_245
timestamp 1586364061
transform 1 0 23644 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_257
timestamp 1586364061
transform 1 0 24748 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_269
timestamp 1586364061
transform 1 0 25852 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_281
timestamp 1586364061
transform 1 0 26956 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_293
timestamp 1586364061
transform 1 0 28060 0 1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_522
timestamp 1586364061
transform 1 0 29164 0 1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_43_306
timestamp 1586364061
transform 1 0 29256 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_318
timestamp 1586364061
transform 1 0 30360 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_330
timestamp 1586364061
transform 1 0 31464 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_342
timestamp 1586364061
transform 1 0 32568 0 1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_523
timestamp 1586364061
transform 1 0 34776 0 1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_43_354
timestamp 1586364061
transform 1 0 33672 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_43_367
timestamp 1586364061
transform 1 0 34868 0 1 25568
box -38 -48 774 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 36616 0 1 25568
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 36432 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 35880 0 1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_43_375
timestamp 1586364061
transform 1 0 35604 0 1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_43_380
timestamp 1586364061
transform 1 0 36064 0 1 25568
box -38 -48 406 592
use scs8hd_conb_1  _63_
timestamp 1586364061
transform 1 0 39192 0 1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 38548 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 38916 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 39836 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_405
timestamp 1586364061
transform 1 0 38364 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_409
timestamp 1586364061
transform 1 0 38732 0 1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_43_413
timestamp 1586364061
transform 1 0 39100 0 1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_43_417
timestamp 1586364061
transform 1 0 39468 0 1 25568
box -38 -48 406 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 40480 0 1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_524
timestamp 1586364061
transform 1 0 40388 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 42136 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 40204 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 41492 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_423
timestamp 1586364061
transform 1 0 40020 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_437
timestamp 1586364061
transform 1 0 41308 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_441
timestamp 1586364061
transform 1 0 41676 0 1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_43_445
timestamp 1586364061
transform 1 0 42044 0 1 25568
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 42320 0 1 25568
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_43_467
timestamp 1586364061
transform 1 0 44068 0 1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_43_471
timestamp 1586364061
transform 1 0 44436 0 1 25568
box -38 -48 130 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1586364061
transform 1 0 46092 0 1 25568
box -38 -48 866 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_3_
timestamp 1586364061
transform 1 0 44804 0 1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_525
timestamp 1586364061
transform 1 0 46000 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 45816 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 45448 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 44528 0 1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_43_474
timestamp 1586364061
transform 1 0 44712 0 1 25568
box -38 -48 130 592
use scs8hd_decap_3  FILLER_43_479
timestamp 1586364061
transform 1 0 45172 0 1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_43_484
timestamp 1586364061
transform 1 0 45632 0 1 25568
box -38 -48 222 592
use scs8hd_decap_3  PHY_87
timestamp 1586364061
transform -1 0 48852 0 1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 47104 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 47472 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_498
timestamp 1586364061
transform 1 0 46920 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_502
timestamp 1586364061
transform 1 0 47288 0 1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_43_506
timestamp 1586364061
transform 1 0 47656 0 1 25568
box -38 -48 774 592
use scs8hd_fill_2  FILLER_43_514
timestamp 1586364061
transform 1 0 48392 0 1 25568
box -38 -48 222 592
use scs8hd_decap_3  PHY_88
timestamp 1586364061
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_44_3
timestamp 1586364061
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_15
timestamp 1586364061
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_526
timestamp 1586364061
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_4  FILLER_44_27
timestamp 1586364061
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use scs8hd_decap_12  FILLER_44_32
timestamp 1586364061
transform 1 0 4048 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_44
timestamp 1586364061
transform 1 0 5152 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_56
timestamp 1586364061
transform 1 0 6256 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_68
timestamp 1586364061
transform 1 0 7360 0 -1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_527
timestamp 1586364061
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_44_80
timestamp 1586364061
transform 1 0 8464 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_93
timestamp 1586364061
transform 1 0 9660 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_105
timestamp 1586364061
transform 1 0 10764 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_117
timestamp 1586364061
transform 1 0 11868 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_129
timestamp 1586364061
transform 1 0 12972 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_141
timestamp 1586364061
transform 1 0 14076 0 -1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_528
timestamp 1586364061
transform 1 0 15180 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_44_154
timestamp 1586364061
transform 1 0 15272 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_166
timestamp 1586364061
transform 1 0 16376 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_178
timestamp 1586364061
transform 1 0 17480 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_190
timestamp 1586364061
transform 1 0 18584 0 -1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_529
timestamp 1586364061
transform 1 0 20792 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_44_202
timestamp 1586364061
transform 1 0 19688 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_215
timestamp 1586364061
transform 1 0 20884 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_227
timestamp 1586364061
transform 1 0 21988 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_239
timestamp 1586364061
transform 1 0 23092 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_251
timestamp 1586364061
transform 1 0 24196 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_263
timestamp 1586364061
transform 1 0 25300 0 -1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_530
timestamp 1586364061
transform 1 0 26404 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_44_276
timestamp 1586364061
transform 1 0 26496 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_288
timestamp 1586364061
transform 1 0 27600 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_300
timestamp 1586364061
transform 1 0 28704 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_312
timestamp 1586364061
transform 1 0 29808 0 -1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_531
timestamp 1586364061
transform 1 0 32016 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_44_324
timestamp 1586364061
transform 1 0 30912 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_337
timestamp 1586364061
transform 1 0 32108 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_349
timestamp 1586364061
transform 1 0 33212 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_361
timestamp 1586364061
transform 1 0 34316 0 -1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_532
timestamp 1586364061
transform 1 0 37628 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 35788 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 36616 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_373
timestamp 1586364061
transform 1 0 35420 0 -1 26656
box -38 -48 406 592
use scs8hd_decap_6  FILLER_44_379
timestamp 1586364061
transform 1 0 35972 0 -1 26656
box -38 -48 590 592
use scs8hd_fill_1  FILLER_44_385
timestamp 1586364061
transform 1 0 36524 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_8  FILLER_44_388
timestamp 1586364061
transform 1 0 36800 0 -1 26656
box -38 -48 774 592
use scs8hd_fill_1  FILLER_44_396
timestamp 1586364061
transform 1 0 37536 0 -1 26656
box -38 -48 130 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 38456 0 -1 26656
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 38272 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_6  FILLER_44_398
timestamp 1586364061
transform 1 0 37720 0 -1 26656
box -38 -48 590 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 41308 0 -1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 40480 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 41124 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_3  FILLER_44_425
timestamp 1586364061
transform 1 0 40204 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_4  FILLER_44_430
timestamp 1586364061
transform 1 0 40664 0 -1 26656
box -38 -48 406 592
use scs8hd_fill_1  FILLER_44_434
timestamp 1586364061
transform 1 0 41032 0 -1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_44_446
timestamp 1586364061
transform 1 0 42136 0 -1 26656
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0_
timestamp 1586364061
transform 1 0 43332 0 -1 26656
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_533
timestamp 1586364061
transform 1 0 43240 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 42320 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_0__A
timestamp 1586364061
transform 1 0 43884 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 44344 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_8  FILLER_44_450
timestamp 1586364061
transform 1 0 42504 0 -1 26656
box -38 -48 774 592
use scs8hd_fill_2  FILLER_44_463
timestamp 1586364061
transform 1 0 43700 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_3  FILLER_44_467
timestamp 1586364061
transform 1 0 44068 0 -1 26656
box -38 -48 314 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1586364061
transform 1 0 44528 0 -1 26656
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 46092 0 -1 26656
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_44_481
timestamp 1586364061
transform 1 0 45356 0 -1 26656
box -38 -48 774 592
use scs8hd_decap_3  PHY_89
timestamp 1586364061
transform -1 0 48852 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_8  FILLER_44_508
timestamp 1586364061
transform 1 0 47840 0 -1 26656
box -38 -48 774 592
use scs8hd_decap_3  PHY_90
timestamp 1586364061
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_45_3
timestamp 1586364061
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_15
timestamp 1586364061
transform 1 0 2484 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_27
timestamp 1586364061
transform 1 0 3588 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_39
timestamp 1586364061
transform 1 0 4692 0 1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_534
timestamp 1586364061
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use scs8hd_decap_8  FILLER_45_51
timestamp 1586364061
transform 1 0 5796 0 1 26656
box -38 -48 774 592
use scs8hd_fill_2  FILLER_45_59
timestamp 1586364061
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_45_62
timestamp 1586364061
transform 1 0 6808 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_74
timestamp 1586364061
transform 1 0 7912 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_86
timestamp 1586364061
transform 1 0 9016 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_98
timestamp 1586364061
transform 1 0 10120 0 1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_535
timestamp 1586364061
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_45_110
timestamp 1586364061
transform 1 0 11224 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_123
timestamp 1586364061
transform 1 0 12420 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_135
timestamp 1586364061
transform 1 0 13524 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_147
timestamp 1586364061
transform 1 0 14628 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_159
timestamp 1586364061
transform 1 0 15732 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_171
timestamp 1586364061
transform 1 0 16836 0 1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_536
timestamp 1586364061
transform 1 0 17940 0 1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_45_184
timestamp 1586364061
transform 1 0 18032 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_196
timestamp 1586364061
transform 1 0 19136 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_208
timestamp 1586364061
transform 1 0 20240 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_220
timestamp 1586364061
transform 1 0 21344 0 1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_537
timestamp 1586364061
transform 1 0 23552 0 1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_45_232
timestamp 1586364061
transform 1 0 22448 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_245
timestamp 1586364061
transform 1 0 23644 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_257
timestamp 1586364061
transform 1 0 24748 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_269
timestamp 1586364061
transform 1 0 25852 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_281
timestamp 1586364061
transform 1 0 26956 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_293
timestamp 1586364061
transform 1 0 28060 0 1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_538
timestamp 1586364061
transform 1 0 29164 0 1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_45_306
timestamp 1586364061
transform 1 0 29256 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_318
timestamp 1586364061
transform 1 0 30360 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_330
timestamp 1586364061
transform 1 0 31464 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_342
timestamp 1586364061
transform 1 0 32568 0 1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_539
timestamp 1586364061
transform 1 0 34776 0 1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_45_354
timestamp 1586364061
transform 1 0 33672 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_45_367
timestamp 1586364061
transform 1 0 34868 0 1 26656
box -38 -48 774 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 35788 0 1 26656
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 35604 0 1 26656
box -38 -48 222 592
use scs8hd_decap_6  FILLER_45_396
timestamp 1586364061
transform 1 0 37536 0 1 26656
box -38 -48 590 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 38272 0 1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__CLK
timestamp 1586364061
transform 1 0 39284 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 38088 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14__D
timestamp 1586364061
transform 1 0 39652 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_413
timestamp 1586364061
transform 1 0 39100 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_417
timestamp 1586364061
transform 1 0 39468 0 1 26656
box -38 -48 222 592
use scs8hd_decap_6  FILLER_45_421
timestamp 1586364061
transform 1 0 39836 0 1 26656
box -38 -48 590 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16_
timestamp 1586364061
transform 1 0 41308 0 1 26656
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_540
timestamp 1586364061
transform 1 0 40388 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__CLK
timestamp 1586364061
transform 1 0 41124 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_16__D
timestamp 1586364061
transform 1 0 40756 0 1 26656
box -38 -48 222 592
use scs8hd_decap_3  FILLER_45_428
timestamp 1586364061
transform 1 0 40480 0 1 26656
box -38 -48 314 592
use scs8hd_fill_2  FILLER_45_433
timestamp 1586364061
transform 1 0 40940 0 1 26656
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1586364061
transform 1 0 43792 0 1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 43608 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 43240 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_456
timestamp 1586364061
transform 1 0 43056 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_460
timestamp 1586364061
transform 1 0 43424 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_481
timestamp 1586364061
transform 1 0 45356 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_477
timestamp 1586364061
transform 1 0 44988 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_473
timestamp 1586364061
transform 1 0 44620 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 45172 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4__A
timestamp 1586364061
transform 1 0 44804 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__CLK
timestamp 1586364061
transform 1 0 45540 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_489
timestamp 1586364061
transform 1 0 46092 0 1 26656
box -38 -48 222 592
use scs8hd_decap_3  FILLER_45_485
timestamp 1586364061
transform 1 0 45724 0 1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4__D
timestamp 1586364061
transform 1 0 46276 0 1 26656
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_541
timestamp 1586364061
transform 1 0 46000 0 1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_45_493
timestamp 1586364061
transform 1 0 46460 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_3  PHY_91
timestamp 1586364061
transform -1 0 48852 0 1 26656
box -38 -48 314 592
use scs8hd_decap_8  FILLER_45_505
timestamp 1586364061
transform 1 0 47564 0 1 26656
box -38 -48 774 592
use scs8hd_decap_3  FILLER_45_513
timestamp 1586364061
transform 1 0 48300 0 1 26656
box -38 -48 314 592
use scs8hd_decap_3  PHY_92
timestamp 1586364061
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_94
timestamp 1586364061
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use scs8hd_decap_12  FILLER_46_3
timestamp 1586364061
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_15
timestamp 1586364061
transform 1 0 2484 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_3
timestamp 1586364061
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_15
timestamp 1586364061
transform 1 0 2484 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_542
timestamp 1586364061
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_46_27
timestamp 1586364061
transform 1 0 3588 0 -1 27744
box -38 -48 406 592
use scs8hd_decap_12  FILLER_46_32
timestamp 1586364061
transform 1 0 4048 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_44
timestamp 1586364061
transform 1 0 5152 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_27
timestamp 1586364061
transform 1 0 3588 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_39
timestamp 1586364061
transform 1 0 4692 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_550
timestamp 1586364061
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_56
timestamp 1586364061
transform 1 0 6256 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_68
timestamp 1586364061
transform 1 0 7360 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_47_51
timestamp 1586364061
transform 1 0 5796 0 1 27744
box -38 -48 774 592
use scs8hd_fill_2  FILLER_47_59
timestamp 1586364061
transform 1 0 6532 0 1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_47_62
timestamp 1586364061
transform 1 0 6808 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_74
timestamp 1586364061
transform 1 0 7912 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_543
timestamp 1586364061
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_80
timestamp 1586364061
transform 1 0 8464 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_93
timestamp 1586364061
transform 1 0 9660 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_86
timestamp 1586364061
transform 1 0 9016 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_98
timestamp 1586364061
transform 1 0 10120 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_551
timestamp 1586364061
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_105
timestamp 1586364061
transform 1 0 10764 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_117
timestamp 1586364061
transform 1 0 11868 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_110
timestamp 1586364061
transform 1 0 11224 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_123
timestamp 1586364061
transform 1 0 12420 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_129
timestamp 1586364061
transform 1 0 12972 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_141
timestamp 1586364061
transform 1 0 14076 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_135
timestamp 1586364061
transform 1 0 13524 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_147
timestamp 1586364061
transform 1 0 14628 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_544
timestamp 1586364061
transform 1 0 15180 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_154
timestamp 1586364061
transform 1 0 15272 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_166
timestamp 1586364061
transform 1 0 16376 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_159
timestamp 1586364061
transform 1 0 15732 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_171
timestamp 1586364061
transform 1 0 16836 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_552
timestamp 1586364061
transform 1 0 17940 0 1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_178
timestamp 1586364061
transform 1 0 17480 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_190
timestamp 1586364061
transform 1 0 18584 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_184
timestamp 1586364061
transform 1 0 18032 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_196
timestamp 1586364061
transform 1 0 19136 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_545
timestamp 1586364061
transform 1 0 20792 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_202
timestamp 1586364061
transform 1 0 19688 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_215
timestamp 1586364061
transform 1 0 20884 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_208
timestamp 1586364061
transform 1 0 20240 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_220
timestamp 1586364061
transform 1 0 21344 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_553
timestamp 1586364061
transform 1 0 23552 0 1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_227
timestamp 1586364061
transform 1 0 21988 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_239
timestamp 1586364061
transform 1 0 23092 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_232
timestamp 1586364061
transform 1 0 22448 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_245
timestamp 1586364061
transform 1 0 23644 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_251
timestamp 1586364061
transform 1 0 24196 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_263
timestamp 1586364061
transform 1 0 25300 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_257
timestamp 1586364061
transform 1 0 24748 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_269
timestamp 1586364061
transform 1 0 25852 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_546
timestamp 1586364061
transform 1 0 26404 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_276
timestamp 1586364061
transform 1 0 26496 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_288
timestamp 1586364061
transform 1 0 27600 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_281
timestamp 1586364061
transform 1 0 26956 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_293
timestamp 1586364061
transform 1 0 28060 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_554
timestamp 1586364061
transform 1 0 29164 0 1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_300
timestamp 1586364061
transform 1 0 28704 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_312
timestamp 1586364061
transform 1 0 29808 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_306
timestamp 1586364061
transform 1 0 29256 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_318
timestamp 1586364061
transform 1 0 30360 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_547
timestamp 1586364061
transform 1 0 32016 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_324
timestamp 1586364061
transform 1 0 30912 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_337
timestamp 1586364061
transform 1 0 32108 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_330
timestamp 1586364061
transform 1 0 31464 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_342
timestamp 1586364061
transform 1 0 32568 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_555
timestamp 1586364061
transform 1 0 34776 0 1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_349
timestamp 1586364061
transform 1 0 33212 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_361
timestamp 1586364061
transform 1 0 34316 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_354
timestamp 1586364061
transform 1 0 33672 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_367
timestamp 1586364061
transform 1 0 34868 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_548
timestamp 1586364061
transform 1 0 37628 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_373
timestamp 1586364061
transform 1 0 35420 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_385
timestamp 1586364061
transform 1 0 36524 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_379
timestamp 1586364061
transform 1 0 35972 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_391
timestamp 1586364061
transform 1 0 37076 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_47_403
timestamp 1586364061
transform 1 0 38180 0 1 27744
box -38 -48 774 592
use scs8hd_decap_6  FILLER_46_406
timestamp 1586364061
transform 1 0 38456 0 -1 27744
box -38 -48 590 592
use scs8hd_decap_3  FILLER_46_401
timestamp 1586364061
transform 1 0 37996 0 -1 27744
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 38272 0 -1 27744
box -38 -48 222 592
use scs8hd_conb_1  _32_
timestamp 1586364061
transform 1 0 37720 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_4  FILLER_47_417
timestamp 1586364061
transform 1 0 39468 0 1 27744
box -38 -48 406 592
use scs8hd_fill_2  FILLER_47_413
timestamp 1586364061
transform 1 0 39100 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_46_412
timestamp 1586364061
transform 1 0 39008 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__D
timestamp 1586364061
transform 1 0 39836 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__D
timestamp 1586364061
transform 1 0 39284 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13__CLK
timestamp 1586364061
transform 1 0 38916 0 1 27744
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_14_
timestamp 1586364061
transform 1 0 39100 0 -1 27744
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_47_423
timestamp 1586364061
transform 1 0 40020 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_432
timestamp 1586364061
transform 1 0 40848 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 41032 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15__CLK
timestamp 1586364061
transform 1 0 40204 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_556
timestamp 1586364061
transform 1 0 40388 0 1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_47_447
timestamp 1586364061
transform 1 0 42228 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_436
timestamp 1586364061
transform 1 0 41216 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1586364061
transform 1 0 41400 0 -1 27744
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1586364061
transform 1 0 41584 0 -1 27744
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_15_
timestamp 1586364061
transform 1 0 40480 0 1 27744
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_47_451
timestamp 1586364061
transform 1 0 42596 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_453
timestamp 1586364061
transform 1 0 42780 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_449
timestamp 1586364061
transform 1 0 42412 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 42596 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 42964 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 42780 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1586364061
transform 1 0 42412 0 1 27744
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1586364061
transform 1 0 42964 0 1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_47_464
timestamp 1586364061
transform 1 0 43792 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_46_466
timestamp 1586364061
transform 1 0 43976 0 -1 27744
box -38 -48 130 592
use scs8hd_fill_1  FILLER_46_463
timestamp 1586364061
transform 1 0 43700 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_46_459
timestamp 1586364061
transform 1 0 43332 0 -1 27744
box -38 -48 406 592
use scs8hd_fill_1  FILLER_46_457
timestamp 1586364061
transform 1 0 43148 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5__A
timestamp 1586364061
transform 1 0 43976 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 43792 0 -1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_549
timestamp 1586364061
transform 1 0 43240 0 -1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_47_468
timestamp 1586364061
transform 1 0 44160 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_471
timestamp 1586364061
transform 1 0 44436 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 44344 0 1 27744
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_4_
timestamp 1586364061
transform 1 0 44068 0 -1 27744
box -38 -48 406 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6_
timestamp 1586364061
transform 1 0 44528 0 1 27744
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 44620 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_475
timestamp 1586364061
transform 1 0 44804 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_476
timestamp 1586364061
transform 1 0 44896 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_6__A
timestamp 1586364061
transform 1 0 45080 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 44988 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_4  FILLER_46_479
timestamp 1586364061
transform 1 0 45172 0 -1 27744
box -38 -48 406 592
use scs8hd_fill_2  FILLER_47_480
timestamp 1586364061
transform 1 0 45264 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__D
timestamp 1586364061
transform 1 0 45448 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_484
timestamp 1586364061
transform 1 0 45632 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5__CLK
timestamp 1586364061
transform 1 0 45816 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_557
timestamp 1586364061
transform 1 0 46000 0 1 27744
box -38 -48 130 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1586364061
transform 1 0 46092 0 1 27744
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_4_
timestamp 1586364061
transform 1 0 45540 0 -1 27744
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_47_506
timestamp 1586364061
transform 1 0 47656 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_502
timestamp 1586364061
transform 1 0 47288 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_498
timestamp 1586364061
transform 1 0 46920 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 47840 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 47472 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 47104 0 1 27744
box -38 -48 222 592
use scs8hd_decap_6  FILLER_47_510
timestamp 1586364061
transform 1 0 48024 0 1 27744
box -38 -48 590 592
use scs8hd_fill_2  FILLER_46_514
timestamp 1586364061
transform 1 0 48392 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_3  PHY_95
timestamp 1586364061
transform -1 0 48852 0 1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_93
timestamp 1586364061
transform -1 0 48852 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_12  FILLER_46_502
timestamp 1586364061
transform 1 0 47288 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_3  PHY_96
timestamp 1586364061
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_48_3
timestamp 1586364061
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_15
timestamp 1586364061
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_558
timestamp 1586364061
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_4  FILLER_48_27
timestamp 1586364061
transform 1 0 3588 0 -1 28832
box -38 -48 406 592
use scs8hd_decap_12  FILLER_48_32
timestamp 1586364061
transform 1 0 4048 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_44
timestamp 1586364061
transform 1 0 5152 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_56
timestamp 1586364061
transform 1 0 6256 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_68
timestamp 1586364061
transform 1 0 7360 0 -1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_559
timestamp 1586364061
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_48_80
timestamp 1586364061
transform 1 0 8464 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_93
timestamp 1586364061
transform 1 0 9660 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_105
timestamp 1586364061
transform 1 0 10764 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_117
timestamp 1586364061
transform 1 0 11868 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_129
timestamp 1586364061
transform 1 0 12972 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_141
timestamp 1586364061
transform 1 0 14076 0 -1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_560
timestamp 1586364061
transform 1 0 15180 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_48_154
timestamp 1586364061
transform 1 0 15272 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_166
timestamp 1586364061
transform 1 0 16376 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_178
timestamp 1586364061
transform 1 0 17480 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_190
timestamp 1586364061
transform 1 0 18584 0 -1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_561
timestamp 1586364061
transform 1 0 20792 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_48_202
timestamp 1586364061
transform 1 0 19688 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_215
timestamp 1586364061
transform 1 0 20884 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_227
timestamp 1586364061
transform 1 0 21988 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_239
timestamp 1586364061
transform 1 0 23092 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_251
timestamp 1586364061
transform 1 0 24196 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_263
timestamp 1586364061
transform 1 0 25300 0 -1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_562
timestamp 1586364061
transform 1 0 26404 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_48_276
timestamp 1586364061
transform 1 0 26496 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_288
timestamp 1586364061
transform 1 0 27600 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_300
timestamp 1586364061
transform 1 0 28704 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_312
timestamp 1586364061
transform 1 0 29808 0 -1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_563
timestamp 1586364061
transform 1 0 32016 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_48_324
timestamp 1586364061
transform 1 0 30912 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_337
timestamp 1586364061
transform 1 0 32108 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_349
timestamp 1586364061
transform 1 0 33212 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_361
timestamp 1586364061
transform 1 0 34316 0 -1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_564
timestamp 1586364061
transform 1 0 37628 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_48_373
timestamp 1586364061
transform 1 0 35420 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_385
timestamp 1586364061
transform 1 0 36524 0 -1 28832
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_13_
timestamp 1586364061
transform 1 0 38916 0 -1 28832
box -38 -48 1786 592
use scs8hd_decap_12  FILLER_48_398
timestamp 1586364061
transform 1 0 37720 0 -1 28832
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_48_410
timestamp 1586364061
transform 1 0 38824 0 -1 28832
box -38 -48 130 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1586364061
transform 1 0 41400 0 -1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1586364061
transform 1 0 41216 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1586364061
transform 1 0 40848 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_430
timestamp 1586364061
transform 1 0 40664 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_434
timestamp 1586364061
transform 1 0 41032 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_447
timestamp 1586364061
transform 1 0 42228 0 -1 28832
box -38 -48 222 592
use scs8hd_buf_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.scs8hd_buf_2_5_
timestamp 1586364061
transform 1 0 43332 0 -1 28832
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_565
timestamp 1586364061
transform 1 0 43240 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1586364061
transform 1 0 42412 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 42780 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_451
timestamp 1586364061
transform 1 0 42596 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_48_455
timestamp 1586364061
transform 1 0 42964 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_8  FILLER_48_463
timestamp 1586364061
transform 1 0 43700 0 -1 28832
box -38 -48 774 592
use scs8hd_fill_1  FILLER_48_471
timestamp 1586364061
transform 1 0 44436 0 -1 28832
box -38 -48 130 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1586364061
transform 1 0 44528 0 -1 28832
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_5_
timestamp 1586364061
transform 1 0 46092 0 -1 28832
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_48_481
timestamp 1586364061
transform 1 0 45356 0 -1 28832
box -38 -48 774 592
use scs8hd_decap_3  PHY_97
timestamp 1586364061
transform -1 0 48852 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_8  FILLER_48_508
timestamp 1586364061
transform 1 0 47840 0 -1 28832
box -38 -48 774 592
use scs8hd_decap_3  PHY_98
timestamp 1586364061
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_49_3
timestamp 1586364061
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_15
timestamp 1586364061
transform 1 0 2484 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_27
timestamp 1586364061
transform 1 0 3588 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_39
timestamp 1586364061
transform 1 0 4692 0 1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_566
timestamp 1586364061
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use scs8hd_decap_8  FILLER_49_51
timestamp 1586364061
transform 1 0 5796 0 1 28832
box -38 -48 774 592
use scs8hd_fill_2  FILLER_49_59
timestamp 1586364061
transform 1 0 6532 0 1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_49_62
timestamp 1586364061
transform 1 0 6808 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_74
timestamp 1586364061
transform 1 0 7912 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_86
timestamp 1586364061
transform 1 0 9016 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_98
timestamp 1586364061
transform 1 0 10120 0 1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_567
timestamp 1586364061
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_49_110
timestamp 1586364061
transform 1 0 11224 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_123
timestamp 1586364061
transform 1 0 12420 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_135
timestamp 1586364061
transform 1 0 13524 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_147
timestamp 1586364061
transform 1 0 14628 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_159
timestamp 1586364061
transform 1 0 15732 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_171
timestamp 1586364061
transform 1 0 16836 0 1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_568
timestamp 1586364061
transform 1 0 17940 0 1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_49_184
timestamp 1586364061
transform 1 0 18032 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_196
timestamp 1586364061
transform 1 0 19136 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_208
timestamp 1586364061
transform 1 0 20240 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_220
timestamp 1586364061
transform 1 0 21344 0 1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_569
timestamp 1586364061
transform 1 0 23552 0 1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_49_232
timestamp 1586364061
transform 1 0 22448 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_245
timestamp 1586364061
transform 1 0 23644 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_257
timestamp 1586364061
transform 1 0 24748 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_269
timestamp 1586364061
transform 1 0 25852 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_281
timestamp 1586364061
transform 1 0 26956 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_293
timestamp 1586364061
transform 1 0 28060 0 1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_570
timestamp 1586364061
transform 1 0 29164 0 1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_49_306
timestamp 1586364061
transform 1 0 29256 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_318
timestamp 1586364061
transform 1 0 30360 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_330
timestamp 1586364061
transform 1 0 31464 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_342
timestamp 1586364061
transform 1 0 32568 0 1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_571
timestamp 1586364061
transform 1 0 34776 0 1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_49_354
timestamp 1586364061
transform 1 0 33672 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_367
timestamp 1586364061
transform 1 0 34868 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_379
timestamp 1586364061
transform 1 0 35972 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_391
timestamp 1586364061
transform 1 0 37076 0 1 28832
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__CLK
timestamp 1586364061
transform 1 0 39100 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12__D
timestamp 1586364061
transform 1 0 39468 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1586364061
transform 1 0 39836 0 1 28832
box -38 -48 222 592
use scs8hd_decap_8  FILLER_49_403
timestamp 1586364061
transform 1 0 38180 0 1 28832
box -38 -48 774 592
use scs8hd_fill_2  FILLER_49_411
timestamp 1586364061
transform 1 0 38916 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_415
timestamp 1586364061
transform 1 0 39284 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_419
timestamp 1586364061
transform 1 0 39652 0 1 28832
box -38 -48 222 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1586364061
transform 1 0 40480 0 1 28832
box -38 -48 866 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1586364061
transform 1 0 42136 0 1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_572
timestamp 1586364061
transform 1 0 40388 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1586364061
transform 1 0 41676 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1586364061
transform 1 0 40204 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_423
timestamp 1586364061
transform 1 0 40020 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_437
timestamp 1586364061
transform 1 0 41308 0 1 28832
box -38 -48 406 592
use scs8hd_decap_3  FILLER_49_443
timestamp 1586364061
transform 1 0 41860 0 1 28832
box -38 -48 314 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1586364061
transform 1 0 44436 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 44252 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 43148 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 43884 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 43516 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_455
timestamp 1586364061
transform 1 0 42964 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_459
timestamp 1586364061
transform 1 0 43332 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_463
timestamp 1586364061
transform 1 0 43700 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_467
timestamp 1586364061
transform 1 0 44068 0 1 28832
box -38 -48 222 592
use scs8hd_buf_2  _74_
timestamp 1586364061
transform 1 0 46736 0 1 28832
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_573
timestamp 1586364061
transform 1 0 46000 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__CLK
timestamp 1586364061
transform 1 0 45448 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7__D
timestamp 1586364061
transform 1 0 45816 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_480
timestamp 1586364061
transform 1 0 45264 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_484
timestamp 1586364061
transform 1 0 45632 0 1 28832
box -38 -48 222 592
use scs8hd_decap_6  FILLER_49_489
timestamp 1586364061
transform 1 0 46092 0 1 28832
box -38 -48 590 592
use scs8hd_fill_1  FILLER_49_495
timestamp 1586364061
transform 1 0 46644 0 1 28832
box -38 -48 130 592
use scs8hd_decap_3  PHY_99
timestamp 1586364061
transform -1 0 48852 0 1 28832
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__74__A
timestamp 1586364061
transform 1 0 47288 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_500
timestamp 1586364061
transform 1 0 47104 0 1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_49_504
timestamp 1586364061
transform 1 0 47472 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_3  PHY_100
timestamp 1586364061
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_50_3
timestamp 1586364061
transform 1 0 1380 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_15
timestamp 1586364061
transform 1 0 2484 0 -1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_574
timestamp 1586364061
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_4  FILLER_50_27
timestamp 1586364061
transform 1 0 3588 0 -1 29920
box -38 -48 406 592
use scs8hd_decap_12  FILLER_50_32
timestamp 1586364061
transform 1 0 4048 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_44
timestamp 1586364061
transform 1 0 5152 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_56
timestamp 1586364061
transform 1 0 6256 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_68
timestamp 1586364061
transform 1 0 7360 0 -1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_575
timestamp 1586364061
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_50_80
timestamp 1586364061
transform 1 0 8464 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_93
timestamp 1586364061
transform 1 0 9660 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_105
timestamp 1586364061
transform 1 0 10764 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_117
timestamp 1586364061
transform 1 0 11868 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_129
timestamp 1586364061
transform 1 0 12972 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_141
timestamp 1586364061
transform 1 0 14076 0 -1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_576
timestamp 1586364061
transform 1 0 15180 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_50_154
timestamp 1586364061
transform 1 0 15272 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_166
timestamp 1586364061
transform 1 0 16376 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_178
timestamp 1586364061
transform 1 0 17480 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_190
timestamp 1586364061
transform 1 0 18584 0 -1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_577
timestamp 1586364061
transform 1 0 20792 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_50_202
timestamp 1586364061
transform 1 0 19688 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_215
timestamp 1586364061
transform 1 0 20884 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_227
timestamp 1586364061
transform 1 0 21988 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_239
timestamp 1586364061
transform 1 0 23092 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_251
timestamp 1586364061
transform 1 0 24196 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_263
timestamp 1586364061
transform 1 0 25300 0 -1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_578
timestamp 1586364061
transform 1 0 26404 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_50_276
timestamp 1586364061
transform 1 0 26496 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_288
timestamp 1586364061
transform 1 0 27600 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_300
timestamp 1586364061
transform 1 0 28704 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_312
timestamp 1586364061
transform 1 0 29808 0 -1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_579
timestamp 1586364061
transform 1 0 32016 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_50_324
timestamp 1586364061
transform 1 0 30912 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_337
timestamp 1586364061
transform 1 0 32108 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_349
timestamp 1586364061
transform 1 0 33212 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_361
timestamp 1586364061
transform 1 0 34316 0 -1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_580
timestamp 1586364061
transform 1 0 37628 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_50_373
timestamp 1586364061
transform 1 0 35420 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_385
timestamp 1586364061
transform 1 0 36524 0 -1 29920
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_12_
timestamp 1586364061
transform 1 0 39100 0 -1 29920
box -38 -48 1786 592
use scs8hd_decap_12  FILLER_50_398
timestamp 1586364061
transform 1 0 37720 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_50_410
timestamp 1586364061
transform 1 0 38824 0 -1 29920
box -38 -48 314 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1586364061
transform 1 0 41676 0 -1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1586364061
transform 1 0 41492 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_6  FILLER_50_432
timestamp 1586364061
transform 1 0 40848 0 -1 29920
box -38 -48 590 592
use scs8hd_fill_1  FILLER_50_438
timestamp 1586364061
transform 1 0 41400 0 -1 29920
box -38 -48 130 592
use scs8hd_fill_2  FILLER_50_450
timestamp 1586364061
transform 1 0 42504 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_50_454
timestamp 1586364061
transform 1 0 42872 0 -1 29920
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__D
timestamp 1586364061
transform 1 0 42688 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_459
timestamp 1586364061
transform 1 0 43332 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__CLK
timestamp 1586364061
transform 1 0 43516 0 -1 29920
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_581
timestamp 1586364061
transform 1 0 43240 0 -1 29920
box -38 -48 130 592
use scs8hd_fill_2  FILLER_50_463
timestamp 1586364061
transform 1 0 43700 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9__D
timestamp 1586364061
transform 1 0 43884 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_50_467
timestamp 1586364061
transform 1 0 44068 0 -1 29920
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 44436 0 -1 29920
box -38 -48 222 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_7_
timestamp 1586364061
transform 1 0 45172 0 -1 29920
box -38 -48 1786 592
use scs8hd_decap_6  FILLER_50_473
timestamp 1586364061
transform 1 0 44620 0 -1 29920
box -38 -48 590 592
use scs8hd_decap_3  PHY_101
timestamp 1586364061
transform -1 0 48852 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_50_498
timestamp 1586364061
transform 1 0 46920 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_50_510
timestamp 1586364061
transform 1 0 48024 0 -1 29920
box -38 -48 590 592
use scs8hd_decap_3  PHY_102
timestamp 1586364061
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_51_3
timestamp 1586364061
transform 1 0 1380 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_15
timestamp 1586364061
transform 1 0 2484 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_27
timestamp 1586364061
transform 1 0 3588 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_39
timestamp 1586364061
transform 1 0 4692 0 1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_582
timestamp 1586364061
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use scs8hd_decap_8  FILLER_51_51
timestamp 1586364061
transform 1 0 5796 0 1 29920
box -38 -48 774 592
use scs8hd_fill_2  FILLER_51_59
timestamp 1586364061
transform 1 0 6532 0 1 29920
box -38 -48 222 592
use scs8hd_decap_12  FILLER_51_62
timestamp 1586364061
transform 1 0 6808 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_74
timestamp 1586364061
transform 1 0 7912 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_86
timestamp 1586364061
transform 1 0 9016 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_98
timestamp 1586364061
transform 1 0 10120 0 1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_583
timestamp 1586364061
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_51_110
timestamp 1586364061
transform 1 0 11224 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_123
timestamp 1586364061
transform 1 0 12420 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_135
timestamp 1586364061
transform 1 0 13524 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_147
timestamp 1586364061
transform 1 0 14628 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_159
timestamp 1586364061
transform 1 0 15732 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_171
timestamp 1586364061
transform 1 0 16836 0 1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_584
timestamp 1586364061
transform 1 0 17940 0 1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_51_184
timestamp 1586364061
transform 1 0 18032 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_196
timestamp 1586364061
transform 1 0 19136 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_208
timestamp 1586364061
transform 1 0 20240 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_220
timestamp 1586364061
transform 1 0 21344 0 1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_585
timestamp 1586364061
transform 1 0 23552 0 1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_51_232
timestamp 1586364061
transform 1 0 22448 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_245
timestamp 1586364061
transform 1 0 23644 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_257
timestamp 1586364061
transform 1 0 24748 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_269
timestamp 1586364061
transform 1 0 25852 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_281
timestamp 1586364061
transform 1 0 26956 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_293
timestamp 1586364061
transform 1 0 28060 0 1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_586
timestamp 1586364061
transform 1 0 29164 0 1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_51_306
timestamp 1586364061
transform 1 0 29256 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_318
timestamp 1586364061
transform 1 0 30360 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_330
timestamp 1586364061
transform 1 0 31464 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_342
timestamp 1586364061
transform 1 0 32568 0 1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_587
timestamp 1586364061
transform 1 0 34776 0 1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_51_354
timestamp 1586364061
transform 1 0 33672 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_367
timestamp 1586364061
transform 1 0 34868 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_379
timestamp 1586364061
transform 1 0 35972 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_391
timestamp 1586364061
transform 1 0 37076 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_403
timestamp 1586364061
transform 1 0 38180 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_415
timestamp 1586364061
transform 1 0 39284 0 1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_588
timestamp 1586364061
transform 1 0 40388 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1586364061
transform 1 0 41676 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1586364061
transform 1 0 42044 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1586364061
transform 1 0 41308 0 1 29920
box -38 -48 222 592
use scs8hd_decap_8  FILLER_51_428
timestamp 1586364061
transform 1 0 40480 0 1 29920
box -38 -48 774 592
use scs8hd_fill_1  FILLER_51_436
timestamp 1586364061
transform 1 0 41216 0 1 29920
box -38 -48 130 592
use scs8hd_fill_2  FILLER_51_439
timestamp 1586364061
transform 1 0 41492 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_443
timestamp 1586364061
transform 1 0 41860 0 1 29920
box -38 -48 222 592
use scs8hd_decap_3  FILLER_51_447
timestamp 1586364061
transform 1 0 42228 0 1 29920
box -38 -48 314 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11_
timestamp 1586364061
transform 1 0 42688 0 1 29920
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_11__CLK
timestamp 1586364061
transform 1 0 42504 0 1 29920
box -38 -48 222 592
use scs8hd_decap_6  FILLER_51_471
timestamp 1586364061
transform 1 0 44436 0 1 29920
box -38 -48 590 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6_
timestamp 1586364061
transform 1 0 46092 0 1 29920
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_589
timestamp 1586364061
transform 1 0 46000 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__CLK
timestamp 1586364061
transform 1 0 45816 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__CLK
timestamp 1586364061
transform 1 0 45448 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8__D
timestamp 1586364061
transform 1 0 45080 0 1 29920
box -38 -48 222 592
use scs8hd_fill_1  FILLER_51_477
timestamp 1586364061
transform 1 0 44988 0 1 29920
box -38 -48 130 592
use scs8hd_fill_2  FILLER_51_480
timestamp 1586364061
transform 1 0 45264 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_484
timestamp 1586364061
transform 1 0 45632 0 1 29920
box -38 -48 222 592
use scs8hd_decap_3  PHY_103
timestamp 1586364061
transform -1 0 48852 0 1 29920
box -38 -48 314 592
use scs8hd_decap_8  FILLER_51_508
timestamp 1586364061
transform 1 0 47840 0 1 29920
box -38 -48 774 592
use scs8hd_decap_3  PHY_104
timestamp 1586364061
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_106
timestamp 1586364061
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use scs8hd_decap_12  FILLER_52_3
timestamp 1586364061
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_15
timestamp 1586364061
transform 1 0 2484 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_3
timestamp 1586364061
transform 1 0 1380 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_15
timestamp 1586364061
transform 1 0 2484 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_590
timestamp 1586364061
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_52_27
timestamp 1586364061
transform 1 0 3588 0 -1 31008
box -38 -48 406 592
use scs8hd_decap_12  FILLER_52_32
timestamp 1586364061
transform 1 0 4048 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_44
timestamp 1586364061
transform 1 0 5152 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_27
timestamp 1586364061
transform 1 0 3588 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_39
timestamp 1586364061
transform 1 0 4692 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_598
timestamp 1586364061
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_56
timestamp 1586364061
transform 1 0 6256 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_68
timestamp 1586364061
transform 1 0 7360 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_53_51
timestamp 1586364061
transform 1 0 5796 0 1 31008
box -38 -48 774 592
use scs8hd_fill_2  FILLER_53_59
timestamp 1586364061
transform 1 0 6532 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_53_62
timestamp 1586364061
transform 1 0 6808 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_74
timestamp 1586364061
transform 1 0 7912 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_591
timestamp 1586364061
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_80
timestamp 1586364061
transform 1 0 8464 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_93
timestamp 1586364061
transform 1 0 9660 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_86
timestamp 1586364061
transform 1 0 9016 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_98
timestamp 1586364061
transform 1 0 10120 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_599
timestamp 1586364061
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_105
timestamp 1586364061
transform 1 0 10764 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_117
timestamp 1586364061
transform 1 0 11868 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_110
timestamp 1586364061
transform 1 0 11224 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_123
timestamp 1586364061
transform 1 0 12420 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_129
timestamp 1586364061
transform 1 0 12972 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_141
timestamp 1586364061
transform 1 0 14076 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_135
timestamp 1586364061
transform 1 0 13524 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_147
timestamp 1586364061
transform 1 0 14628 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_592
timestamp 1586364061
transform 1 0 15180 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_154
timestamp 1586364061
transform 1 0 15272 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_166
timestamp 1586364061
transform 1 0 16376 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_159
timestamp 1586364061
transform 1 0 15732 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_171
timestamp 1586364061
transform 1 0 16836 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_600
timestamp 1586364061
transform 1 0 17940 0 1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_178
timestamp 1586364061
transform 1 0 17480 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_190
timestamp 1586364061
transform 1 0 18584 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_184
timestamp 1586364061
transform 1 0 18032 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_196
timestamp 1586364061
transform 1 0 19136 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_593
timestamp 1586364061
transform 1 0 20792 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_202
timestamp 1586364061
transform 1 0 19688 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_215
timestamp 1586364061
transform 1 0 20884 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_208
timestamp 1586364061
transform 1 0 20240 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_220
timestamp 1586364061
transform 1 0 21344 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_601
timestamp 1586364061
transform 1 0 23552 0 1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_227
timestamp 1586364061
transform 1 0 21988 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_239
timestamp 1586364061
transform 1 0 23092 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_232
timestamp 1586364061
transform 1 0 22448 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_245
timestamp 1586364061
transform 1 0 23644 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_251
timestamp 1586364061
transform 1 0 24196 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_263
timestamp 1586364061
transform 1 0 25300 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_257
timestamp 1586364061
transform 1 0 24748 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_269
timestamp 1586364061
transform 1 0 25852 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_594
timestamp 1586364061
transform 1 0 26404 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_276
timestamp 1586364061
transform 1 0 26496 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_288
timestamp 1586364061
transform 1 0 27600 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_281
timestamp 1586364061
transform 1 0 26956 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_293
timestamp 1586364061
transform 1 0 28060 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_602
timestamp 1586364061
transform 1 0 29164 0 1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_300
timestamp 1586364061
transform 1 0 28704 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_312
timestamp 1586364061
transform 1 0 29808 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_306
timestamp 1586364061
transform 1 0 29256 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_318
timestamp 1586364061
transform 1 0 30360 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_595
timestamp 1586364061
transform 1 0 32016 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_324
timestamp 1586364061
transform 1 0 30912 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_337
timestamp 1586364061
transform 1 0 32108 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_330
timestamp 1586364061
transform 1 0 31464 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_342
timestamp 1586364061
transform 1 0 32568 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_603
timestamp 1586364061
transform 1 0 34776 0 1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_349
timestamp 1586364061
transform 1 0 33212 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_361
timestamp 1586364061
transform 1 0 34316 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_354
timestamp 1586364061
transform 1 0 33672 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_367
timestamp 1586364061
transform 1 0 34868 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_596
timestamp 1586364061
transform 1 0 37628 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_373
timestamp 1586364061
transform 1 0 35420 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_385
timestamp 1586364061
transform 1 0 36524 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_379
timestamp 1586364061
transform 1 0 35972 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_391
timestamp 1586364061
transform 1 0 37076 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_398
timestamp 1586364061
transform 1 0 37720 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_410
timestamp 1586364061
transform 1 0 38824 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_422
timestamp 1586364061
transform 1 0 39928 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_403
timestamp 1586364061
transform 1 0 38180 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_415
timestamp 1586364061
transform 1 0 39284 0 1 31008
box -38 -48 1142 592
use scs8hd_mux2_2  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1586364061
transform 1 0 41676 0 -1 31008
box -38 -48 866 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10_
timestamp 1586364061
transform 1 0 42044 0 1 31008
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_604
timestamp 1586364061
transform 1 0 40388 0 1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__CLK
timestamp 1586364061
transform 1 0 41860 0 1 31008
box -38 -48 222 592
use scs8hd_decap_6  FILLER_52_434
timestamp 1586364061
transform 1 0 41032 0 -1 31008
box -38 -48 590 592
use scs8hd_fill_1  FILLER_52_440
timestamp 1586364061
transform 1 0 41584 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_53_428
timestamp 1586364061
transform 1 0 40480 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_53_440
timestamp 1586364061
transform 1 0 41584 0 1 31008
box -38 -48 314 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_9_
timestamp 1586364061
transform 1 0 43332 0 -1 31008
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_597
timestamp 1586364061
transform 1 0 43240 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_8  FILLER_52_450
timestamp 1586364061
transform 1 0 42504 0 -1 31008
box -38 -48 774 592
use scs8hd_decap_12  FILLER_53_464
timestamp 1586364061
transform 1 0 43792 0 1 31008
box -38 -48 1142 592
use scs8hd_dfxbp_1  ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_8_
timestamp 1586364061
transform 1 0 45816 0 -1 31008
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_605
timestamp 1586364061
transform 1 0 46000 0 1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__75__A
timestamp 1586364061
transform 1 0 46736 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_6__D
timestamp 1586364061
transform 1 0 45632 0 -1 31008
box -38 -48 222 592
use scs8hd_decap_6  FILLER_52_478
timestamp 1586364061
transform 1 0 45080 0 -1 31008
box -38 -48 590 592
use scs8hd_decap_12  FILLER_53_476
timestamp 1586364061
transform 1 0 44896 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_53_489
timestamp 1586364061
transform 1 0 46092 0 1 31008
box -38 -48 590 592
use scs8hd_fill_1  FILLER_53_495
timestamp 1586364061
transform 1 0 46644 0 1 31008
box -38 -48 130 592
use scs8hd_decap_3  PHY_105
timestamp 1586364061
transform -1 0 48852 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_107
timestamp 1586364061
transform -1 0 48852 0 1 31008
box -38 -48 314 592
use scs8hd_decap_8  FILLER_52_505
timestamp 1586364061
transform 1 0 47564 0 -1 31008
box -38 -48 774 592
use scs8hd_decap_3  FILLER_52_513
timestamp 1586364061
transform 1 0 48300 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_12  FILLER_53_498
timestamp 1586364061
transform 1 0 46920 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_53_510
timestamp 1586364061
transform 1 0 48024 0 1 31008
box -38 -48 590 592
use scs8hd_decap_3  PHY_108
timestamp 1586364061
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_54_3
timestamp 1586364061
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_15
timestamp 1586364061
transform 1 0 2484 0 -1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_606
timestamp 1586364061
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_4  FILLER_54_27
timestamp 1586364061
transform 1 0 3588 0 -1 32096
box -38 -48 406 592
use scs8hd_decap_12  FILLER_54_32
timestamp 1586364061
transform 1 0 4048 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_44
timestamp 1586364061
transform 1 0 5152 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_56
timestamp 1586364061
transform 1 0 6256 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_68
timestamp 1586364061
transform 1 0 7360 0 -1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_607
timestamp 1586364061
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_54_80
timestamp 1586364061
transform 1 0 8464 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_93
timestamp 1586364061
transform 1 0 9660 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_105
timestamp 1586364061
transform 1 0 10764 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_117
timestamp 1586364061
transform 1 0 11868 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_129
timestamp 1586364061
transform 1 0 12972 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_141
timestamp 1586364061
transform 1 0 14076 0 -1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_608
timestamp 1586364061
transform 1 0 15180 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_54_154
timestamp 1586364061
transform 1 0 15272 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_166
timestamp 1586364061
transform 1 0 16376 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_178
timestamp 1586364061
transform 1 0 17480 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_190
timestamp 1586364061
transform 1 0 18584 0 -1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_609
timestamp 1586364061
transform 1 0 20792 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_54_202
timestamp 1586364061
transform 1 0 19688 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_215
timestamp 1586364061
transform 1 0 20884 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_227
timestamp 1586364061
transform 1 0 21988 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_239
timestamp 1586364061
transform 1 0 23092 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_251
timestamp 1586364061
transform 1 0 24196 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_263
timestamp 1586364061
transform 1 0 25300 0 -1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_610
timestamp 1586364061
transform 1 0 26404 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_54_276
timestamp 1586364061
transform 1 0 26496 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_288
timestamp 1586364061
transform 1 0 27600 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_300
timestamp 1586364061
transform 1 0 28704 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_312
timestamp 1586364061
transform 1 0 29808 0 -1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_611
timestamp 1586364061
transform 1 0 32016 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_54_324
timestamp 1586364061
transform 1 0 30912 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_337
timestamp 1586364061
transform 1 0 32108 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_349
timestamp 1586364061
transform 1 0 33212 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_361
timestamp 1586364061
transform 1 0 34316 0 -1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_612
timestamp 1586364061
transform 1 0 37628 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_54_373
timestamp 1586364061
transform 1 0 35420 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_385
timestamp 1586364061
transform 1 0 36524 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_398
timestamp 1586364061
transform 1 0 37720 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_410
timestamp 1586364061
transform 1 0 38824 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_422
timestamp 1586364061
transform 1 0 39928 0 -1 32096
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_md_fle_mp_fab_md_flogic_md_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.scs8hd_dfxbp_1_10__D
timestamp 1586364061
transform 1 0 42044 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_8  FILLER_54_434
timestamp 1586364061
transform 1 0 41032 0 -1 32096
box -38 -48 774 592
use scs8hd_decap_3  FILLER_54_442
timestamp 1586364061
transform 1 0 41768 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_8  FILLER_54_447
timestamp 1586364061
transform 1 0 42228 0 -1 32096
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_613
timestamp 1586364061
transform 1 0 43240 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_3  FILLER_54_455
timestamp 1586364061
transform 1 0 42964 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_54_459
timestamp 1586364061
transform 1 0 43332 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_471
timestamp 1586364061
transform 1 0 44436 0 -1 32096
box -38 -48 1142 592
use scs8hd_buf_2  _75_
timestamp 1586364061
transform 1 0 46736 0 -1 32096
box -38 -48 406 592
use scs8hd_decap_12  FILLER_54_483
timestamp 1586364061
transform 1 0 45540 0 -1 32096
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_54_495
timestamp 1586364061
transform 1 0 46644 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_3  PHY_109
timestamp 1586364061
transform -1 0 48852 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_54_500
timestamp 1586364061
transform 1 0 47104 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_54_512
timestamp 1586364061
transform 1 0 48208 0 -1 32096
box -38 -48 406 592
use scs8hd_decap_3  PHY_110
timestamp 1586364061
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_55_3
timestamp 1586364061
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_15
timestamp 1586364061
transform 1 0 2484 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_27
timestamp 1586364061
transform 1 0 3588 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_39
timestamp 1586364061
transform 1 0 4692 0 1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_614
timestamp 1586364061
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use scs8hd_decap_8  FILLER_55_51
timestamp 1586364061
transform 1 0 5796 0 1 32096
box -38 -48 774 592
use scs8hd_fill_2  FILLER_55_59
timestamp 1586364061
transform 1 0 6532 0 1 32096
box -38 -48 222 592
use scs8hd_decap_12  FILLER_55_62
timestamp 1586364061
transform 1 0 6808 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_74
timestamp 1586364061
transform 1 0 7912 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_86
timestamp 1586364061
transform 1 0 9016 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_98
timestamp 1586364061
transform 1 0 10120 0 1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_615
timestamp 1586364061
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_55_110
timestamp 1586364061
transform 1 0 11224 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_123
timestamp 1586364061
transform 1 0 12420 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_135
timestamp 1586364061
transform 1 0 13524 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_147
timestamp 1586364061
transform 1 0 14628 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_159
timestamp 1586364061
transform 1 0 15732 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_171
timestamp 1586364061
transform 1 0 16836 0 1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_616
timestamp 1586364061
transform 1 0 17940 0 1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_55_184
timestamp 1586364061
transform 1 0 18032 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_196
timestamp 1586364061
transform 1 0 19136 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_208
timestamp 1586364061
transform 1 0 20240 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_220
timestamp 1586364061
transform 1 0 21344 0 1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_617
timestamp 1586364061
transform 1 0 23552 0 1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_55_232
timestamp 1586364061
transform 1 0 22448 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_245
timestamp 1586364061
transform 1 0 23644 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_257
timestamp 1586364061
transform 1 0 24748 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_269
timestamp 1586364061
transform 1 0 25852 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_281
timestamp 1586364061
transform 1 0 26956 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_293
timestamp 1586364061
transform 1 0 28060 0 1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_618
timestamp 1586364061
transform 1 0 29164 0 1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_55_306
timestamp 1586364061
transform 1 0 29256 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_318
timestamp 1586364061
transform 1 0 30360 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_330
timestamp 1586364061
transform 1 0 31464 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_342
timestamp 1586364061
transform 1 0 32568 0 1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_619
timestamp 1586364061
transform 1 0 34776 0 1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_55_354
timestamp 1586364061
transform 1 0 33672 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_367
timestamp 1586364061
transform 1 0 34868 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_379
timestamp 1586364061
transform 1 0 35972 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_391
timestamp 1586364061
transform 1 0 37076 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_403
timestamp 1586364061
transform 1 0 38180 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_415
timestamp 1586364061
transform 1 0 39284 0 1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_620
timestamp 1586364061
transform 1 0 40388 0 1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_55_428
timestamp 1586364061
transform 1 0 40480 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_440
timestamp 1586364061
transform 1 0 41584 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_452
timestamp 1586364061
transform 1 0 42688 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_464
timestamp 1586364061
transform 1 0 43792 0 1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_621
timestamp 1586364061
transform 1 0 46000 0 1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_55_476
timestamp 1586364061
transform 1 0 44896 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_489
timestamp 1586364061
transform 1 0 46092 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_3  PHY_111
timestamp 1586364061
transform -1 0 48852 0 1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_55_501
timestamp 1586364061
transform 1 0 47196 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_55_513
timestamp 1586364061
transform 1 0 48300 0 1 32096
box -38 -48 314 592
use scs8hd_decap_3  PHY_112
timestamp 1586364061
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_56_3
timestamp 1586364061
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_15
timestamp 1586364061
transform 1 0 2484 0 -1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_622
timestamp 1586364061
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_4  FILLER_56_27
timestamp 1586364061
transform 1 0 3588 0 -1 33184
box -38 -48 406 592
use scs8hd_decap_12  FILLER_56_32
timestamp 1586364061
transform 1 0 4048 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_44
timestamp 1586364061
transform 1 0 5152 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_56
timestamp 1586364061
transform 1 0 6256 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_68
timestamp 1586364061
transform 1 0 7360 0 -1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_623
timestamp 1586364061
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_56_80
timestamp 1586364061
transform 1 0 8464 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_93
timestamp 1586364061
transform 1 0 9660 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_105
timestamp 1586364061
transform 1 0 10764 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_117
timestamp 1586364061
transform 1 0 11868 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_129
timestamp 1586364061
transform 1 0 12972 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_141
timestamp 1586364061
transform 1 0 14076 0 -1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_624
timestamp 1586364061
transform 1 0 15180 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_56_154
timestamp 1586364061
transform 1 0 15272 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_166
timestamp 1586364061
transform 1 0 16376 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_178
timestamp 1586364061
transform 1 0 17480 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_190
timestamp 1586364061
transform 1 0 18584 0 -1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_625
timestamp 1586364061
transform 1 0 20792 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_56_202
timestamp 1586364061
transform 1 0 19688 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_215
timestamp 1586364061
transform 1 0 20884 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_227
timestamp 1586364061
transform 1 0 21988 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_239
timestamp 1586364061
transform 1 0 23092 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_251
timestamp 1586364061
transform 1 0 24196 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_263
timestamp 1586364061
transform 1 0 25300 0 -1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_626
timestamp 1586364061
transform 1 0 26404 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_56_276
timestamp 1586364061
transform 1 0 26496 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_288
timestamp 1586364061
transform 1 0 27600 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_300
timestamp 1586364061
transform 1 0 28704 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_312
timestamp 1586364061
transform 1 0 29808 0 -1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_627
timestamp 1586364061
transform 1 0 32016 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_56_324
timestamp 1586364061
transform 1 0 30912 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_337
timestamp 1586364061
transform 1 0 32108 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_349
timestamp 1586364061
transform 1 0 33212 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_361
timestamp 1586364061
transform 1 0 34316 0 -1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_628
timestamp 1586364061
transform 1 0 37628 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_56_373
timestamp 1586364061
transform 1 0 35420 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_385
timestamp 1586364061
transform 1 0 36524 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_398
timestamp 1586364061
transform 1 0 37720 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_410
timestamp 1586364061
transform 1 0 38824 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_422
timestamp 1586364061
transform 1 0 39928 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_434
timestamp 1586364061
transform 1 0 41032 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_446
timestamp 1586364061
transform 1 0 42136 0 -1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_629
timestamp 1586364061
transform 1 0 43240 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_56_459
timestamp 1586364061
transform 1 0 43332 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_471
timestamp 1586364061
transform 1 0 44436 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_483
timestamp 1586364061
transform 1 0 45540 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_495
timestamp 1586364061
transform 1 0 46644 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_3  PHY_113
timestamp 1586364061
transform -1 0 48852 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_8  FILLER_56_507
timestamp 1586364061
transform 1 0 47748 0 -1 33184
box -38 -48 774 592
use scs8hd_fill_1  FILLER_56_515
timestamp 1586364061
transform 1 0 48484 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_3  PHY_114
timestamp 1586364061
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_57_3
timestamp 1586364061
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_15
timestamp 1586364061
transform 1 0 2484 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_27
timestamp 1586364061
transform 1 0 3588 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_39
timestamp 1586364061
transform 1 0 4692 0 1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_630
timestamp 1586364061
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use scs8hd_decap_8  FILLER_57_51
timestamp 1586364061
transform 1 0 5796 0 1 33184
box -38 -48 774 592
use scs8hd_fill_2  FILLER_57_59
timestamp 1586364061
transform 1 0 6532 0 1 33184
box -38 -48 222 592
use scs8hd_decap_12  FILLER_57_62
timestamp 1586364061
transform 1 0 6808 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_74
timestamp 1586364061
transform 1 0 7912 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_86
timestamp 1586364061
transform 1 0 9016 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_98
timestamp 1586364061
transform 1 0 10120 0 1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_631
timestamp 1586364061
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_57_110
timestamp 1586364061
transform 1 0 11224 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_123
timestamp 1586364061
transform 1 0 12420 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_135
timestamp 1586364061
transform 1 0 13524 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_147
timestamp 1586364061
transform 1 0 14628 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_159
timestamp 1586364061
transform 1 0 15732 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_171
timestamp 1586364061
transform 1 0 16836 0 1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_632
timestamp 1586364061
transform 1 0 17940 0 1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_57_184
timestamp 1586364061
transform 1 0 18032 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_196
timestamp 1586364061
transform 1 0 19136 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_208
timestamp 1586364061
transform 1 0 20240 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_220
timestamp 1586364061
transform 1 0 21344 0 1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_633
timestamp 1586364061
transform 1 0 23552 0 1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_57_232
timestamp 1586364061
transform 1 0 22448 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_245
timestamp 1586364061
transform 1 0 23644 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_257
timestamp 1586364061
transform 1 0 24748 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_269
timestamp 1586364061
transform 1 0 25852 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_281
timestamp 1586364061
transform 1 0 26956 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_293
timestamp 1586364061
transform 1 0 28060 0 1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_634
timestamp 1586364061
transform 1 0 29164 0 1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_57_306
timestamp 1586364061
transform 1 0 29256 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_318
timestamp 1586364061
transform 1 0 30360 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_330
timestamp 1586364061
transform 1 0 31464 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_342
timestamp 1586364061
transform 1 0 32568 0 1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_635
timestamp 1586364061
transform 1 0 34776 0 1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_57_354
timestamp 1586364061
transform 1 0 33672 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_367
timestamp 1586364061
transform 1 0 34868 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_379
timestamp 1586364061
transform 1 0 35972 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_391
timestamp 1586364061
transform 1 0 37076 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_403
timestamp 1586364061
transform 1 0 38180 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_415
timestamp 1586364061
transform 1 0 39284 0 1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_636
timestamp 1586364061
transform 1 0 40388 0 1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_57_428
timestamp 1586364061
transform 1 0 40480 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_440
timestamp 1586364061
transform 1 0 41584 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_452
timestamp 1586364061
transform 1 0 42688 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_464
timestamp 1586364061
transform 1 0 43792 0 1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_637
timestamp 1586364061
transform 1 0 46000 0 1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_57_476
timestamp 1586364061
transform 1 0 44896 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_489
timestamp 1586364061
transform 1 0 46092 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_3  PHY_115
timestamp 1586364061
transform -1 0 48852 0 1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_57_501
timestamp 1586364061
transform 1 0 47196 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_57_513
timestamp 1586364061
transform 1 0 48300 0 1 33184
box -38 -48 314 592
use scs8hd_decap_3  PHY_116
timestamp 1586364061
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_12  FILLER_58_3
timestamp 1586364061
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_15
timestamp 1586364061
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_638
timestamp 1586364061
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_4  FILLER_58_27
timestamp 1586364061
transform 1 0 3588 0 -1 34272
box -38 -48 406 592
use scs8hd_decap_12  FILLER_58_32
timestamp 1586364061
transform 1 0 4048 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_44
timestamp 1586364061
transform 1 0 5152 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_56
timestamp 1586364061
transform 1 0 6256 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_68
timestamp 1586364061
transform 1 0 7360 0 -1 34272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_639
timestamp 1586364061
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_58_80
timestamp 1586364061
transform 1 0 8464 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_93
timestamp 1586364061
transform 1 0 9660 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_105
timestamp 1586364061
transform 1 0 10764 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_117
timestamp 1586364061
transform 1 0 11868 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_129
timestamp 1586364061
transform 1 0 12972 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_141
timestamp 1586364061
transform 1 0 14076 0 -1 34272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_640
timestamp 1586364061
transform 1 0 15180 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_58_154
timestamp 1586364061
transform 1 0 15272 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_166
timestamp 1586364061
transform 1 0 16376 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_178
timestamp 1586364061
transform 1 0 17480 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_190
timestamp 1586364061
transform 1 0 18584 0 -1 34272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_641
timestamp 1586364061
transform 1 0 20792 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_58_202
timestamp 1586364061
transform 1 0 19688 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_215
timestamp 1586364061
transform 1 0 20884 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_227
timestamp 1586364061
transform 1 0 21988 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_239
timestamp 1586364061
transform 1 0 23092 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_251
timestamp 1586364061
transform 1 0 24196 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_263
timestamp 1586364061
transform 1 0 25300 0 -1 34272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_642
timestamp 1586364061
transform 1 0 26404 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_58_276
timestamp 1586364061
transform 1 0 26496 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_288
timestamp 1586364061
transform 1 0 27600 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_300
timestamp 1586364061
transform 1 0 28704 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_312
timestamp 1586364061
transform 1 0 29808 0 -1 34272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_643
timestamp 1586364061
transform 1 0 32016 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_58_324
timestamp 1586364061
transform 1 0 30912 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_337
timestamp 1586364061
transform 1 0 32108 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_349
timestamp 1586364061
transform 1 0 33212 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_361
timestamp 1586364061
transform 1 0 34316 0 -1 34272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_644
timestamp 1586364061
transform 1 0 37628 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_58_373
timestamp 1586364061
transform 1 0 35420 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_385
timestamp 1586364061
transform 1 0 36524 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_398
timestamp 1586364061
transform 1 0 37720 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_410
timestamp 1586364061
transform 1 0 38824 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_422
timestamp 1586364061
transform 1 0 39928 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_434
timestamp 1586364061
transform 1 0 41032 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_446
timestamp 1586364061
transform 1 0 42136 0 -1 34272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_645
timestamp 1586364061
transform 1 0 43240 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_58_459
timestamp 1586364061
transform 1 0 43332 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_471
timestamp 1586364061
transform 1 0 44436 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_483
timestamp 1586364061
transform 1 0 45540 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_495
timestamp 1586364061
transform 1 0 46644 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_3  PHY_117
timestamp 1586364061
transform -1 0 48852 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_8  FILLER_58_507
timestamp 1586364061
transform 1 0 47748 0 -1 34272
box -38 -48 774 592
use scs8hd_fill_1  FILLER_58_515
timestamp 1586364061
transform 1 0 48484 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_3  PHY_118
timestamp 1586364061
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_120
timestamp 1586364061
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_59_3
timestamp 1586364061
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_15
timestamp 1586364061
transform 1 0 2484 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_3
timestamp 1586364061
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_15
timestamp 1586364061
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_654
timestamp 1586364061
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_27
timestamp 1586364061
transform 1 0 3588 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_39
timestamp 1586364061
transform 1 0 4692 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_60_27
timestamp 1586364061
transform 1 0 3588 0 -1 35360
box -38 -48 406 592
use scs8hd_decap_12  FILLER_60_32
timestamp 1586364061
transform 1 0 4048 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_44
timestamp 1586364061
transform 1 0 5152 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_646
timestamp 1586364061
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use scs8hd_decap_8  FILLER_59_51
timestamp 1586364061
transform 1 0 5796 0 1 34272
box -38 -48 774 592
use scs8hd_fill_2  FILLER_59_59
timestamp 1586364061
transform 1 0 6532 0 1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_59_62
timestamp 1586364061
transform 1 0 6808 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_74
timestamp 1586364061
transform 1 0 7912 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_56
timestamp 1586364061
transform 1 0 6256 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_68
timestamp 1586364061
transform 1 0 7360 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_655
timestamp 1586364061
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_86
timestamp 1586364061
transform 1 0 9016 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_98
timestamp 1586364061
transform 1 0 10120 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_80
timestamp 1586364061
transform 1 0 8464 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_93
timestamp 1586364061
transform 1 0 9660 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_647
timestamp 1586364061
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_110
timestamp 1586364061
transform 1 0 11224 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_123
timestamp 1586364061
transform 1 0 12420 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_105
timestamp 1586364061
transform 1 0 10764 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_117
timestamp 1586364061
transform 1 0 11868 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_135
timestamp 1586364061
transform 1 0 13524 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_147
timestamp 1586364061
transform 1 0 14628 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_129
timestamp 1586364061
transform 1 0 12972 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_141
timestamp 1586364061
transform 1 0 14076 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_656
timestamp 1586364061
transform 1 0 15180 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_159
timestamp 1586364061
transform 1 0 15732 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_171
timestamp 1586364061
transform 1 0 16836 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_154
timestamp 1586364061
transform 1 0 15272 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_166
timestamp 1586364061
transform 1 0 16376 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_648
timestamp 1586364061
transform 1 0 17940 0 1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_184
timestamp 1586364061
transform 1 0 18032 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_196
timestamp 1586364061
transform 1 0 19136 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_178
timestamp 1586364061
transform 1 0 17480 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_190
timestamp 1586364061
transform 1 0 18584 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_657
timestamp 1586364061
transform 1 0 20792 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_208
timestamp 1586364061
transform 1 0 20240 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_220
timestamp 1586364061
transform 1 0 21344 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_202
timestamp 1586364061
transform 1 0 19688 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_215
timestamp 1586364061
transform 1 0 20884 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_649
timestamp 1586364061
transform 1 0 23552 0 1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_232
timestamp 1586364061
transform 1 0 22448 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_245
timestamp 1586364061
transform 1 0 23644 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_227
timestamp 1586364061
transform 1 0 21988 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_239
timestamp 1586364061
transform 1 0 23092 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_257
timestamp 1586364061
transform 1 0 24748 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_269
timestamp 1586364061
transform 1 0 25852 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_251
timestamp 1586364061
transform 1 0 24196 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_263
timestamp 1586364061
transform 1 0 25300 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_658
timestamp 1586364061
transform 1 0 26404 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_281
timestamp 1586364061
transform 1 0 26956 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_293
timestamp 1586364061
transform 1 0 28060 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_276
timestamp 1586364061
transform 1 0 26496 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_288
timestamp 1586364061
transform 1 0 27600 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_650
timestamp 1586364061
transform 1 0 29164 0 1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_306
timestamp 1586364061
transform 1 0 29256 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_318
timestamp 1586364061
transform 1 0 30360 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_300
timestamp 1586364061
transform 1 0 28704 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_312
timestamp 1586364061
transform 1 0 29808 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_659
timestamp 1586364061
transform 1 0 32016 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_330
timestamp 1586364061
transform 1 0 31464 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_342
timestamp 1586364061
transform 1 0 32568 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_324
timestamp 1586364061
transform 1 0 30912 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_337
timestamp 1586364061
transform 1 0 32108 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_651
timestamp 1586364061
transform 1 0 34776 0 1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_354
timestamp 1586364061
transform 1 0 33672 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_367
timestamp 1586364061
transform 1 0 34868 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_349
timestamp 1586364061
transform 1 0 33212 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_361
timestamp 1586364061
transform 1 0 34316 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_660
timestamp 1586364061
transform 1 0 37628 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_379
timestamp 1586364061
transform 1 0 35972 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_391
timestamp 1586364061
transform 1 0 37076 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_373
timestamp 1586364061
transform 1 0 35420 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_385
timestamp 1586364061
transform 1 0 36524 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_403
timestamp 1586364061
transform 1 0 38180 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_415
timestamp 1586364061
transform 1 0 39284 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_398
timestamp 1586364061
transform 1 0 37720 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_410
timestamp 1586364061
transform 1 0 38824 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_422
timestamp 1586364061
transform 1 0 39928 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_652
timestamp 1586364061
transform 1 0 40388 0 1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_428
timestamp 1586364061
transform 1 0 40480 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_440
timestamp 1586364061
transform 1 0 41584 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_434
timestamp 1586364061
transform 1 0 41032 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_446
timestamp 1586364061
transform 1 0 42136 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_661
timestamp 1586364061
transform 1 0 43240 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_452
timestamp 1586364061
transform 1 0 42688 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_464
timestamp 1586364061
transform 1 0 43792 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_459
timestamp 1586364061
transform 1 0 43332 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_471
timestamp 1586364061
transform 1 0 44436 0 -1 35360
box -38 -48 1142 592
use scs8hd_buf_2  _76_
timestamp 1586364061
transform 1 0 46736 0 -1 35360
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_653
timestamp 1586364061
transform 1 0 46000 0 1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__76__A
timestamp 1586364061
transform 1 0 46736 0 1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_59_476
timestamp 1586364061
transform 1 0 44896 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_59_489
timestamp 1586364061
transform 1 0 46092 0 1 34272
box -38 -48 590 592
use scs8hd_fill_1  FILLER_59_495
timestamp 1586364061
transform 1 0 46644 0 1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_60_483
timestamp 1586364061
transform 1 0 45540 0 -1 35360
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_60_495
timestamp 1586364061
transform 1 0 46644 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_3  PHY_119
timestamp 1586364061
transform -1 0 48852 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_121
timestamp 1586364061
transform -1 0 48852 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_59_498
timestamp 1586364061
transform 1 0 46920 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_59_510
timestamp 1586364061
transform 1 0 48024 0 1 34272
box -38 -48 590 592
use scs8hd_decap_12  FILLER_60_500
timestamp 1586364061
transform 1 0 47104 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_60_512
timestamp 1586364061
transform 1 0 48208 0 -1 35360
box -38 -48 406 592
use scs8hd_decap_3  PHY_122
timestamp 1586364061
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_61_3
timestamp 1586364061
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_15
timestamp 1586364061
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_27
timestamp 1586364061
transform 1 0 3588 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_39
timestamp 1586364061
transform 1 0 4692 0 1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_662
timestamp 1586364061
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use scs8hd_decap_8  FILLER_61_51
timestamp 1586364061
transform 1 0 5796 0 1 35360
box -38 -48 774 592
use scs8hd_fill_2  FILLER_61_59
timestamp 1586364061
transform 1 0 6532 0 1 35360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_61_62
timestamp 1586364061
transform 1 0 6808 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_74
timestamp 1586364061
transform 1 0 7912 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_86
timestamp 1586364061
transform 1 0 9016 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_98
timestamp 1586364061
transform 1 0 10120 0 1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_663
timestamp 1586364061
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_61_110
timestamp 1586364061
transform 1 0 11224 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_123
timestamp 1586364061
transform 1 0 12420 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_135
timestamp 1586364061
transform 1 0 13524 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_147
timestamp 1586364061
transform 1 0 14628 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_159
timestamp 1586364061
transform 1 0 15732 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_171
timestamp 1586364061
transform 1 0 16836 0 1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_664
timestamp 1586364061
transform 1 0 17940 0 1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_61_184
timestamp 1586364061
transform 1 0 18032 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_196
timestamp 1586364061
transform 1 0 19136 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_208
timestamp 1586364061
transform 1 0 20240 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_220
timestamp 1586364061
transform 1 0 21344 0 1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_665
timestamp 1586364061
transform 1 0 23552 0 1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_61_232
timestamp 1586364061
transform 1 0 22448 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_245
timestamp 1586364061
transform 1 0 23644 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_257
timestamp 1586364061
transform 1 0 24748 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_269
timestamp 1586364061
transform 1 0 25852 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_281
timestamp 1586364061
transform 1 0 26956 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_293
timestamp 1586364061
transform 1 0 28060 0 1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_666
timestamp 1586364061
transform 1 0 29164 0 1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_61_306
timestamp 1586364061
transform 1 0 29256 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_318
timestamp 1586364061
transform 1 0 30360 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_330
timestamp 1586364061
transform 1 0 31464 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_342
timestamp 1586364061
transform 1 0 32568 0 1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_667
timestamp 1586364061
transform 1 0 34776 0 1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_61_354
timestamp 1586364061
transform 1 0 33672 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_367
timestamp 1586364061
transform 1 0 34868 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_379
timestamp 1586364061
transform 1 0 35972 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_391
timestamp 1586364061
transform 1 0 37076 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_403
timestamp 1586364061
transform 1 0 38180 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_415
timestamp 1586364061
transform 1 0 39284 0 1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_668
timestamp 1586364061
transform 1 0 40388 0 1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_61_428
timestamp 1586364061
transform 1 0 40480 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_440
timestamp 1586364061
transform 1 0 41584 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_452
timestamp 1586364061
transform 1 0 42688 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_464
timestamp 1586364061
transform 1 0 43792 0 1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_669
timestamp 1586364061
transform 1 0 46000 0 1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_61_476
timestamp 1586364061
transform 1 0 44896 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_489
timestamp 1586364061
transform 1 0 46092 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_3  PHY_123
timestamp 1586364061
transform -1 0 48852 0 1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_61_501
timestamp 1586364061
transform 1 0 47196 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_61_513
timestamp 1586364061
transform 1 0 48300 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  PHY_124
timestamp 1586364061
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_62_3
timestamp 1586364061
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_15
timestamp 1586364061
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_670
timestamp 1586364061
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_4  FILLER_62_27
timestamp 1586364061
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use scs8hd_decap_12  FILLER_62_32
timestamp 1586364061
transform 1 0 4048 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_44
timestamp 1586364061
transform 1 0 5152 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_56
timestamp 1586364061
transform 1 0 6256 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_68
timestamp 1586364061
transform 1 0 7360 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_671
timestamp 1586364061
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_80
timestamp 1586364061
transform 1 0 8464 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_93
timestamp 1586364061
transform 1 0 9660 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_105
timestamp 1586364061
transform 1 0 10764 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_117
timestamp 1586364061
transform 1 0 11868 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_129
timestamp 1586364061
transform 1 0 12972 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_141
timestamp 1586364061
transform 1 0 14076 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_672
timestamp 1586364061
transform 1 0 15180 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_154
timestamp 1586364061
transform 1 0 15272 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_166
timestamp 1586364061
transform 1 0 16376 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_178
timestamp 1586364061
transform 1 0 17480 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_190
timestamp 1586364061
transform 1 0 18584 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_673
timestamp 1586364061
transform 1 0 20792 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_202
timestamp 1586364061
transform 1 0 19688 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_215
timestamp 1586364061
transform 1 0 20884 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_227
timestamp 1586364061
transform 1 0 21988 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_239
timestamp 1586364061
transform 1 0 23092 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_251
timestamp 1586364061
transform 1 0 24196 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_263
timestamp 1586364061
transform 1 0 25300 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_674
timestamp 1586364061
transform 1 0 26404 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_276
timestamp 1586364061
transform 1 0 26496 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_288
timestamp 1586364061
transform 1 0 27600 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_300
timestamp 1586364061
transform 1 0 28704 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_312
timestamp 1586364061
transform 1 0 29808 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_675
timestamp 1586364061
transform 1 0 32016 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_324
timestamp 1586364061
transform 1 0 30912 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_337
timestamp 1586364061
transform 1 0 32108 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_349
timestamp 1586364061
transform 1 0 33212 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_361
timestamp 1586364061
transform 1 0 34316 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_676
timestamp 1586364061
transform 1 0 37628 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_373
timestamp 1586364061
transform 1 0 35420 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_385
timestamp 1586364061
transform 1 0 36524 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_398
timestamp 1586364061
transform 1 0 37720 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_410
timestamp 1586364061
transform 1 0 38824 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_422
timestamp 1586364061
transform 1 0 39928 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_434
timestamp 1586364061
transform 1 0 41032 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_446
timestamp 1586364061
transform 1 0 42136 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_677
timestamp 1586364061
transform 1 0 43240 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_459
timestamp 1586364061
transform 1 0 43332 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_471
timestamp 1586364061
transform 1 0 44436 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_483
timestamp 1586364061
transform 1 0 45540 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_495
timestamp 1586364061
transform 1 0 46644 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_3  PHY_125
timestamp 1586364061
transform -1 0 48852 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_8  FILLER_62_507
timestamp 1586364061
transform 1 0 47748 0 -1 36448
box -38 -48 774 592
use scs8hd_fill_1  FILLER_62_515
timestamp 1586364061
transform 1 0 48484 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_3  PHY_126
timestamp 1586364061
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_63_3
timestamp 1586364061
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_15
timestamp 1586364061
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_27
timestamp 1586364061
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_39
timestamp 1586364061
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_678
timestamp 1586364061
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use scs8hd_decap_8  FILLER_63_51
timestamp 1586364061
transform 1 0 5796 0 1 36448
box -38 -48 774 592
use scs8hd_fill_2  FILLER_63_59
timestamp 1586364061
transform 1 0 6532 0 1 36448
box -38 -48 222 592
use scs8hd_decap_12  FILLER_63_62
timestamp 1586364061
transform 1 0 6808 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_74
timestamp 1586364061
transform 1 0 7912 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_86
timestamp 1586364061
transform 1 0 9016 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_98
timestamp 1586364061
transform 1 0 10120 0 1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_679
timestamp 1586364061
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_63_110
timestamp 1586364061
transform 1 0 11224 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_123
timestamp 1586364061
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_135
timestamp 1586364061
transform 1 0 13524 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_147
timestamp 1586364061
transform 1 0 14628 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_159
timestamp 1586364061
transform 1 0 15732 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_171
timestamp 1586364061
transform 1 0 16836 0 1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_680
timestamp 1586364061
transform 1 0 17940 0 1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_63_184
timestamp 1586364061
transform 1 0 18032 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_196
timestamp 1586364061
transform 1 0 19136 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_208
timestamp 1586364061
transform 1 0 20240 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_220
timestamp 1586364061
transform 1 0 21344 0 1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_681
timestamp 1586364061
transform 1 0 23552 0 1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_63_232
timestamp 1586364061
transform 1 0 22448 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_245
timestamp 1586364061
transform 1 0 23644 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_257
timestamp 1586364061
transform 1 0 24748 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_269
timestamp 1586364061
transform 1 0 25852 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_281
timestamp 1586364061
transform 1 0 26956 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_293
timestamp 1586364061
transform 1 0 28060 0 1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_682
timestamp 1586364061
transform 1 0 29164 0 1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_63_306
timestamp 1586364061
transform 1 0 29256 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_318
timestamp 1586364061
transform 1 0 30360 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_330
timestamp 1586364061
transform 1 0 31464 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_342
timestamp 1586364061
transform 1 0 32568 0 1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_683
timestamp 1586364061
transform 1 0 34776 0 1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_63_354
timestamp 1586364061
transform 1 0 33672 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_367
timestamp 1586364061
transform 1 0 34868 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_379
timestamp 1586364061
transform 1 0 35972 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_391
timestamp 1586364061
transform 1 0 37076 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_403
timestamp 1586364061
transform 1 0 38180 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_415
timestamp 1586364061
transform 1 0 39284 0 1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_684
timestamp 1586364061
transform 1 0 40388 0 1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_63_428
timestamp 1586364061
transform 1 0 40480 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_440
timestamp 1586364061
transform 1 0 41584 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_452
timestamp 1586364061
transform 1 0 42688 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_464
timestamp 1586364061
transform 1 0 43792 0 1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_685
timestamp 1586364061
transform 1 0 46000 0 1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_63_476
timestamp 1586364061
transform 1 0 44896 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_489
timestamp 1586364061
transform 1 0 46092 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_3  PHY_127
timestamp 1586364061
transform -1 0 48852 0 1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_63_501
timestamp 1586364061
transform 1 0 47196 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_63_513
timestamp 1586364061
transform 1 0 48300 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  PHY_128
timestamp 1586364061
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_64_3
timestamp 1586364061
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_15
timestamp 1586364061
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_686
timestamp 1586364061
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_4  FILLER_64_27
timestamp 1586364061
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use scs8hd_decap_12  FILLER_64_32
timestamp 1586364061
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_44
timestamp 1586364061
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_56
timestamp 1586364061
transform 1 0 6256 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_68
timestamp 1586364061
transform 1 0 7360 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_687
timestamp 1586364061
transform 1 0 9568 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_80
timestamp 1586364061
transform 1 0 8464 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_93
timestamp 1586364061
transform 1 0 9660 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_105
timestamp 1586364061
transform 1 0 10764 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_117
timestamp 1586364061
transform 1 0 11868 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_129
timestamp 1586364061
transform 1 0 12972 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_141
timestamp 1586364061
transform 1 0 14076 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_688
timestamp 1586364061
transform 1 0 15180 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_154
timestamp 1586364061
transform 1 0 15272 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_166
timestamp 1586364061
transform 1 0 16376 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_178
timestamp 1586364061
transform 1 0 17480 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_190
timestamp 1586364061
transform 1 0 18584 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_689
timestamp 1586364061
transform 1 0 20792 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_202
timestamp 1586364061
transform 1 0 19688 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_215
timestamp 1586364061
transform 1 0 20884 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_227
timestamp 1586364061
transform 1 0 21988 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_239
timestamp 1586364061
transform 1 0 23092 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_251
timestamp 1586364061
transform 1 0 24196 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_263
timestamp 1586364061
transform 1 0 25300 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_690
timestamp 1586364061
transform 1 0 26404 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_276
timestamp 1586364061
transform 1 0 26496 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_288
timestamp 1586364061
transform 1 0 27600 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_300
timestamp 1586364061
transform 1 0 28704 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_312
timestamp 1586364061
transform 1 0 29808 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_691
timestamp 1586364061
transform 1 0 32016 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_324
timestamp 1586364061
transform 1 0 30912 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_337
timestamp 1586364061
transform 1 0 32108 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_349
timestamp 1586364061
transform 1 0 33212 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_361
timestamp 1586364061
transform 1 0 34316 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_692
timestamp 1586364061
transform 1 0 37628 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_373
timestamp 1586364061
transform 1 0 35420 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_385
timestamp 1586364061
transform 1 0 36524 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_398
timestamp 1586364061
transform 1 0 37720 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_410
timestamp 1586364061
transform 1 0 38824 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_422
timestamp 1586364061
transform 1 0 39928 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_434
timestamp 1586364061
transform 1 0 41032 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_446
timestamp 1586364061
transform 1 0 42136 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_693
timestamp 1586364061
transform 1 0 43240 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_459
timestamp 1586364061
transform 1 0 43332 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_471
timestamp 1586364061
transform 1 0 44436 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_483
timestamp 1586364061
transform 1 0 45540 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_495
timestamp 1586364061
transform 1 0 46644 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_3  PHY_129
timestamp 1586364061
transform -1 0 48852 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_8  FILLER_64_507
timestamp 1586364061
transform 1 0 47748 0 -1 37536
box -38 -48 774 592
use scs8hd_fill_1  FILLER_64_515
timestamp 1586364061
transform 1 0 48484 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_3  PHY_130
timestamp 1586364061
transform 1 0 1104 0 1 37536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_65_3
timestamp 1586364061
transform 1 0 1380 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_15
timestamp 1586364061
transform 1 0 2484 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_27
timestamp 1586364061
transform 1 0 3588 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_39
timestamp 1586364061
transform 1 0 4692 0 1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_694
timestamp 1586364061
transform 1 0 6716 0 1 37536
box -38 -48 130 592
use scs8hd_decap_8  FILLER_65_51
timestamp 1586364061
transform 1 0 5796 0 1 37536
box -38 -48 774 592
use scs8hd_fill_2  FILLER_65_59
timestamp 1586364061
transform 1 0 6532 0 1 37536
box -38 -48 222 592
use scs8hd_decap_12  FILLER_65_62
timestamp 1586364061
transform 1 0 6808 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_74
timestamp 1586364061
transform 1 0 7912 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_86
timestamp 1586364061
transform 1 0 9016 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_98
timestamp 1586364061
transform 1 0 10120 0 1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_695
timestamp 1586364061
transform 1 0 12328 0 1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_65_110
timestamp 1586364061
transform 1 0 11224 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_123
timestamp 1586364061
transform 1 0 12420 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_135
timestamp 1586364061
transform 1 0 13524 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_147
timestamp 1586364061
transform 1 0 14628 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_159
timestamp 1586364061
transform 1 0 15732 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_171
timestamp 1586364061
transform 1 0 16836 0 1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_696
timestamp 1586364061
transform 1 0 17940 0 1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_65_184
timestamp 1586364061
transform 1 0 18032 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_196
timestamp 1586364061
transform 1 0 19136 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_208
timestamp 1586364061
transform 1 0 20240 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_220
timestamp 1586364061
transform 1 0 21344 0 1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_697
timestamp 1586364061
transform 1 0 23552 0 1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_65_232
timestamp 1586364061
transform 1 0 22448 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_245
timestamp 1586364061
transform 1 0 23644 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_257
timestamp 1586364061
transform 1 0 24748 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_269
timestamp 1586364061
transform 1 0 25852 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_281
timestamp 1586364061
transform 1 0 26956 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_293
timestamp 1586364061
transform 1 0 28060 0 1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_698
timestamp 1586364061
transform 1 0 29164 0 1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_65_306
timestamp 1586364061
transform 1 0 29256 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_318
timestamp 1586364061
transform 1 0 30360 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_330
timestamp 1586364061
transform 1 0 31464 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_342
timestamp 1586364061
transform 1 0 32568 0 1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_699
timestamp 1586364061
transform 1 0 34776 0 1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_65_354
timestamp 1586364061
transform 1 0 33672 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_367
timestamp 1586364061
transform 1 0 34868 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_379
timestamp 1586364061
transform 1 0 35972 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_391
timestamp 1586364061
transform 1 0 37076 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_403
timestamp 1586364061
transform 1 0 38180 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_415
timestamp 1586364061
transform 1 0 39284 0 1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_700
timestamp 1586364061
transform 1 0 40388 0 1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_65_428
timestamp 1586364061
transform 1 0 40480 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_440
timestamp 1586364061
transform 1 0 41584 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_452
timestamp 1586364061
transform 1 0 42688 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_464
timestamp 1586364061
transform 1 0 43792 0 1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_701
timestamp 1586364061
transform 1 0 46000 0 1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__77__A
timestamp 1586364061
transform 1 0 46736 0 1 37536
box -38 -48 222 592
use scs8hd_decap_12  FILLER_65_476
timestamp 1586364061
transform 1 0 44896 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_65_489
timestamp 1586364061
transform 1 0 46092 0 1 37536
box -38 -48 590 592
use scs8hd_fill_1  FILLER_65_495
timestamp 1586364061
transform 1 0 46644 0 1 37536
box -38 -48 130 592
use scs8hd_decap_3  PHY_131
timestamp 1586364061
transform -1 0 48852 0 1 37536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_65_498
timestamp 1586364061
transform 1 0 46920 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_65_510
timestamp 1586364061
transform 1 0 48024 0 1 37536
box -38 -48 590 592
use scs8hd_decap_3  PHY_132
timestamp 1586364061
transform 1 0 1104 0 -1 38624
box -38 -48 314 592
use scs8hd_decap_3  PHY_134
timestamp 1586364061
transform 1 0 1104 0 1 38624
box -38 -48 314 592
use scs8hd_decap_12  FILLER_66_3
timestamp 1586364061
transform 1 0 1380 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_15
timestamp 1586364061
transform 1 0 2484 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_3
timestamp 1586364061
transform 1 0 1380 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_15
timestamp 1586364061
transform 1 0 2484 0 1 38624
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_702
timestamp 1586364061
transform 1 0 3956 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_4  FILLER_66_27
timestamp 1586364061
transform 1 0 3588 0 -1 38624
box -38 -48 406 592
use scs8hd_decap_12  FILLER_66_32
timestamp 1586364061
transform 1 0 4048 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_44
timestamp 1586364061
transform 1 0 5152 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_27
timestamp 1586364061
transform 1 0 3588 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_39
timestamp 1586364061
transform 1 0 4692 0 1 38624
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_710
timestamp 1586364061
transform 1 0 6716 0 1 38624
box -38 -48 130 592
use scs8hd_decap_12  FILLER_66_56
timestamp 1586364061
transform 1 0 6256 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_68
timestamp 1586364061
transform 1 0 7360 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_67_51
timestamp 1586364061
transform 1 0 5796 0 1 38624
box -38 -48 774 592
use scs8hd_fill_2  FILLER_67_59
timestamp 1586364061
transform 1 0 6532 0 1 38624
box -38 -48 222 592
use scs8hd_decap_12  FILLER_67_62
timestamp 1586364061
transform 1 0 6808 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_74
timestamp 1586364061
transform 1 0 7912 0 1 38624
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_703
timestamp 1586364061
transform 1 0 9568 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_12  FILLER_66_80
timestamp 1586364061
transform 1 0 8464 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_93
timestamp 1586364061
transform 1 0 9660 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_86
timestamp 1586364061
transform 1 0 9016 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_98
timestamp 1586364061
transform 1 0 10120 0 1 38624
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_711
timestamp 1586364061
transform 1 0 12328 0 1 38624
box -38 -48 130 592
use scs8hd_decap_12  FILLER_66_105
timestamp 1586364061
transform 1 0 10764 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_117
timestamp 1586364061
transform 1 0 11868 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_110
timestamp 1586364061
transform 1 0 11224 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_123
timestamp 1586364061
transform 1 0 12420 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_129
timestamp 1586364061
transform 1 0 12972 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_141
timestamp 1586364061
transform 1 0 14076 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_135
timestamp 1586364061
transform 1 0 13524 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_147
timestamp 1586364061
transform 1 0 14628 0 1 38624
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_704
timestamp 1586364061
transform 1 0 15180 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_12  FILLER_66_154
timestamp 1586364061
transform 1 0 15272 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_166
timestamp 1586364061
transform 1 0 16376 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_159
timestamp 1586364061
transform 1 0 15732 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_171
timestamp 1586364061
transform 1 0 16836 0 1 38624
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_712
timestamp 1586364061
transform 1 0 17940 0 1 38624
box -38 -48 130 592
use scs8hd_decap_12  FILLER_66_178
timestamp 1586364061
transform 1 0 17480 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_190
timestamp 1586364061
transform 1 0 18584 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_184
timestamp 1586364061
transform 1 0 18032 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_196
timestamp 1586364061
transform 1 0 19136 0 1 38624
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_705
timestamp 1586364061
transform 1 0 20792 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_12  FILLER_66_202
timestamp 1586364061
transform 1 0 19688 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_215
timestamp 1586364061
transform 1 0 20884 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_208
timestamp 1586364061
transform 1 0 20240 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_220
timestamp 1586364061
transform 1 0 21344 0 1 38624
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_713
timestamp 1586364061
transform 1 0 23552 0 1 38624
box -38 -48 130 592
use scs8hd_decap_12  FILLER_66_227
timestamp 1586364061
transform 1 0 21988 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_239
timestamp 1586364061
transform 1 0 23092 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_232
timestamp 1586364061
transform 1 0 22448 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_245
timestamp 1586364061
transform 1 0 23644 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_251
timestamp 1586364061
transform 1 0 24196 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_263
timestamp 1586364061
transform 1 0 25300 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_257
timestamp 1586364061
transform 1 0 24748 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_269
timestamp 1586364061
transform 1 0 25852 0 1 38624
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_706
timestamp 1586364061
transform 1 0 26404 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_12  FILLER_66_276
timestamp 1586364061
transform 1 0 26496 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_288
timestamp 1586364061
transform 1 0 27600 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_281
timestamp 1586364061
transform 1 0 26956 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_293
timestamp 1586364061
transform 1 0 28060 0 1 38624
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_714
timestamp 1586364061
transform 1 0 29164 0 1 38624
box -38 -48 130 592
use scs8hd_decap_12  FILLER_66_300
timestamp 1586364061
transform 1 0 28704 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_312
timestamp 1586364061
transform 1 0 29808 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_306
timestamp 1586364061
transform 1 0 29256 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_318
timestamp 1586364061
transform 1 0 30360 0 1 38624
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_707
timestamp 1586364061
transform 1 0 32016 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_12  FILLER_66_324
timestamp 1586364061
transform 1 0 30912 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_337
timestamp 1586364061
transform 1 0 32108 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_330
timestamp 1586364061
transform 1 0 31464 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_342
timestamp 1586364061
transform 1 0 32568 0 1 38624
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_715
timestamp 1586364061
transform 1 0 34776 0 1 38624
box -38 -48 130 592
use scs8hd_decap_12  FILLER_66_349
timestamp 1586364061
transform 1 0 33212 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_361
timestamp 1586364061
transform 1 0 34316 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_354
timestamp 1586364061
transform 1 0 33672 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_367
timestamp 1586364061
transform 1 0 34868 0 1 38624
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_708
timestamp 1586364061
transform 1 0 37628 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_12  FILLER_66_373
timestamp 1586364061
transform 1 0 35420 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_385
timestamp 1586364061
transform 1 0 36524 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_379
timestamp 1586364061
transform 1 0 35972 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_391
timestamp 1586364061
transform 1 0 37076 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_398
timestamp 1586364061
transform 1 0 37720 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_410
timestamp 1586364061
transform 1 0 38824 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_422
timestamp 1586364061
transform 1 0 39928 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_403
timestamp 1586364061
transform 1 0 38180 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_415
timestamp 1586364061
transform 1 0 39284 0 1 38624
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_716
timestamp 1586364061
transform 1 0 40388 0 1 38624
box -38 -48 130 592
use scs8hd_decap_12  FILLER_66_434
timestamp 1586364061
transform 1 0 41032 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_446
timestamp 1586364061
transform 1 0 42136 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_428
timestamp 1586364061
transform 1 0 40480 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_440
timestamp 1586364061
transform 1 0 41584 0 1 38624
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_709
timestamp 1586364061
transform 1 0 43240 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_12  FILLER_66_459
timestamp 1586364061
transform 1 0 43332 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_471
timestamp 1586364061
transform 1 0 44436 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_452
timestamp 1586364061
transform 1 0 42688 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_464
timestamp 1586364061
transform 1 0 43792 0 1 38624
box -38 -48 1142 592
use scs8hd_buf_2  _77_
timestamp 1586364061
transform 1 0 46736 0 -1 38624
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_717
timestamp 1586364061
transform 1 0 46000 0 1 38624
box -38 -48 130 592
use scs8hd_decap_12  FILLER_66_483
timestamp 1586364061
transform 1 0 45540 0 -1 38624
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_66_495
timestamp 1586364061
transform 1 0 46644 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_12  FILLER_67_476
timestamp 1586364061
transform 1 0 44896 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_489
timestamp 1586364061
transform 1 0 46092 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_3  PHY_133
timestamp 1586364061
transform -1 0 48852 0 -1 38624
box -38 -48 314 592
use scs8hd_decap_3  PHY_135
timestamp 1586364061
transform -1 0 48852 0 1 38624
box -38 -48 314 592
use scs8hd_decap_12  FILLER_66_500
timestamp 1586364061
transform 1 0 47104 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_66_512
timestamp 1586364061
transform 1 0 48208 0 -1 38624
box -38 -48 406 592
use scs8hd_decap_12  FILLER_67_501
timestamp 1586364061
transform 1 0 47196 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_67_513
timestamp 1586364061
transform 1 0 48300 0 1 38624
box -38 -48 314 592
use scs8hd_decap_3  PHY_136
timestamp 1586364061
transform 1 0 1104 0 -1 39712
box -38 -48 314 592
use scs8hd_decap_12  FILLER_68_3
timestamp 1586364061
transform 1 0 1380 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_15
timestamp 1586364061
transform 1 0 2484 0 -1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_718
timestamp 1586364061
transform 1 0 3956 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_4  FILLER_68_27
timestamp 1586364061
transform 1 0 3588 0 -1 39712
box -38 -48 406 592
use scs8hd_decap_12  FILLER_68_32
timestamp 1586364061
transform 1 0 4048 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_44
timestamp 1586364061
transform 1 0 5152 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_56
timestamp 1586364061
transform 1 0 6256 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_68
timestamp 1586364061
transform 1 0 7360 0 -1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_719
timestamp 1586364061
transform 1 0 9568 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_68_80
timestamp 1586364061
transform 1 0 8464 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_93
timestamp 1586364061
transform 1 0 9660 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_105
timestamp 1586364061
transform 1 0 10764 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_117
timestamp 1586364061
transform 1 0 11868 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_129
timestamp 1586364061
transform 1 0 12972 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_141
timestamp 1586364061
transform 1 0 14076 0 -1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_720
timestamp 1586364061
transform 1 0 15180 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_68_154
timestamp 1586364061
transform 1 0 15272 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_166
timestamp 1586364061
transform 1 0 16376 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_178
timestamp 1586364061
transform 1 0 17480 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_190
timestamp 1586364061
transform 1 0 18584 0 -1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_721
timestamp 1586364061
transform 1 0 20792 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_68_202
timestamp 1586364061
transform 1 0 19688 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_215
timestamp 1586364061
transform 1 0 20884 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_227
timestamp 1586364061
transform 1 0 21988 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_239
timestamp 1586364061
transform 1 0 23092 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_251
timestamp 1586364061
transform 1 0 24196 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_263
timestamp 1586364061
transform 1 0 25300 0 -1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_722
timestamp 1586364061
transform 1 0 26404 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_68_276
timestamp 1586364061
transform 1 0 26496 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_288
timestamp 1586364061
transform 1 0 27600 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_300
timestamp 1586364061
transform 1 0 28704 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_312
timestamp 1586364061
transform 1 0 29808 0 -1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_723
timestamp 1586364061
transform 1 0 32016 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_68_324
timestamp 1586364061
transform 1 0 30912 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_337
timestamp 1586364061
transform 1 0 32108 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_349
timestamp 1586364061
transform 1 0 33212 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_361
timestamp 1586364061
transform 1 0 34316 0 -1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_724
timestamp 1586364061
transform 1 0 37628 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_68_373
timestamp 1586364061
transform 1 0 35420 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_385
timestamp 1586364061
transform 1 0 36524 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_398
timestamp 1586364061
transform 1 0 37720 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_410
timestamp 1586364061
transform 1 0 38824 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_422
timestamp 1586364061
transform 1 0 39928 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_434
timestamp 1586364061
transform 1 0 41032 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_446
timestamp 1586364061
transform 1 0 42136 0 -1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_725
timestamp 1586364061
transform 1 0 43240 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_68_459
timestamp 1586364061
transform 1 0 43332 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_471
timestamp 1586364061
transform 1 0 44436 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_483
timestamp 1586364061
transform 1 0 45540 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_495
timestamp 1586364061
transform 1 0 46644 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_3  PHY_137
timestamp 1586364061
transform -1 0 48852 0 -1 39712
box -38 -48 314 592
use scs8hd_decap_8  FILLER_68_507
timestamp 1586364061
transform 1 0 47748 0 -1 39712
box -38 -48 774 592
use scs8hd_fill_1  FILLER_68_515
timestamp 1586364061
transform 1 0 48484 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_3  PHY_138
timestamp 1586364061
transform 1 0 1104 0 1 39712
box -38 -48 314 592
use scs8hd_decap_12  FILLER_69_3
timestamp 1586364061
transform 1 0 1380 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_15
timestamp 1586364061
transform 1 0 2484 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_27
timestamp 1586364061
transform 1 0 3588 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_39
timestamp 1586364061
transform 1 0 4692 0 1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_726
timestamp 1586364061
transform 1 0 6716 0 1 39712
box -38 -48 130 592
use scs8hd_decap_8  FILLER_69_51
timestamp 1586364061
transform 1 0 5796 0 1 39712
box -38 -48 774 592
use scs8hd_fill_2  FILLER_69_59
timestamp 1586364061
transform 1 0 6532 0 1 39712
box -38 -48 222 592
use scs8hd_decap_12  FILLER_69_62
timestamp 1586364061
transform 1 0 6808 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_74
timestamp 1586364061
transform 1 0 7912 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_86
timestamp 1586364061
transform 1 0 9016 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_98
timestamp 1586364061
transform 1 0 10120 0 1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_727
timestamp 1586364061
transform 1 0 12328 0 1 39712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_69_110
timestamp 1586364061
transform 1 0 11224 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_123
timestamp 1586364061
transform 1 0 12420 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_135
timestamp 1586364061
transform 1 0 13524 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_147
timestamp 1586364061
transform 1 0 14628 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_159
timestamp 1586364061
transform 1 0 15732 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_171
timestamp 1586364061
transform 1 0 16836 0 1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_728
timestamp 1586364061
transform 1 0 17940 0 1 39712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_69_184
timestamp 1586364061
transform 1 0 18032 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_196
timestamp 1586364061
transform 1 0 19136 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_208
timestamp 1586364061
transform 1 0 20240 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_220
timestamp 1586364061
transform 1 0 21344 0 1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_729
timestamp 1586364061
transform 1 0 23552 0 1 39712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_69_232
timestamp 1586364061
transform 1 0 22448 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_245
timestamp 1586364061
transform 1 0 23644 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_257
timestamp 1586364061
transform 1 0 24748 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_269
timestamp 1586364061
transform 1 0 25852 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_281
timestamp 1586364061
transform 1 0 26956 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_293
timestamp 1586364061
transform 1 0 28060 0 1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_730
timestamp 1586364061
transform 1 0 29164 0 1 39712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_69_306
timestamp 1586364061
transform 1 0 29256 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_318
timestamp 1586364061
transform 1 0 30360 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_330
timestamp 1586364061
transform 1 0 31464 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_342
timestamp 1586364061
transform 1 0 32568 0 1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_731
timestamp 1586364061
transform 1 0 34776 0 1 39712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_69_354
timestamp 1586364061
transform 1 0 33672 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_367
timestamp 1586364061
transform 1 0 34868 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_379
timestamp 1586364061
transform 1 0 35972 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_391
timestamp 1586364061
transform 1 0 37076 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_403
timestamp 1586364061
transform 1 0 38180 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_415
timestamp 1586364061
transform 1 0 39284 0 1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_732
timestamp 1586364061
transform 1 0 40388 0 1 39712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_69_428
timestamp 1586364061
transform 1 0 40480 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_440
timestamp 1586364061
transform 1 0 41584 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_452
timestamp 1586364061
transform 1 0 42688 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_464
timestamp 1586364061
transform 1 0 43792 0 1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_733
timestamp 1586364061
transform 1 0 46000 0 1 39712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_69_476
timestamp 1586364061
transform 1 0 44896 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_489
timestamp 1586364061
transform 1 0 46092 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_3  PHY_139
timestamp 1586364061
transform -1 0 48852 0 1 39712
box -38 -48 314 592
use scs8hd_decap_12  FILLER_69_501
timestamp 1586364061
transform 1 0 47196 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_69_513
timestamp 1586364061
transform 1 0 48300 0 1 39712
box -38 -48 314 592
use scs8hd_decap_3  PHY_140
timestamp 1586364061
transform 1 0 1104 0 -1 40800
box -38 -48 314 592
use scs8hd_decap_12  FILLER_70_3
timestamp 1586364061
transform 1 0 1380 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_15
timestamp 1586364061
transform 1 0 2484 0 -1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_734
timestamp 1586364061
transform 1 0 3956 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_4  FILLER_70_27
timestamp 1586364061
transform 1 0 3588 0 -1 40800
box -38 -48 406 592
use scs8hd_decap_12  FILLER_70_32
timestamp 1586364061
transform 1 0 4048 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_44
timestamp 1586364061
transform 1 0 5152 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_56
timestamp 1586364061
transform 1 0 6256 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_68
timestamp 1586364061
transform 1 0 7360 0 -1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_735
timestamp 1586364061
transform 1 0 9568 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_70_80
timestamp 1586364061
transform 1 0 8464 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_93
timestamp 1586364061
transform 1 0 9660 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_105
timestamp 1586364061
transform 1 0 10764 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_117
timestamp 1586364061
transform 1 0 11868 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_129
timestamp 1586364061
transform 1 0 12972 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_141
timestamp 1586364061
transform 1 0 14076 0 -1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_736
timestamp 1586364061
transform 1 0 15180 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_70_154
timestamp 1586364061
transform 1 0 15272 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_166
timestamp 1586364061
transform 1 0 16376 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_178
timestamp 1586364061
transform 1 0 17480 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_190
timestamp 1586364061
transform 1 0 18584 0 -1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_737
timestamp 1586364061
transform 1 0 20792 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_70_202
timestamp 1586364061
transform 1 0 19688 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_215
timestamp 1586364061
transform 1 0 20884 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_227
timestamp 1586364061
transform 1 0 21988 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_239
timestamp 1586364061
transform 1 0 23092 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_251
timestamp 1586364061
transform 1 0 24196 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_263
timestamp 1586364061
transform 1 0 25300 0 -1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_738
timestamp 1586364061
transform 1 0 26404 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_70_276
timestamp 1586364061
transform 1 0 26496 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_288
timestamp 1586364061
transform 1 0 27600 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_300
timestamp 1586364061
transform 1 0 28704 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_312
timestamp 1586364061
transform 1 0 29808 0 -1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_739
timestamp 1586364061
transform 1 0 32016 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_70_324
timestamp 1586364061
transform 1 0 30912 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_337
timestamp 1586364061
transform 1 0 32108 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_349
timestamp 1586364061
transform 1 0 33212 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_361
timestamp 1586364061
transform 1 0 34316 0 -1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_740
timestamp 1586364061
transform 1 0 37628 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_70_373
timestamp 1586364061
transform 1 0 35420 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_385
timestamp 1586364061
transform 1 0 36524 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_398
timestamp 1586364061
transform 1 0 37720 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_410
timestamp 1586364061
transform 1 0 38824 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_422
timestamp 1586364061
transform 1 0 39928 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_434
timestamp 1586364061
transform 1 0 41032 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_446
timestamp 1586364061
transform 1 0 42136 0 -1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_741
timestamp 1586364061
transform 1 0 43240 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_70_459
timestamp 1586364061
transform 1 0 43332 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_471
timestamp 1586364061
transform 1 0 44436 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_483
timestamp 1586364061
transform 1 0 45540 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_495
timestamp 1586364061
transform 1 0 46644 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_3  PHY_141
timestamp 1586364061
transform -1 0 48852 0 -1 40800
box -38 -48 314 592
use scs8hd_decap_8  FILLER_70_507
timestamp 1586364061
transform 1 0 47748 0 -1 40800
box -38 -48 774 592
use scs8hd_fill_1  FILLER_70_515
timestamp 1586364061
transform 1 0 48484 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_3  PHY_142
timestamp 1586364061
transform 1 0 1104 0 1 40800
box -38 -48 314 592
use scs8hd_decap_12  FILLER_71_3
timestamp 1586364061
transform 1 0 1380 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_15
timestamp 1586364061
transform 1 0 2484 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_27
timestamp 1586364061
transform 1 0 3588 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_39
timestamp 1586364061
transform 1 0 4692 0 1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_742
timestamp 1586364061
transform 1 0 6716 0 1 40800
box -38 -48 130 592
use scs8hd_decap_8  FILLER_71_51
timestamp 1586364061
transform 1 0 5796 0 1 40800
box -38 -48 774 592
use scs8hd_fill_2  FILLER_71_59
timestamp 1586364061
transform 1 0 6532 0 1 40800
box -38 -48 222 592
use scs8hd_decap_12  FILLER_71_62
timestamp 1586364061
transform 1 0 6808 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_74
timestamp 1586364061
transform 1 0 7912 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_86
timestamp 1586364061
transform 1 0 9016 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_98
timestamp 1586364061
transform 1 0 10120 0 1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_743
timestamp 1586364061
transform 1 0 12328 0 1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_71_110
timestamp 1586364061
transform 1 0 11224 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_123
timestamp 1586364061
transform 1 0 12420 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_135
timestamp 1586364061
transform 1 0 13524 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_147
timestamp 1586364061
transform 1 0 14628 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_159
timestamp 1586364061
transform 1 0 15732 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_171
timestamp 1586364061
transform 1 0 16836 0 1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_744
timestamp 1586364061
transform 1 0 17940 0 1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_71_184
timestamp 1586364061
transform 1 0 18032 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_196
timestamp 1586364061
transform 1 0 19136 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_208
timestamp 1586364061
transform 1 0 20240 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_220
timestamp 1586364061
transform 1 0 21344 0 1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_745
timestamp 1586364061
transform 1 0 23552 0 1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_71_232
timestamp 1586364061
transform 1 0 22448 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_245
timestamp 1586364061
transform 1 0 23644 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_257
timestamp 1586364061
transform 1 0 24748 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_269
timestamp 1586364061
transform 1 0 25852 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_281
timestamp 1586364061
transform 1 0 26956 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_293
timestamp 1586364061
transform 1 0 28060 0 1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_746
timestamp 1586364061
transform 1 0 29164 0 1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_71_306
timestamp 1586364061
transform 1 0 29256 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_318
timestamp 1586364061
transform 1 0 30360 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_330
timestamp 1586364061
transform 1 0 31464 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_342
timestamp 1586364061
transform 1 0 32568 0 1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_747
timestamp 1586364061
transform 1 0 34776 0 1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_71_354
timestamp 1586364061
transform 1 0 33672 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_367
timestamp 1586364061
transform 1 0 34868 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_379
timestamp 1586364061
transform 1 0 35972 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_391
timestamp 1586364061
transform 1 0 37076 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_403
timestamp 1586364061
transform 1 0 38180 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_415
timestamp 1586364061
transform 1 0 39284 0 1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_748
timestamp 1586364061
transform 1 0 40388 0 1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_71_428
timestamp 1586364061
transform 1 0 40480 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_440
timestamp 1586364061
transform 1 0 41584 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_452
timestamp 1586364061
transform 1 0 42688 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_464
timestamp 1586364061
transform 1 0 43792 0 1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_749
timestamp 1586364061
transform 1 0 46000 0 1 40800
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__78__A
timestamp 1586364061
transform 1 0 46736 0 1 40800
box -38 -48 222 592
use scs8hd_decap_12  FILLER_71_476
timestamp 1586364061
transform 1 0 44896 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_71_489
timestamp 1586364061
transform 1 0 46092 0 1 40800
box -38 -48 590 592
use scs8hd_fill_1  FILLER_71_495
timestamp 1586364061
transform 1 0 46644 0 1 40800
box -38 -48 130 592
use scs8hd_decap_3  PHY_143
timestamp 1586364061
transform -1 0 48852 0 1 40800
box -38 -48 314 592
use scs8hd_decap_12  FILLER_71_498
timestamp 1586364061
transform 1 0 46920 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_71_510
timestamp 1586364061
transform 1 0 48024 0 1 40800
box -38 -48 590 592
use scs8hd_decap_3  PHY_144
timestamp 1586364061
transform 1 0 1104 0 -1 41888
box -38 -48 314 592
use scs8hd_decap_3  PHY_146
timestamp 1586364061
transform 1 0 1104 0 1 41888
box -38 -48 314 592
use scs8hd_decap_12  FILLER_72_3
timestamp 1586364061
transform 1 0 1380 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_15
timestamp 1586364061
transform 1 0 2484 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_3
timestamp 1586364061
transform 1 0 1380 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_15
timestamp 1586364061
transform 1 0 2484 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_750
timestamp 1586364061
transform 1 0 3956 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_4  FILLER_72_27
timestamp 1586364061
transform 1 0 3588 0 -1 41888
box -38 -48 406 592
use scs8hd_decap_12  FILLER_72_32
timestamp 1586364061
transform 1 0 4048 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_44
timestamp 1586364061
transform 1 0 5152 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_27
timestamp 1586364061
transform 1 0 3588 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_39
timestamp 1586364061
transform 1 0 4692 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_758
timestamp 1586364061
transform 1 0 6716 0 1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_56
timestamp 1586364061
transform 1 0 6256 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_68
timestamp 1586364061
transform 1 0 7360 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_73_51
timestamp 1586364061
transform 1 0 5796 0 1 41888
box -38 -48 774 592
use scs8hd_fill_2  FILLER_73_59
timestamp 1586364061
transform 1 0 6532 0 1 41888
box -38 -48 222 592
use scs8hd_decap_12  FILLER_73_62
timestamp 1586364061
transform 1 0 6808 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_74
timestamp 1586364061
transform 1 0 7912 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_751
timestamp 1586364061
transform 1 0 9568 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_80
timestamp 1586364061
transform 1 0 8464 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_93
timestamp 1586364061
transform 1 0 9660 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_86
timestamp 1586364061
transform 1 0 9016 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_98
timestamp 1586364061
transform 1 0 10120 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_759
timestamp 1586364061
transform 1 0 12328 0 1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_105
timestamp 1586364061
transform 1 0 10764 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_117
timestamp 1586364061
transform 1 0 11868 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_110
timestamp 1586364061
transform 1 0 11224 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_123
timestamp 1586364061
transform 1 0 12420 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_129
timestamp 1586364061
transform 1 0 12972 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_141
timestamp 1586364061
transform 1 0 14076 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_135
timestamp 1586364061
transform 1 0 13524 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_147
timestamp 1586364061
transform 1 0 14628 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_752
timestamp 1586364061
transform 1 0 15180 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_154
timestamp 1586364061
transform 1 0 15272 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_166
timestamp 1586364061
transform 1 0 16376 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_159
timestamp 1586364061
transform 1 0 15732 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_171
timestamp 1586364061
transform 1 0 16836 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_760
timestamp 1586364061
transform 1 0 17940 0 1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_178
timestamp 1586364061
transform 1 0 17480 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_190
timestamp 1586364061
transform 1 0 18584 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_184
timestamp 1586364061
transform 1 0 18032 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_196
timestamp 1586364061
transform 1 0 19136 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_753
timestamp 1586364061
transform 1 0 20792 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_202
timestamp 1586364061
transform 1 0 19688 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_215
timestamp 1586364061
transform 1 0 20884 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_208
timestamp 1586364061
transform 1 0 20240 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_220
timestamp 1586364061
transform 1 0 21344 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_761
timestamp 1586364061
transform 1 0 23552 0 1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_227
timestamp 1586364061
transform 1 0 21988 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_239
timestamp 1586364061
transform 1 0 23092 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_232
timestamp 1586364061
transform 1 0 22448 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_245
timestamp 1586364061
transform 1 0 23644 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_251
timestamp 1586364061
transform 1 0 24196 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_263
timestamp 1586364061
transform 1 0 25300 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_257
timestamp 1586364061
transform 1 0 24748 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_269
timestamp 1586364061
transform 1 0 25852 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_754
timestamp 1586364061
transform 1 0 26404 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_276
timestamp 1586364061
transform 1 0 26496 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_288
timestamp 1586364061
transform 1 0 27600 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_281
timestamp 1586364061
transform 1 0 26956 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_293
timestamp 1586364061
transform 1 0 28060 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_762
timestamp 1586364061
transform 1 0 29164 0 1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_300
timestamp 1586364061
transform 1 0 28704 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_312
timestamp 1586364061
transform 1 0 29808 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_306
timestamp 1586364061
transform 1 0 29256 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_318
timestamp 1586364061
transform 1 0 30360 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_755
timestamp 1586364061
transform 1 0 32016 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_324
timestamp 1586364061
transform 1 0 30912 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_337
timestamp 1586364061
transform 1 0 32108 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_330
timestamp 1586364061
transform 1 0 31464 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_342
timestamp 1586364061
transform 1 0 32568 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_763
timestamp 1586364061
transform 1 0 34776 0 1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_349
timestamp 1586364061
transform 1 0 33212 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_361
timestamp 1586364061
transform 1 0 34316 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_354
timestamp 1586364061
transform 1 0 33672 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_367
timestamp 1586364061
transform 1 0 34868 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_756
timestamp 1586364061
transform 1 0 37628 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_373
timestamp 1586364061
transform 1 0 35420 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_385
timestamp 1586364061
transform 1 0 36524 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_379
timestamp 1586364061
transform 1 0 35972 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_391
timestamp 1586364061
transform 1 0 37076 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_398
timestamp 1586364061
transform 1 0 37720 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_410
timestamp 1586364061
transform 1 0 38824 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_422
timestamp 1586364061
transform 1 0 39928 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_403
timestamp 1586364061
transform 1 0 38180 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_415
timestamp 1586364061
transform 1 0 39284 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_764
timestamp 1586364061
transform 1 0 40388 0 1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_434
timestamp 1586364061
transform 1 0 41032 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_446
timestamp 1586364061
transform 1 0 42136 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_428
timestamp 1586364061
transform 1 0 40480 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_440
timestamp 1586364061
transform 1 0 41584 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_757
timestamp 1586364061
transform 1 0 43240 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_459
timestamp 1586364061
transform 1 0 43332 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_471
timestamp 1586364061
transform 1 0 44436 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_452
timestamp 1586364061
transform 1 0 42688 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_464
timestamp 1586364061
transform 1 0 43792 0 1 41888
box -38 -48 1142 592
use scs8hd_buf_2  _78_
timestamp 1586364061
transform 1 0 46736 0 -1 41888
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_765
timestamp 1586364061
transform 1 0 46000 0 1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_483
timestamp 1586364061
transform 1 0 45540 0 -1 41888
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_72_495
timestamp 1586364061
transform 1 0 46644 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_73_476
timestamp 1586364061
transform 1 0 44896 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_489
timestamp 1586364061
transform 1 0 46092 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_3  PHY_145
timestamp 1586364061
transform -1 0 48852 0 -1 41888
box -38 -48 314 592
use scs8hd_decap_3  PHY_147
timestamp 1586364061
transform -1 0 48852 0 1 41888
box -38 -48 314 592
use scs8hd_decap_12  FILLER_72_500
timestamp 1586364061
transform 1 0 47104 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_72_512
timestamp 1586364061
transform 1 0 48208 0 -1 41888
box -38 -48 406 592
use scs8hd_decap_12  FILLER_73_501
timestamp 1586364061
transform 1 0 47196 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_73_513
timestamp 1586364061
transform 1 0 48300 0 1 41888
box -38 -48 314 592
use scs8hd_decap_3  PHY_148
timestamp 1586364061
transform 1 0 1104 0 -1 42976
box -38 -48 314 592
use scs8hd_decap_12  FILLER_74_3
timestamp 1586364061
transform 1 0 1380 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_15
timestamp 1586364061
transform 1 0 2484 0 -1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_766
timestamp 1586364061
transform 1 0 3956 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_4  FILLER_74_27
timestamp 1586364061
transform 1 0 3588 0 -1 42976
box -38 -48 406 592
use scs8hd_decap_12  FILLER_74_32
timestamp 1586364061
transform 1 0 4048 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_44
timestamp 1586364061
transform 1 0 5152 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_56
timestamp 1586364061
transform 1 0 6256 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_68
timestamp 1586364061
transform 1 0 7360 0 -1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_767
timestamp 1586364061
transform 1 0 9568 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_74_80
timestamp 1586364061
transform 1 0 8464 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_93
timestamp 1586364061
transform 1 0 9660 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_105
timestamp 1586364061
transform 1 0 10764 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_117
timestamp 1586364061
transform 1 0 11868 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_129
timestamp 1586364061
transform 1 0 12972 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_141
timestamp 1586364061
transform 1 0 14076 0 -1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_768
timestamp 1586364061
transform 1 0 15180 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_74_154
timestamp 1586364061
transform 1 0 15272 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_166
timestamp 1586364061
transform 1 0 16376 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_178
timestamp 1586364061
transform 1 0 17480 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_190
timestamp 1586364061
transform 1 0 18584 0 -1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_769
timestamp 1586364061
transform 1 0 20792 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_74_202
timestamp 1586364061
transform 1 0 19688 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_215
timestamp 1586364061
transform 1 0 20884 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_227
timestamp 1586364061
transform 1 0 21988 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_239
timestamp 1586364061
transform 1 0 23092 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_251
timestamp 1586364061
transform 1 0 24196 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_263
timestamp 1586364061
transform 1 0 25300 0 -1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_770
timestamp 1586364061
transform 1 0 26404 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_74_276
timestamp 1586364061
transform 1 0 26496 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_288
timestamp 1586364061
transform 1 0 27600 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_300
timestamp 1586364061
transform 1 0 28704 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_312
timestamp 1586364061
transform 1 0 29808 0 -1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_771
timestamp 1586364061
transform 1 0 32016 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_74_324
timestamp 1586364061
transform 1 0 30912 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_337
timestamp 1586364061
transform 1 0 32108 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_349
timestamp 1586364061
transform 1 0 33212 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_361
timestamp 1586364061
transform 1 0 34316 0 -1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_772
timestamp 1586364061
transform 1 0 37628 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_74_373
timestamp 1586364061
transform 1 0 35420 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_385
timestamp 1586364061
transform 1 0 36524 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_398
timestamp 1586364061
transform 1 0 37720 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_410
timestamp 1586364061
transform 1 0 38824 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_422
timestamp 1586364061
transform 1 0 39928 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_434
timestamp 1586364061
transform 1 0 41032 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_446
timestamp 1586364061
transform 1 0 42136 0 -1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_773
timestamp 1586364061
transform 1 0 43240 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_74_459
timestamp 1586364061
transform 1 0 43332 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_471
timestamp 1586364061
transform 1 0 44436 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_483
timestamp 1586364061
transform 1 0 45540 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_495
timestamp 1586364061
transform 1 0 46644 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_3  PHY_149
timestamp 1586364061
transform -1 0 48852 0 -1 42976
box -38 -48 314 592
use scs8hd_decap_8  FILLER_74_507
timestamp 1586364061
transform 1 0 47748 0 -1 42976
box -38 -48 774 592
use scs8hd_fill_1  FILLER_74_515
timestamp 1586364061
transform 1 0 48484 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_3  PHY_150
timestamp 1586364061
transform 1 0 1104 0 1 42976
box -38 -48 314 592
use scs8hd_decap_12  FILLER_75_3
timestamp 1586364061
transform 1 0 1380 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_15
timestamp 1586364061
transform 1 0 2484 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_27
timestamp 1586364061
transform 1 0 3588 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_39
timestamp 1586364061
transform 1 0 4692 0 1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_774
timestamp 1586364061
transform 1 0 6716 0 1 42976
box -38 -48 130 592
use scs8hd_decap_8  FILLER_75_51
timestamp 1586364061
transform 1 0 5796 0 1 42976
box -38 -48 774 592
use scs8hd_fill_2  FILLER_75_59
timestamp 1586364061
transform 1 0 6532 0 1 42976
box -38 -48 222 592
use scs8hd_decap_12  FILLER_75_62
timestamp 1586364061
transform 1 0 6808 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_74
timestamp 1586364061
transform 1 0 7912 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_86
timestamp 1586364061
transform 1 0 9016 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_98
timestamp 1586364061
transform 1 0 10120 0 1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_775
timestamp 1586364061
transform 1 0 12328 0 1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_75_110
timestamp 1586364061
transform 1 0 11224 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_123
timestamp 1586364061
transform 1 0 12420 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_135
timestamp 1586364061
transform 1 0 13524 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_147
timestamp 1586364061
transform 1 0 14628 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_159
timestamp 1586364061
transform 1 0 15732 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_171
timestamp 1586364061
transform 1 0 16836 0 1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_776
timestamp 1586364061
transform 1 0 17940 0 1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_75_184
timestamp 1586364061
transform 1 0 18032 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_196
timestamp 1586364061
transform 1 0 19136 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_208
timestamp 1586364061
transform 1 0 20240 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_220
timestamp 1586364061
transform 1 0 21344 0 1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_777
timestamp 1586364061
transform 1 0 23552 0 1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_75_232
timestamp 1586364061
transform 1 0 22448 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_245
timestamp 1586364061
transform 1 0 23644 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_257
timestamp 1586364061
transform 1 0 24748 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_269
timestamp 1586364061
transform 1 0 25852 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_281
timestamp 1586364061
transform 1 0 26956 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_293
timestamp 1586364061
transform 1 0 28060 0 1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_778
timestamp 1586364061
transform 1 0 29164 0 1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_75_306
timestamp 1586364061
transform 1 0 29256 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_318
timestamp 1586364061
transform 1 0 30360 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_330
timestamp 1586364061
transform 1 0 31464 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_342
timestamp 1586364061
transform 1 0 32568 0 1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_779
timestamp 1586364061
transform 1 0 34776 0 1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_75_354
timestamp 1586364061
transform 1 0 33672 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_367
timestamp 1586364061
transform 1 0 34868 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_379
timestamp 1586364061
transform 1 0 35972 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_391
timestamp 1586364061
transform 1 0 37076 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_403
timestamp 1586364061
transform 1 0 38180 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_415
timestamp 1586364061
transform 1 0 39284 0 1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_780
timestamp 1586364061
transform 1 0 40388 0 1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_75_428
timestamp 1586364061
transform 1 0 40480 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_440
timestamp 1586364061
transform 1 0 41584 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_452
timestamp 1586364061
transform 1 0 42688 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_464
timestamp 1586364061
transform 1 0 43792 0 1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_781
timestamp 1586364061
transform 1 0 46000 0 1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_75_476
timestamp 1586364061
transform 1 0 44896 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_489
timestamp 1586364061
transform 1 0 46092 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_3  PHY_151
timestamp 1586364061
transform -1 0 48852 0 1 42976
box -38 -48 314 592
use scs8hd_decap_12  FILLER_75_501
timestamp 1586364061
transform 1 0 47196 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_75_513
timestamp 1586364061
transform 1 0 48300 0 1 42976
box -38 -48 314 592
use scs8hd_decap_3  PHY_152
timestamp 1586364061
transform 1 0 1104 0 -1 44064
box -38 -48 314 592
use scs8hd_decap_12  FILLER_76_3
timestamp 1586364061
transform 1 0 1380 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_15
timestamp 1586364061
transform 1 0 2484 0 -1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_782
timestamp 1586364061
transform 1 0 3956 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_4  FILLER_76_27
timestamp 1586364061
transform 1 0 3588 0 -1 44064
box -38 -48 406 592
use scs8hd_decap_12  FILLER_76_32
timestamp 1586364061
transform 1 0 4048 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_44
timestamp 1586364061
transform 1 0 5152 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_56
timestamp 1586364061
transform 1 0 6256 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_68
timestamp 1586364061
transform 1 0 7360 0 -1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_783
timestamp 1586364061
transform 1 0 9568 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_76_80
timestamp 1586364061
transform 1 0 8464 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_93
timestamp 1586364061
transform 1 0 9660 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_105
timestamp 1586364061
transform 1 0 10764 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_117
timestamp 1586364061
transform 1 0 11868 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_129
timestamp 1586364061
transform 1 0 12972 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_141
timestamp 1586364061
transform 1 0 14076 0 -1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_784
timestamp 1586364061
transform 1 0 15180 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_76_154
timestamp 1586364061
transform 1 0 15272 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_166
timestamp 1586364061
transform 1 0 16376 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_178
timestamp 1586364061
transform 1 0 17480 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_190
timestamp 1586364061
transform 1 0 18584 0 -1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_785
timestamp 1586364061
transform 1 0 20792 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_76_202
timestamp 1586364061
transform 1 0 19688 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_215
timestamp 1586364061
transform 1 0 20884 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_227
timestamp 1586364061
transform 1 0 21988 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_239
timestamp 1586364061
transform 1 0 23092 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_251
timestamp 1586364061
transform 1 0 24196 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_263
timestamp 1586364061
transform 1 0 25300 0 -1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_786
timestamp 1586364061
transform 1 0 26404 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_76_276
timestamp 1586364061
transform 1 0 26496 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_288
timestamp 1586364061
transform 1 0 27600 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_300
timestamp 1586364061
transform 1 0 28704 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_312
timestamp 1586364061
transform 1 0 29808 0 -1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_787
timestamp 1586364061
transform 1 0 32016 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_76_324
timestamp 1586364061
transform 1 0 30912 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_337
timestamp 1586364061
transform 1 0 32108 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_349
timestamp 1586364061
transform 1 0 33212 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_361
timestamp 1586364061
transform 1 0 34316 0 -1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_788
timestamp 1586364061
transform 1 0 37628 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_76_373
timestamp 1586364061
transform 1 0 35420 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_385
timestamp 1586364061
transform 1 0 36524 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_398
timestamp 1586364061
transform 1 0 37720 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_410
timestamp 1586364061
transform 1 0 38824 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_422
timestamp 1586364061
transform 1 0 39928 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_434
timestamp 1586364061
transform 1 0 41032 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_446
timestamp 1586364061
transform 1 0 42136 0 -1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_789
timestamp 1586364061
transform 1 0 43240 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_76_459
timestamp 1586364061
transform 1 0 43332 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_471
timestamp 1586364061
transform 1 0 44436 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_483
timestamp 1586364061
transform 1 0 45540 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_495
timestamp 1586364061
transform 1 0 46644 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_3  PHY_153
timestamp 1586364061
transform -1 0 48852 0 -1 44064
box -38 -48 314 592
use scs8hd_decap_8  FILLER_76_507
timestamp 1586364061
transform 1 0 47748 0 -1 44064
box -38 -48 774 592
use scs8hd_fill_1  FILLER_76_515
timestamp 1586364061
transform 1 0 48484 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_3  PHY_154
timestamp 1586364061
transform 1 0 1104 0 1 44064
box -38 -48 314 592
use scs8hd_decap_12  FILLER_77_3
timestamp 1586364061
transform 1 0 1380 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_15
timestamp 1586364061
transform 1 0 2484 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_27
timestamp 1586364061
transform 1 0 3588 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_39
timestamp 1586364061
transform 1 0 4692 0 1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_790
timestamp 1586364061
transform 1 0 6716 0 1 44064
box -38 -48 130 592
use scs8hd_decap_8  FILLER_77_51
timestamp 1586364061
transform 1 0 5796 0 1 44064
box -38 -48 774 592
use scs8hd_fill_2  FILLER_77_59
timestamp 1586364061
transform 1 0 6532 0 1 44064
box -38 -48 222 592
use scs8hd_decap_12  FILLER_77_62
timestamp 1586364061
transform 1 0 6808 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_74
timestamp 1586364061
transform 1 0 7912 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_86
timestamp 1586364061
transform 1 0 9016 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_98
timestamp 1586364061
transform 1 0 10120 0 1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_791
timestamp 1586364061
transform 1 0 12328 0 1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_77_110
timestamp 1586364061
transform 1 0 11224 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_123
timestamp 1586364061
transform 1 0 12420 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_135
timestamp 1586364061
transform 1 0 13524 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_147
timestamp 1586364061
transform 1 0 14628 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_159
timestamp 1586364061
transform 1 0 15732 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_171
timestamp 1586364061
transform 1 0 16836 0 1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_792
timestamp 1586364061
transform 1 0 17940 0 1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_77_184
timestamp 1586364061
transform 1 0 18032 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_196
timestamp 1586364061
transform 1 0 19136 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_208
timestamp 1586364061
transform 1 0 20240 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_220
timestamp 1586364061
transform 1 0 21344 0 1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_793
timestamp 1586364061
transform 1 0 23552 0 1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_77_232
timestamp 1586364061
transform 1 0 22448 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_245
timestamp 1586364061
transform 1 0 23644 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_257
timestamp 1586364061
transform 1 0 24748 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_269
timestamp 1586364061
transform 1 0 25852 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_281
timestamp 1586364061
transform 1 0 26956 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_293
timestamp 1586364061
transform 1 0 28060 0 1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_794
timestamp 1586364061
transform 1 0 29164 0 1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_77_306
timestamp 1586364061
transform 1 0 29256 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_318
timestamp 1586364061
transform 1 0 30360 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_330
timestamp 1586364061
transform 1 0 31464 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_342
timestamp 1586364061
transform 1 0 32568 0 1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_795
timestamp 1586364061
transform 1 0 34776 0 1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_77_354
timestamp 1586364061
transform 1 0 33672 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_367
timestamp 1586364061
transform 1 0 34868 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_379
timestamp 1586364061
transform 1 0 35972 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_391
timestamp 1586364061
transform 1 0 37076 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_403
timestamp 1586364061
transform 1 0 38180 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_415
timestamp 1586364061
transform 1 0 39284 0 1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_796
timestamp 1586364061
transform 1 0 40388 0 1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_77_428
timestamp 1586364061
transform 1 0 40480 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_440
timestamp 1586364061
transform 1 0 41584 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_452
timestamp 1586364061
transform 1 0 42688 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_464
timestamp 1586364061
transform 1 0 43792 0 1 44064
box -38 -48 1142 592
use scs8hd_buf_2  _79_
timestamp 1586364061
transform 1 0 46736 0 1 44064
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_797
timestamp 1586364061
transform 1 0 46000 0 1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_77_476
timestamp 1586364061
transform 1 0 44896 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_77_489
timestamp 1586364061
transform 1 0 46092 0 1 44064
box -38 -48 590 592
use scs8hd_fill_1  FILLER_77_495
timestamp 1586364061
transform 1 0 46644 0 1 44064
box -38 -48 130 592
use scs8hd_decap_3  PHY_155
timestamp 1586364061
transform -1 0 48852 0 1 44064
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__79__A
timestamp 1586364061
transform 1 0 47288 0 1 44064
box -38 -48 222 592
use scs8hd_fill_2  FILLER_77_500
timestamp 1586364061
transform 1 0 47104 0 1 44064
box -38 -48 222 592
use scs8hd_decap_12  FILLER_77_504
timestamp 1586364061
transform 1 0 47472 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_3  PHY_156
timestamp 1586364061
transform 1 0 1104 0 -1 45152
box -38 -48 314 592
use scs8hd_decap_12  FILLER_78_3
timestamp 1586364061
transform 1 0 1380 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_15
timestamp 1586364061
transform 1 0 2484 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_798
timestamp 1586364061
transform 1 0 3956 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_4  FILLER_78_27
timestamp 1586364061
transform 1 0 3588 0 -1 45152
box -38 -48 406 592
use scs8hd_decap_12  FILLER_78_32
timestamp 1586364061
transform 1 0 4048 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_44
timestamp 1586364061
transform 1 0 5152 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_56
timestamp 1586364061
transform 1 0 6256 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_68
timestamp 1586364061
transform 1 0 7360 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_799
timestamp 1586364061
transform 1 0 9568 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_78_80
timestamp 1586364061
transform 1 0 8464 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_93
timestamp 1586364061
transform 1 0 9660 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_105
timestamp 1586364061
transform 1 0 10764 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_117
timestamp 1586364061
transform 1 0 11868 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_129
timestamp 1586364061
transform 1 0 12972 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_141
timestamp 1586364061
transform 1 0 14076 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_800
timestamp 1586364061
transform 1 0 15180 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_78_154
timestamp 1586364061
transform 1 0 15272 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_166
timestamp 1586364061
transform 1 0 16376 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_178
timestamp 1586364061
transform 1 0 17480 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_190
timestamp 1586364061
transform 1 0 18584 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_801
timestamp 1586364061
transform 1 0 20792 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_78_202
timestamp 1586364061
transform 1 0 19688 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_215
timestamp 1586364061
transform 1 0 20884 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_227
timestamp 1586364061
transform 1 0 21988 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_239
timestamp 1586364061
transform 1 0 23092 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_251
timestamp 1586364061
transform 1 0 24196 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_263
timestamp 1586364061
transform 1 0 25300 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_802
timestamp 1586364061
transform 1 0 26404 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_78_276
timestamp 1586364061
transform 1 0 26496 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_288
timestamp 1586364061
transform 1 0 27600 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_300
timestamp 1586364061
transform 1 0 28704 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_312
timestamp 1586364061
transform 1 0 29808 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_803
timestamp 1586364061
transform 1 0 32016 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_78_324
timestamp 1586364061
transform 1 0 30912 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_337
timestamp 1586364061
transform 1 0 32108 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_349
timestamp 1586364061
transform 1 0 33212 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_361
timestamp 1586364061
transform 1 0 34316 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_804
timestamp 1586364061
transform 1 0 37628 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_78_373
timestamp 1586364061
transform 1 0 35420 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_385
timestamp 1586364061
transform 1 0 36524 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_398
timestamp 1586364061
transform 1 0 37720 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_410
timestamp 1586364061
transform 1 0 38824 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_422
timestamp 1586364061
transform 1 0 39928 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_434
timestamp 1586364061
transform 1 0 41032 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_446
timestamp 1586364061
transform 1 0 42136 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_805
timestamp 1586364061
transform 1 0 43240 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_78_459
timestamp 1586364061
transform 1 0 43332 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_471
timestamp 1586364061
transform 1 0 44436 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_483
timestamp 1586364061
transform 1 0 45540 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_495
timestamp 1586364061
transform 1 0 46644 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_3  PHY_157
timestamp 1586364061
transform -1 0 48852 0 -1 45152
box -38 -48 314 592
use scs8hd_decap_8  FILLER_78_507
timestamp 1586364061
transform 1 0 47748 0 -1 45152
box -38 -48 774 592
use scs8hd_fill_1  FILLER_78_515
timestamp 1586364061
transform 1 0 48484 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_3  PHY_158
timestamp 1586364061
transform 1 0 1104 0 1 45152
box -38 -48 314 592
use scs8hd_decap_3  PHY_160
timestamp 1586364061
transform 1 0 1104 0 -1 46240
box -38 -48 314 592
use scs8hd_decap_12  FILLER_79_3
timestamp 1586364061
transform 1 0 1380 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_15
timestamp 1586364061
transform 1 0 2484 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_3
timestamp 1586364061
transform 1 0 1380 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_15
timestamp 1586364061
transform 1 0 2484 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_814
timestamp 1586364061
transform 1 0 3956 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_27
timestamp 1586364061
transform 1 0 3588 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_39
timestamp 1586364061
transform 1 0 4692 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_80_27
timestamp 1586364061
transform 1 0 3588 0 -1 46240
box -38 -48 406 592
use scs8hd_decap_12  FILLER_80_32
timestamp 1586364061
transform 1 0 4048 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_44
timestamp 1586364061
transform 1 0 5152 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_806
timestamp 1586364061
transform 1 0 6716 0 1 45152
box -38 -48 130 592
use scs8hd_decap_8  FILLER_79_51
timestamp 1586364061
transform 1 0 5796 0 1 45152
box -38 -48 774 592
use scs8hd_fill_2  FILLER_79_59
timestamp 1586364061
transform 1 0 6532 0 1 45152
box -38 -48 222 592
use scs8hd_decap_12  FILLER_79_62
timestamp 1586364061
transform 1 0 6808 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_74
timestamp 1586364061
transform 1 0 7912 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_56
timestamp 1586364061
transform 1 0 6256 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_68
timestamp 1586364061
transform 1 0 7360 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_815
timestamp 1586364061
transform 1 0 9568 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_86
timestamp 1586364061
transform 1 0 9016 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_98
timestamp 1586364061
transform 1 0 10120 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_80
timestamp 1586364061
transform 1 0 8464 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_93
timestamp 1586364061
transform 1 0 9660 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_807
timestamp 1586364061
transform 1 0 12328 0 1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_110
timestamp 1586364061
transform 1 0 11224 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_123
timestamp 1586364061
transform 1 0 12420 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_105
timestamp 1586364061
transform 1 0 10764 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_117
timestamp 1586364061
transform 1 0 11868 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_135
timestamp 1586364061
transform 1 0 13524 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_147
timestamp 1586364061
transform 1 0 14628 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_129
timestamp 1586364061
transform 1 0 12972 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_141
timestamp 1586364061
transform 1 0 14076 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_816
timestamp 1586364061
transform 1 0 15180 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_159
timestamp 1586364061
transform 1 0 15732 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_171
timestamp 1586364061
transform 1 0 16836 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_154
timestamp 1586364061
transform 1 0 15272 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_166
timestamp 1586364061
transform 1 0 16376 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_808
timestamp 1586364061
transform 1 0 17940 0 1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_184
timestamp 1586364061
transform 1 0 18032 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_196
timestamp 1586364061
transform 1 0 19136 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_178
timestamp 1586364061
transform 1 0 17480 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_190
timestamp 1586364061
transform 1 0 18584 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_817
timestamp 1586364061
transform 1 0 20792 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_208
timestamp 1586364061
transform 1 0 20240 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_220
timestamp 1586364061
transform 1 0 21344 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_202
timestamp 1586364061
transform 1 0 19688 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_215
timestamp 1586364061
transform 1 0 20884 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_809
timestamp 1586364061
transform 1 0 23552 0 1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_232
timestamp 1586364061
transform 1 0 22448 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_245
timestamp 1586364061
transform 1 0 23644 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_227
timestamp 1586364061
transform 1 0 21988 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_239
timestamp 1586364061
transform 1 0 23092 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_257
timestamp 1586364061
transform 1 0 24748 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_269
timestamp 1586364061
transform 1 0 25852 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_251
timestamp 1586364061
transform 1 0 24196 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_263
timestamp 1586364061
transform 1 0 25300 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_818
timestamp 1586364061
transform 1 0 26404 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_281
timestamp 1586364061
transform 1 0 26956 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_293
timestamp 1586364061
transform 1 0 28060 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_276
timestamp 1586364061
transform 1 0 26496 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_288
timestamp 1586364061
transform 1 0 27600 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_810
timestamp 1586364061
transform 1 0 29164 0 1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_306
timestamp 1586364061
transform 1 0 29256 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_318
timestamp 1586364061
transform 1 0 30360 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_300
timestamp 1586364061
transform 1 0 28704 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_312
timestamp 1586364061
transform 1 0 29808 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_819
timestamp 1586364061
transform 1 0 32016 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_330
timestamp 1586364061
transform 1 0 31464 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_342
timestamp 1586364061
transform 1 0 32568 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_324
timestamp 1586364061
transform 1 0 30912 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_337
timestamp 1586364061
transform 1 0 32108 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_811
timestamp 1586364061
transform 1 0 34776 0 1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_354
timestamp 1586364061
transform 1 0 33672 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_367
timestamp 1586364061
transform 1 0 34868 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_349
timestamp 1586364061
transform 1 0 33212 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_361
timestamp 1586364061
transform 1 0 34316 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_820
timestamp 1586364061
transform 1 0 37628 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_379
timestamp 1586364061
transform 1 0 35972 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_391
timestamp 1586364061
transform 1 0 37076 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_373
timestamp 1586364061
transform 1 0 35420 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_385
timestamp 1586364061
transform 1 0 36524 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_403
timestamp 1586364061
transform 1 0 38180 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_415
timestamp 1586364061
transform 1 0 39284 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_398
timestamp 1586364061
transform 1 0 37720 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_410
timestamp 1586364061
transform 1 0 38824 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_422
timestamp 1586364061
transform 1 0 39928 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_812
timestamp 1586364061
transform 1 0 40388 0 1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_428
timestamp 1586364061
transform 1 0 40480 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_440
timestamp 1586364061
transform 1 0 41584 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_434
timestamp 1586364061
transform 1 0 41032 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_446
timestamp 1586364061
transform 1 0 42136 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_821
timestamp 1586364061
transform 1 0 43240 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_452
timestamp 1586364061
transform 1 0 42688 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_464
timestamp 1586364061
transform 1 0 43792 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_459
timestamp 1586364061
transform 1 0 43332 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_471
timestamp 1586364061
transform 1 0 44436 0 -1 46240
box -38 -48 1142 592
use scs8hd_buf_2  _80_
timestamp 1586364061
transform 1 0 46736 0 1 45152
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_813
timestamp 1586364061
transform 1 0 46000 0 1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_476
timestamp 1586364061
transform 1 0 44896 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_79_489
timestamp 1586364061
transform 1 0 46092 0 1 45152
box -38 -48 590 592
use scs8hd_fill_1  FILLER_79_495
timestamp 1586364061
transform 1 0 46644 0 1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_80_483
timestamp 1586364061
transform 1 0 45540 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_495
timestamp 1586364061
transform 1 0 46644 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_3  PHY_159
timestamp 1586364061
transform -1 0 48852 0 1 45152
box -38 -48 314 592
use scs8hd_decap_3  PHY_161
timestamp 1586364061
transform -1 0 48852 0 -1 46240
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__80__A
timestamp 1586364061
transform 1 0 47288 0 1 45152
box -38 -48 222 592
use scs8hd_fill_2  FILLER_79_500
timestamp 1586364061
transform 1 0 47104 0 1 45152
box -38 -48 222 592
use scs8hd_decap_12  FILLER_79_504
timestamp 1586364061
transform 1 0 47472 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_80_507
timestamp 1586364061
transform 1 0 47748 0 -1 46240
box -38 -48 774 592
use scs8hd_fill_1  FILLER_80_515
timestamp 1586364061
transform 1 0 48484 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_3  PHY_162
timestamp 1586364061
transform 1 0 1104 0 1 46240
box -38 -48 314 592
use scs8hd_decap_12  FILLER_81_3
timestamp 1586364061
transform 1 0 1380 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_15
timestamp 1586364061
transform 1 0 2484 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_27
timestamp 1586364061
transform 1 0 3588 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_39
timestamp 1586364061
transform 1 0 4692 0 1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_822
timestamp 1586364061
transform 1 0 6716 0 1 46240
box -38 -48 130 592
use scs8hd_decap_8  FILLER_81_51
timestamp 1586364061
transform 1 0 5796 0 1 46240
box -38 -48 774 592
use scs8hd_fill_2  FILLER_81_59
timestamp 1586364061
transform 1 0 6532 0 1 46240
box -38 -48 222 592
use scs8hd_decap_12  FILLER_81_62
timestamp 1586364061
transform 1 0 6808 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_74
timestamp 1586364061
transform 1 0 7912 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_86
timestamp 1586364061
transform 1 0 9016 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_98
timestamp 1586364061
transform 1 0 10120 0 1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_823
timestamp 1586364061
transform 1 0 12328 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_110
timestamp 1586364061
transform 1 0 11224 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_123
timestamp 1586364061
transform 1 0 12420 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_135
timestamp 1586364061
transform 1 0 13524 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_147
timestamp 1586364061
transform 1 0 14628 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_159
timestamp 1586364061
transform 1 0 15732 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_171
timestamp 1586364061
transform 1 0 16836 0 1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_824
timestamp 1586364061
transform 1 0 17940 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_184
timestamp 1586364061
transform 1 0 18032 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_196
timestamp 1586364061
transform 1 0 19136 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_208
timestamp 1586364061
transform 1 0 20240 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_220
timestamp 1586364061
transform 1 0 21344 0 1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_825
timestamp 1586364061
transform 1 0 23552 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_232
timestamp 1586364061
transform 1 0 22448 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_245
timestamp 1586364061
transform 1 0 23644 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_257
timestamp 1586364061
transform 1 0 24748 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_269
timestamp 1586364061
transform 1 0 25852 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_281
timestamp 1586364061
transform 1 0 26956 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_293
timestamp 1586364061
transform 1 0 28060 0 1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_826
timestamp 1586364061
transform 1 0 29164 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_306
timestamp 1586364061
transform 1 0 29256 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_318
timestamp 1586364061
transform 1 0 30360 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_330
timestamp 1586364061
transform 1 0 31464 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_342
timestamp 1586364061
transform 1 0 32568 0 1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_827
timestamp 1586364061
transform 1 0 34776 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_354
timestamp 1586364061
transform 1 0 33672 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_367
timestamp 1586364061
transform 1 0 34868 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_379
timestamp 1586364061
transform 1 0 35972 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_391
timestamp 1586364061
transform 1 0 37076 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_403
timestamp 1586364061
transform 1 0 38180 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_415
timestamp 1586364061
transform 1 0 39284 0 1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_828
timestamp 1586364061
transform 1 0 40388 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_428
timestamp 1586364061
transform 1 0 40480 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_440
timestamp 1586364061
transform 1 0 41584 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_452
timestamp 1586364061
transform 1 0 42688 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_464
timestamp 1586364061
transform 1 0 43792 0 1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_829
timestamp 1586364061
transform 1 0 46000 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_476
timestamp 1586364061
transform 1 0 44896 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_489
timestamp 1586364061
transform 1 0 46092 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_3  PHY_163
timestamp 1586364061
transform -1 0 48852 0 1 46240
box -38 -48 314 592
use scs8hd_decap_12  FILLER_81_501
timestamp 1586364061
transform 1 0 47196 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_81_513
timestamp 1586364061
transform 1 0 48300 0 1 46240
box -38 -48 314 592
use scs8hd_decap_3  PHY_164
timestamp 1586364061
transform 1 0 1104 0 -1 47328
box -38 -48 314 592
use scs8hd_decap_12  FILLER_82_3
timestamp 1586364061
transform 1 0 1380 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_15
timestamp 1586364061
transform 1 0 2484 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_830
timestamp 1586364061
transform 1 0 3956 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_4  FILLER_82_27
timestamp 1586364061
transform 1 0 3588 0 -1 47328
box -38 -48 406 592
use scs8hd_decap_12  FILLER_82_32
timestamp 1586364061
transform 1 0 4048 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_44
timestamp 1586364061
transform 1 0 5152 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_831
timestamp 1586364061
transform 1 0 6808 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_6  FILLER_82_56
timestamp 1586364061
transform 1 0 6256 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_63
timestamp 1586364061
transform 1 0 6900 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_832
timestamp 1586364061
transform 1 0 9660 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_75
timestamp 1586364061
transform 1 0 8004 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_87
timestamp 1586364061
transform 1 0 9108 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_94
timestamp 1586364061
transform 1 0 9752 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_833
timestamp 1586364061
transform 1 0 12512 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_106
timestamp 1586364061
transform 1 0 10856 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_118
timestamp 1586364061
transform 1 0 11960 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_125
timestamp 1586364061
transform 1 0 12604 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_137
timestamp 1586364061
transform 1 0 13708 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_149
timestamp 1586364061
transform 1 0 14812 0 -1 47328
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_834
timestamp 1586364061
transform 1 0 15364 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_156
timestamp 1586364061
transform 1 0 15456 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_168
timestamp 1586364061
transform 1 0 16560 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_835
timestamp 1586364061
transform 1 0 18216 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_6  FILLER_82_180
timestamp 1586364061
transform 1 0 17664 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_187
timestamp 1586364061
transform 1 0 18308 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_836
timestamp 1586364061
transform 1 0 21068 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_199
timestamp 1586364061
transform 1 0 19412 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_211
timestamp 1586364061
transform 1 0 20516 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_218
timestamp 1586364061
transform 1 0 21160 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_837
timestamp 1586364061
transform 1 0 23920 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_230
timestamp 1586364061
transform 1 0 22264 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_242
timestamp 1586364061
transform 1 0 23368 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_249
timestamp 1586364061
transform 1 0 24012 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_261
timestamp 1586364061
transform 1 0 25116 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_273
timestamp 1586364061
transform 1 0 26220 0 -1 47328
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_838
timestamp 1586364061
transform 1 0 26772 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_280
timestamp 1586364061
transform 1 0 26864 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_292
timestamp 1586364061
transform 1 0 27968 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_839
timestamp 1586364061
transform 1 0 29624 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_6  FILLER_82_304
timestamp 1586364061
transform 1 0 29072 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_311
timestamp 1586364061
transform 1 0 29716 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_840
timestamp 1586364061
transform 1 0 32476 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_323
timestamp 1586364061
transform 1 0 30820 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_335
timestamp 1586364061
transform 1 0 31924 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_342
timestamp 1586364061
transform 1 0 32568 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_841
timestamp 1586364061
transform 1 0 35328 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_354
timestamp 1586364061
transform 1 0 33672 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_366
timestamp 1586364061
transform 1 0 34776 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_373
timestamp 1586364061
transform 1 0 35420 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_385
timestamp 1586364061
transform 1 0 36524 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_397
timestamp 1586364061
transform 1 0 37628 0 -1 47328
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_842
timestamp 1586364061
transform 1 0 38180 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_404
timestamp 1586364061
transform 1 0 38272 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_416
timestamp 1586364061
transform 1 0 39376 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_843
timestamp 1586364061
transform 1 0 41032 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_6  FILLER_82_428
timestamp 1586364061
transform 1 0 40480 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_435
timestamp 1586364061
transform 1 0 41124 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_447
timestamp 1586364061
transform 1 0 42228 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_844
timestamp 1586364061
transform 1 0 43884 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_6  FILLER_82_459
timestamp 1586364061
transform 1 0 43332 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_466
timestamp 1586364061
transform 1 0 43976 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_845
timestamp 1586364061
transform 1 0 46736 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_478
timestamp 1586364061
transform 1 0 45080 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_490
timestamp 1586364061
transform 1 0 46184 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_3  PHY_165
timestamp 1586364061
transform -1 0 48852 0 -1 47328
box -38 -48 314 592
use scs8hd_decap_12  FILLER_82_497
timestamp 1586364061
transform 1 0 46828 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_509
timestamp 1586364061
transform 1 0 47932 0 -1 47328
box -38 -48 590 592
use scs8hd_fill_1  FILLER_82_515
timestamp 1586364061
transform 1 0 48484 0 -1 47328
box -38 -48 130 592
<< labels >>
rlabel metal2 s 47858 0 47914 480 6 Test_en
port 0 nsew default input
rlabel metal2 s 1950 0 2006 480 6 bottom_width_0_height_0__pin_16_
port 1 nsew default input
rlabel metal2 s 3330 0 3386 480 6 bottom_width_0_height_0__pin_17_
port 2 nsew default input
rlabel metal2 s 4710 0 4766 480 6 bottom_width_0_height_0__pin_18_
port 3 nsew default input
rlabel metal2 s 5998 0 6054 480 6 bottom_width_0_height_0__pin_19_
port 4 nsew default input
rlabel metal2 s 7378 0 7434 480 6 bottom_width_0_height_0__pin_20_
port 5 nsew default input
rlabel metal2 s 8758 0 8814 480 6 bottom_width_0_height_0__pin_21_
port 6 nsew default input
rlabel metal2 s 10046 0 10102 480 6 bottom_width_0_height_0__pin_22_
port 7 nsew default input
rlabel metal2 s 11426 0 11482 480 6 bottom_width_0_height_0__pin_23_
port 8 nsew default input
rlabel metal2 s 12806 0 12862 480 6 bottom_width_0_height_0__pin_24_
port 9 nsew default input
rlabel metal2 s 14094 0 14150 480 6 bottom_width_0_height_0__pin_25_
port 10 nsew default input
rlabel metal2 s 15474 0 15530 480 6 bottom_width_0_height_0__pin_26_
port 11 nsew default input
rlabel metal2 s 16854 0 16910 480 6 bottom_width_0_height_0__pin_27_
port 12 nsew default input
rlabel metal2 s 18142 0 18198 480 6 bottom_width_0_height_0__pin_28_
port 13 nsew default input
rlabel metal2 s 19522 0 19578 480 6 bottom_width_0_height_0__pin_29_
port 14 nsew default input
rlabel metal2 s 20902 0 20958 480 6 bottom_width_0_height_0__pin_30_
port 15 nsew default input
rlabel metal2 s 22190 0 22246 480 6 bottom_width_0_height_0__pin_31_
port 16 nsew default input
rlabel metal2 s 23570 0 23626 480 6 bottom_width_0_height_0__pin_42_lower
port 17 nsew default tristate
rlabel metal2 s 24950 0 25006 480 6 bottom_width_0_height_0__pin_42_upper
port 18 nsew default tristate
rlabel metal2 s 26238 0 26294 480 6 bottom_width_0_height_0__pin_43_lower
port 19 nsew default tristate
rlabel metal2 s 27618 0 27674 480 6 bottom_width_0_height_0__pin_43_upper
port 20 nsew default tristate
rlabel metal2 s 28998 0 29054 480 6 bottom_width_0_height_0__pin_44_lower
port 21 nsew default tristate
rlabel metal2 s 30286 0 30342 480 6 bottom_width_0_height_0__pin_44_upper
port 22 nsew default tristate
rlabel metal2 s 31666 0 31722 480 6 bottom_width_0_height_0__pin_45_lower
port 23 nsew default tristate
rlabel metal2 s 33046 0 33102 480 6 bottom_width_0_height_0__pin_45_upper
port 24 nsew default tristate
rlabel metal2 s 34334 0 34390 480 6 bottom_width_0_height_0__pin_46_lower
port 25 nsew default tristate
rlabel metal2 s 35714 0 35770 480 6 bottom_width_0_height_0__pin_46_upper
port 26 nsew default tristate
rlabel metal2 s 37094 0 37150 480 6 bottom_width_0_height_0__pin_47_lower
port 27 nsew default tristate
rlabel metal2 s 38382 0 38438 480 6 bottom_width_0_height_0__pin_47_upper
port 28 nsew default tristate
rlabel metal2 s 39762 0 39818 480 6 bottom_width_0_height_0__pin_48_lower
port 29 nsew default tristate
rlabel metal2 s 41142 0 41198 480 6 bottom_width_0_height_0__pin_48_upper
port 30 nsew default tristate
rlabel metal2 s 42430 0 42486 480 6 bottom_width_0_height_0__pin_49_lower
port 31 nsew default tristate
rlabel metal2 s 43810 0 43866 480 6 bottom_width_0_height_0__pin_49_upper
port 32 nsew default tristate
rlabel metal2 s 45190 0 45246 480 6 bottom_width_0_height_0__pin_50_
port 33 nsew default tristate
rlabel metal2 s 46478 0 46534 480 6 bottom_width_0_height_0__pin_51_
port 34 nsew default tristate
rlabel metal3 s 0 37544 480 37664 6 ccff_head
port 35 nsew default input
rlabel metal2 s 41602 49520 41658 50000 6 ccff_tail
port 36 nsew default tristate
rlabel metal2 s 662 0 718 480 6 clk
port 37 nsew default input
rlabel metal3 s 0 12520 480 12640 6 left_width_0_height_0__pin_52_
port 38 nsew default input
rlabel metal2 s 49238 0 49294 480 6 prog_clk
port 39 nsew default input
rlabel metal3 s 49520 688 50000 808 6 right_width_0_height_0__pin_0_
port 40 nsew default input
rlabel metal3 s 49520 16328 50000 16448 6 right_width_0_height_0__pin_10_
port 41 nsew default input
rlabel metal3 s 49520 17824 50000 17944 6 right_width_0_height_0__pin_11_
port 42 nsew default input
rlabel metal3 s 49520 19456 50000 19576 6 right_width_0_height_0__pin_12_
port 43 nsew default input
rlabel metal3 s 49520 20952 50000 21072 6 right_width_0_height_0__pin_13_
port 44 nsew default input
rlabel metal3 s 49520 22584 50000 22704 6 right_width_0_height_0__pin_14_
port 45 nsew default input
rlabel metal3 s 49520 24080 50000 24200 6 right_width_0_height_0__pin_15_
port 46 nsew default input
rlabel metal3 s 49520 2184 50000 2304 6 right_width_0_height_0__pin_1_
port 47 nsew default input
rlabel metal3 s 49520 3816 50000 3936 6 right_width_0_height_0__pin_2_
port 48 nsew default input
rlabel metal3 s 49520 25712 50000 25832 6 right_width_0_height_0__pin_34_lower
port 49 nsew default tristate
rlabel metal3 s 49520 27208 50000 27328 6 right_width_0_height_0__pin_34_upper
port 50 nsew default tristate
rlabel metal3 s 49520 28840 50000 28960 6 right_width_0_height_0__pin_35_lower
port 51 nsew default tristate
rlabel metal3 s 49520 30336 50000 30456 6 right_width_0_height_0__pin_35_upper
port 52 nsew default tristate
rlabel metal3 s 49520 31968 50000 32088 6 right_width_0_height_0__pin_36_lower
port 53 nsew default tristate
rlabel metal3 s 49520 33464 50000 33584 6 right_width_0_height_0__pin_36_upper
port 54 nsew default tristate
rlabel metal3 s 49520 35096 50000 35216 6 right_width_0_height_0__pin_37_lower
port 55 nsew default tristate
rlabel metal3 s 49520 36592 50000 36712 6 right_width_0_height_0__pin_37_upper
port 56 nsew default tristate
rlabel metal3 s 49520 38224 50000 38344 6 right_width_0_height_0__pin_38_lower
port 57 nsew default tristate
rlabel metal3 s 49520 39720 50000 39840 6 right_width_0_height_0__pin_38_upper
port 58 nsew default tristate
rlabel metal3 s 49520 41352 50000 41472 6 right_width_0_height_0__pin_39_lower
port 59 nsew default tristate
rlabel metal3 s 49520 42848 50000 42968 6 right_width_0_height_0__pin_39_upper
port 60 nsew default tristate
rlabel metal3 s 49520 5312 50000 5432 6 right_width_0_height_0__pin_3_
port 61 nsew default input
rlabel metal3 s 49520 44480 50000 44600 6 right_width_0_height_0__pin_40_lower
port 62 nsew default tristate
rlabel metal3 s 49520 45976 50000 46096 6 right_width_0_height_0__pin_40_upper
port 63 nsew default tristate
rlabel metal3 s 49520 47608 50000 47728 6 right_width_0_height_0__pin_41_lower
port 64 nsew default tristate
rlabel metal3 s 49520 49104 50000 49224 6 right_width_0_height_0__pin_41_upper
port 65 nsew default tristate
rlabel metal3 s 49520 6944 50000 7064 6 right_width_0_height_0__pin_4_
port 66 nsew default input
rlabel metal3 s 49520 8440 50000 8560 6 right_width_0_height_0__pin_5_
port 67 nsew default input
rlabel metal3 s 49520 10072 50000 10192 6 right_width_0_height_0__pin_6_
port 68 nsew default input
rlabel metal3 s 49520 11568 50000 11688 6 right_width_0_height_0__pin_7_
port 69 nsew default input
rlabel metal3 s 49520 13200 50000 13320 6 right_width_0_height_0__pin_8_
port 70 nsew default input
rlabel metal3 s 49520 14696 50000 14816 6 right_width_0_height_0__pin_9_
port 71 nsew default input
rlabel metal2 s 8298 49520 8354 50000 6 top_width_0_height_0__pin_32_
port 72 nsew default input
rlabel metal2 s 24950 49520 25006 50000 6 top_width_0_height_0__pin_33_
port 73 nsew default input
rlabel metal4 s 4208 2128 4528 47376 6 vpwr
port 74 nsew default input
rlabel metal4 s 19568 2128 19888 47376 6 vgnd
port 75 nsew default input
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
