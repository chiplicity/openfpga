magic
tech EFS8A
magscale 1 2
timestamp 1602540333
<< locali >>
rect 222761 3995 222795 4165
rect 225337 3927 225371 4029
rect 218529 3451 218563 3553
<< viali >>
rect 215309 7497 215343 7531
rect 238125 7497 238159 7531
rect 239229 7497 239263 7531
rect 215125 7293 215159 7327
rect 237941 7293 237975 7327
rect 239045 7293 239079 7327
rect 404185 7293 404219 7327
rect 404737 7293 404771 7327
rect 239689 7225 239723 7259
rect 215769 7157 215803 7191
rect 238585 7157 238619 7191
rect 404369 7157 404403 7191
rect 219535 6885 219569 6919
rect 212825 6817 212859 6851
rect 215769 6817 215803 6851
rect 216229 6817 216263 6851
rect 215585 6749 215619 6783
rect 219173 6749 219207 6783
rect 220093 6681 220127 6715
rect 213009 6613 213043 6647
rect 215033 6409 215067 6443
rect 215309 6409 215343 6443
rect 238125 6409 238159 6443
rect 400045 6409 400079 6443
rect 216413 6341 216447 6375
rect 215493 6273 215527 6307
rect 215677 6205 215711 6239
rect 237481 6205 237515 6239
rect 237665 6205 237699 6239
rect 399493 6205 399527 6239
rect 399677 6205 399711 6239
rect 399861 6205 399895 6239
rect 219265 6137 219299 6171
rect 212917 6069 212951 6103
rect 216137 6069 216171 6103
rect 219633 6069 219667 6103
rect 237389 6069 237423 6103
rect 216229 5865 216263 5899
rect 220645 5865 220679 5899
rect 220046 5797 220080 5831
rect 234490 5797 234524 5831
rect 209329 5729 209363 5763
rect 215309 5729 215343 5763
rect 215493 5661 215527 5695
rect 219725 5661 219759 5695
rect 234169 5661 234203 5695
rect 209513 5525 209547 5559
rect 215953 5525 215987 5559
rect 220921 5525 220955 5559
rect 232421 5525 232455 5559
rect 235089 5525 235123 5559
rect 237481 5525 237515 5559
rect 399677 5525 399711 5559
rect 215309 5321 215343 5355
rect 233341 5321 233375 5355
rect 239137 5321 239171 5355
rect 290105 5321 290139 5355
rect 219449 5185 219483 5219
rect 221105 5185 221139 5219
rect 217609 5117 217643 5151
rect 220369 5117 220403 5151
rect 220553 5117 220587 5151
rect 221381 5117 221415 5151
rect 232421 5117 232455 5151
rect 238493 5117 238527 5151
rect 238677 5117 238711 5151
rect 289461 5117 289495 5151
rect 217517 5049 217551 5083
rect 217930 5049 217964 5083
rect 220737 5049 220771 5083
rect 232742 5049 232776 5083
rect 234169 5049 234203 5083
rect 209421 4981 209455 5015
rect 215769 4981 215803 5015
rect 218529 4981 218563 5015
rect 219817 4981 219851 5015
rect 220645 4981 220679 5015
rect 221841 4981 221875 5015
rect 232237 4981 232271 5015
rect 234537 4981 234571 5015
rect 238401 4981 238435 5015
rect 289645 4981 289679 5015
rect 219357 4777 219391 4811
rect 220645 4777 220679 4811
rect 218799 4709 218833 4743
rect 232650 4709 232684 4743
rect 213009 4641 213043 4675
rect 220553 4641 220587 4675
rect 221197 4641 221231 4675
rect 221381 4641 221415 4675
rect 221841 4641 221875 4675
rect 233249 4641 233283 4675
rect 238493 4641 238527 4675
rect 212365 4573 212399 4607
rect 212549 4573 212583 4607
rect 218437 4573 218471 4607
rect 232329 4573 232363 4607
rect 217701 4437 217735 4471
rect 218253 4437 218287 4471
rect 220461 4437 220495 4471
rect 223221 4437 223255 4471
rect 225797 4437 225831 4471
rect 212825 4233 212859 4267
rect 218161 4233 218195 4267
rect 219541 4233 219575 4267
rect 232329 4233 232363 4267
rect 232697 4233 232731 4267
rect 221473 4165 221507 4199
rect 222761 4165 222795 4199
rect 217793 4097 217827 4131
rect 220829 4097 220863 4131
rect 216413 4029 216447 4063
rect 218253 4029 218287 4063
rect 219173 4029 219207 4063
rect 222577 4029 222611 4063
rect 224601 4097 224635 4131
rect 226441 4097 226475 4131
rect 223129 4029 223163 4063
rect 223589 4029 223623 4063
rect 223957 4029 223991 4063
rect 224509 4029 224543 4063
rect 225337 4029 225371 4063
rect 225705 4029 225739 4063
rect 217057 3961 217091 3995
rect 218574 3961 218608 3995
rect 220093 3961 220127 3995
rect 220461 3961 220495 3995
rect 222761 3961 222795 3995
rect 225153 3961 225187 3995
rect 226073 3961 226107 3995
rect 212365 3893 212399 3927
rect 216137 3893 216171 3927
rect 219909 3893 219943 3927
rect 220277 3893 220311 3927
rect 220369 3893 220403 3927
rect 221105 3893 221139 3927
rect 221841 3893 221875 3927
rect 222209 3893 222243 3927
rect 222945 3893 222979 3927
rect 225337 3893 225371 3927
rect 225429 3893 225463 3927
rect 225889 3893 225923 3927
rect 225981 3893 226015 3927
rect 217701 3689 217735 3723
rect 218253 3689 218287 3723
rect 218713 3689 218747 3723
rect 223129 3689 223163 3723
rect 220369 3621 220403 3655
rect 221565 3621 221599 3655
rect 225153 3621 225187 3655
rect 225245 3621 225279 3655
rect 218529 3553 218563 3587
rect 218621 3553 218655 3587
rect 219081 3553 219115 3587
rect 219541 3553 219575 3587
rect 219817 3553 219851 3587
rect 221105 3553 221139 3587
rect 222945 3553 222979 3587
rect 225061 3553 225095 3587
rect 225613 3553 225647 3587
rect 220737 3485 220771 3519
rect 220921 3485 220955 3519
rect 223405 3485 223439 3519
rect 224877 3485 224911 3519
rect 218529 3417 218563 3451
rect 225889 3349 225923 3383
rect 219449 3145 219483 3179
rect 221473 3145 221507 3179
rect 224877 3145 224911 3179
rect 225245 3145 225279 3179
rect 224601 3077 224635 3111
rect 216873 3009 216907 3043
rect 220093 3009 220127 3043
rect 223037 3009 223071 3043
rect 217793 2941 217827 2975
rect 218161 2941 218195 2975
rect 218529 2941 218563 2975
rect 218989 2941 219023 2975
rect 219909 2941 219943 2975
rect 220461 2941 220495 2975
rect 217609 2873 217643 2907
rect 217241 2805 217275 2839
rect 217977 2805 218011 2839
rect 221105 2805 221139 2839
rect 208685 2601 208719 2635
rect 217793 2601 217827 2635
rect 219817 2601 219851 2635
rect 224877 2601 224911 2635
rect 218437 2533 218471 2567
rect 219449 2533 219483 2567
rect 208041 2465 208075 2499
rect 218345 2465 218379 2499
rect 218989 2465 219023 2499
rect 208225 2329 208259 2363
<< metal1 >>
rect 79778 8236 79784 8288
rect 79836 8276 79842 8288
rect 239214 8276 239220 8288
rect 79836 8248 239220 8276
rect 79836 8236 79842 8248
rect 239214 8236 239220 8248
rect 239272 8236 239278 8288
rect 106 7760 112 7812
rect 164 7800 170 7812
rect 215294 7800 215300 7812
rect 164 7772 215300 7800
rect 164 7760 170 7772
rect 215294 7760 215300 7772
rect 215352 7760 215358 7812
rect 14 7692 20 7744
rect 72 7732 78 7744
rect 215202 7732 215208 7744
rect 72 7704 215208 7732
rect 72 7692 78 7704
rect 215202 7692 215208 7704
rect 215260 7692 215266 7744
rect 1104 7642 422832 7664
rect 1104 7590 71648 7642
rect 71700 7590 71712 7642
rect 71764 7590 71776 7642
rect 71828 7590 71840 7642
rect 71892 7590 212982 7642
rect 213034 7590 213046 7642
rect 213098 7590 213110 7642
rect 213162 7590 213174 7642
rect 213226 7590 354315 7642
rect 354367 7590 354379 7642
rect 354431 7590 354443 7642
rect 354495 7590 354507 7642
rect 354559 7590 422832 7642
rect 1104 7568 422832 7590
rect 215294 7528 215300 7540
rect 215255 7500 215300 7528
rect 215294 7488 215300 7500
rect 215352 7488 215358 7540
rect 238113 7531 238171 7537
rect 238113 7497 238125 7531
rect 238159 7528 238171 7531
rect 238202 7528 238208 7540
rect 238159 7500 238208 7528
rect 238159 7497 238171 7500
rect 238113 7491 238171 7497
rect 238202 7488 238208 7500
rect 238260 7488 238266 7540
rect 239214 7528 239220 7540
rect 239175 7500 239220 7528
rect 239214 7488 239220 7500
rect 239272 7488 239278 7540
rect 215113 7327 215171 7333
rect 215113 7293 215125 7327
rect 215159 7324 215171 7327
rect 237929 7327 237987 7333
rect 215159 7296 215800 7324
rect 215159 7293 215171 7296
rect 215113 7287 215171 7293
rect 215772 7197 215800 7296
rect 237929 7293 237941 7327
rect 237975 7324 237987 7327
rect 239033 7327 239091 7333
rect 237975 7296 238616 7324
rect 237975 7293 237987 7296
rect 237929 7287 237987 7293
rect 238588 7200 238616 7296
rect 239033 7293 239045 7327
rect 239079 7324 239091 7327
rect 239122 7324 239128 7336
rect 239079 7296 239128 7324
rect 239079 7293 239091 7296
rect 239033 7287 239091 7293
rect 239122 7284 239128 7296
rect 239180 7324 239186 7336
rect 404170 7324 404176 7336
rect 239180 7296 239720 7324
rect 404131 7296 404176 7324
rect 239180 7284 239186 7296
rect 239692 7265 239720 7296
rect 404170 7284 404176 7296
rect 404228 7324 404234 7336
rect 404725 7327 404783 7333
rect 404725 7324 404737 7327
rect 404228 7296 404737 7324
rect 404228 7284 404234 7296
rect 404725 7293 404737 7296
rect 404771 7293 404783 7327
rect 404725 7287 404783 7293
rect 239677 7259 239735 7265
rect 239677 7225 239689 7259
rect 239723 7256 239735 7259
rect 423582 7256 423588 7268
rect 239723 7228 423588 7256
rect 239723 7225 239735 7228
rect 239677 7219 239735 7225
rect 423582 7216 423588 7228
rect 423640 7216 423646 7268
rect 215757 7191 215815 7197
rect 215757 7157 215769 7191
rect 215803 7188 215815 7191
rect 216214 7188 216220 7200
rect 215803 7160 216220 7188
rect 215803 7157 215815 7160
rect 215757 7151 215815 7157
rect 216214 7148 216220 7160
rect 216272 7148 216278 7200
rect 238570 7188 238576 7200
rect 238531 7160 238576 7188
rect 238570 7148 238576 7160
rect 238628 7148 238634 7200
rect 404357 7191 404415 7197
rect 404357 7157 404369 7191
rect 404403 7188 404415 7191
rect 423674 7188 423680 7200
rect 404403 7160 423680 7188
rect 404403 7157 404415 7160
rect 404357 7151 404415 7157
rect 423674 7148 423680 7160
rect 423732 7148 423738 7200
rect 1104 7098 422832 7120
rect 1104 7046 142315 7098
rect 142367 7046 142379 7098
rect 142431 7046 142443 7098
rect 142495 7046 142507 7098
rect 142559 7046 283648 7098
rect 283700 7046 283712 7098
rect 283764 7046 283776 7098
rect 283828 7046 283840 7098
rect 283892 7046 422832 7098
rect 1104 7024 422832 7046
rect 238570 6944 238576 6996
rect 238628 6984 238634 6996
rect 423490 6984 423496 6996
rect 238628 6956 423496 6984
rect 238628 6944 238634 6956
rect 423490 6944 423496 6956
rect 423548 6944 423554 6996
rect 219523 6919 219581 6925
rect 219523 6885 219535 6919
rect 219569 6916 219581 6919
rect 219802 6916 219808 6928
rect 219569 6888 219808 6916
rect 219569 6885 219581 6888
rect 219523 6879 219581 6885
rect 219802 6876 219808 6888
rect 219860 6876 219866 6928
rect 212810 6848 212816 6860
rect 212771 6820 212816 6848
rect 212810 6808 212816 6820
rect 212868 6808 212874 6860
rect 215018 6808 215024 6860
rect 215076 6848 215082 6860
rect 215757 6851 215815 6857
rect 215757 6848 215769 6851
rect 215076 6820 215769 6848
rect 215076 6808 215082 6820
rect 215757 6817 215769 6820
rect 215803 6817 215815 6851
rect 216214 6848 216220 6860
rect 216175 6820 216220 6848
rect 215757 6811 215815 6817
rect 215570 6780 215576 6792
rect 215531 6752 215576 6780
rect 215570 6740 215576 6752
rect 215628 6740 215634 6792
rect 215772 6712 215800 6811
rect 216214 6808 216220 6820
rect 216272 6808 216278 6860
rect 219161 6783 219219 6789
rect 219161 6749 219173 6783
rect 219207 6780 219219 6783
rect 219618 6780 219624 6792
rect 219207 6752 219624 6780
rect 219207 6749 219219 6752
rect 219161 6743 219219 6749
rect 219618 6740 219624 6752
rect 219676 6740 219682 6792
rect 220081 6715 220139 6721
rect 220081 6712 220093 6715
rect 215772 6684 220093 6712
rect 220081 6681 220093 6684
rect 220127 6681 220139 6715
rect 220081 6675 220139 6681
rect 202138 6604 202144 6656
rect 202196 6644 202202 6656
rect 212997 6647 213055 6653
rect 212997 6644 213009 6647
rect 202196 6616 213009 6644
rect 202196 6604 202202 6616
rect 212997 6613 213009 6616
rect 213043 6613 213055 6647
rect 212997 6607 213055 6613
rect 1104 6554 422832 6576
rect 1104 6502 71648 6554
rect 71700 6502 71712 6554
rect 71764 6502 71776 6554
rect 71828 6502 71840 6554
rect 71892 6502 212982 6554
rect 213034 6502 213046 6554
rect 213098 6502 213110 6554
rect 213162 6502 213174 6554
rect 213226 6502 354315 6554
rect 354367 6502 354379 6554
rect 354431 6502 354443 6554
rect 354495 6502 354507 6554
rect 354559 6502 422832 6554
rect 1104 6480 422832 6502
rect 215018 6440 215024 6452
rect 214979 6412 215024 6440
rect 215018 6400 215024 6412
rect 215076 6400 215082 6452
rect 215294 6440 215300 6452
rect 215255 6412 215300 6440
rect 215294 6400 215300 6412
rect 215352 6440 215358 6452
rect 238113 6443 238171 6449
rect 215352 6412 215524 6440
rect 215352 6400 215358 6412
rect 215496 6313 215524 6412
rect 238113 6409 238125 6443
rect 238159 6440 238171 6443
rect 238570 6440 238576 6452
rect 238159 6412 238576 6440
rect 238159 6409 238171 6412
rect 238113 6403 238171 6409
rect 238570 6400 238576 6412
rect 238628 6400 238634 6452
rect 397730 6400 397736 6452
rect 397788 6440 397794 6452
rect 400033 6443 400091 6449
rect 400033 6440 400045 6443
rect 397788 6412 400045 6440
rect 397788 6400 397794 6412
rect 400033 6409 400045 6412
rect 400079 6440 400091 6443
rect 404170 6440 404176 6452
rect 400079 6412 404176 6440
rect 400079 6409 400091 6412
rect 400033 6403 400091 6409
rect 404170 6400 404176 6412
rect 404228 6400 404234 6452
rect 215570 6332 215576 6384
rect 215628 6372 215634 6384
rect 216401 6375 216459 6381
rect 216401 6372 216413 6375
rect 215628 6344 216413 6372
rect 215628 6332 215634 6344
rect 216401 6341 216413 6344
rect 216447 6341 216459 6375
rect 216401 6335 216459 6341
rect 215481 6307 215539 6313
rect 215481 6273 215493 6307
rect 215527 6273 215539 6307
rect 215481 6267 215539 6273
rect 215665 6239 215723 6245
rect 215665 6205 215677 6239
rect 215711 6236 215723 6239
rect 216214 6236 216220 6248
rect 215711 6208 216220 6236
rect 215711 6205 215723 6208
rect 215665 6199 215723 6205
rect 216214 6196 216220 6208
rect 216272 6196 216278 6248
rect 237469 6239 237527 6245
rect 237469 6205 237481 6239
rect 237515 6205 237527 6239
rect 237469 6199 237527 6205
rect 219253 6171 219311 6177
rect 219253 6137 219265 6171
rect 219299 6168 219311 6171
rect 219802 6168 219808 6180
rect 219299 6140 219808 6168
rect 219299 6137 219311 6140
rect 219253 6131 219311 6137
rect 219802 6128 219808 6140
rect 219860 6128 219866 6180
rect 212810 6060 212816 6112
rect 212868 6100 212874 6112
rect 212905 6103 212963 6109
rect 212905 6100 212917 6103
rect 212868 6072 212917 6100
rect 212868 6060 212874 6072
rect 212905 6069 212917 6072
rect 212951 6100 212963 6103
rect 216122 6100 216128 6112
rect 212951 6072 216128 6100
rect 212951 6069 212963 6072
rect 212905 6063 212963 6069
rect 216122 6060 216128 6072
rect 216180 6060 216186 6112
rect 219618 6100 219624 6112
rect 219579 6072 219624 6100
rect 219618 6060 219624 6072
rect 219676 6060 219682 6112
rect 237374 6100 237380 6112
rect 237335 6072 237380 6100
rect 237374 6060 237380 6072
rect 237432 6100 237438 6112
rect 237484 6100 237512 6199
rect 237558 6196 237564 6248
rect 237616 6236 237622 6248
rect 237653 6239 237711 6245
rect 237653 6236 237665 6239
rect 237616 6208 237665 6236
rect 237616 6196 237622 6208
rect 237653 6205 237665 6208
rect 237699 6205 237711 6239
rect 237653 6199 237711 6205
rect 399481 6239 399539 6245
rect 399481 6205 399493 6239
rect 399527 6236 399539 6239
rect 399662 6236 399668 6248
rect 399527 6208 399668 6236
rect 399527 6205 399539 6208
rect 399481 6199 399539 6205
rect 399662 6196 399668 6208
rect 399720 6196 399726 6248
rect 399754 6196 399760 6248
rect 399812 6236 399818 6248
rect 399849 6239 399907 6245
rect 399849 6236 399861 6239
rect 399812 6208 399861 6236
rect 399812 6196 399818 6208
rect 399849 6205 399861 6208
rect 399895 6205 399907 6239
rect 399849 6199 399907 6205
rect 237432 6072 237512 6100
rect 237432 6060 237438 6072
rect 1104 6010 422832 6032
rect 1104 5958 142315 6010
rect 142367 5958 142379 6010
rect 142431 5958 142443 6010
rect 142495 5958 142507 6010
rect 142559 5958 283648 6010
rect 283700 5958 283712 6010
rect 283764 5958 283776 6010
rect 283828 5958 283840 6010
rect 283892 5958 422832 6010
rect 1104 5936 422832 5958
rect 216214 5896 216220 5908
rect 216175 5868 216220 5896
rect 216214 5856 216220 5868
rect 216272 5896 216278 5908
rect 220633 5899 220691 5905
rect 220633 5896 220645 5899
rect 216272 5868 220645 5896
rect 216272 5856 216278 5868
rect 220633 5865 220645 5868
rect 220679 5865 220691 5899
rect 220633 5859 220691 5865
rect 219802 5788 219808 5840
rect 219860 5828 219866 5840
rect 220034 5831 220092 5837
rect 220034 5828 220046 5831
rect 219860 5800 220046 5828
rect 219860 5788 219866 5800
rect 220034 5797 220046 5800
rect 220080 5797 220092 5831
rect 220034 5791 220092 5797
rect 234246 5788 234252 5840
rect 234304 5828 234310 5840
rect 234478 5831 234536 5837
rect 234478 5828 234490 5831
rect 234304 5800 234490 5828
rect 234304 5788 234310 5800
rect 234478 5797 234490 5800
rect 234524 5797 234536 5831
rect 234478 5791 234536 5797
rect 209314 5760 209320 5772
rect 209275 5732 209320 5760
rect 209314 5720 209320 5732
rect 209372 5720 209378 5772
rect 215202 5720 215208 5772
rect 215260 5760 215266 5772
rect 215297 5763 215355 5769
rect 215297 5760 215309 5763
rect 215260 5732 215309 5760
rect 215260 5720 215266 5732
rect 215297 5729 215309 5732
rect 215343 5729 215355 5763
rect 215297 5723 215355 5729
rect 215481 5695 215539 5701
rect 215481 5661 215493 5695
rect 215527 5692 215539 5695
rect 215754 5692 215760 5704
rect 215527 5664 215760 5692
rect 215527 5661 215539 5664
rect 215481 5655 215539 5661
rect 215754 5652 215760 5664
rect 215812 5652 215818 5704
rect 219710 5692 219716 5704
rect 219671 5664 219716 5692
rect 219710 5652 219716 5664
rect 219768 5652 219774 5704
rect 234157 5695 234215 5701
rect 234157 5661 234169 5695
rect 234203 5692 234215 5695
rect 234522 5692 234528 5704
rect 234203 5664 234528 5692
rect 234203 5661 234215 5664
rect 234157 5655 234215 5661
rect 234522 5652 234528 5664
rect 234580 5652 234586 5704
rect 209498 5556 209504 5568
rect 209459 5528 209504 5556
rect 209498 5516 209504 5528
rect 209556 5516 209562 5568
rect 215938 5556 215944 5568
rect 215899 5528 215944 5556
rect 215938 5516 215944 5528
rect 215996 5516 216002 5568
rect 220354 5516 220360 5568
rect 220412 5556 220418 5568
rect 220909 5559 220967 5565
rect 220909 5556 220921 5559
rect 220412 5528 220921 5556
rect 220412 5516 220418 5528
rect 220909 5525 220921 5528
rect 220955 5525 220967 5559
rect 232406 5556 232412 5568
rect 232367 5528 232412 5556
rect 220909 5519 220967 5525
rect 232406 5516 232412 5528
rect 232464 5516 232470 5568
rect 235074 5556 235080 5568
rect 235035 5528 235080 5556
rect 235074 5516 235080 5528
rect 235132 5516 235138 5568
rect 237466 5556 237472 5568
rect 237427 5528 237472 5556
rect 237466 5516 237472 5528
rect 237524 5516 237530 5568
rect 399662 5556 399668 5568
rect 399623 5528 399668 5556
rect 399662 5516 399668 5528
rect 399720 5516 399726 5568
rect 1104 5466 422832 5488
rect 1104 5414 71648 5466
rect 71700 5414 71712 5466
rect 71764 5414 71776 5466
rect 71828 5414 71840 5466
rect 71892 5414 212982 5466
rect 213034 5414 213046 5466
rect 213098 5414 213110 5466
rect 213162 5414 213174 5466
rect 213226 5414 354315 5466
rect 354367 5414 354379 5466
rect 354431 5414 354443 5466
rect 354495 5414 354507 5466
rect 354559 5414 422832 5466
rect 1104 5392 422832 5414
rect 215202 5312 215208 5364
rect 215260 5352 215266 5364
rect 215297 5355 215355 5361
rect 215297 5352 215309 5355
rect 215260 5324 215309 5352
rect 215260 5312 215266 5324
rect 215297 5321 215309 5324
rect 215343 5321 215355 5355
rect 215297 5315 215355 5321
rect 233329 5355 233387 5361
rect 233329 5321 233341 5355
rect 233375 5352 233387 5355
rect 237466 5352 237472 5364
rect 233375 5324 237472 5352
rect 233375 5321 233387 5324
rect 233329 5315 233387 5321
rect 237466 5312 237472 5324
rect 237524 5312 237530 5364
rect 239122 5352 239128 5364
rect 239083 5324 239128 5352
rect 239122 5312 239128 5324
rect 239180 5312 239186 5364
rect 290093 5355 290151 5361
rect 290093 5321 290105 5355
rect 290139 5352 290151 5355
rect 291102 5352 291108 5364
rect 290139 5324 291108 5352
rect 290139 5321 290151 5324
rect 290093 5315 290151 5321
rect 219437 5219 219495 5225
rect 219437 5185 219449 5219
rect 219483 5216 219495 5219
rect 219710 5216 219716 5228
rect 219483 5188 219716 5216
rect 219483 5185 219495 5188
rect 219437 5179 219495 5185
rect 219710 5176 219716 5188
rect 219768 5216 219774 5228
rect 221093 5219 221151 5225
rect 221093 5216 221105 5219
rect 219768 5188 221105 5216
rect 219768 5176 219774 5188
rect 221093 5185 221105 5188
rect 221139 5185 221151 5219
rect 221093 5179 221151 5185
rect 217597 5151 217655 5157
rect 217597 5117 217609 5151
rect 217643 5148 217655 5151
rect 217686 5148 217692 5160
rect 217643 5120 217692 5148
rect 217643 5117 217655 5120
rect 217597 5111 217655 5117
rect 217686 5108 217692 5120
rect 217744 5108 217750 5160
rect 220354 5148 220360 5160
rect 220315 5120 220360 5148
rect 220354 5108 220360 5120
rect 220412 5108 220418 5160
rect 220446 5108 220452 5160
rect 220504 5148 220510 5160
rect 220541 5151 220599 5157
rect 220541 5148 220553 5151
rect 220504 5120 220553 5148
rect 220504 5108 220510 5120
rect 220541 5117 220553 5120
rect 220587 5148 220599 5151
rect 221369 5151 221427 5157
rect 221369 5148 221381 5151
rect 220587 5120 221381 5148
rect 220587 5117 220599 5120
rect 220541 5111 220599 5117
rect 221369 5117 221381 5120
rect 221415 5117 221427 5151
rect 221369 5111 221427 5117
rect 226426 5108 226432 5160
rect 226484 5148 226490 5160
rect 232406 5148 232412 5160
rect 226484 5120 232412 5148
rect 226484 5108 226490 5120
rect 232406 5108 232412 5120
rect 232464 5108 232470 5160
rect 238481 5151 238539 5157
rect 238481 5117 238493 5151
rect 238527 5117 238539 5151
rect 238662 5148 238668 5160
rect 238623 5120 238668 5148
rect 238481 5111 238539 5117
rect 217502 5080 217508 5092
rect 217463 5052 217508 5080
rect 217502 5040 217508 5052
rect 217560 5080 217566 5092
rect 217918 5083 217976 5089
rect 217918 5080 217930 5083
rect 217560 5052 217930 5080
rect 217560 5040 217566 5052
rect 217918 5049 217930 5052
rect 217964 5049 217976 5083
rect 217918 5043 217976 5049
rect 220725 5083 220783 5089
rect 220725 5049 220737 5083
rect 220771 5080 220783 5083
rect 232730 5083 232788 5089
rect 232730 5080 232742 5083
rect 220771 5052 221872 5080
rect 220771 5049 220783 5052
rect 220725 5043 220783 5049
rect 221844 5024 221872 5052
rect 232240 5052 232742 5080
rect 232240 5024 232268 5052
rect 232730 5049 232742 5052
rect 232776 5080 232788 5083
rect 234157 5083 234215 5089
rect 234157 5080 234169 5083
rect 232776 5052 234169 5080
rect 232776 5049 232788 5052
rect 232730 5043 232788 5049
rect 234157 5049 234169 5052
rect 234203 5080 234215 5083
rect 234246 5080 234252 5092
rect 234203 5052 234252 5080
rect 234203 5049 234215 5052
rect 234157 5043 234215 5049
rect 234246 5040 234252 5052
rect 234304 5040 234310 5092
rect 209314 4972 209320 5024
rect 209372 5012 209378 5024
rect 209409 5015 209467 5021
rect 209409 5012 209421 5015
rect 209372 4984 209421 5012
rect 209372 4972 209378 4984
rect 209409 4981 209421 4984
rect 209455 5012 209467 5015
rect 212994 5012 213000 5024
rect 209455 4984 213000 5012
rect 209455 4981 209467 4984
rect 209409 4975 209467 4981
rect 212994 4972 213000 4984
rect 213052 4972 213058 5024
rect 215754 5012 215760 5024
rect 215715 4984 215760 5012
rect 215754 4972 215760 4984
rect 215812 4972 215818 5024
rect 217594 4972 217600 5024
rect 217652 5012 217658 5024
rect 218517 5015 218575 5021
rect 218517 5012 218529 5015
rect 217652 4984 218529 5012
rect 217652 4972 217658 4984
rect 218517 4981 218529 4984
rect 218563 4981 218575 5015
rect 219802 5012 219808 5024
rect 219763 4984 219808 5012
rect 218517 4975 218575 4981
rect 219802 4972 219808 4984
rect 219860 4972 219866 5024
rect 220630 5012 220636 5024
rect 220591 4984 220636 5012
rect 220630 4972 220636 4984
rect 220688 4972 220694 5024
rect 221826 5012 221832 5024
rect 221787 4984 221832 5012
rect 221826 4972 221832 4984
rect 221884 4972 221890 5024
rect 232222 5012 232228 5024
rect 232183 4984 232228 5012
rect 232222 4972 232228 4984
rect 232280 4972 232286 5024
rect 234522 5012 234528 5024
rect 234483 4984 234528 5012
rect 234522 4972 234528 4984
rect 234580 4972 234586 5024
rect 238386 5012 238392 5024
rect 238347 4984 238392 5012
rect 238386 4972 238392 4984
rect 238444 5012 238450 5024
rect 238496 5012 238524 5111
rect 238662 5108 238668 5120
rect 238720 5108 238726 5160
rect 289446 5148 289452 5160
rect 289359 5120 289452 5148
rect 289446 5108 289452 5120
rect 289504 5148 289510 5160
rect 290108 5148 290136 5315
rect 291102 5312 291108 5324
rect 291160 5312 291166 5364
rect 289504 5120 290136 5148
rect 289504 5108 289510 5120
rect 289630 5012 289636 5024
rect 238444 4984 238524 5012
rect 289591 4984 289636 5012
rect 238444 4972 238450 4984
rect 289630 4972 289636 4984
rect 289688 4972 289694 5024
rect 1104 4922 422832 4944
rect 1104 4870 142315 4922
rect 142367 4870 142379 4922
rect 142431 4870 142443 4922
rect 142495 4870 142507 4922
rect 142559 4870 283648 4922
rect 283700 4870 283712 4922
rect 283764 4870 283776 4922
rect 283828 4870 283840 4922
rect 283892 4870 422832 4922
rect 1104 4848 422832 4870
rect 215754 4768 215760 4820
rect 215812 4808 215818 4820
rect 219345 4811 219403 4817
rect 219345 4808 219357 4811
rect 215812 4780 219357 4808
rect 215812 4768 215818 4780
rect 219345 4777 219357 4780
rect 219391 4777 219403 4811
rect 219345 4771 219403 4777
rect 219618 4768 219624 4820
rect 219676 4808 219682 4820
rect 220633 4811 220691 4817
rect 220633 4808 220645 4811
rect 219676 4780 220645 4808
rect 219676 4768 219682 4780
rect 220633 4777 220645 4780
rect 220679 4777 220691 4811
rect 220633 4771 220691 4777
rect 217502 4700 217508 4752
rect 217560 4740 217566 4752
rect 218146 4740 218152 4752
rect 217560 4712 218152 4740
rect 217560 4700 217566 4712
rect 218146 4700 218152 4712
rect 218204 4740 218210 4752
rect 218787 4743 218845 4749
rect 218787 4740 218799 4743
rect 218204 4712 218799 4740
rect 218204 4700 218210 4712
rect 218787 4709 218799 4712
rect 218833 4740 218845 4743
rect 219802 4740 219808 4752
rect 218833 4712 219808 4740
rect 218833 4709 218845 4712
rect 218787 4703 218845 4709
rect 219802 4700 219808 4712
rect 219860 4700 219866 4752
rect 221918 4740 221924 4752
rect 221200 4712 221924 4740
rect 212994 4672 213000 4684
rect 212955 4644 213000 4672
rect 212994 4632 213000 4644
rect 213052 4632 213058 4684
rect 220354 4632 220360 4684
rect 220412 4672 220418 4684
rect 221200 4681 221228 4712
rect 221918 4700 221924 4712
rect 221976 4700 221982 4752
rect 232222 4700 232228 4752
rect 232280 4740 232286 4752
rect 232638 4743 232696 4749
rect 232638 4740 232650 4743
rect 232280 4712 232650 4740
rect 232280 4700 232286 4712
rect 232638 4709 232650 4712
rect 232684 4709 232696 4743
rect 232638 4703 232696 4709
rect 220541 4675 220599 4681
rect 220541 4672 220553 4675
rect 220412 4644 220553 4672
rect 220412 4632 220418 4644
rect 220541 4641 220553 4644
rect 220587 4641 220599 4675
rect 220541 4635 220599 4641
rect 221185 4675 221243 4681
rect 221185 4641 221197 4675
rect 221231 4641 221243 4675
rect 221366 4672 221372 4684
rect 221327 4644 221372 4672
rect 221185 4635 221243 4641
rect 221366 4632 221372 4644
rect 221424 4632 221430 4684
rect 221826 4672 221832 4684
rect 221787 4644 221832 4672
rect 221826 4632 221832 4644
rect 221884 4632 221890 4684
rect 233237 4675 233295 4681
rect 233237 4641 233249 4675
rect 233283 4672 233295 4675
rect 238481 4675 238539 4681
rect 238481 4672 238493 4675
rect 233283 4644 238493 4672
rect 233283 4641 233295 4644
rect 233237 4635 233295 4641
rect 238481 4641 238493 4644
rect 238527 4672 238539 4675
rect 238662 4672 238668 4684
rect 238527 4644 238668 4672
rect 238527 4641 238539 4644
rect 238481 4635 238539 4641
rect 238662 4632 238668 4644
rect 238720 4632 238726 4684
rect 212350 4604 212356 4616
rect 212311 4576 212356 4604
rect 212350 4564 212356 4576
rect 212408 4564 212414 4616
rect 212537 4607 212595 4613
rect 212537 4573 212549 4607
rect 212583 4604 212595 4607
rect 212810 4604 212816 4616
rect 212583 4576 212816 4604
rect 212583 4573 212595 4576
rect 212537 4567 212595 4573
rect 212810 4564 212816 4576
rect 212868 4604 212874 4616
rect 217594 4604 217600 4616
rect 212868 4576 217600 4604
rect 212868 4564 212874 4576
rect 217594 4564 217600 4576
rect 217652 4564 217658 4616
rect 218422 4604 218428 4616
rect 218383 4576 218428 4604
rect 218422 4564 218428 4576
rect 218480 4564 218486 4616
rect 224586 4564 224592 4616
rect 224644 4604 224650 4616
rect 232317 4607 232375 4613
rect 232317 4604 232329 4607
rect 224644 4576 232329 4604
rect 224644 4564 224650 4576
rect 232317 4573 232329 4576
rect 232363 4604 232375 4607
rect 232682 4604 232688 4616
rect 232363 4576 232688 4604
rect 232363 4573 232375 4576
rect 232317 4567 232375 4573
rect 232682 4564 232688 4576
rect 232740 4564 232746 4616
rect 217686 4468 217692 4480
rect 217647 4440 217692 4468
rect 217686 4428 217692 4440
rect 217744 4428 217750 4480
rect 217962 4428 217968 4480
rect 218020 4468 218026 4480
rect 218241 4471 218299 4477
rect 218241 4468 218253 4471
rect 218020 4440 218253 4468
rect 218020 4428 218026 4440
rect 218241 4437 218253 4440
rect 218287 4437 218299 4471
rect 218241 4431 218299 4437
rect 220449 4471 220507 4477
rect 220449 4437 220461 4471
rect 220495 4468 220507 4471
rect 220630 4468 220636 4480
rect 220495 4440 220636 4468
rect 220495 4437 220507 4440
rect 220449 4431 220507 4437
rect 220630 4428 220636 4440
rect 220688 4468 220694 4480
rect 221182 4468 221188 4480
rect 220688 4440 221188 4468
rect 220688 4428 220694 4440
rect 221182 4428 221188 4440
rect 221240 4428 221246 4480
rect 223206 4468 223212 4480
rect 223167 4440 223212 4468
rect 223206 4428 223212 4440
rect 223264 4468 223270 4480
rect 224494 4468 224500 4480
rect 223264 4440 224500 4468
rect 223264 4428 223270 4440
rect 224494 4428 224500 4440
rect 224552 4428 224558 4480
rect 225785 4471 225843 4477
rect 225785 4437 225797 4471
rect 225831 4468 225843 4471
rect 226150 4468 226156 4480
rect 225831 4440 226156 4468
rect 225831 4437 225843 4440
rect 225785 4431 225843 4437
rect 226150 4428 226156 4440
rect 226208 4428 226214 4480
rect 1104 4378 422832 4400
rect 1104 4326 71648 4378
rect 71700 4326 71712 4378
rect 71764 4326 71776 4378
rect 71828 4326 71840 4378
rect 71892 4326 212982 4378
rect 213034 4326 213046 4378
rect 213098 4326 213110 4378
rect 213162 4326 213174 4378
rect 213226 4326 354315 4378
rect 354367 4326 354379 4378
rect 354431 4326 354443 4378
rect 354495 4326 354507 4378
rect 354559 4326 422832 4378
rect 1104 4304 422832 4326
rect 212810 4264 212816 4276
rect 212771 4236 212816 4264
rect 212810 4224 212816 4236
rect 212868 4224 212874 4276
rect 218146 4264 218152 4276
rect 218107 4236 218152 4264
rect 218146 4224 218152 4236
rect 218204 4224 218210 4276
rect 219529 4267 219587 4273
rect 219529 4233 219541 4267
rect 219575 4264 219587 4267
rect 220446 4264 220452 4276
rect 219575 4236 220452 4264
rect 219575 4233 219587 4236
rect 219529 4227 219587 4233
rect 220446 4224 220452 4236
rect 220504 4224 220510 4276
rect 232222 4224 232228 4276
rect 232280 4264 232286 4276
rect 232317 4267 232375 4273
rect 232317 4264 232329 4267
rect 232280 4236 232329 4264
rect 232280 4224 232286 4236
rect 232317 4233 232329 4236
rect 232363 4233 232375 4267
rect 232682 4264 232688 4276
rect 232643 4236 232688 4264
rect 232317 4227 232375 4233
rect 232682 4224 232688 4236
rect 232740 4224 232746 4276
rect 220354 4156 220360 4208
rect 220412 4196 220418 4208
rect 221461 4199 221519 4205
rect 221461 4196 221473 4199
rect 220412 4168 221473 4196
rect 220412 4156 220418 4168
rect 221461 4165 221473 4168
rect 221507 4165 221519 4199
rect 221461 4159 221519 4165
rect 222749 4199 222807 4205
rect 222749 4165 222761 4199
rect 222795 4196 222807 4199
rect 222795 4168 225184 4196
rect 222795 4165 222807 4168
rect 222749 4159 222807 4165
rect 217781 4131 217839 4137
rect 217781 4097 217793 4131
rect 217827 4128 217839 4131
rect 218422 4128 218428 4140
rect 217827 4100 218428 4128
rect 217827 4097 217839 4100
rect 217781 4091 217839 4097
rect 218422 4088 218428 4100
rect 218480 4128 218486 4140
rect 220817 4131 220875 4137
rect 220817 4128 220829 4131
rect 218480 4100 220829 4128
rect 218480 4088 218486 4100
rect 220817 4097 220829 4100
rect 220863 4097 220875 4131
rect 224586 4128 224592 4140
rect 220817 4091 220875 4097
rect 222580 4100 223988 4128
rect 224547 4100 224592 4128
rect 222580 4072 222608 4100
rect 223960 4072 223988 4100
rect 224586 4088 224592 4100
rect 224644 4088 224650 4140
rect 216401 4063 216459 4069
rect 216401 4060 216413 4063
rect 216140 4032 216413 4060
rect 216140 3936 216168 4032
rect 216401 4029 216413 4032
rect 216447 4029 216459 4063
rect 216401 4023 216459 4029
rect 217962 4020 217968 4072
rect 218020 4060 218026 4072
rect 218241 4063 218299 4069
rect 218241 4060 218253 4063
rect 218020 4032 218253 4060
rect 218020 4020 218026 4032
rect 218241 4029 218253 4032
rect 218287 4029 218299 4063
rect 218241 4023 218299 4029
rect 219161 4063 219219 4069
rect 219161 4029 219173 4063
rect 219207 4060 219219 4063
rect 221090 4060 221096 4072
rect 219207 4032 221096 4060
rect 219207 4029 219219 4032
rect 219161 4023 219219 4029
rect 221090 4020 221096 4032
rect 221148 4020 221154 4072
rect 221366 4020 221372 4072
rect 221424 4060 221430 4072
rect 222562 4060 222568 4072
rect 221424 4032 222568 4060
rect 221424 4020 221430 4032
rect 222562 4020 222568 4032
rect 222620 4020 222626 4072
rect 223117 4063 223175 4069
rect 223117 4060 223129 4063
rect 222948 4032 223129 4060
rect 217042 3992 217048 4004
rect 217003 3964 217048 3992
rect 217042 3952 217048 3964
rect 217100 3952 217106 4004
rect 218146 3952 218152 4004
rect 218204 3992 218210 4004
rect 218562 3995 218620 4001
rect 218562 3992 218574 3995
rect 218204 3964 218574 3992
rect 218204 3952 218210 3964
rect 218562 3961 218574 3964
rect 218608 3961 218620 3995
rect 220078 3992 220084 4004
rect 220039 3964 220084 3992
rect 218562 3955 218620 3961
rect 220078 3952 220084 3964
rect 220136 3952 220142 4004
rect 220446 3992 220452 4004
rect 220359 3964 220452 3992
rect 220446 3952 220452 3964
rect 220504 3992 220510 4004
rect 222749 3995 222807 4001
rect 222749 3992 222761 3995
rect 220504 3964 222761 3992
rect 220504 3952 220510 3964
rect 222749 3961 222761 3964
rect 222795 3961 222807 3995
rect 222749 3955 222807 3961
rect 212350 3924 212356 3936
rect 212311 3896 212356 3924
rect 212350 3884 212356 3896
rect 212408 3884 212414 3936
rect 216122 3924 216128 3936
rect 216083 3896 216128 3924
rect 216122 3884 216128 3896
rect 216180 3884 216186 3936
rect 218974 3884 218980 3936
rect 219032 3924 219038 3936
rect 219897 3927 219955 3933
rect 219897 3924 219909 3927
rect 219032 3896 219909 3924
rect 219032 3884 219038 3896
rect 219897 3893 219909 3896
rect 219943 3924 219955 3927
rect 220262 3924 220268 3936
rect 219943 3896 220268 3924
rect 219943 3893 219955 3896
rect 219897 3887 219955 3893
rect 220262 3884 220268 3896
rect 220320 3884 220326 3936
rect 220354 3884 220360 3936
rect 220412 3924 220418 3936
rect 220412 3896 220457 3924
rect 220412 3884 220418 3896
rect 220998 3884 221004 3936
rect 221056 3924 221062 3936
rect 221093 3927 221151 3933
rect 221093 3924 221105 3927
rect 221056 3896 221105 3924
rect 221056 3884 221062 3896
rect 221093 3893 221105 3896
rect 221139 3924 221151 3927
rect 221366 3924 221372 3936
rect 221139 3896 221372 3924
rect 221139 3893 221151 3896
rect 221093 3887 221151 3893
rect 221366 3884 221372 3896
rect 221424 3884 221430 3936
rect 221826 3924 221832 3936
rect 221787 3896 221832 3924
rect 221826 3884 221832 3896
rect 221884 3884 221890 3936
rect 221918 3884 221924 3936
rect 221976 3924 221982 3936
rect 222197 3927 222255 3933
rect 222197 3924 222209 3927
rect 221976 3896 222209 3924
rect 221976 3884 221982 3896
rect 222197 3893 222209 3896
rect 222243 3893 222255 3927
rect 222197 3887 222255 3893
rect 222838 3884 222844 3936
rect 222896 3924 222902 3936
rect 222948 3933 222976 4032
rect 223117 4029 223129 4032
rect 223163 4029 223175 4063
rect 223574 4060 223580 4072
rect 223535 4032 223580 4060
rect 223117 4023 223175 4029
rect 223574 4020 223580 4032
rect 223632 4020 223638 4072
rect 223942 4060 223948 4072
rect 223855 4032 223948 4060
rect 223942 4020 223948 4032
rect 224000 4020 224006 4072
rect 224494 4060 224500 4072
rect 224407 4032 224500 4060
rect 224494 4020 224500 4032
rect 224552 4060 224558 4072
rect 225046 4060 225052 4072
rect 224552 4032 225052 4060
rect 224552 4020 224558 4032
rect 225046 4020 225052 4032
rect 225104 4020 225110 4072
rect 225156 4001 225184 4168
rect 226426 4128 226432 4140
rect 226387 4100 226432 4128
rect 226426 4088 226432 4100
rect 226484 4088 226490 4140
rect 225325 4063 225383 4069
rect 225325 4029 225337 4063
rect 225371 4060 225383 4063
rect 225693 4063 225751 4069
rect 225693 4060 225705 4063
rect 225371 4032 225705 4060
rect 225371 4029 225383 4032
rect 225325 4023 225383 4029
rect 225693 4029 225705 4032
rect 225739 4029 225751 4063
rect 225693 4023 225751 4029
rect 225141 3995 225199 4001
rect 225141 3961 225153 3995
rect 225187 3992 225199 3995
rect 225187 3964 225552 3992
rect 225187 3961 225199 3964
rect 225141 3955 225199 3961
rect 222933 3927 222991 3933
rect 222933 3924 222945 3927
rect 222896 3896 222945 3924
rect 222896 3884 222902 3896
rect 222933 3893 222945 3896
rect 222979 3893 222991 3927
rect 222933 3887 222991 3893
rect 224954 3884 224960 3936
rect 225012 3924 225018 3936
rect 225325 3927 225383 3933
rect 225325 3924 225337 3927
rect 225012 3896 225337 3924
rect 225012 3884 225018 3896
rect 225325 3893 225337 3896
rect 225371 3924 225383 3927
rect 225417 3927 225475 3933
rect 225417 3924 225429 3927
rect 225371 3896 225429 3924
rect 225371 3893 225383 3896
rect 225325 3887 225383 3893
rect 225417 3893 225429 3896
rect 225463 3893 225475 3927
rect 225524 3924 225552 3964
rect 225782 3952 225788 4004
rect 225840 3992 225846 4004
rect 226061 3995 226119 4001
rect 226061 3992 226073 3995
rect 225840 3964 226073 3992
rect 225840 3952 225846 3964
rect 226061 3961 226073 3964
rect 226107 3961 226119 3995
rect 226061 3955 226119 3961
rect 225874 3924 225880 3936
rect 225524 3896 225880 3924
rect 225417 3887 225475 3893
rect 225874 3884 225880 3896
rect 225932 3884 225938 3936
rect 225969 3927 226027 3933
rect 225969 3893 225981 3927
rect 226015 3924 226027 3927
rect 226150 3924 226156 3936
rect 226015 3896 226156 3924
rect 226015 3893 226027 3896
rect 225969 3887 226027 3893
rect 226150 3884 226156 3896
rect 226208 3884 226214 3936
rect 1104 3834 422832 3856
rect 1104 3782 142315 3834
rect 142367 3782 142379 3834
rect 142431 3782 142443 3834
rect 142495 3782 142507 3834
rect 142559 3782 283648 3834
rect 283700 3782 283712 3834
rect 283764 3782 283776 3834
rect 283828 3782 283840 3834
rect 283892 3782 422832 3834
rect 1104 3760 422832 3782
rect 217042 3680 217048 3732
rect 217100 3720 217106 3732
rect 217689 3723 217747 3729
rect 217689 3720 217701 3723
rect 217100 3692 217701 3720
rect 217100 3680 217106 3692
rect 217689 3689 217701 3692
rect 217735 3720 217747 3723
rect 217778 3720 217784 3732
rect 217735 3692 217784 3720
rect 217735 3689 217747 3692
rect 217689 3683 217747 3689
rect 217778 3680 217784 3692
rect 217836 3680 217842 3732
rect 218146 3680 218152 3732
rect 218204 3720 218210 3732
rect 218241 3723 218299 3729
rect 218241 3720 218253 3723
rect 218204 3692 218253 3720
rect 218204 3680 218210 3692
rect 218241 3689 218253 3692
rect 218287 3689 218299 3723
rect 218701 3723 218759 3729
rect 218701 3720 218713 3723
rect 218241 3683 218299 3689
rect 218348 3692 218713 3720
rect 217686 3544 217692 3596
rect 217744 3584 217750 3596
rect 218348 3584 218376 3692
rect 218701 3689 218713 3692
rect 218747 3689 218759 3723
rect 218701 3683 218759 3689
rect 219802 3680 219808 3732
rect 219860 3720 219866 3732
rect 221826 3720 221832 3732
rect 219860 3692 221832 3720
rect 219860 3680 219866 3692
rect 221826 3680 221832 3692
rect 221884 3680 221890 3732
rect 222562 3680 222568 3732
rect 222620 3720 222626 3732
rect 223117 3723 223175 3729
rect 223117 3720 223129 3723
rect 222620 3692 223129 3720
rect 222620 3680 222626 3692
rect 223117 3689 223129 3692
rect 223163 3689 223175 3723
rect 223117 3683 223175 3689
rect 220078 3652 220084 3664
rect 219544 3624 220084 3652
rect 219544 3596 219572 3624
rect 220078 3612 220084 3624
rect 220136 3652 220142 3664
rect 220357 3655 220415 3661
rect 220357 3652 220369 3655
rect 220136 3624 220369 3652
rect 220136 3612 220142 3624
rect 220357 3621 220369 3624
rect 220403 3652 220415 3655
rect 220998 3652 221004 3664
rect 220403 3624 221004 3652
rect 220403 3621 220415 3624
rect 220357 3615 220415 3621
rect 220998 3612 221004 3624
rect 221056 3612 221062 3664
rect 221553 3655 221611 3661
rect 221553 3621 221565 3655
rect 221599 3652 221611 3655
rect 224862 3652 224868 3664
rect 221599 3624 224868 3652
rect 221599 3621 221611 3624
rect 221553 3615 221611 3621
rect 224862 3612 224868 3624
rect 224920 3612 224926 3664
rect 224954 3612 224960 3664
rect 225012 3652 225018 3664
rect 225141 3655 225199 3661
rect 225141 3652 225153 3655
rect 225012 3624 225153 3652
rect 225012 3612 225018 3624
rect 225141 3621 225153 3624
rect 225187 3621 225199 3655
rect 225141 3615 225199 3621
rect 225233 3655 225291 3661
rect 225233 3621 225245 3655
rect 225279 3652 225291 3655
rect 225874 3652 225880 3664
rect 225279 3624 225880 3652
rect 225279 3621 225291 3624
rect 225233 3615 225291 3621
rect 225874 3612 225880 3624
rect 225932 3612 225938 3664
rect 217744 3556 218376 3584
rect 218517 3587 218575 3593
rect 217744 3544 217750 3556
rect 218517 3553 218529 3587
rect 218563 3584 218575 3587
rect 218609 3587 218667 3593
rect 218609 3584 218621 3587
rect 218563 3556 218621 3584
rect 218563 3553 218575 3556
rect 218517 3547 218575 3553
rect 218609 3553 218621 3556
rect 218655 3553 218667 3587
rect 219066 3584 219072 3596
rect 219027 3556 219072 3584
rect 218609 3547 218667 3553
rect 219066 3544 219072 3556
rect 219124 3544 219130 3596
rect 219526 3584 219532 3596
rect 219487 3556 219532 3584
rect 219526 3544 219532 3556
rect 219584 3544 219590 3596
rect 219802 3584 219808 3596
rect 219763 3556 219808 3584
rect 219802 3544 219808 3556
rect 219860 3544 219866 3596
rect 221090 3584 221096 3596
rect 221051 3556 221096 3584
rect 221090 3544 221096 3556
rect 221148 3544 221154 3596
rect 221182 3544 221188 3596
rect 221240 3584 221246 3596
rect 222930 3584 222936 3596
rect 221240 3556 222936 3584
rect 221240 3544 221246 3556
rect 222930 3544 222936 3556
rect 222988 3544 222994 3596
rect 225046 3584 225052 3596
rect 225007 3556 225052 3584
rect 225046 3544 225052 3556
rect 225104 3544 225110 3596
rect 225601 3587 225659 3593
rect 225601 3553 225613 3587
rect 225647 3584 225659 3587
rect 226058 3584 226064 3596
rect 225647 3556 226064 3584
rect 225647 3553 225659 3556
rect 225601 3547 225659 3553
rect 226058 3544 226064 3556
rect 226116 3544 226122 3596
rect 214006 3476 214012 3528
rect 214064 3516 214070 3528
rect 216122 3516 216128 3528
rect 214064 3488 216128 3516
rect 214064 3476 214070 3488
rect 216122 3476 216128 3488
rect 216180 3516 216186 3528
rect 216180 3488 216674 3516
rect 216180 3476 216186 3488
rect 216646 3448 216674 3488
rect 217778 3476 217784 3528
rect 217836 3516 217842 3528
rect 220354 3516 220360 3528
rect 217836 3488 220360 3516
rect 217836 3476 217842 3488
rect 220354 3476 220360 3488
rect 220412 3516 220418 3528
rect 220725 3519 220783 3525
rect 220725 3516 220737 3519
rect 220412 3488 220737 3516
rect 220412 3476 220418 3488
rect 220725 3485 220737 3488
rect 220771 3485 220783 3519
rect 220725 3479 220783 3485
rect 220909 3519 220967 3525
rect 220909 3485 220921 3519
rect 220955 3516 220967 3519
rect 220998 3516 221004 3528
rect 220955 3488 221004 3516
rect 220955 3485 220967 3488
rect 220909 3479 220967 3485
rect 220998 3476 221004 3488
rect 221056 3476 221062 3528
rect 221918 3476 221924 3528
rect 221976 3516 221982 3528
rect 223393 3519 223451 3525
rect 223393 3516 223405 3519
rect 221976 3488 223405 3516
rect 221976 3476 221982 3488
rect 223393 3485 223405 3488
rect 223439 3516 223451 3519
rect 223574 3516 223580 3528
rect 223439 3488 223580 3516
rect 223439 3485 223451 3488
rect 223393 3479 223451 3485
rect 223574 3476 223580 3488
rect 223632 3476 223638 3528
rect 223942 3476 223948 3528
rect 224000 3516 224006 3528
rect 224865 3519 224923 3525
rect 224865 3516 224877 3519
rect 224000 3488 224877 3516
rect 224000 3476 224006 3488
rect 224865 3485 224877 3488
rect 224911 3485 224923 3519
rect 224865 3479 224923 3485
rect 218517 3451 218575 3457
rect 218517 3448 218529 3451
rect 216646 3420 218529 3448
rect 218517 3417 218529 3420
rect 218563 3448 218575 3451
rect 219434 3448 219440 3460
rect 218563 3420 219440 3448
rect 218563 3417 218575 3420
rect 218517 3411 218575 3417
rect 219434 3408 219440 3420
rect 219492 3448 219498 3460
rect 222838 3448 222844 3460
rect 219492 3420 222844 3448
rect 219492 3408 219498 3420
rect 222838 3408 222844 3420
rect 222896 3408 222902 3460
rect 221826 3340 221832 3392
rect 221884 3380 221890 3392
rect 225782 3380 225788 3392
rect 221884 3352 225788 3380
rect 221884 3340 221890 3352
rect 225782 3340 225788 3352
rect 225840 3380 225846 3392
rect 225877 3383 225935 3389
rect 225877 3380 225889 3383
rect 225840 3352 225889 3380
rect 225840 3340 225846 3352
rect 225877 3349 225889 3352
rect 225923 3349 225935 3383
rect 225877 3343 225935 3349
rect 1104 3290 422832 3312
rect 1104 3238 71648 3290
rect 71700 3238 71712 3290
rect 71764 3238 71776 3290
rect 71828 3238 71840 3290
rect 71892 3238 212982 3290
rect 213034 3238 213046 3290
rect 213098 3238 213110 3290
rect 213162 3238 213174 3290
rect 213226 3238 354315 3290
rect 354367 3238 354379 3290
rect 354431 3238 354443 3290
rect 354495 3238 354507 3290
rect 354559 3238 422832 3290
rect 1104 3216 422832 3238
rect 219434 3176 219440 3188
rect 219395 3148 219440 3176
rect 219434 3136 219440 3148
rect 219492 3136 219498 3188
rect 221090 3136 221096 3188
rect 221148 3176 221154 3188
rect 221461 3179 221519 3185
rect 221461 3176 221473 3179
rect 221148 3148 221473 3176
rect 221148 3136 221154 3148
rect 221461 3145 221473 3148
rect 221507 3145 221519 3179
rect 221461 3139 221519 3145
rect 222838 3136 222844 3188
rect 222896 3176 222902 3188
rect 224865 3179 224923 3185
rect 224865 3176 224877 3179
rect 222896 3148 224877 3176
rect 222896 3136 222902 3148
rect 224865 3145 224877 3148
rect 224911 3176 224923 3179
rect 224954 3176 224960 3188
rect 224911 3148 224960 3176
rect 224911 3145 224923 3148
rect 224865 3139 224923 3145
rect 224954 3136 224960 3148
rect 225012 3136 225018 3188
rect 225046 3136 225052 3188
rect 225104 3176 225110 3188
rect 225233 3179 225291 3185
rect 225233 3176 225245 3179
rect 225104 3148 225245 3176
rect 225104 3136 225110 3148
rect 225233 3145 225245 3148
rect 225279 3145 225291 3179
rect 225233 3139 225291 3145
rect 224589 3111 224647 3117
rect 224589 3077 224601 3111
rect 224635 3108 224647 3111
rect 225874 3108 225880 3120
rect 224635 3080 225880 3108
rect 224635 3077 224647 3080
rect 224589 3071 224647 3077
rect 225874 3068 225880 3080
rect 225932 3068 225938 3120
rect 216861 3043 216919 3049
rect 216861 3009 216873 3043
rect 216907 3040 216919 3043
rect 219066 3040 219072 3052
rect 216907 3012 219072 3040
rect 216907 3009 216919 3012
rect 216861 3003 216919 3009
rect 217778 2972 217784 2984
rect 217739 2944 217784 2972
rect 217778 2932 217784 2944
rect 217836 2932 217842 2984
rect 218164 2981 218192 3012
rect 219066 3000 219072 3012
rect 219124 3040 219130 3052
rect 220081 3043 220139 3049
rect 220081 3040 220093 3043
rect 219124 3012 220093 3040
rect 219124 3000 219130 3012
rect 220081 3009 220093 3012
rect 220127 3040 220139 3043
rect 221918 3040 221924 3052
rect 220127 3012 221924 3040
rect 220127 3009 220139 3012
rect 220081 3003 220139 3009
rect 221918 3000 221924 3012
rect 221976 3000 221982 3052
rect 222930 3000 222936 3052
rect 222988 3040 222994 3052
rect 223025 3043 223083 3049
rect 223025 3040 223037 3043
rect 222988 3012 223037 3040
rect 222988 3000 222994 3012
rect 223025 3009 223037 3012
rect 223071 3040 223083 3043
rect 226150 3040 226156 3052
rect 223071 3012 226156 3040
rect 223071 3009 223083 3012
rect 223025 3003 223083 3009
rect 226150 3000 226156 3012
rect 226208 3000 226214 3052
rect 218149 2975 218207 2981
rect 218149 2941 218161 2975
rect 218195 2941 218207 2975
rect 218514 2972 218520 2984
rect 218475 2944 218520 2972
rect 218149 2935 218207 2941
rect 218514 2932 218520 2944
rect 218572 2932 218578 2984
rect 218974 2972 218980 2984
rect 218935 2944 218980 2972
rect 218974 2932 218980 2944
rect 219032 2932 219038 2984
rect 219897 2975 219955 2981
rect 219897 2941 219909 2975
rect 219943 2972 219955 2975
rect 220446 2972 220452 2984
rect 219943 2944 220452 2972
rect 219943 2941 219955 2944
rect 219897 2935 219955 2941
rect 220446 2932 220452 2944
rect 220504 2932 220510 2984
rect 217594 2904 217600 2916
rect 217507 2876 217600 2904
rect 217594 2864 217600 2876
rect 217652 2904 217658 2916
rect 218992 2904 219020 2932
rect 217652 2876 219020 2904
rect 217652 2864 217658 2876
rect 217226 2836 217232 2848
rect 217187 2808 217232 2836
rect 217226 2796 217232 2808
rect 217284 2796 217290 2848
rect 217962 2836 217968 2848
rect 217923 2808 217968 2836
rect 217962 2796 217968 2808
rect 218020 2796 218026 2848
rect 221090 2836 221096 2848
rect 221051 2808 221096 2836
rect 221090 2796 221096 2808
rect 221148 2796 221154 2848
rect 1104 2746 422832 2768
rect 1104 2694 142315 2746
rect 142367 2694 142379 2746
rect 142431 2694 142443 2746
rect 142495 2694 142507 2746
rect 142559 2694 283648 2746
rect 283700 2694 283712 2746
rect 283764 2694 283776 2746
rect 283828 2694 283840 2746
rect 283892 2694 422832 2746
rect 1104 2672 422832 2694
rect 208673 2635 208731 2641
rect 208673 2601 208685 2635
rect 208719 2632 208731 2635
rect 215938 2632 215944 2644
rect 208719 2604 215944 2632
rect 208719 2601 208731 2604
rect 208673 2595 208731 2601
rect 208029 2499 208087 2505
rect 208029 2465 208041 2499
rect 208075 2496 208087 2499
rect 208688 2496 208716 2595
rect 215938 2592 215944 2604
rect 215996 2592 216002 2644
rect 217781 2635 217839 2641
rect 217781 2601 217793 2635
rect 217827 2632 217839 2635
rect 218514 2632 218520 2644
rect 217827 2604 218520 2632
rect 217827 2601 217839 2604
rect 217781 2595 217839 2601
rect 218514 2592 218520 2604
rect 218572 2592 218578 2644
rect 219066 2592 219072 2644
rect 219124 2632 219130 2644
rect 219805 2635 219863 2641
rect 219805 2632 219817 2635
rect 219124 2604 219817 2632
rect 219124 2592 219130 2604
rect 219805 2601 219817 2604
rect 219851 2601 219863 2635
rect 219805 2595 219863 2601
rect 223942 2592 223948 2644
rect 224000 2632 224006 2644
rect 224865 2635 224923 2641
rect 224865 2632 224877 2635
rect 224000 2604 224877 2632
rect 224000 2592 224006 2604
rect 224865 2601 224877 2604
rect 224911 2601 224923 2635
rect 224865 2595 224923 2601
rect 217226 2524 217232 2576
rect 217284 2564 217290 2576
rect 218425 2567 218483 2573
rect 218425 2564 218437 2567
rect 217284 2536 218437 2564
rect 217284 2524 217290 2536
rect 208075 2468 208716 2496
rect 208075 2465 208087 2468
rect 208029 2459 208087 2465
rect 218256 2428 218284 2536
rect 218425 2533 218437 2536
rect 218471 2533 218483 2567
rect 218532 2564 218560 2592
rect 219437 2567 219495 2573
rect 219437 2564 219449 2567
rect 218532 2536 219449 2564
rect 218425 2527 218483 2533
rect 219437 2533 219449 2536
rect 219483 2564 219495 2567
rect 219526 2564 219532 2576
rect 219483 2536 219532 2564
rect 219483 2533 219495 2536
rect 219437 2527 219495 2533
rect 219526 2524 219532 2536
rect 219584 2524 219590 2576
rect 218333 2499 218391 2505
rect 218333 2465 218345 2499
rect 218379 2496 218391 2499
rect 218974 2496 218980 2508
rect 218379 2468 218980 2496
rect 218379 2465 218391 2468
rect 218333 2459 218391 2465
rect 218974 2456 218980 2468
rect 219032 2456 219038 2508
rect 219802 2428 219808 2440
rect 218256 2400 219808 2428
rect 219802 2388 219808 2400
rect 219860 2388 219866 2440
rect 208213 2363 208271 2369
rect 208213 2329 208225 2363
rect 208259 2360 208271 2363
rect 211614 2360 211620 2372
rect 208259 2332 211620 2360
rect 208259 2329 208271 2332
rect 208213 2323 208271 2329
rect 211614 2320 211620 2332
rect 211672 2320 211678 2372
rect 1104 2202 422832 2224
rect 1104 2150 71648 2202
rect 71700 2150 71712 2202
rect 71764 2150 71776 2202
rect 71828 2150 71840 2202
rect 71892 2150 212982 2202
rect 213034 2150 213046 2202
rect 213098 2150 213110 2202
rect 213162 2150 213174 2202
rect 213226 2150 354315 2202
rect 354367 2150 354379 2202
rect 354431 2150 354443 2202
rect 354495 2150 354507 2202
rect 354559 2150 422832 2202
rect 1104 2128 422832 2150
<< via1 >>
rect 79784 8236 79836 8288
rect 239220 8236 239272 8288
rect 112 7760 164 7812
rect 215300 7760 215352 7812
rect 20 7692 72 7744
rect 215208 7692 215260 7744
rect 71648 7590 71700 7642
rect 71712 7590 71764 7642
rect 71776 7590 71828 7642
rect 71840 7590 71892 7642
rect 212982 7590 213034 7642
rect 213046 7590 213098 7642
rect 213110 7590 213162 7642
rect 213174 7590 213226 7642
rect 354315 7590 354367 7642
rect 354379 7590 354431 7642
rect 354443 7590 354495 7642
rect 354507 7590 354559 7642
rect 215300 7531 215352 7540
rect 215300 7497 215309 7531
rect 215309 7497 215343 7531
rect 215343 7497 215352 7531
rect 215300 7488 215352 7497
rect 238208 7488 238260 7540
rect 239220 7531 239272 7540
rect 239220 7497 239229 7531
rect 239229 7497 239263 7531
rect 239263 7497 239272 7531
rect 239220 7488 239272 7497
rect 239128 7284 239180 7336
rect 404176 7327 404228 7336
rect 404176 7293 404185 7327
rect 404185 7293 404219 7327
rect 404219 7293 404228 7327
rect 404176 7284 404228 7293
rect 423588 7216 423640 7268
rect 216220 7148 216272 7200
rect 238576 7191 238628 7200
rect 238576 7157 238585 7191
rect 238585 7157 238619 7191
rect 238619 7157 238628 7191
rect 238576 7148 238628 7157
rect 423680 7148 423732 7200
rect 142315 7046 142367 7098
rect 142379 7046 142431 7098
rect 142443 7046 142495 7098
rect 142507 7046 142559 7098
rect 283648 7046 283700 7098
rect 283712 7046 283764 7098
rect 283776 7046 283828 7098
rect 283840 7046 283892 7098
rect 238576 6944 238628 6996
rect 423496 6944 423548 6996
rect 219808 6876 219860 6928
rect 212816 6851 212868 6860
rect 212816 6817 212825 6851
rect 212825 6817 212859 6851
rect 212859 6817 212868 6851
rect 212816 6808 212868 6817
rect 215024 6808 215076 6860
rect 216220 6851 216272 6860
rect 215576 6783 215628 6792
rect 215576 6749 215585 6783
rect 215585 6749 215619 6783
rect 215619 6749 215628 6783
rect 215576 6740 215628 6749
rect 216220 6817 216229 6851
rect 216229 6817 216263 6851
rect 216263 6817 216272 6851
rect 216220 6808 216272 6817
rect 219624 6740 219676 6792
rect 202144 6604 202196 6656
rect 71648 6502 71700 6554
rect 71712 6502 71764 6554
rect 71776 6502 71828 6554
rect 71840 6502 71892 6554
rect 212982 6502 213034 6554
rect 213046 6502 213098 6554
rect 213110 6502 213162 6554
rect 213174 6502 213226 6554
rect 354315 6502 354367 6554
rect 354379 6502 354431 6554
rect 354443 6502 354495 6554
rect 354507 6502 354559 6554
rect 215024 6443 215076 6452
rect 215024 6409 215033 6443
rect 215033 6409 215067 6443
rect 215067 6409 215076 6443
rect 215024 6400 215076 6409
rect 215300 6443 215352 6452
rect 215300 6409 215309 6443
rect 215309 6409 215343 6443
rect 215343 6409 215352 6443
rect 215300 6400 215352 6409
rect 238576 6400 238628 6452
rect 397736 6400 397788 6452
rect 404176 6400 404228 6452
rect 215576 6332 215628 6384
rect 216220 6196 216272 6248
rect 219808 6128 219860 6180
rect 212816 6060 212868 6112
rect 216128 6103 216180 6112
rect 216128 6069 216137 6103
rect 216137 6069 216171 6103
rect 216171 6069 216180 6103
rect 216128 6060 216180 6069
rect 219624 6103 219676 6112
rect 219624 6069 219633 6103
rect 219633 6069 219667 6103
rect 219667 6069 219676 6103
rect 219624 6060 219676 6069
rect 237380 6103 237432 6112
rect 237380 6069 237389 6103
rect 237389 6069 237423 6103
rect 237423 6069 237432 6103
rect 237564 6196 237616 6248
rect 399668 6239 399720 6248
rect 399668 6205 399677 6239
rect 399677 6205 399711 6239
rect 399711 6205 399720 6239
rect 399668 6196 399720 6205
rect 399760 6196 399812 6248
rect 237380 6060 237432 6069
rect 142315 5958 142367 6010
rect 142379 5958 142431 6010
rect 142443 5958 142495 6010
rect 142507 5958 142559 6010
rect 283648 5958 283700 6010
rect 283712 5958 283764 6010
rect 283776 5958 283828 6010
rect 283840 5958 283892 6010
rect 216220 5899 216272 5908
rect 216220 5865 216229 5899
rect 216229 5865 216263 5899
rect 216263 5865 216272 5899
rect 216220 5856 216272 5865
rect 219808 5788 219860 5840
rect 234252 5788 234304 5840
rect 209320 5763 209372 5772
rect 209320 5729 209329 5763
rect 209329 5729 209363 5763
rect 209363 5729 209372 5763
rect 209320 5720 209372 5729
rect 215208 5720 215260 5772
rect 215760 5652 215812 5704
rect 219716 5695 219768 5704
rect 219716 5661 219725 5695
rect 219725 5661 219759 5695
rect 219759 5661 219768 5695
rect 219716 5652 219768 5661
rect 234528 5652 234580 5704
rect 209504 5559 209556 5568
rect 209504 5525 209513 5559
rect 209513 5525 209547 5559
rect 209547 5525 209556 5559
rect 209504 5516 209556 5525
rect 215944 5559 215996 5568
rect 215944 5525 215953 5559
rect 215953 5525 215987 5559
rect 215987 5525 215996 5559
rect 215944 5516 215996 5525
rect 220360 5516 220412 5568
rect 232412 5559 232464 5568
rect 232412 5525 232421 5559
rect 232421 5525 232455 5559
rect 232455 5525 232464 5559
rect 232412 5516 232464 5525
rect 235080 5559 235132 5568
rect 235080 5525 235089 5559
rect 235089 5525 235123 5559
rect 235123 5525 235132 5559
rect 235080 5516 235132 5525
rect 237472 5559 237524 5568
rect 237472 5525 237481 5559
rect 237481 5525 237515 5559
rect 237515 5525 237524 5559
rect 237472 5516 237524 5525
rect 399668 5559 399720 5568
rect 399668 5525 399677 5559
rect 399677 5525 399711 5559
rect 399711 5525 399720 5559
rect 399668 5516 399720 5525
rect 71648 5414 71700 5466
rect 71712 5414 71764 5466
rect 71776 5414 71828 5466
rect 71840 5414 71892 5466
rect 212982 5414 213034 5466
rect 213046 5414 213098 5466
rect 213110 5414 213162 5466
rect 213174 5414 213226 5466
rect 354315 5414 354367 5466
rect 354379 5414 354431 5466
rect 354443 5414 354495 5466
rect 354507 5414 354559 5466
rect 215208 5312 215260 5364
rect 237472 5312 237524 5364
rect 239128 5355 239180 5364
rect 239128 5321 239137 5355
rect 239137 5321 239171 5355
rect 239171 5321 239180 5355
rect 239128 5312 239180 5321
rect 219716 5176 219768 5228
rect 217692 5108 217744 5160
rect 220360 5151 220412 5160
rect 220360 5117 220369 5151
rect 220369 5117 220403 5151
rect 220403 5117 220412 5151
rect 220360 5108 220412 5117
rect 220452 5108 220504 5160
rect 226432 5108 226484 5160
rect 232412 5151 232464 5160
rect 232412 5117 232421 5151
rect 232421 5117 232455 5151
rect 232455 5117 232464 5151
rect 232412 5108 232464 5117
rect 238668 5151 238720 5160
rect 217508 5083 217560 5092
rect 217508 5049 217517 5083
rect 217517 5049 217551 5083
rect 217551 5049 217560 5083
rect 217508 5040 217560 5049
rect 234252 5040 234304 5092
rect 209320 4972 209372 5024
rect 213000 4972 213052 5024
rect 215760 5015 215812 5024
rect 215760 4981 215769 5015
rect 215769 4981 215803 5015
rect 215803 4981 215812 5015
rect 215760 4972 215812 4981
rect 217600 4972 217652 5024
rect 219808 5015 219860 5024
rect 219808 4981 219817 5015
rect 219817 4981 219851 5015
rect 219851 4981 219860 5015
rect 219808 4972 219860 4981
rect 220636 5015 220688 5024
rect 220636 4981 220645 5015
rect 220645 4981 220679 5015
rect 220679 4981 220688 5015
rect 220636 4972 220688 4981
rect 221832 5015 221884 5024
rect 221832 4981 221841 5015
rect 221841 4981 221875 5015
rect 221875 4981 221884 5015
rect 221832 4972 221884 4981
rect 232228 5015 232280 5024
rect 232228 4981 232237 5015
rect 232237 4981 232271 5015
rect 232271 4981 232280 5015
rect 232228 4972 232280 4981
rect 234528 5015 234580 5024
rect 234528 4981 234537 5015
rect 234537 4981 234571 5015
rect 234571 4981 234580 5015
rect 234528 4972 234580 4981
rect 238392 5015 238444 5024
rect 238392 4981 238401 5015
rect 238401 4981 238435 5015
rect 238435 4981 238444 5015
rect 238668 5117 238677 5151
rect 238677 5117 238711 5151
rect 238711 5117 238720 5151
rect 238668 5108 238720 5117
rect 289452 5151 289504 5160
rect 289452 5117 289461 5151
rect 289461 5117 289495 5151
rect 289495 5117 289504 5151
rect 291108 5312 291160 5364
rect 289452 5108 289504 5117
rect 289636 5015 289688 5024
rect 238392 4972 238444 4981
rect 289636 4981 289645 5015
rect 289645 4981 289679 5015
rect 289679 4981 289688 5015
rect 289636 4972 289688 4981
rect 142315 4870 142367 4922
rect 142379 4870 142431 4922
rect 142443 4870 142495 4922
rect 142507 4870 142559 4922
rect 283648 4870 283700 4922
rect 283712 4870 283764 4922
rect 283776 4870 283828 4922
rect 283840 4870 283892 4922
rect 215760 4768 215812 4820
rect 219624 4768 219676 4820
rect 217508 4700 217560 4752
rect 218152 4700 218204 4752
rect 219808 4700 219860 4752
rect 213000 4675 213052 4684
rect 213000 4641 213009 4675
rect 213009 4641 213043 4675
rect 213043 4641 213052 4675
rect 213000 4632 213052 4641
rect 220360 4632 220412 4684
rect 221924 4700 221976 4752
rect 232228 4700 232280 4752
rect 221372 4675 221424 4684
rect 221372 4641 221381 4675
rect 221381 4641 221415 4675
rect 221415 4641 221424 4675
rect 221372 4632 221424 4641
rect 221832 4675 221884 4684
rect 221832 4641 221841 4675
rect 221841 4641 221875 4675
rect 221875 4641 221884 4675
rect 221832 4632 221884 4641
rect 238668 4632 238720 4684
rect 212356 4607 212408 4616
rect 212356 4573 212365 4607
rect 212365 4573 212399 4607
rect 212399 4573 212408 4607
rect 212356 4564 212408 4573
rect 212816 4564 212868 4616
rect 217600 4564 217652 4616
rect 218428 4607 218480 4616
rect 218428 4573 218437 4607
rect 218437 4573 218471 4607
rect 218471 4573 218480 4607
rect 218428 4564 218480 4573
rect 224592 4564 224644 4616
rect 232688 4564 232740 4616
rect 217692 4471 217744 4480
rect 217692 4437 217701 4471
rect 217701 4437 217735 4471
rect 217735 4437 217744 4471
rect 217692 4428 217744 4437
rect 217968 4428 218020 4480
rect 220636 4428 220688 4480
rect 221188 4428 221240 4480
rect 223212 4471 223264 4480
rect 223212 4437 223221 4471
rect 223221 4437 223255 4471
rect 223255 4437 223264 4471
rect 223212 4428 223264 4437
rect 224500 4428 224552 4480
rect 226156 4428 226208 4480
rect 71648 4326 71700 4378
rect 71712 4326 71764 4378
rect 71776 4326 71828 4378
rect 71840 4326 71892 4378
rect 212982 4326 213034 4378
rect 213046 4326 213098 4378
rect 213110 4326 213162 4378
rect 213174 4326 213226 4378
rect 354315 4326 354367 4378
rect 354379 4326 354431 4378
rect 354443 4326 354495 4378
rect 354507 4326 354559 4378
rect 212816 4267 212868 4276
rect 212816 4233 212825 4267
rect 212825 4233 212859 4267
rect 212859 4233 212868 4267
rect 212816 4224 212868 4233
rect 218152 4267 218204 4276
rect 218152 4233 218161 4267
rect 218161 4233 218195 4267
rect 218195 4233 218204 4267
rect 218152 4224 218204 4233
rect 220452 4224 220504 4276
rect 232228 4224 232280 4276
rect 232688 4267 232740 4276
rect 232688 4233 232697 4267
rect 232697 4233 232731 4267
rect 232731 4233 232740 4267
rect 232688 4224 232740 4233
rect 220360 4156 220412 4208
rect 218428 4088 218480 4140
rect 224592 4131 224644 4140
rect 224592 4097 224601 4131
rect 224601 4097 224635 4131
rect 224635 4097 224644 4131
rect 224592 4088 224644 4097
rect 217968 4020 218020 4072
rect 221096 4020 221148 4072
rect 221372 4020 221424 4072
rect 222568 4063 222620 4072
rect 222568 4029 222577 4063
rect 222577 4029 222611 4063
rect 222611 4029 222620 4063
rect 222568 4020 222620 4029
rect 217048 3995 217100 4004
rect 217048 3961 217057 3995
rect 217057 3961 217091 3995
rect 217091 3961 217100 3995
rect 217048 3952 217100 3961
rect 218152 3952 218204 4004
rect 220084 3995 220136 4004
rect 220084 3961 220093 3995
rect 220093 3961 220127 3995
rect 220127 3961 220136 3995
rect 220084 3952 220136 3961
rect 220452 3995 220504 4004
rect 220452 3961 220461 3995
rect 220461 3961 220495 3995
rect 220495 3961 220504 3995
rect 220452 3952 220504 3961
rect 212356 3927 212408 3936
rect 212356 3893 212365 3927
rect 212365 3893 212399 3927
rect 212399 3893 212408 3927
rect 212356 3884 212408 3893
rect 216128 3927 216180 3936
rect 216128 3893 216137 3927
rect 216137 3893 216171 3927
rect 216171 3893 216180 3927
rect 216128 3884 216180 3893
rect 218980 3884 219032 3936
rect 220268 3927 220320 3936
rect 220268 3893 220277 3927
rect 220277 3893 220311 3927
rect 220311 3893 220320 3927
rect 220268 3884 220320 3893
rect 220360 3927 220412 3936
rect 220360 3893 220369 3927
rect 220369 3893 220403 3927
rect 220403 3893 220412 3927
rect 220360 3884 220412 3893
rect 221004 3884 221056 3936
rect 221372 3884 221424 3936
rect 221832 3927 221884 3936
rect 221832 3893 221841 3927
rect 221841 3893 221875 3927
rect 221875 3893 221884 3927
rect 221832 3884 221884 3893
rect 221924 3884 221976 3936
rect 222844 3884 222896 3936
rect 223580 4063 223632 4072
rect 223580 4029 223589 4063
rect 223589 4029 223623 4063
rect 223623 4029 223632 4063
rect 223580 4020 223632 4029
rect 223948 4063 224000 4072
rect 223948 4029 223957 4063
rect 223957 4029 223991 4063
rect 223991 4029 224000 4063
rect 223948 4020 224000 4029
rect 224500 4063 224552 4072
rect 224500 4029 224509 4063
rect 224509 4029 224543 4063
rect 224543 4029 224552 4063
rect 224500 4020 224552 4029
rect 225052 4020 225104 4072
rect 226432 4131 226484 4140
rect 226432 4097 226441 4131
rect 226441 4097 226475 4131
rect 226475 4097 226484 4131
rect 226432 4088 226484 4097
rect 224960 3884 225012 3936
rect 225788 3952 225840 4004
rect 225880 3927 225932 3936
rect 225880 3893 225889 3927
rect 225889 3893 225923 3927
rect 225923 3893 225932 3927
rect 225880 3884 225932 3893
rect 226156 3884 226208 3936
rect 142315 3782 142367 3834
rect 142379 3782 142431 3834
rect 142443 3782 142495 3834
rect 142507 3782 142559 3834
rect 283648 3782 283700 3834
rect 283712 3782 283764 3834
rect 283776 3782 283828 3834
rect 283840 3782 283892 3834
rect 217048 3680 217100 3732
rect 217784 3680 217836 3732
rect 218152 3680 218204 3732
rect 217692 3544 217744 3596
rect 219808 3680 219860 3732
rect 221832 3680 221884 3732
rect 222568 3680 222620 3732
rect 220084 3612 220136 3664
rect 221004 3612 221056 3664
rect 224868 3612 224920 3664
rect 224960 3612 225012 3664
rect 225880 3612 225932 3664
rect 219072 3587 219124 3596
rect 219072 3553 219081 3587
rect 219081 3553 219115 3587
rect 219115 3553 219124 3587
rect 219072 3544 219124 3553
rect 219532 3587 219584 3596
rect 219532 3553 219541 3587
rect 219541 3553 219575 3587
rect 219575 3553 219584 3587
rect 219532 3544 219584 3553
rect 219808 3587 219860 3596
rect 219808 3553 219817 3587
rect 219817 3553 219851 3587
rect 219851 3553 219860 3587
rect 219808 3544 219860 3553
rect 221096 3587 221148 3596
rect 221096 3553 221105 3587
rect 221105 3553 221139 3587
rect 221139 3553 221148 3587
rect 221096 3544 221148 3553
rect 221188 3544 221240 3596
rect 222936 3587 222988 3596
rect 222936 3553 222945 3587
rect 222945 3553 222979 3587
rect 222979 3553 222988 3587
rect 222936 3544 222988 3553
rect 225052 3587 225104 3596
rect 225052 3553 225061 3587
rect 225061 3553 225095 3587
rect 225095 3553 225104 3587
rect 225052 3544 225104 3553
rect 226064 3544 226116 3596
rect 214012 3476 214064 3528
rect 216128 3476 216180 3528
rect 217784 3476 217836 3528
rect 220360 3476 220412 3528
rect 221004 3476 221056 3528
rect 221924 3476 221976 3528
rect 223580 3476 223632 3528
rect 223948 3476 224000 3528
rect 219440 3408 219492 3460
rect 222844 3408 222896 3460
rect 221832 3340 221884 3392
rect 225788 3340 225840 3392
rect 71648 3238 71700 3290
rect 71712 3238 71764 3290
rect 71776 3238 71828 3290
rect 71840 3238 71892 3290
rect 212982 3238 213034 3290
rect 213046 3238 213098 3290
rect 213110 3238 213162 3290
rect 213174 3238 213226 3290
rect 354315 3238 354367 3290
rect 354379 3238 354431 3290
rect 354443 3238 354495 3290
rect 354507 3238 354559 3290
rect 219440 3179 219492 3188
rect 219440 3145 219449 3179
rect 219449 3145 219483 3179
rect 219483 3145 219492 3179
rect 219440 3136 219492 3145
rect 221096 3136 221148 3188
rect 222844 3136 222896 3188
rect 224960 3136 225012 3188
rect 225052 3136 225104 3188
rect 225880 3068 225932 3120
rect 217784 2975 217836 2984
rect 217784 2941 217793 2975
rect 217793 2941 217827 2975
rect 217827 2941 217836 2975
rect 217784 2932 217836 2941
rect 219072 3000 219124 3052
rect 221924 3000 221976 3052
rect 222936 3000 222988 3052
rect 226156 3000 226208 3052
rect 218520 2975 218572 2984
rect 218520 2941 218529 2975
rect 218529 2941 218563 2975
rect 218563 2941 218572 2975
rect 218520 2932 218572 2941
rect 218980 2975 219032 2984
rect 218980 2941 218989 2975
rect 218989 2941 219023 2975
rect 219023 2941 219032 2975
rect 218980 2932 219032 2941
rect 220452 2975 220504 2984
rect 220452 2941 220461 2975
rect 220461 2941 220495 2975
rect 220495 2941 220504 2975
rect 220452 2932 220504 2941
rect 217600 2907 217652 2916
rect 217600 2873 217609 2907
rect 217609 2873 217643 2907
rect 217643 2873 217652 2907
rect 217600 2864 217652 2873
rect 217232 2839 217284 2848
rect 217232 2805 217241 2839
rect 217241 2805 217275 2839
rect 217275 2805 217284 2839
rect 217232 2796 217284 2805
rect 217968 2839 218020 2848
rect 217968 2805 217977 2839
rect 217977 2805 218011 2839
rect 218011 2805 218020 2839
rect 217968 2796 218020 2805
rect 221096 2839 221148 2848
rect 221096 2805 221105 2839
rect 221105 2805 221139 2839
rect 221139 2805 221148 2839
rect 221096 2796 221148 2805
rect 142315 2694 142367 2746
rect 142379 2694 142431 2746
rect 142443 2694 142495 2746
rect 142507 2694 142559 2746
rect 283648 2694 283700 2746
rect 283712 2694 283764 2746
rect 283776 2694 283828 2746
rect 283840 2694 283892 2746
rect 215944 2592 215996 2644
rect 218520 2592 218572 2644
rect 219072 2592 219124 2644
rect 223948 2592 224000 2644
rect 217232 2524 217284 2576
rect 219532 2524 219584 2576
rect 218980 2499 219032 2508
rect 218980 2465 218989 2499
rect 218989 2465 219023 2499
rect 219023 2465 219032 2499
rect 218980 2456 219032 2465
rect 219808 2388 219860 2440
rect 211620 2320 211672 2372
rect 71648 2150 71700 2202
rect 71712 2150 71764 2202
rect 71776 2150 71828 2202
rect 71840 2150 71892 2202
rect 212982 2150 213034 2202
rect 213046 2150 213098 2202
rect 213110 2150 213162 2202
rect 213174 2150 213226 2202
rect 354315 2150 354367 2202
rect 354379 2150 354431 2202
rect 354443 2150 354495 2202
rect 354507 2150 354559 2202
<< metal2 >>
rect 26514 9520 26570 10000
rect 79506 9602 79562 10000
rect 132498 9602 132554 10000
rect 185490 9602 185546 10000
rect 238482 9602 238538 10000
rect 291474 9602 291530 10000
rect 79506 9574 79824 9602
rect 79506 9520 79562 9574
rect 18 9208 74 9217
rect 18 9143 74 9152
rect 32 7750 60 9143
rect 79796 8294 79824 9574
rect 132498 9574 132816 9602
rect 132498 9520 132554 9574
rect 79784 8288 79836 8294
rect 79784 8230 79836 8236
rect 112 7812 164 7818
rect 112 7754 164 7760
rect 20 7744 72 7750
rect 20 7686 72 7692
rect 124 7585 152 7754
rect 71622 7644 71918 7664
rect 71678 7642 71702 7644
rect 71758 7642 71782 7644
rect 71838 7642 71862 7644
rect 71700 7590 71702 7642
rect 71764 7590 71776 7642
rect 71838 7590 71840 7642
rect 71678 7588 71702 7590
rect 71758 7588 71782 7590
rect 71838 7588 71862 7590
rect 110 7576 166 7585
rect 71622 7568 71918 7588
rect 110 7511 166 7520
rect 132788 6905 132816 9574
rect 185490 9574 185808 9602
rect 185490 9520 185546 9574
rect 142289 7100 142585 7120
rect 142345 7098 142369 7100
rect 142425 7098 142449 7100
rect 142505 7098 142529 7100
rect 142367 7046 142369 7098
rect 142431 7046 142443 7098
rect 142505 7046 142507 7098
rect 142345 7044 142369 7046
rect 142425 7044 142449 7046
rect 142505 7044 142529 7046
rect 142289 7024 142585 7044
rect 132774 6896 132830 6905
rect 132774 6831 132830 6840
rect 185780 6769 185808 9574
rect 238220 9574 238538 9602
rect 215300 7812 215352 7818
rect 215300 7754 215352 7760
rect 215208 7744 215260 7750
rect 215208 7686 215260 7692
rect 212956 7644 213252 7664
rect 213012 7642 213036 7644
rect 213092 7642 213116 7644
rect 213172 7642 213196 7644
rect 213034 7590 213036 7642
rect 213098 7590 213110 7642
rect 213172 7590 213174 7642
rect 213012 7588 213036 7590
rect 213092 7588 213116 7590
rect 213172 7588 213196 7590
rect 212956 7568 213252 7588
rect 212816 6860 212868 6866
rect 212816 6802 212868 6808
rect 215024 6860 215076 6866
rect 215024 6802 215076 6808
rect 185766 6760 185822 6769
rect 185766 6695 185822 6704
rect 202142 6760 202198 6769
rect 202142 6695 202198 6704
rect 202156 6662 202184 6695
rect 202144 6656 202196 6662
rect 202144 6598 202196 6604
rect 71622 6556 71918 6576
rect 71678 6554 71702 6556
rect 71758 6554 71782 6556
rect 71838 6554 71862 6556
rect 71700 6502 71702 6554
rect 71764 6502 71776 6554
rect 71838 6502 71840 6554
rect 71678 6500 71702 6502
rect 71758 6500 71782 6502
rect 71838 6500 71862 6502
rect 71622 6480 71918 6500
rect 212828 6118 212856 6802
rect 212956 6556 213252 6576
rect 213012 6554 213036 6556
rect 213092 6554 213116 6556
rect 213172 6554 213196 6556
rect 213034 6502 213036 6554
rect 213098 6502 213110 6554
rect 213172 6502 213174 6554
rect 213012 6500 213036 6502
rect 213092 6500 213116 6502
rect 213172 6500 213196 6502
rect 212956 6480 213252 6500
rect 215036 6458 215064 6802
rect 215024 6452 215076 6458
rect 215024 6394 215076 6400
rect 212816 6112 212868 6118
rect 212816 6054 212868 6060
rect 142289 6012 142585 6032
rect 142345 6010 142369 6012
rect 142425 6010 142449 6012
rect 142505 6010 142529 6012
rect 142367 5958 142369 6010
rect 142431 5958 142443 6010
rect 142505 5958 142507 6010
rect 142345 5956 142369 5958
rect 142425 5956 142449 5958
rect 142505 5956 142529 5958
rect 142289 5936 142585 5956
rect 215220 5778 215248 7686
rect 215312 7546 215340 7754
rect 238220 7546 238248 9574
rect 238482 9520 238538 9574
rect 291120 9574 291530 9602
rect 239220 8288 239272 8294
rect 239220 8230 239272 8236
rect 239232 7546 239260 8230
rect 215300 7540 215352 7546
rect 215300 7482 215352 7488
rect 238208 7540 238260 7546
rect 238208 7482 238260 7488
rect 239220 7540 239272 7546
rect 239220 7482 239272 7488
rect 239128 7336 239180 7342
rect 239128 7278 239180 7284
rect 216220 7200 216272 7206
rect 216220 7142 216272 7148
rect 238576 7200 238628 7206
rect 238576 7142 238628 7148
rect 215298 6896 215354 6905
rect 216232 6866 216260 7142
rect 238588 7002 238616 7142
rect 238576 6996 238628 7002
rect 238576 6938 238628 6944
rect 219808 6928 219860 6934
rect 219808 6870 219860 6876
rect 215298 6831 215354 6840
rect 216220 6860 216272 6866
rect 215312 6458 215340 6831
rect 216220 6802 216272 6808
rect 215576 6792 215628 6798
rect 216232 6769 216260 6802
rect 219624 6792 219676 6798
rect 215576 6734 215628 6740
rect 216218 6760 216274 6769
rect 215300 6452 215352 6458
rect 215300 6394 215352 6400
rect 215588 6390 215616 6734
rect 219624 6734 219676 6740
rect 216218 6695 216274 6704
rect 215576 6384 215628 6390
rect 215576 6326 215628 6332
rect 215588 6225 215616 6326
rect 216220 6248 216272 6254
rect 215574 6216 215630 6225
rect 216220 6190 216272 6196
rect 215574 6151 215630 6160
rect 216128 6112 216180 6118
rect 216128 6054 216180 6060
rect 209320 5772 209372 5778
rect 209320 5714 209372 5720
rect 215208 5772 215260 5778
rect 215208 5714 215260 5720
rect 71622 5468 71918 5488
rect 71678 5466 71702 5468
rect 71758 5466 71782 5468
rect 71838 5466 71862 5468
rect 71700 5414 71702 5466
rect 71764 5414 71776 5466
rect 71838 5414 71840 5466
rect 71678 5412 71702 5414
rect 71758 5412 71782 5414
rect 71838 5412 71862 5414
rect 71622 5392 71918 5412
rect 110 5264 166 5273
rect 110 5199 166 5208
rect 124 4185 152 5199
rect 209332 5030 209360 5714
rect 209504 5568 209556 5574
rect 209504 5510 209556 5516
rect 209516 5273 209544 5510
rect 212956 5468 213252 5488
rect 213012 5466 213036 5468
rect 213092 5466 213116 5468
rect 213172 5466 213196 5468
rect 213034 5414 213036 5466
rect 213098 5414 213110 5466
rect 213172 5414 213174 5466
rect 213012 5412 213036 5414
rect 213092 5412 213116 5414
rect 213172 5412 213196 5414
rect 212956 5392 213252 5412
rect 215220 5370 215248 5714
rect 215760 5704 215812 5710
rect 215760 5646 215812 5652
rect 215208 5364 215260 5370
rect 215208 5306 215260 5312
rect 209502 5264 209558 5273
rect 209502 5199 209558 5208
rect 215772 5030 215800 5646
rect 215944 5568 215996 5574
rect 215944 5510 215996 5516
rect 209320 5024 209372 5030
rect 209320 4966 209372 4972
rect 213000 5024 213052 5030
rect 213000 4966 213052 4972
rect 215760 5024 215812 5030
rect 215760 4966 215812 4972
rect 142289 4924 142585 4944
rect 142345 4922 142369 4924
rect 142425 4922 142449 4924
rect 142505 4922 142529 4924
rect 142367 4870 142369 4922
rect 142431 4870 142443 4922
rect 142505 4870 142507 4922
rect 142345 4868 142369 4870
rect 142425 4868 142449 4870
rect 142505 4868 142529 4870
rect 142289 4848 142585 4868
rect 213012 4690 213040 4966
rect 215772 4826 215800 4966
rect 215760 4820 215812 4826
rect 215760 4762 215812 4768
rect 213000 4684 213052 4690
rect 213000 4626 213052 4632
rect 212356 4616 212408 4622
rect 212356 4558 212408 4564
rect 212816 4616 212868 4622
rect 213012 4593 213040 4626
rect 212816 4558 212868 4564
rect 212998 4584 213054 4593
rect 71622 4380 71918 4400
rect 71678 4378 71702 4380
rect 71758 4378 71782 4380
rect 71838 4378 71862 4380
rect 71700 4326 71702 4378
rect 71764 4326 71776 4378
rect 71838 4326 71840 4378
rect 71678 4324 71702 4326
rect 71758 4324 71782 4326
rect 71838 4324 71862 4326
rect 71622 4304 71918 4324
rect 110 4176 166 4185
rect 110 4111 166 4120
rect 212368 3942 212396 4558
rect 212828 4282 212856 4558
rect 212998 4519 213054 4528
rect 212956 4380 213252 4400
rect 213012 4378 213036 4380
rect 213092 4378 213116 4380
rect 213172 4378 213196 4380
rect 213034 4326 213036 4378
rect 213098 4326 213110 4378
rect 213172 4326 213174 4378
rect 213012 4324 213036 4326
rect 213092 4324 213116 4326
rect 213172 4324 213196 4326
rect 212956 4304 213252 4324
rect 212816 4276 212868 4282
rect 212816 4218 212868 4224
rect 212356 3936 212408 3942
rect 212356 3878 212408 3884
rect 142289 3836 142585 3856
rect 142345 3834 142369 3836
rect 142425 3834 142449 3836
rect 142505 3834 142529 3836
rect 142367 3782 142369 3834
rect 142431 3782 142443 3834
rect 142505 3782 142507 3834
rect 142345 3780 142369 3782
rect 142425 3780 142449 3782
rect 142505 3780 142529 3782
rect 142289 3760 142585 3780
rect 71622 3292 71918 3312
rect 71678 3290 71702 3292
rect 71758 3290 71782 3292
rect 71838 3290 71862 3292
rect 71700 3238 71702 3290
rect 71764 3238 71776 3290
rect 71838 3238 71840 3290
rect 71678 3236 71702 3238
rect 71758 3236 71782 3238
rect 71838 3236 71862 3238
rect 71622 3216 71918 3236
rect 142289 2748 142585 2768
rect 142345 2746 142369 2748
rect 142425 2746 142449 2748
rect 142505 2746 142529 2748
rect 142367 2694 142369 2746
rect 142431 2694 142443 2746
rect 142505 2694 142507 2746
rect 142345 2692 142369 2694
rect 142425 2692 142449 2694
rect 142505 2692 142529 2694
rect 142289 2672 142585 2692
rect 211620 2372 211672 2378
rect 211620 2314 211672 2320
rect 71622 2204 71918 2224
rect 71678 2202 71702 2204
rect 71758 2202 71782 2204
rect 71838 2202 71862 2204
rect 71700 2150 71702 2202
rect 71764 2150 71776 2202
rect 71838 2150 71840 2202
rect 71678 2148 71702 2150
rect 71758 2148 71782 2150
rect 71838 2148 71862 2150
rect 71622 2128 71918 2148
rect 42522 1592 42578 1601
rect 42522 1527 42578 1536
rect 42338 82 42394 480
rect 42536 82 42564 1527
rect 42338 54 42564 82
rect 127070 96 127126 480
rect 42338 0 42394 54
rect 211632 82 211660 2314
rect 212368 1737 212396 3878
rect 214012 3528 214064 3534
rect 214012 3470 214064 3476
rect 212956 3292 213252 3312
rect 213012 3290 213036 3292
rect 213092 3290 213116 3292
rect 213172 3290 213196 3292
rect 213034 3238 213036 3290
rect 213098 3238 213110 3290
rect 213172 3238 213174 3290
rect 213012 3236 213036 3238
rect 213092 3236 213116 3238
rect 213172 3236 213196 3238
rect 212956 3216 213252 3236
rect 212956 2204 213252 2224
rect 213012 2202 213036 2204
rect 213092 2202 213116 2204
rect 213172 2202 213196 2204
rect 213034 2150 213036 2202
rect 213098 2150 213110 2202
rect 213172 2150 213174 2202
rect 213012 2148 213036 2150
rect 213092 2148 213116 2150
rect 213172 2148 213196 2150
rect 212956 2128 213252 2148
rect 212354 1728 212410 1737
rect 212354 1663 212410 1672
rect 214024 1193 214052 3470
rect 215956 2650 215984 5510
rect 216140 4154 216168 6054
rect 216232 5914 216260 6190
rect 219636 6118 219664 6734
rect 219820 6186 219848 6870
rect 238588 6458 238616 6938
rect 238576 6452 238628 6458
rect 238576 6394 238628 6400
rect 237564 6248 237616 6254
rect 237484 6208 237564 6236
rect 219808 6180 219860 6186
rect 219808 6122 219860 6128
rect 219624 6112 219676 6118
rect 219624 6054 219676 6060
rect 216220 5908 216272 5914
rect 216220 5850 216272 5856
rect 217692 5160 217744 5166
rect 217692 5102 217744 5108
rect 217508 5092 217560 5098
rect 217508 5034 217560 5040
rect 217520 4758 217548 5034
rect 217600 5024 217652 5030
rect 217600 4966 217652 4972
rect 217508 4752 217560 4758
rect 217508 4694 217560 4700
rect 217612 4622 217640 4966
rect 217600 4616 217652 4622
rect 217600 4558 217652 4564
rect 217704 4486 217732 5102
rect 219636 4826 219664 6054
rect 219820 5846 219848 6122
rect 237380 6112 237432 6118
rect 237380 6054 237432 6060
rect 219808 5840 219860 5846
rect 219808 5782 219860 5788
rect 234252 5840 234304 5846
rect 234252 5782 234304 5788
rect 219716 5704 219768 5710
rect 219716 5646 219768 5652
rect 219728 5234 219756 5646
rect 219716 5228 219768 5234
rect 219716 5170 219768 5176
rect 219820 5137 219848 5782
rect 220360 5568 220412 5574
rect 220360 5510 220412 5516
rect 232412 5568 232464 5574
rect 232412 5510 232464 5516
rect 220372 5166 220400 5510
rect 232424 5166 232452 5510
rect 220360 5160 220412 5166
rect 219806 5128 219862 5137
rect 220360 5102 220412 5108
rect 220452 5160 220504 5166
rect 220452 5102 220504 5108
rect 226432 5160 226484 5166
rect 232412 5160 232464 5166
rect 226432 5102 226484 5108
rect 232226 5128 232282 5137
rect 219806 5063 219862 5072
rect 219820 5030 219848 5063
rect 219808 5024 219860 5030
rect 219808 4966 219860 4972
rect 219624 4820 219676 4826
rect 219624 4762 219676 4768
rect 219820 4758 219848 4966
rect 218152 4752 218204 4758
rect 218152 4694 218204 4700
rect 219808 4752 219860 4758
rect 219808 4694 219860 4700
rect 217692 4480 217744 4486
rect 217692 4422 217744 4428
rect 217968 4480 218020 4486
rect 217968 4422 218020 4428
rect 216140 4126 216260 4154
rect 216128 3936 216180 3942
rect 216128 3878 216180 3884
rect 216140 3534 216168 3878
rect 216128 3528 216180 3534
rect 216128 3470 216180 3476
rect 216232 3369 216260 4126
rect 217048 4004 217100 4010
rect 217048 3946 217100 3952
rect 217060 3738 217088 3946
rect 217048 3732 217100 3738
rect 217048 3674 217100 3680
rect 217704 3602 217732 4422
rect 217980 4078 218008 4422
rect 218164 4282 218192 4694
rect 220372 4690 220400 5102
rect 220360 4684 220412 4690
rect 220360 4626 220412 4632
rect 218428 4616 218480 4622
rect 218428 4558 218480 4564
rect 218152 4276 218204 4282
rect 218152 4218 218204 4224
rect 217968 4072 218020 4078
rect 217968 4014 218020 4020
rect 217784 3732 217836 3738
rect 217784 3674 217836 3680
rect 217692 3596 217744 3602
rect 217692 3538 217744 3544
rect 217796 3534 217824 3674
rect 217784 3528 217836 3534
rect 217784 3470 217836 3476
rect 216218 3360 216274 3369
rect 216218 3295 216274 3304
rect 217796 2990 217824 3470
rect 217784 2984 217836 2990
rect 217784 2926 217836 2932
rect 217600 2916 217652 2922
rect 217600 2858 217652 2864
rect 217232 2848 217284 2854
rect 217232 2790 217284 2796
rect 215944 2644 215996 2650
rect 215944 2586 215996 2592
rect 215956 2009 215984 2586
rect 217244 2582 217272 2790
rect 217232 2576 217284 2582
rect 217232 2518 217284 2524
rect 215942 2000 215998 2009
rect 215942 1935 215998 1944
rect 217612 1601 217640 2858
rect 217980 2854 218008 4014
rect 218164 4010 218192 4218
rect 218440 4146 218468 4558
rect 220372 4214 220400 4626
rect 220464 4282 220492 5102
rect 220636 5024 220688 5030
rect 220636 4966 220688 4972
rect 221832 5024 221884 5030
rect 221832 4966 221884 4972
rect 220648 4486 220676 4966
rect 221844 4690 221872 4966
rect 221924 4752 221976 4758
rect 221924 4694 221976 4700
rect 221372 4684 221424 4690
rect 221372 4626 221424 4632
rect 221832 4684 221884 4690
rect 221832 4626 221884 4632
rect 220636 4480 220688 4486
rect 220636 4422 220688 4428
rect 221188 4480 221240 4486
rect 221188 4422 221240 4428
rect 220452 4276 220504 4282
rect 220452 4218 220504 4224
rect 220360 4208 220412 4214
rect 220360 4150 220412 4156
rect 218428 4140 218480 4146
rect 218428 4082 218480 4088
rect 220266 4040 220322 4049
rect 218152 4004 218204 4010
rect 218152 3946 218204 3952
rect 220084 4004 220136 4010
rect 220266 3975 220322 3984
rect 220084 3946 220136 3952
rect 218164 3738 218192 3946
rect 218980 3936 219032 3942
rect 218980 3878 219032 3884
rect 218152 3732 218204 3738
rect 218152 3674 218204 3680
rect 218992 2990 219020 3878
rect 219808 3732 219860 3738
rect 219808 3674 219860 3680
rect 219820 3602 219848 3674
rect 220096 3670 220124 3946
rect 220280 3942 220308 3975
rect 220372 3942 220400 4150
rect 220464 4010 220492 4218
rect 221096 4072 221148 4078
rect 221096 4014 221148 4020
rect 220452 4004 220504 4010
rect 220452 3946 220504 3952
rect 220268 3936 220320 3942
rect 220268 3878 220320 3884
rect 220360 3936 220412 3942
rect 220360 3878 220412 3884
rect 220084 3664 220136 3670
rect 220084 3606 220136 3612
rect 219072 3596 219124 3602
rect 219072 3538 219124 3544
rect 219532 3596 219584 3602
rect 219532 3538 219584 3544
rect 219808 3596 219860 3602
rect 219808 3538 219860 3544
rect 219084 3058 219112 3538
rect 219440 3460 219492 3466
rect 219440 3402 219492 3408
rect 219452 3194 219480 3402
rect 219440 3188 219492 3194
rect 219440 3130 219492 3136
rect 219072 3052 219124 3058
rect 219072 2994 219124 3000
rect 218520 2984 218572 2990
rect 218520 2926 218572 2932
rect 218980 2984 219032 2990
rect 218980 2926 219032 2932
rect 217968 2848 218020 2854
rect 217968 2790 218020 2796
rect 218532 2650 218560 2926
rect 218520 2644 218572 2650
rect 218520 2586 218572 2592
rect 218992 2514 219020 2926
rect 219084 2650 219112 2994
rect 219072 2644 219124 2650
rect 219072 2586 219124 2592
rect 219544 2582 219572 3538
rect 219532 2576 219584 2582
rect 219532 2518 219584 2524
rect 218980 2508 219032 2514
rect 218980 2450 219032 2456
rect 219820 2446 219848 3538
rect 220372 3534 220400 3878
rect 220360 3528 220412 3534
rect 220360 3470 220412 3476
rect 220464 2990 220492 3946
rect 221004 3936 221056 3942
rect 221004 3878 221056 3884
rect 221016 3670 221044 3878
rect 221004 3664 221056 3670
rect 221004 3606 221056 3612
rect 221108 3602 221136 4014
rect 221200 3602 221228 4422
rect 221384 4078 221412 4626
rect 221372 4072 221424 4078
rect 221372 4014 221424 4020
rect 221384 3942 221412 4014
rect 221844 3942 221872 4626
rect 221936 3942 221964 4694
rect 224592 4616 224644 4622
rect 224592 4558 224644 4564
rect 223212 4480 223264 4486
rect 223212 4422 223264 4428
rect 224500 4480 224552 4486
rect 224500 4422 224552 4428
rect 222568 4072 222620 4078
rect 223224 4049 223252 4422
rect 224512 4078 224540 4422
rect 224604 4146 224632 4558
rect 226156 4480 226208 4486
rect 226156 4422 226208 4428
rect 224592 4140 224644 4146
rect 224592 4082 224644 4088
rect 223580 4072 223632 4078
rect 222568 4014 222620 4020
rect 223210 4040 223266 4049
rect 221372 3936 221424 3942
rect 221372 3878 221424 3884
rect 221832 3936 221884 3942
rect 221832 3878 221884 3884
rect 221924 3936 221976 3942
rect 221924 3878 221976 3884
rect 221844 3738 221872 3878
rect 221832 3732 221884 3738
rect 221832 3674 221884 3680
rect 221096 3596 221148 3602
rect 221096 3538 221148 3544
rect 221188 3596 221240 3602
rect 221188 3538 221240 3544
rect 221004 3528 221056 3534
rect 221004 3470 221056 3476
rect 220452 2984 220504 2990
rect 220452 2926 220504 2932
rect 221016 2836 221044 3470
rect 221108 3194 221136 3538
rect 221844 3398 221872 3674
rect 221936 3534 221964 3878
rect 222580 3738 222608 4014
rect 223580 4014 223632 4020
rect 223948 4072 224000 4078
rect 223948 4014 224000 4020
rect 224500 4072 224552 4078
rect 224500 4014 224552 4020
rect 225052 4072 225104 4078
rect 225052 4014 225104 4020
rect 223210 3975 223266 3984
rect 222844 3936 222896 3942
rect 222844 3878 222896 3884
rect 222568 3732 222620 3738
rect 222568 3674 222620 3680
rect 221924 3528 221976 3534
rect 221924 3470 221976 3476
rect 221832 3392 221884 3398
rect 221832 3334 221884 3340
rect 221096 3188 221148 3194
rect 221096 3130 221148 3136
rect 221936 3058 221964 3470
rect 222856 3466 222884 3878
rect 222936 3596 222988 3602
rect 222936 3538 222988 3544
rect 222844 3460 222896 3466
rect 222844 3402 222896 3408
rect 222856 3194 222884 3402
rect 222844 3188 222896 3194
rect 222844 3130 222896 3136
rect 222948 3058 222976 3538
rect 223592 3534 223620 4014
rect 223960 3534 223988 4014
rect 224960 3936 225012 3942
rect 224960 3878 225012 3884
rect 224972 3670 225000 3878
rect 224868 3664 224920 3670
rect 224868 3606 224920 3612
rect 224960 3664 225012 3670
rect 224960 3606 225012 3612
rect 223580 3528 223632 3534
rect 223580 3470 223632 3476
rect 223948 3528 224000 3534
rect 224880 3505 224908 3606
rect 223948 3470 224000 3476
rect 224866 3496 224922 3505
rect 221924 3052 221976 3058
rect 221924 2994 221976 3000
rect 222936 3052 222988 3058
rect 222936 2994 222988 3000
rect 221096 2848 221148 2854
rect 221016 2808 221096 2836
rect 221096 2790 221148 2796
rect 219808 2440 219860 2446
rect 221108 2417 221136 2790
rect 223960 2650 223988 3470
rect 224866 3431 224922 3440
rect 224972 3194 225000 3606
rect 225064 3602 225092 4014
rect 225788 4004 225840 4010
rect 225788 3946 225840 3952
rect 225052 3596 225104 3602
rect 225052 3538 225104 3544
rect 225064 3194 225092 3538
rect 225800 3398 225828 3946
rect 226168 3942 226196 4422
rect 226444 4146 226472 5102
rect 232412 5102 232464 5108
rect 234264 5098 234292 5782
rect 234528 5704 234580 5710
rect 234528 5646 234580 5652
rect 232226 5063 232282 5072
rect 234252 5092 234304 5098
rect 232240 5030 232268 5063
rect 234252 5034 234304 5040
rect 232228 5024 232280 5030
rect 232228 4966 232280 4972
rect 232240 4758 232268 4966
rect 232228 4752 232280 4758
rect 232228 4694 232280 4700
rect 232240 4282 232268 4694
rect 232688 4616 232740 4622
rect 232688 4558 232740 4564
rect 232700 4282 232728 4558
rect 232228 4276 232280 4282
rect 232228 4218 232280 4224
rect 232688 4276 232740 4282
rect 232688 4218 232740 4224
rect 226432 4140 226484 4146
rect 226432 4082 226484 4088
rect 225880 3936 225932 3942
rect 225880 3878 225932 3884
rect 226156 3936 226208 3942
rect 226156 3878 226208 3884
rect 225892 3670 225920 3878
rect 225880 3664 225932 3670
rect 225880 3606 225932 3612
rect 225970 3632 226026 3641
rect 225788 3392 225840 3398
rect 225788 3334 225840 3340
rect 224960 3188 225012 3194
rect 224960 3130 225012 3136
rect 225052 3188 225104 3194
rect 225052 3130 225104 3136
rect 225892 3126 225920 3606
rect 226026 3602 226104 3618
rect 226026 3596 226116 3602
rect 226026 3590 226064 3596
rect 225970 3567 226026 3576
rect 226064 3538 226116 3544
rect 225880 3120 225932 3126
rect 225880 3062 225932 3068
rect 223948 2644 224000 2650
rect 223948 2586 224000 2592
rect 219808 2382 219860 2388
rect 221094 2408 221150 2417
rect 221094 2343 221150 2352
rect 217598 1592 217654 1601
rect 217598 1527 217654 1536
rect 214010 1184 214066 1193
rect 214010 1119 214066 1128
rect 211894 82 211950 480
rect 225892 105 225920 3062
rect 226168 3058 226196 3878
rect 226156 3052 226208 3058
rect 226156 2994 226208 3000
rect 226168 1601 226196 2994
rect 226154 1592 226210 1601
rect 226154 1527 226210 1536
rect 234264 241 234292 5034
rect 234540 5030 234568 5646
rect 235080 5568 235132 5574
rect 235080 5510 235132 5516
rect 235092 5273 235120 5510
rect 235078 5264 235134 5273
rect 235078 5199 235134 5208
rect 234528 5024 234580 5030
rect 234528 4966 234580 4972
rect 234540 3641 234568 4966
rect 237392 4185 237420 6054
rect 237484 5574 237512 6208
rect 237564 6190 237616 6196
rect 237472 5568 237524 5574
rect 237472 5510 237524 5516
rect 237484 5370 237512 5510
rect 239140 5370 239168 7278
rect 283622 7100 283918 7120
rect 283678 7098 283702 7100
rect 283758 7098 283782 7100
rect 283838 7098 283862 7100
rect 283700 7046 283702 7098
rect 283764 7046 283776 7098
rect 283838 7046 283840 7098
rect 283678 7044 283702 7046
rect 283758 7044 283782 7046
rect 283838 7044 283862 7046
rect 283622 7024 283918 7044
rect 283622 6012 283918 6032
rect 283678 6010 283702 6012
rect 283758 6010 283782 6012
rect 283838 6010 283862 6012
rect 283700 5958 283702 6010
rect 283764 5958 283776 6010
rect 283838 5958 283840 6010
rect 283678 5956 283702 5958
rect 283758 5956 283782 5958
rect 283838 5956 283862 5958
rect 283622 5936 283918 5956
rect 291120 5370 291148 9574
rect 291474 9520 291530 9574
rect 344466 9602 344522 10000
rect 397458 9602 397514 10000
rect 423586 9616 423642 9625
rect 344466 9574 344600 9602
rect 344466 9520 344522 9574
rect 344572 6769 344600 9574
rect 397458 9574 397776 9602
rect 397458 9520 397514 9574
rect 354289 7644 354585 7664
rect 354345 7642 354369 7644
rect 354425 7642 354449 7644
rect 354505 7642 354529 7644
rect 354367 7590 354369 7642
rect 354431 7590 354443 7642
rect 354505 7590 354507 7642
rect 354345 7588 354369 7590
rect 354425 7588 354449 7590
rect 354505 7588 354529 7590
rect 354289 7568 354585 7588
rect 344558 6760 344614 6769
rect 344558 6695 344614 6704
rect 354289 6556 354585 6576
rect 354345 6554 354369 6556
rect 354425 6554 354449 6556
rect 354505 6554 354529 6556
rect 354367 6502 354369 6554
rect 354431 6502 354443 6554
rect 354505 6502 354507 6554
rect 354345 6500 354369 6502
rect 354425 6500 354449 6502
rect 354505 6500 354529 6502
rect 354289 6480 354585 6500
rect 397748 6458 397776 9574
rect 423508 9574 423586 9602
rect 404176 7336 404228 7342
rect 404176 7278 404228 7284
rect 404188 6458 404216 7278
rect 423508 7002 423536 9574
rect 423586 9551 423642 9560
rect 423586 7712 423642 7721
rect 423586 7647 423642 7656
rect 423600 7274 423628 7647
rect 423588 7268 423640 7274
rect 423588 7210 423640 7216
rect 423680 7200 423732 7206
rect 423680 7142 423732 7148
rect 423496 6996 423548 7002
rect 423496 6938 423548 6944
rect 423692 6905 423720 7142
rect 423678 6896 423734 6905
rect 423678 6831 423734 6840
rect 397736 6452 397788 6458
rect 397736 6394 397788 6400
rect 404176 6452 404228 6458
rect 404176 6394 404228 6400
rect 399666 6352 399722 6361
rect 399666 6287 399722 6296
rect 399680 6254 399708 6287
rect 399668 6248 399720 6254
rect 399668 6190 399720 6196
rect 399760 6248 399812 6254
rect 399760 6190 399812 6196
rect 399668 5568 399720 5574
rect 399772 5556 399800 6190
rect 399720 5528 399800 5556
rect 399668 5510 399720 5516
rect 354289 5468 354585 5488
rect 354345 5466 354369 5468
rect 354425 5466 354449 5468
rect 354505 5466 354529 5468
rect 354367 5414 354369 5466
rect 354431 5414 354443 5466
rect 354505 5414 354507 5466
rect 354345 5412 354369 5414
rect 354425 5412 354449 5414
rect 354505 5412 354529 5414
rect 354289 5392 354585 5412
rect 237472 5364 237524 5370
rect 237472 5306 237524 5312
rect 239128 5364 239180 5370
rect 239128 5306 239180 5312
rect 291108 5364 291160 5370
rect 291108 5306 291160 5312
rect 399680 5273 399708 5510
rect 399666 5264 399722 5273
rect 399666 5199 399722 5208
rect 238668 5160 238720 5166
rect 238668 5102 238720 5108
rect 289452 5160 289504 5166
rect 289452 5102 289504 5108
rect 238392 5024 238444 5030
rect 238392 4966 238444 4972
rect 237378 4176 237434 4185
rect 237378 4111 237434 4120
rect 234526 3632 234582 3641
rect 234526 3567 234582 3576
rect 238404 2961 238432 4966
rect 238680 4690 238708 5102
rect 283622 4924 283918 4944
rect 283678 4922 283702 4924
rect 283758 4922 283782 4924
rect 283838 4922 283862 4924
rect 283700 4870 283702 4922
rect 283764 4870 283776 4922
rect 283838 4870 283840 4922
rect 283678 4868 283702 4870
rect 283758 4868 283782 4870
rect 283838 4868 283862 4870
rect 283622 4848 283918 4868
rect 238668 4684 238720 4690
rect 238668 4626 238720 4632
rect 283622 3836 283918 3856
rect 283678 3834 283702 3836
rect 283758 3834 283782 3836
rect 283838 3834 283862 3836
rect 283700 3782 283702 3834
rect 283764 3782 283776 3834
rect 283838 3782 283840 3834
rect 283678 3780 283702 3782
rect 283758 3780 283782 3782
rect 283838 3780 283862 3782
rect 283622 3760 283918 3780
rect 289464 3505 289492 5102
rect 289636 5024 289688 5030
rect 289636 4966 289688 4972
rect 289450 3496 289506 3505
rect 289450 3431 289506 3440
rect 289648 3097 289676 4966
rect 354289 4380 354585 4400
rect 354345 4378 354369 4380
rect 354425 4378 354449 4380
rect 354505 4378 354529 4380
rect 354367 4326 354369 4378
rect 354431 4326 354443 4378
rect 354505 4326 354507 4378
rect 354345 4324 354369 4326
rect 354425 4324 354449 4326
rect 354505 4324 354529 4326
rect 354289 4304 354585 4324
rect 296442 3360 296498 3369
rect 296442 3295 296498 3304
rect 289634 3088 289690 3097
rect 289634 3023 289690 3032
rect 238390 2952 238446 2961
rect 238390 2887 238446 2896
rect 283622 2748 283918 2768
rect 283678 2746 283702 2748
rect 283758 2746 283782 2748
rect 283838 2746 283862 2748
rect 283700 2694 283702 2746
rect 283764 2694 283776 2746
rect 283838 2694 283840 2746
rect 283678 2692 283702 2694
rect 283758 2692 283782 2694
rect 283838 2692 283862 2694
rect 283622 2672 283918 2692
rect 234250 232 234306 241
rect 234250 167 234306 176
rect 211632 54 211950 82
rect 127070 0 127126 40
rect 211894 0 211950 54
rect 225878 96 225934 105
rect 296456 82 296484 3295
rect 354289 3292 354585 3312
rect 354345 3290 354369 3292
rect 354425 3290 354449 3292
rect 354505 3290 354529 3292
rect 354367 3238 354369 3290
rect 354431 3238 354443 3290
rect 354505 3238 354507 3290
rect 354345 3236 354369 3238
rect 354425 3236 354449 3238
rect 354505 3236 354529 3238
rect 354289 3216 354585 3236
rect 354289 2204 354585 2224
rect 354345 2202 354369 2204
rect 354425 2202 354449 2204
rect 354505 2202 354529 2204
rect 354367 2150 354369 2202
rect 354431 2150 354443 2202
rect 354505 2150 354507 2202
rect 354345 2148 354369 2150
rect 354425 2148 354449 2150
rect 354505 2148 354529 2150
rect 354289 2128 354585 2148
rect 381266 2000 381322 2009
rect 381266 1935 381322 1944
rect 296718 82 296774 480
rect 296456 54 296774 82
rect 381280 82 381308 1935
rect 423586 1320 423642 1329
rect 423508 1278 423586 1306
rect 381542 82 381598 480
rect 423508 241 423536 1278
rect 423586 1255 423642 1264
rect 423494 232 423550 241
rect 423494 167 423550 176
rect 381280 54 381598 82
rect 225878 31 225934 40
rect 296718 0 296774 54
rect 381542 0 381598 54
<< via2 >>
rect 18 9152 74 9208
rect 71622 7642 71678 7644
rect 71702 7642 71758 7644
rect 71782 7642 71838 7644
rect 71862 7642 71918 7644
rect 71622 7590 71648 7642
rect 71648 7590 71678 7642
rect 71702 7590 71712 7642
rect 71712 7590 71758 7642
rect 71782 7590 71828 7642
rect 71828 7590 71838 7642
rect 71862 7590 71892 7642
rect 71892 7590 71918 7642
rect 71622 7588 71678 7590
rect 71702 7588 71758 7590
rect 71782 7588 71838 7590
rect 71862 7588 71918 7590
rect 110 7520 166 7576
rect 142289 7098 142345 7100
rect 142369 7098 142425 7100
rect 142449 7098 142505 7100
rect 142529 7098 142585 7100
rect 142289 7046 142315 7098
rect 142315 7046 142345 7098
rect 142369 7046 142379 7098
rect 142379 7046 142425 7098
rect 142449 7046 142495 7098
rect 142495 7046 142505 7098
rect 142529 7046 142559 7098
rect 142559 7046 142585 7098
rect 142289 7044 142345 7046
rect 142369 7044 142425 7046
rect 142449 7044 142505 7046
rect 142529 7044 142585 7046
rect 132774 6840 132830 6896
rect 212956 7642 213012 7644
rect 213036 7642 213092 7644
rect 213116 7642 213172 7644
rect 213196 7642 213252 7644
rect 212956 7590 212982 7642
rect 212982 7590 213012 7642
rect 213036 7590 213046 7642
rect 213046 7590 213092 7642
rect 213116 7590 213162 7642
rect 213162 7590 213172 7642
rect 213196 7590 213226 7642
rect 213226 7590 213252 7642
rect 212956 7588 213012 7590
rect 213036 7588 213092 7590
rect 213116 7588 213172 7590
rect 213196 7588 213252 7590
rect 185766 6704 185822 6760
rect 202142 6704 202198 6760
rect 71622 6554 71678 6556
rect 71702 6554 71758 6556
rect 71782 6554 71838 6556
rect 71862 6554 71918 6556
rect 71622 6502 71648 6554
rect 71648 6502 71678 6554
rect 71702 6502 71712 6554
rect 71712 6502 71758 6554
rect 71782 6502 71828 6554
rect 71828 6502 71838 6554
rect 71862 6502 71892 6554
rect 71892 6502 71918 6554
rect 71622 6500 71678 6502
rect 71702 6500 71758 6502
rect 71782 6500 71838 6502
rect 71862 6500 71918 6502
rect 212956 6554 213012 6556
rect 213036 6554 213092 6556
rect 213116 6554 213172 6556
rect 213196 6554 213252 6556
rect 212956 6502 212982 6554
rect 212982 6502 213012 6554
rect 213036 6502 213046 6554
rect 213046 6502 213092 6554
rect 213116 6502 213162 6554
rect 213162 6502 213172 6554
rect 213196 6502 213226 6554
rect 213226 6502 213252 6554
rect 212956 6500 213012 6502
rect 213036 6500 213092 6502
rect 213116 6500 213172 6502
rect 213196 6500 213252 6502
rect 142289 6010 142345 6012
rect 142369 6010 142425 6012
rect 142449 6010 142505 6012
rect 142529 6010 142585 6012
rect 142289 5958 142315 6010
rect 142315 5958 142345 6010
rect 142369 5958 142379 6010
rect 142379 5958 142425 6010
rect 142449 5958 142495 6010
rect 142495 5958 142505 6010
rect 142529 5958 142559 6010
rect 142559 5958 142585 6010
rect 142289 5956 142345 5958
rect 142369 5956 142425 5958
rect 142449 5956 142505 5958
rect 142529 5956 142585 5958
rect 215298 6840 215354 6896
rect 216218 6704 216274 6760
rect 215574 6160 215630 6216
rect 71622 5466 71678 5468
rect 71702 5466 71758 5468
rect 71782 5466 71838 5468
rect 71862 5466 71918 5468
rect 71622 5414 71648 5466
rect 71648 5414 71678 5466
rect 71702 5414 71712 5466
rect 71712 5414 71758 5466
rect 71782 5414 71828 5466
rect 71828 5414 71838 5466
rect 71862 5414 71892 5466
rect 71892 5414 71918 5466
rect 71622 5412 71678 5414
rect 71702 5412 71758 5414
rect 71782 5412 71838 5414
rect 71862 5412 71918 5414
rect 110 5208 166 5264
rect 212956 5466 213012 5468
rect 213036 5466 213092 5468
rect 213116 5466 213172 5468
rect 213196 5466 213252 5468
rect 212956 5414 212982 5466
rect 212982 5414 213012 5466
rect 213036 5414 213046 5466
rect 213046 5414 213092 5466
rect 213116 5414 213162 5466
rect 213162 5414 213172 5466
rect 213196 5414 213226 5466
rect 213226 5414 213252 5466
rect 212956 5412 213012 5414
rect 213036 5412 213092 5414
rect 213116 5412 213172 5414
rect 213196 5412 213252 5414
rect 209502 5208 209558 5264
rect 142289 4922 142345 4924
rect 142369 4922 142425 4924
rect 142449 4922 142505 4924
rect 142529 4922 142585 4924
rect 142289 4870 142315 4922
rect 142315 4870 142345 4922
rect 142369 4870 142379 4922
rect 142379 4870 142425 4922
rect 142449 4870 142495 4922
rect 142495 4870 142505 4922
rect 142529 4870 142559 4922
rect 142559 4870 142585 4922
rect 142289 4868 142345 4870
rect 142369 4868 142425 4870
rect 142449 4868 142505 4870
rect 142529 4868 142585 4870
rect 71622 4378 71678 4380
rect 71702 4378 71758 4380
rect 71782 4378 71838 4380
rect 71862 4378 71918 4380
rect 71622 4326 71648 4378
rect 71648 4326 71678 4378
rect 71702 4326 71712 4378
rect 71712 4326 71758 4378
rect 71782 4326 71828 4378
rect 71828 4326 71838 4378
rect 71862 4326 71892 4378
rect 71892 4326 71918 4378
rect 71622 4324 71678 4326
rect 71702 4324 71758 4326
rect 71782 4324 71838 4326
rect 71862 4324 71918 4326
rect 110 4120 166 4176
rect 212998 4528 213054 4584
rect 212956 4378 213012 4380
rect 213036 4378 213092 4380
rect 213116 4378 213172 4380
rect 213196 4378 213252 4380
rect 212956 4326 212982 4378
rect 212982 4326 213012 4378
rect 213036 4326 213046 4378
rect 213046 4326 213092 4378
rect 213116 4326 213162 4378
rect 213162 4326 213172 4378
rect 213196 4326 213226 4378
rect 213226 4326 213252 4378
rect 212956 4324 213012 4326
rect 213036 4324 213092 4326
rect 213116 4324 213172 4326
rect 213196 4324 213252 4326
rect 142289 3834 142345 3836
rect 142369 3834 142425 3836
rect 142449 3834 142505 3836
rect 142529 3834 142585 3836
rect 142289 3782 142315 3834
rect 142315 3782 142345 3834
rect 142369 3782 142379 3834
rect 142379 3782 142425 3834
rect 142449 3782 142495 3834
rect 142495 3782 142505 3834
rect 142529 3782 142559 3834
rect 142559 3782 142585 3834
rect 142289 3780 142345 3782
rect 142369 3780 142425 3782
rect 142449 3780 142505 3782
rect 142529 3780 142585 3782
rect 71622 3290 71678 3292
rect 71702 3290 71758 3292
rect 71782 3290 71838 3292
rect 71862 3290 71918 3292
rect 71622 3238 71648 3290
rect 71648 3238 71678 3290
rect 71702 3238 71712 3290
rect 71712 3238 71758 3290
rect 71782 3238 71828 3290
rect 71828 3238 71838 3290
rect 71862 3238 71892 3290
rect 71892 3238 71918 3290
rect 71622 3236 71678 3238
rect 71702 3236 71758 3238
rect 71782 3236 71838 3238
rect 71862 3236 71918 3238
rect 142289 2746 142345 2748
rect 142369 2746 142425 2748
rect 142449 2746 142505 2748
rect 142529 2746 142585 2748
rect 142289 2694 142315 2746
rect 142315 2694 142345 2746
rect 142369 2694 142379 2746
rect 142379 2694 142425 2746
rect 142449 2694 142495 2746
rect 142495 2694 142505 2746
rect 142529 2694 142559 2746
rect 142559 2694 142585 2746
rect 142289 2692 142345 2694
rect 142369 2692 142425 2694
rect 142449 2692 142505 2694
rect 142529 2692 142585 2694
rect 71622 2202 71678 2204
rect 71702 2202 71758 2204
rect 71782 2202 71838 2204
rect 71862 2202 71918 2204
rect 71622 2150 71648 2202
rect 71648 2150 71678 2202
rect 71702 2150 71712 2202
rect 71712 2150 71758 2202
rect 71782 2150 71828 2202
rect 71828 2150 71838 2202
rect 71862 2150 71892 2202
rect 71892 2150 71918 2202
rect 71622 2148 71678 2150
rect 71702 2148 71758 2150
rect 71782 2148 71838 2150
rect 71862 2148 71918 2150
rect 42522 1536 42578 1592
rect 127070 40 127126 96
rect 212956 3290 213012 3292
rect 213036 3290 213092 3292
rect 213116 3290 213172 3292
rect 213196 3290 213252 3292
rect 212956 3238 212982 3290
rect 212982 3238 213012 3290
rect 213036 3238 213046 3290
rect 213046 3238 213092 3290
rect 213116 3238 213162 3290
rect 213162 3238 213172 3290
rect 213196 3238 213226 3290
rect 213226 3238 213252 3290
rect 212956 3236 213012 3238
rect 213036 3236 213092 3238
rect 213116 3236 213172 3238
rect 213196 3236 213252 3238
rect 212956 2202 213012 2204
rect 213036 2202 213092 2204
rect 213116 2202 213172 2204
rect 213196 2202 213252 2204
rect 212956 2150 212982 2202
rect 212982 2150 213012 2202
rect 213036 2150 213046 2202
rect 213046 2150 213092 2202
rect 213116 2150 213162 2202
rect 213162 2150 213172 2202
rect 213196 2150 213226 2202
rect 213226 2150 213252 2202
rect 212956 2148 213012 2150
rect 213036 2148 213092 2150
rect 213116 2148 213172 2150
rect 213196 2148 213252 2150
rect 212354 1672 212410 1728
rect 219806 5072 219862 5128
rect 216218 3304 216274 3360
rect 215942 1944 215998 2000
rect 220266 3984 220322 4040
rect 223210 3984 223266 4040
rect 224866 3440 224922 3496
rect 232226 5072 232282 5128
rect 225970 3576 226026 3632
rect 221094 2352 221150 2408
rect 217598 1536 217654 1592
rect 214010 1128 214066 1184
rect 226154 1536 226210 1592
rect 235078 5208 235134 5264
rect 283622 7098 283678 7100
rect 283702 7098 283758 7100
rect 283782 7098 283838 7100
rect 283862 7098 283918 7100
rect 283622 7046 283648 7098
rect 283648 7046 283678 7098
rect 283702 7046 283712 7098
rect 283712 7046 283758 7098
rect 283782 7046 283828 7098
rect 283828 7046 283838 7098
rect 283862 7046 283892 7098
rect 283892 7046 283918 7098
rect 283622 7044 283678 7046
rect 283702 7044 283758 7046
rect 283782 7044 283838 7046
rect 283862 7044 283918 7046
rect 283622 6010 283678 6012
rect 283702 6010 283758 6012
rect 283782 6010 283838 6012
rect 283862 6010 283918 6012
rect 283622 5958 283648 6010
rect 283648 5958 283678 6010
rect 283702 5958 283712 6010
rect 283712 5958 283758 6010
rect 283782 5958 283828 6010
rect 283828 5958 283838 6010
rect 283862 5958 283892 6010
rect 283892 5958 283918 6010
rect 283622 5956 283678 5958
rect 283702 5956 283758 5958
rect 283782 5956 283838 5958
rect 283862 5956 283918 5958
rect 354289 7642 354345 7644
rect 354369 7642 354425 7644
rect 354449 7642 354505 7644
rect 354529 7642 354585 7644
rect 354289 7590 354315 7642
rect 354315 7590 354345 7642
rect 354369 7590 354379 7642
rect 354379 7590 354425 7642
rect 354449 7590 354495 7642
rect 354495 7590 354505 7642
rect 354529 7590 354559 7642
rect 354559 7590 354585 7642
rect 354289 7588 354345 7590
rect 354369 7588 354425 7590
rect 354449 7588 354505 7590
rect 354529 7588 354585 7590
rect 344558 6704 344614 6760
rect 354289 6554 354345 6556
rect 354369 6554 354425 6556
rect 354449 6554 354505 6556
rect 354529 6554 354585 6556
rect 354289 6502 354315 6554
rect 354315 6502 354345 6554
rect 354369 6502 354379 6554
rect 354379 6502 354425 6554
rect 354449 6502 354495 6554
rect 354495 6502 354505 6554
rect 354529 6502 354559 6554
rect 354559 6502 354585 6554
rect 354289 6500 354345 6502
rect 354369 6500 354425 6502
rect 354449 6500 354505 6502
rect 354529 6500 354585 6502
rect 423586 9560 423642 9616
rect 423586 7656 423642 7712
rect 423678 6840 423734 6896
rect 399666 6296 399722 6352
rect 354289 5466 354345 5468
rect 354369 5466 354425 5468
rect 354449 5466 354505 5468
rect 354529 5466 354585 5468
rect 354289 5414 354315 5466
rect 354315 5414 354345 5466
rect 354369 5414 354379 5466
rect 354379 5414 354425 5466
rect 354449 5414 354495 5466
rect 354495 5414 354505 5466
rect 354529 5414 354559 5466
rect 354559 5414 354585 5466
rect 354289 5412 354345 5414
rect 354369 5412 354425 5414
rect 354449 5412 354505 5414
rect 354529 5412 354585 5414
rect 399666 5208 399722 5264
rect 237378 4120 237434 4176
rect 234526 3576 234582 3632
rect 283622 4922 283678 4924
rect 283702 4922 283758 4924
rect 283782 4922 283838 4924
rect 283862 4922 283918 4924
rect 283622 4870 283648 4922
rect 283648 4870 283678 4922
rect 283702 4870 283712 4922
rect 283712 4870 283758 4922
rect 283782 4870 283828 4922
rect 283828 4870 283838 4922
rect 283862 4870 283892 4922
rect 283892 4870 283918 4922
rect 283622 4868 283678 4870
rect 283702 4868 283758 4870
rect 283782 4868 283838 4870
rect 283862 4868 283918 4870
rect 283622 3834 283678 3836
rect 283702 3834 283758 3836
rect 283782 3834 283838 3836
rect 283862 3834 283918 3836
rect 283622 3782 283648 3834
rect 283648 3782 283678 3834
rect 283702 3782 283712 3834
rect 283712 3782 283758 3834
rect 283782 3782 283828 3834
rect 283828 3782 283838 3834
rect 283862 3782 283892 3834
rect 283892 3782 283918 3834
rect 283622 3780 283678 3782
rect 283702 3780 283758 3782
rect 283782 3780 283838 3782
rect 283862 3780 283918 3782
rect 289450 3440 289506 3496
rect 354289 4378 354345 4380
rect 354369 4378 354425 4380
rect 354449 4378 354505 4380
rect 354529 4378 354585 4380
rect 354289 4326 354315 4378
rect 354315 4326 354345 4378
rect 354369 4326 354379 4378
rect 354379 4326 354425 4378
rect 354449 4326 354495 4378
rect 354495 4326 354505 4378
rect 354529 4326 354559 4378
rect 354559 4326 354585 4378
rect 354289 4324 354345 4326
rect 354369 4324 354425 4326
rect 354449 4324 354505 4326
rect 354529 4324 354585 4326
rect 296442 3304 296498 3360
rect 289634 3032 289690 3088
rect 238390 2896 238446 2952
rect 283622 2746 283678 2748
rect 283702 2746 283758 2748
rect 283782 2746 283838 2748
rect 283862 2746 283918 2748
rect 283622 2694 283648 2746
rect 283648 2694 283678 2746
rect 283702 2694 283712 2746
rect 283712 2694 283758 2746
rect 283782 2694 283828 2746
rect 283828 2694 283838 2746
rect 283862 2694 283892 2746
rect 283892 2694 283918 2746
rect 283622 2692 283678 2694
rect 283702 2692 283758 2694
rect 283782 2692 283838 2694
rect 283862 2692 283918 2694
rect 234250 176 234306 232
rect 225878 40 225934 96
rect 354289 3290 354345 3292
rect 354369 3290 354425 3292
rect 354449 3290 354505 3292
rect 354529 3290 354585 3292
rect 354289 3238 354315 3290
rect 354315 3238 354345 3290
rect 354369 3238 354379 3290
rect 354379 3238 354425 3290
rect 354449 3238 354495 3290
rect 354495 3238 354505 3290
rect 354529 3238 354559 3290
rect 354559 3238 354585 3290
rect 354289 3236 354345 3238
rect 354369 3236 354425 3238
rect 354449 3236 354505 3238
rect 354529 3236 354585 3238
rect 354289 2202 354345 2204
rect 354369 2202 354425 2204
rect 354449 2202 354505 2204
rect 354529 2202 354585 2204
rect 354289 2150 354315 2202
rect 354315 2150 354345 2202
rect 354369 2150 354379 2202
rect 354379 2150 354425 2202
rect 354449 2150 354495 2202
rect 354495 2150 354505 2202
rect 354529 2150 354559 2202
rect 354559 2150 354585 2202
rect 354289 2148 354345 2150
rect 354369 2148 354425 2150
rect 354449 2148 354505 2150
rect 354529 2148 354585 2150
rect 381266 1944 381322 2000
rect 423586 1264 423642 1320
rect 423494 176 423550 232
<< metal3 >>
rect 423520 9616 424000 9648
rect 423520 9560 423586 9616
rect 423642 9560 424000 9616
rect 423520 9528 424000 9560
rect 0 9208 480 9240
rect 0 9152 18 9208
rect 74 9152 480 9208
rect 0 9120 480 9152
rect 423520 8668 424000 8696
rect 423520 8666 423628 8668
rect 423500 8606 423628 8666
rect 423520 8604 423628 8606
rect 423692 8604 424000 8668
rect 423520 8576 424000 8604
rect 423520 7712 424000 7744
rect 423520 7656 423586 7712
rect 423642 7656 424000 7712
rect 71610 7648 71930 7649
rect 0 7576 480 7608
rect 71610 7584 71618 7648
rect 71682 7584 71698 7648
rect 71762 7584 71778 7648
rect 71842 7584 71858 7648
rect 71922 7584 71930 7648
rect 71610 7583 71930 7584
rect 212944 7648 213264 7649
rect 212944 7584 212952 7648
rect 213016 7584 213032 7648
rect 213096 7584 213112 7648
rect 213176 7584 213192 7648
rect 213256 7584 213264 7648
rect 212944 7583 213264 7584
rect 354277 7648 354597 7649
rect 354277 7584 354285 7648
rect 354349 7584 354365 7648
rect 354429 7584 354445 7648
rect 354509 7584 354525 7648
rect 354589 7584 354597 7648
rect 423520 7624 424000 7656
rect 354277 7583 354597 7584
rect 0 7520 110 7576
rect 166 7520 480 7576
rect 0 7488 480 7520
rect 142277 7104 142597 7105
rect 142277 7040 142285 7104
rect 142349 7040 142365 7104
rect 142429 7040 142445 7104
rect 142509 7040 142525 7104
rect 142589 7040 142597 7104
rect 142277 7039 142597 7040
rect 283610 7104 283930 7105
rect 283610 7040 283618 7104
rect 283682 7040 283698 7104
rect 283762 7040 283778 7104
rect 283842 7040 283858 7104
rect 283922 7040 283930 7104
rect 283610 7039 283930 7040
rect 132769 6898 132835 6901
rect 215293 6898 215359 6901
rect 132769 6896 215359 6898
rect 132769 6840 132774 6896
rect 132830 6840 215298 6896
rect 215354 6840 215359 6896
rect 132769 6838 215359 6840
rect 132769 6835 132835 6838
rect 215293 6835 215359 6838
rect 423520 6896 424000 6928
rect 423520 6840 423678 6896
rect 423734 6840 424000 6896
rect 423520 6808 424000 6840
rect 185761 6762 185827 6765
rect 202137 6762 202203 6765
rect 185761 6760 202203 6762
rect 185761 6704 185766 6760
rect 185822 6704 202142 6760
rect 202198 6704 202203 6760
rect 185761 6702 202203 6704
rect 185761 6699 185827 6702
rect 202137 6699 202203 6702
rect 216213 6762 216279 6765
rect 344553 6762 344619 6765
rect 216213 6760 344619 6762
rect 216213 6704 216218 6760
rect 216274 6704 344558 6760
rect 344614 6704 344619 6760
rect 216213 6702 344619 6704
rect 216213 6699 216279 6702
rect 344553 6699 344619 6702
rect 71610 6560 71930 6561
rect 71610 6496 71618 6560
rect 71682 6496 71698 6560
rect 71762 6496 71778 6560
rect 71842 6496 71858 6560
rect 71922 6496 71930 6560
rect 71610 6495 71930 6496
rect 212944 6560 213264 6561
rect 212944 6496 212952 6560
rect 213016 6496 213032 6560
rect 213096 6496 213112 6560
rect 213176 6496 213192 6560
rect 213256 6496 213264 6560
rect 212944 6495 213264 6496
rect 354277 6560 354597 6561
rect 354277 6496 354285 6560
rect 354349 6496 354365 6560
rect 354429 6496 354445 6560
rect 354509 6496 354525 6560
rect 354589 6496 354597 6560
rect 354277 6495 354597 6496
rect 399661 6354 399727 6357
rect 399661 6352 423690 6354
rect 399661 6296 399666 6352
rect 399722 6296 423690 6352
rect 399661 6294 423690 6296
rect 399661 6291 399727 6294
rect 215569 6218 215635 6221
rect 62 6216 215635 6218
rect 62 6160 215574 6216
rect 215630 6160 215635 6216
rect 62 6158 215635 6160
rect 62 5976 122 6158
rect 215569 6155 215635 6158
rect 142277 6016 142597 6017
rect 0 5856 480 5976
rect 142277 5952 142285 6016
rect 142349 5952 142365 6016
rect 142429 5952 142445 6016
rect 142509 5952 142525 6016
rect 142589 5952 142597 6016
rect 142277 5951 142597 5952
rect 283610 6016 283930 6017
rect 283610 5952 283618 6016
rect 283682 5952 283698 6016
rect 283762 5952 283778 6016
rect 283842 5952 283858 6016
rect 283922 5952 283930 6016
rect 423630 5976 423690 6294
rect 283610 5951 283930 5952
rect 423520 5856 424000 5976
rect 71610 5472 71930 5473
rect 71610 5408 71618 5472
rect 71682 5408 71698 5472
rect 71762 5408 71778 5472
rect 71842 5408 71858 5472
rect 71922 5408 71930 5472
rect 71610 5407 71930 5408
rect 212944 5472 213264 5473
rect 212944 5408 212952 5472
rect 213016 5408 213032 5472
rect 213096 5408 213112 5472
rect 213176 5408 213192 5472
rect 213256 5408 213264 5472
rect 212944 5407 213264 5408
rect 354277 5472 354597 5473
rect 354277 5408 354285 5472
rect 354349 5408 354365 5472
rect 354429 5408 354445 5472
rect 354509 5408 354525 5472
rect 354589 5408 354597 5472
rect 354277 5407 354597 5408
rect 105 5266 171 5269
rect 209497 5266 209563 5269
rect 105 5264 209563 5266
rect 105 5208 110 5264
rect 166 5208 209502 5264
rect 209558 5208 209563 5264
rect 105 5206 209563 5208
rect 105 5203 171 5206
rect 209497 5203 209563 5206
rect 235073 5266 235139 5269
rect 399661 5266 399727 5269
rect 235073 5264 399727 5266
rect 235073 5208 235078 5264
rect 235134 5208 399666 5264
rect 399722 5208 399727 5264
rect 235073 5206 399727 5208
rect 235073 5203 235139 5206
rect 399661 5203 399727 5206
rect 219801 5130 219867 5133
rect 232221 5130 232287 5133
rect 219801 5128 232287 5130
rect 219801 5072 219806 5128
rect 219862 5072 232226 5128
rect 232282 5072 232287 5128
rect 219801 5070 232287 5072
rect 219801 5067 219867 5070
rect 232221 5067 232287 5070
rect 142277 4928 142597 4929
rect 142277 4864 142285 4928
rect 142349 4864 142365 4928
rect 142429 4864 142445 4928
rect 142509 4864 142525 4928
rect 142589 4864 142597 4928
rect 142277 4863 142597 4864
rect 283610 4928 283930 4929
rect 283610 4864 283618 4928
rect 283682 4864 283698 4928
rect 283762 4864 283778 4928
rect 283842 4864 283858 4928
rect 283922 4864 283930 4928
rect 423520 4904 424000 5024
rect 283610 4863 283930 4864
rect 212993 4586 213059 4589
rect 423438 4586 423444 4588
rect 212993 4584 423444 4586
rect 212993 4528 212998 4584
rect 213054 4528 423444 4584
rect 212993 4526 423444 4528
rect 212993 4523 213059 4526
rect 423438 4524 423444 4526
rect 423508 4524 423514 4588
rect 71610 4384 71930 4385
rect 71610 4320 71618 4384
rect 71682 4320 71698 4384
rect 71762 4320 71778 4384
rect 71842 4320 71858 4384
rect 71922 4320 71930 4384
rect 71610 4319 71930 4320
rect 212944 4384 213264 4385
rect 212944 4320 212952 4384
rect 213016 4320 213032 4384
rect 213096 4320 213112 4384
rect 213176 4320 213192 4384
rect 213256 4320 213264 4384
rect 212944 4319 213264 4320
rect 354277 4384 354597 4385
rect 354277 4320 354285 4384
rect 354349 4320 354365 4384
rect 354429 4320 354445 4384
rect 354509 4320 354525 4384
rect 354589 4320 354597 4384
rect 354277 4319 354597 4320
rect 423630 4314 423690 4904
rect 415350 4254 423690 4314
rect 0 4176 480 4208
rect 0 4120 110 4176
rect 166 4120 480 4176
rect 0 4088 480 4120
rect 237373 4178 237439 4181
rect 415350 4178 415410 4254
rect 237373 4176 415410 4178
rect 237373 4120 237378 4176
rect 237434 4120 415410 4176
rect 237373 4118 415410 4120
rect 237373 4115 237439 4118
rect 220261 4042 220327 4045
rect 223205 4042 223271 4045
rect 220261 4040 223271 4042
rect 220261 3984 220266 4040
rect 220322 3984 223210 4040
rect 223266 3984 223271 4040
rect 220261 3982 223271 3984
rect 220261 3979 220327 3982
rect 223205 3979 223271 3982
rect 423520 3952 424000 4072
rect 142277 3840 142597 3841
rect 142277 3776 142285 3840
rect 142349 3776 142365 3840
rect 142429 3776 142445 3840
rect 142509 3776 142525 3840
rect 142589 3776 142597 3840
rect 142277 3775 142597 3776
rect 283610 3840 283930 3841
rect 283610 3776 283618 3840
rect 283682 3776 283698 3840
rect 283762 3776 283778 3840
rect 283842 3776 283858 3840
rect 283922 3776 283930 3840
rect 283610 3775 283930 3776
rect 225965 3634 226031 3637
rect 234521 3634 234587 3637
rect 225965 3632 234587 3634
rect 225965 3576 225970 3632
rect 226026 3576 234526 3632
rect 234582 3576 234587 3632
rect 225965 3574 234587 3576
rect 225965 3571 226031 3574
rect 234521 3571 234587 3574
rect 224861 3498 224927 3501
rect 289445 3498 289511 3501
rect 423630 3498 423690 3952
rect 224861 3496 289511 3498
rect 224861 3440 224866 3496
rect 224922 3440 289450 3496
rect 289506 3440 289511 3496
rect 224861 3438 289511 3440
rect 224861 3435 224927 3438
rect 289445 3435 289511 3438
rect 415350 3438 423690 3498
rect 216213 3362 216279 3365
rect 296437 3362 296503 3365
rect 415350 3362 415410 3438
rect 216213 3360 296503 3362
rect 216213 3304 216218 3360
rect 216274 3304 296442 3360
rect 296498 3304 296503 3360
rect 216213 3302 296503 3304
rect 216213 3299 216279 3302
rect 296437 3299 296503 3302
rect 409830 3302 415410 3362
rect 71610 3296 71930 3297
rect 71610 3232 71618 3296
rect 71682 3232 71698 3296
rect 71762 3232 71778 3296
rect 71842 3232 71858 3296
rect 71922 3232 71930 3296
rect 71610 3231 71930 3232
rect 212944 3296 213264 3297
rect 212944 3232 212952 3296
rect 213016 3232 213032 3296
rect 213096 3232 213112 3296
rect 213176 3232 213192 3296
rect 213256 3232 213264 3296
rect 212944 3231 213264 3232
rect 354277 3296 354597 3297
rect 354277 3232 354285 3296
rect 354349 3232 354365 3296
rect 354429 3232 354445 3296
rect 354509 3232 354525 3296
rect 354589 3232 354597 3296
rect 354277 3231 354597 3232
rect 289629 3090 289695 3093
rect 409830 3090 409890 3302
rect 423520 3136 424000 3256
rect 289629 3088 409890 3090
rect 289629 3032 289634 3088
rect 289690 3032 409890 3088
rect 289629 3030 409890 3032
rect 289629 3027 289695 3030
rect 238385 2954 238451 2957
rect 423630 2954 423690 3136
rect 238385 2952 423690 2954
rect 238385 2896 238390 2952
rect 238446 2896 423690 2952
rect 238385 2894 423690 2896
rect 238385 2891 238451 2894
rect 142277 2752 142597 2753
rect 142277 2688 142285 2752
rect 142349 2688 142365 2752
rect 142429 2688 142445 2752
rect 142509 2688 142525 2752
rect 142589 2688 142597 2752
rect 142277 2687 142597 2688
rect 283610 2752 283930 2753
rect 283610 2688 283618 2752
rect 283682 2688 283698 2752
rect 283762 2688 283778 2752
rect 283842 2688 283858 2752
rect 283922 2688 283930 2752
rect 283610 2687 283930 2688
rect 0 2456 480 2576
rect 62 1730 122 2456
rect 216622 2348 216628 2412
rect 216692 2410 216698 2412
rect 221089 2410 221155 2413
rect 216692 2408 221155 2410
rect 216692 2352 221094 2408
rect 221150 2352 221155 2408
rect 216692 2350 221155 2352
rect 216692 2348 216698 2350
rect 221089 2347 221155 2350
rect 71610 2208 71930 2209
rect 71610 2144 71618 2208
rect 71682 2144 71698 2208
rect 71762 2144 71778 2208
rect 71842 2144 71858 2208
rect 71922 2144 71930 2208
rect 71610 2143 71930 2144
rect 212944 2208 213264 2209
rect 212944 2144 212952 2208
rect 213016 2144 213032 2208
rect 213096 2144 213112 2208
rect 213176 2144 213192 2208
rect 213256 2144 213264 2208
rect 212944 2143 213264 2144
rect 354277 2208 354597 2209
rect 354277 2144 354285 2208
rect 354349 2144 354365 2208
rect 354429 2144 354445 2208
rect 354509 2144 354525 2208
rect 354589 2144 354597 2208
rect 423520 2184 424000 2304
rect 354277 2143 354597 2144
rect 215937 2002 216003 2005
rect 381261 2002 381327 2005
rect 215937 2000 381327 2002
rect 215937 1944 215942 2000
rect 215998 1944 381266 2000
rect 381322 1944 381327 2000
rect 215937 1942 381327 1944
rect 215937 1939 216003 1942
rect 381261 1939 381327 1942
rect 212349 1730 212415 1733
rect 62 1728 212415 1730
rect 62 1672 212354 1728
rect 212410 1672 212415 1728
rect 62 1670 212415 1672
rect 212349 1667 212415 1670
rect 42517 1594 42583 1597
rect 217593 1594 217659 1597
rect 42517 1592 217659 1594
rect 42517 1536 42522 1592
rect 42578 1536 217598 1592
rect 217654 1536 217659 1592
rect 42517 1534 217659 1536
rect 42517 1531 42583 1534
rect 217593 1531 217659 1534
rect 226149 1594 226215 1597
rect 423630 1594 423690 2184
rect 226149 1592 423690 1594
rect 226149 1536 226154 1592
rect 226210 1536 423690 1592
rect 226149 1534 423690 1536
rect 226149 1531 226215 1534
rect 423520 1320 424000 1352
rect 423520 1264 423586 1320
rect 423642 1264 424000 1320
rect 423520 1232 424000 1264
rect 214005 1186 214071 1189
rect 62 1184 214071 1186
rect 62 1128 214010 1184
rect 214066 1128 214071 1184
rect 62 1126 214071 1128
rect 62 944 122 1126
rect 214005 1123 214071 1126
rect 0 824 480 944
rect 423520 416 424000 536
rect 234245 234 234311 237
rect 423489 234 423555 237
rect 234245 232 423555 234
rect 234245 176 234250 232
rect 234306 176 423494 232
rect 423550 176 423555 232
rect 234245 174 423555 176
rect 234245 171 234311 174
rect 423489 171 423555 174
rect 127065 98 127131 101
rect 127198 98 127204 100
rect 127065 96 127204 98
rect 127065 40 127070 96
rect 127126 40 127204 96
rect 127065 38 127204 40
rect 127065 35 127131 38
rect 127198 36 127204 38
rect 127268 36 127274 100
rect 225873 98 225939 101
rect 423630 98 423690 416
rect 225873 96 423690 98
rect 225873 40 225878 96
rect 225934 40 423690 96
rect 225873 38 423690 40
rect 225873 35 225939 38
<< via3 >>
rect 423628 8604 423692 8668
rect 71618 7644 71682 7648
rect 71618 7588 71622 7644
rect 71622 7588 71678 7644
rect 71678 7588 71682 7644
rect 71618 7584 71682 7588
rect 71698 7644 71762 7648
rect 71698 7588 71702 7644
rect 71702 7588 71758 7644
rect 71758 7588 71762 7644
rect 71698 7584 71762 7588
rect 71778 7644 71842 7648
rect 71778 7588 71782 7644
rect 71782 7588 71838 7644
rect 71838 7588 71842 7644
rect 71778 7584 71842 7588
rect 71858 7644 71922 7648
rect 71858 7588 71862 7644
rect 71862 7588 71918 7644
rect 71918 7588 71922 7644
rect 71858 7584 71922 7588
rect 212952 7644 213016 7648
rect 212952 7588 212956 7644
rect 212956 7588 213012 7644
rect 213012 7588 213016 7644
rect 212952 7584 213016 7588
rect 213032 7644 213096 7648
rect 213032 7588 213036 7644
rect 213036 7588 213092 7644
rect 213092 7588 213096 7644
rect 213032 7584 213096 7588
rect 213112 7644 213176 7648
rect 213112 7588 213116 7644
rect 213116 7588 213172 7644
rect 213172 7588 213176 7644
rect 213112 7584 213176 7588
rect 213192 7644 213256 7648
rect 213192 7588 213196 7644
rect 213196 7588 213252 7644
rect 213252 7588 213256 7644
rect 213192 7584 213256 7588
rect 354285 7644 354349 7648
rect 354285 7588 354289 7644
rect 354289 7588 354345 7644
rect 354345 7588 354349 7644
rect 354285 7584 354349 7588
rect 354365 7644 354429 7648
rect 354365 7588 354369 7644
rect 354369 7588 354425 7644
rect 354425 7588 354429 7644
rect 354365 7584 354429 7588
rect 354445 7644 354509 7648
rect 354445 7588 354449 7644
rect 354449 7588 354505 7644
rect 354505 7588 354509 7644
rect 354445 7584 354509 7588
rect 354525 7644 354589 7648
rect 354525 7588 354529 7644
rect 354529 7588 354585 7644
rect 354585 7588 354589 7644
rect 354525 7584 354589 7588
rect 142285 7100 142349 7104
rect 142285 7044 142289 7100
rect 142289 7044 142345 7100
rect 142345 7044 142349 7100
rect 142285 7040 142349 7044
rect 142365 7100 142429 7104
rect 142365 7044 142369 7100
rect 142369 7044 142425 7100
rect 142425 7044 142429 7100
rect 142365 7040 142429 7044
rect 142445 7100 142509 7104
rect 142445 7044 142449 7100
rect 142449 7044 142505 7100
rect 142505 7044 142509 7100
rect 142445 7040 142509 7044
rect 142525 7100 142589 7104
rect 142525 7044 142529 7100
rect 142529 7044 142585 7100
rect 142585 7044 142589 7100
rect 142525 7040 142589 7044
rect 283618 7100 283682 7104
rect 283618 7044 283622 7100
rect 283622 7044 283678 7100
rect 283678 7044 283682 7100
rect 283618 7040 283682 7044
rect 283698 7100 283762 7104
rect 283698 7044 283702 7100
rect 283702 7044 283758 7100
rect 283758 7044 283762 7100
rect 283698 7040 283762 7044
rect 283778 7100 283842 7104
rect 283778 7044 283782 7100
rect 283782 7044 283838 7100
rect 283838 7044 283842 7100
rect 283778 7040 283842 7044
rect 283858 7100 283922 7104
rect 283858 7044 283862 7100
rect 283862 7044 283918 7100
rect 283918 7044 283922 7100
rect 283858 7040 283922 7044
rect 71618 6556 71682 6560
rect 71618 6500 71622 6556
rect 71622 6500 71678 6556
rect 71678 6500 71682 6556
rect 71618 6496 71682 6500
rect 71698 6556 71762 6560
rect 71698 6500 71702 6556
rect 71702 6500 71758 6556
rect 71758 6500 71762 6556
rect 71698 6496 71762 6500
rect 71778 6556 71842 6560
rect 71778 6500 71782 6556
rect 71782 6500 71838 6556
rect 71838 6500 71842 6556
rect 71778 6496 71842 6500
rect 71858 6556 71922 6560
rect 71858 6500 71862 6556
rect 71862 6500 71918 6556
rect 71918 6500 71922 6556
rect 71858 6496 71922 6500
rect 212952 6556 213016 6560
rect 212952 6500 212956 6556
rect 212956 6500 213012 6556
rect 213012 6500 213016 6556
rect 212952 6496 213016 6500
rect 213032 6556 213096 6560
rect 213032 6500 213036 6556
rect 213036 6500 213092 6556
rect 213092 6500 213096 6556
rect 213032 6496 213096 6500
rect 213112 6556 213176 6560
rect 213112 6500 213116 6556
rect 213116 6500 213172 6556
rect 213172 6500 213176 6556
rect 213112 6496 213176 6500
rect 213192 6556 213256 6560
rect 213192 6500 213196 6556
rect 213196 6500 213252 6556
rect 213252 6500 213256 6556
rect 213192 6496 213256 6500
rect 354285 6556 354349 6560
rect 354285 6500 354289 6556
rect 354289 6500 354345 6556
rect 354345 6500 354349 6556
rect 354285 6496 354349 6500
rect 354365 6556 354429 6560
rect 354365 6500 354369 6556
rect 354369 6500 354425 6556
rect 354425 6500 354429 6556
rect 354365 6496 354429 6500
rect 354445 6556 354509 6560
rect 354445 6500 354449 6556
rect 354449 6500 354505 6556
rect 354505 6500 354509 6556
rect 354445 6496 354509 6500
rect 354525 6556 354589 6560
rect 354525 6500 354529 6556
rect 354529 6500 354585 6556
rect 354585 6500 354589 6556
rect 354525 6496 354589 6500
rect 142285 6012 142349 6016
rect 142285 5956 142289 6012
rect 142289 5956 142345 6012
rect 142345 5956 142349 6012
rect 142285 5952 142349 5956
rect 142365 6012 142429 6016
rect 142365 5956 142369 6012
rect 142369 5956 142425 6012
rect 142425 5956 142429 6012
rect 142365 5952 142429 5956
rect 142445 6012 142509 6016
rect 142445 5956 142449 6012
rect 142449 5956 142505 6012
rect 142505 5956 142509 6012
rect 142445 5952 142509 5956
rect 142525 6012 142589 6016
rect 142525 5956 142529 6012
rect 142529 5956 142585 6012
rect 142585 5956 142589 6012
rect 142525 5952 142589 5956
rect 283618 6012 283682 6016
rect 283618 5956 283622 6012
rect 283622 5956 283678 6012
rect 283678 5956 283682 6012
rect 283618 5952 283682 5956
rect 283698 6012 283762 6016
rect 283698 5956 283702 6012
rect 283702 5956 283758 6012
rect 283758 5956 283762 6012
rect 283698 5952 283762 5956
rect 283778 6012 283842 6016
rect 283778 5956 283782 6012
rect 283782 5956 283838 6012
rect 283838 5956 283842 6012
rect 283778 5952 283842 5956
rect 283858 6012 283922 6016
rect 283858 5956 283862 6012
rect 283862 5956 283918 6012
rect 283918 5956 283922 6012
rect 283858 5952 283922 5956
rect 71618 5468 71682 5472
rect 71618 5412 71622 5468
rect 71622 5412 71678 5468
rect 71678 5412 71682 5468
rect 71618 5408 71682 5412
rect 71698 5468 71762 5472
rect 71698 5412 71702 5468
rect 71702 5412 71758 5468
rect 71758 5412 71762 5468
rect 71698 5408 71762 5412
rect 71778 5468 71842 5472
rect 71778 5412 71782 5468
rect 71782 5412 71838 5468
rect 71838 5412 71842 5468
rect 71778 5408 71842 5412
rect 71858 5468 71922 5472
rect 71858 5412 71862 5468
rect 71862 5412 71918 5468
rect 71918 5412 71922 5468
rect 71858 5408 71922 5412
rect 212952 5468 213016 5472
rect 212952 5412 212956 5468
rect 212956 5412 213012 5468
rect 213012 5412 213016 5468
rect 212952 5408 213016 5412
rect 213032 5468 213096 5472
rect 213032 5412 213036 5468
rect 213036 5412 213092 5468
rect 213092 5412 213096 5468
rect 213032 5408 213096 5412
rect 213112 5468 213176 5472
rect 213112 5412 213116 5468
rect 213116 5412 213172 5468
rect 213172 5412 213176 5468
rect 213112 5408 213176 5412
rect 213192 5468 213256 5472
rect 213192 5412 213196 5468
rect 213196 5412 213252 5468
rect 213252 5412 213256 5468
rect 213192 5408 213256 5412
rect 354285 5468 354349 5472
rect 354285 5412 354289 5468
rect 354289 5412 354345 5468
rect 354345 5412 354349 5468
rect 354285 5408 354349 5412
rect 354365 5468 354429 5472
rect 354365 5412 354369 5468
rect 354369 5412 354425 5468
rect 354425 5412 354429 5468
rect 354365 5408 354429 5412
rect 354445 5468 354509 5472
rect 354445 5412 354449 5468
rect 354449 5412 354505 5468
rect 354505 5412 354509 5468
rect 354445 5408 354509 5412
rect 354525 5468 354589 5472
rect 354525 5412 354529 5468
rect 354529 5412 354585 5468
rect 354585 5412 354589 5468
rect 354525 5408 354589 5412
rect 142285 4924 142349 4928
rect 142285 4868 142289 4924
rect 142289 4868 142345 4924
rect 142345 4868 142349 4924
rect 142285 4864 142349 4868
rect 142365 4924 142429 4928
rect 142365 4868 142369 4924
rect 142369 4868 142425 4924
rect 142425 4868 142429 4924
rect 142365 4864 142429 4868
rect 142445 4924 142509 4928
rect 142445 4868 142449 4924
rect 142449 4868 142505 4924
rect 142505 4868 142509 4924
rect 142445 4864 142509 4868
rect 142525 4924 142589 4928
rect 142525 4868 142529 4924
rect 142529 4868 142585 4924
rect 142585 4868 142589 4924
rect 142525 4864 142589 4868
rect 283618 4924 283682 4928
rect 283618 4868 283622 4924
rect 283622 4868 283678 4924
rect 283678 4868 283682 4924
rect 283618 4864 283682 4868
rect 283698 4924 283762 4928
rect 283698 4868 283702 4924
rect 283702 4868 283758 4924
rect 283758 4868 283762 4924
rect 283698 4864 283762 4868
rect 283778 4924 283842 4928
rect 283778 4868 283782 4924
rect 283782 4868 283838 4924
rect 283838 4868 283842 4924
rect 283778 4864 283842 4868
rect 283858 4924 283922 4928
rect 283858 4868 283862 4924
rect 283862 4868 283918 4924
rect 283918 4868 283922 4924
rect 283858 4864 283922 4868
rect 423444 4524 423508 4588
rect 71618 4380 71682 4384
rect 71618 4324 71622 4380
rect 71622 4324 71678 4380
rect 71678 4324 71682 4380
rect 71618 4320 71682 4324
rect 71698 4380 71762 4384
rect 71698 4324 71702 4380
rect 71702 4324 71758 4380
rect 71758 4324 71762 4380
rect 71698 4320 71762 4324
rect 71778 4380 71842 4384
rect 71778 4324 71782 4380
rect 71782 4324 71838 4380
rect 71838 4324 71842 4380
rect 71778 4320 71842 4324
rect 71858 4380 71922 4384
rect 71858 4324 71862 4380
rect 71862 4324 71918 4380
rect 71918 4324 71922 4380
rect 71858 4320 71922 4324
rect 212952 4380 213016 4384
rect 212952 4324 212956 4380
rect 212956 4324 213012 4380
rect 213012 4324 213016 4380
rect 212952 4320 213016 4324
rect 213032 4380 213096 4384
rect 213032 4324 213036 4380
rect 213036 4324 213092 4380
rect 213092 4324 213096 4380
rect 213032 4320 213096 4324
rect 213112 4380 213176 4384
rect 213112 4324 213116 4380
rect 213116 4324 213172 4380
rect 213172 4324 213176 4380
rect 213112 4320 213176 4324
rect 213192 4380 213256 4384
rect 213192 4324 213196 4380
rect 213196 4324 213252 4380
rect 213252 4324 213256 4380
rect 213192 4320 213256 4324
rect 354285 4380 354349 4384
rect 354285 4324 354289 4380
rect 354289 4324 354345 4380
rect 354345 4324 354349 4380
rect 354285 4320 354349 4324
rect 354365 4380 354429 4384
rect 354365 4324 354369 4380
rect 354369 4324 354425 4380
rect 354425 4324 354429 4380
rect 354365 4320 354429 4324
rect 354445 4380 354509 4384
rect 354445 4324 354449 4380
rect 354449 4324 354505 4380
rect 354505 4324 354509 4380
rect 354445 4320 354509 4324
rect 354525 4380 354589 4384
rect 354525 4324 354529 4380
rect 354529 4324 354585 4380
rect 354585 4324 354589 4380
rect 354525 4320 354589 4324
rect 142285 3836 142349 3840
rect 142285 3780 142289 3836
rect 142289 3780 142345 3836
rect 142345 3780 142349 3836
rect 142285 3776 142349 3780
rect 142365 3836 142429 3840
rect 142365 3780 142369 3836
rect 142369 3780 142425 3836
rect 142425 3780 142429 3836
rect 142365 3776 142429 3780
rect 142445 3836 142509 3840
rect 142445 3780 142449 3836
rect 142449 3780 142505 3836
rect 142505 3780 142509 3836
rect 142445 3776 142509 3780
rect 142525 3836 142589 3840
rect 142525 3780 142529 3836
rect 142529 3780 142585 3836
rect 142585 3780 142589 3836
rect 142525 3776 142589 3780
rect 283618 3836 283682 3840
rect 283618 3780 283622 3836
rect 283622 3780 283678 3836
rect 283678 3780 283682 3836
rect 283618 3776 283682 3780
rect 283698 3836 283762 3840
rect 283698 3780 283702 3836
rect 283702 3780 283758 3836
rect 283758 3780 283762 3836
rect 283698 3776 283762 3780
rect 283778 3836 283842 3840
rect 283778 3780 283782 3836
rect 283782 3780 283838 3836
rect 283838 3780 283842 3836
rect 283778 3776 283842 3780
rect 283858 3836 283922 3840
rect 283858 3780 283862 3836
rect 283862 3780 283918 3836
rect 283918 3780 283922 3836
rect 283858 3776 283922 3780
rect 71618 3292 71682 3296
rect 71618 3236 71622 3292
rect 71622 3236 71678 3292
rect 71678 3236 71682 3292
rect 71618 3232 71682 3236
rect 71698 3292 71762 3296
rect 71698 3236 71702 3292
rect 71702 3236 71758 3292
rect 71758 3236 71762 3292
rect 71698 3232 71762 3236
rect 71778 3292 71842 3296
rect 71778 3236 71782 3292
rect 71782 3236 71838 3292
rect 71838 3236 71842 3292
rect 71778 3232 71842 3236
rect 71858 3292 71922 3296
rect 71858 3236 71862 3292
rect 71862 3236 71918 3292
rect 71918 3236 71922 3292
rect 71858 3232 71922 3236
rect 212952 3292 213016 3296
rect 212952 3236 212956 3292
rect 212956 3236 213012 3292
rect 213012 3236 213016 3292
rect 212952 3232 213016 3236
rect 213032 3292 213096 3296
rect 213032 3236 213036 3292
rect 213036 3236 213092 3292
rect 213092 3236 213096 3292
rect 213032 3232 213096 3236
rect 213112 3292 213176 3296
rect 213112 3236 213116 3292
rect 213116 3236 213172 3292
rect 213172 3236 213176 3292
rect 213112 3232 213176 3236
rect 213192 3292 213256 3296
rect 213192 3236 213196 3292
rect 213196 3236 213252 3292
rect 213252 3236 213256 3292
rect 213192 3232 213256 3236
rect 354285 3292 354349 3296
rect 354285 3236 354289 3292
rect 354289 3236 354345 3292
rect 354345 3236 354349 3292
rect 354285 3232 354349 3236
rect 354365 3292 354429 3296
rect 354365 3236 354369 3292
rect 354369 3236 354425 3292
rect 354425 3236 354429 3292
rect 354365 3232 354429 3236
rect 354445 3292 354509 3296
rect 354445 3236 354449 3292
rect 354449 3236 354505 3292
rect 354505 3236 354509 3292
rect 354445 3232 354509 3236
rect 354525 3292 354589 3296
rect 354525 3236 354529 3292
rect 354529 3236 354585 3292
rect 354585 3236 354589 3292
rect 354525 3232 354589 3236
rect 142285 2748 142349 2752
rect 142285 2692 142289 2748
rect 142289 2692 142345 2748
rect 142345 2692 142349 2748
rect 142285 2688 142349 2692
rect 142365 2748 142429 2752
rect 142365 2692 142369 2748
rect 142369 2692 142425 2748
rect 142425 2692 142429 2748
rect 142365 2688 142429 2692
rect 142445 2748 142509 2752
rect 142445 2692 142449 2748
rect 142449 2692 142505 2748
rect 142505 2692 142509 2748
rect 142445 2688 142509 2692
rect 142525 2748 142589 2752
rect 142525 2692 142529 2748
rect 142529 2692 142585 2748
rect 142585 2692 142589 2748
rect 142525 2688 142589 2692
rect 283618 2748 283682 2752
rect 283618 2692 283622 2748
rect 283622 2692 283678 2748
rect 283678 2692 283682 2748
rect 283618 2688 283682 2692
rect 283698 2748 283762 2752
rect 283698 2692 283702 2748
rect 283702 2692 283758 2748
rect 283758 2692 283762 2748
rect 283698 2688 283762 2692
rect 283778 2748 283842 2752
rect 283778 2692 283782 2748
rect 283782 2692 283838 2748
rect 283838 2692 283842 2748
rect 283778 2688 283842 2692
rect 283858 2748 283922 2752
rect 283858 2692 283862 2748
rect 283862 2692 283918 2748
rect 283918 2692 283922 2748
rect 283858 2688 283922 2692
rect 216628 2348 216692 2412
rect 71618 2204 71682 2208
rect 71618 2148 71622 2204
rect 71622 2148 71678 2204
rect 71678 2148 71682 2204
rect 71618 2144 71682 2148
rect 71698 2204 71762 2208
rect 71698 2148 71702 2204
rect 71702 2148 71758 2204
rect 71758 2148 71762 2204
rect 71698 2144 71762 2148
rect 71778 2204 71842 2208
rect 71778 2148 71782 2204
rect 71782 2148 71838 2204
rect 71838 2148 71842 2204
rect 71778 2144 71842 2148
rect 71858 2204 71922 2208
rect 71858 2148 71862 2204
rect 71862 2148 71918 2204
rect 71918 2148 71922 2204
rect 71858 2144 71922 2148
rect 212952 2204 213016 2208
rect 212952 2148 212956 2204
rect 212956 2148 213012 2204
rect 213012 2148 213016 2204
rect 212952 2144 213016 2148
rect 213032 2204 213096 2208
rect 213032 2148 213036 2204
rect 213036 2148 213092 2204
rect 213092 2148 213096 2204
rect 213032 2144 213096 2148
rect 213112 2204 213176 2208
rect 213112 2148 213116 2204
rect 213116 2148 213172 2204
rect 213172 2148 213176 2204
rect 213112 2144 213176 2148
rect 213192 2204 213256 2208
rect 213192 2148 213196 2204
rect 213196 2148 213252 2204
rect 213252 2148 213256 2204
rect 213192 2144 213256 2148
rect 354285 2204 354349 2208
rect 354285 2148 354289 2204
rect 354289 2148 354345 2204
rect 354345 2148 354349 2204
rect 354285 2144 354349 2148
rect 354365 2204 354429 2208
rect 354365 2148 354369 2204
rect 354369 2148 354425 2204
rect 354425 2148 354429 2204
rect 354365 2144 354429 2148
rect 354445 2204 354509 2208
rect 354445 2148 354449 2204
rect 354449 2148 354505 2204
rect 354505 2148 354509 2204
rect 354445 2144 354509 2148
rect 354525 2204 354589 2208
rect 354525 2148 354529 2204
rect 354529 2148 354585 2204
rect 354585 2148 354589 2204
rect 354525 2144 354589 2148
rect 127204 36 127268 100
<< metal4 >>
rect 423627 8668 423693 8669
rect 423627 8666 423628 8668
rect 423446 8606 423628 8666
rect 71610 7648 71931 7664
rect 71610 7584 71618 7648
rect 71682 7584 71698 7648
rect 71762 7584 71778 7648
rect 71842 7584 71858 7648
rect 71922 7584 71931 7648
rect 71610 6560 71931 7584
rect 71610 6496 71618 6560
rect 71682 6496 71698 6560
rect 71762 6496 71778 6560
rect 71842 6496 71858 6560
rect 71922 6496 71931 6560
rect 71610 5472 71931 6496
rect 71610 5408 71618 5472
rect 71682 5408 71698 5472
rect 71762 5408 71778 5472
rect 71842 5408 71858 5472
rect 71922 5408 71931 5472
rect 71610 4384 71931 5408
rect 71610 4320 71618 4384
rect 71682 4320 71698 4384
rect 71762 4320 71778 4384
rect 71842 4320 71858 4384
rect 71922 4320 71931 4384
rect 71610 3296 71931 4320
rect 71610 3232 71618 3296
rect 71682 3232 71698 3296
rect 71762 3232 71778 3296
rect 71842 3232 71858 3296
rect 71922 3232 71931 3296
rect 71610 2208 71931 3232
rect 142277 7104 142597 7664
rect 142277 7040 142285 7104
rect 142349 7040 142365 7104
rect 142429 7040 142445 7104
rect 142509 7040 142525 7104
rect 142589 7040 142597 7104
rect 142277 6016 142597 7040
rect 142277 5952 142285 6016
rect 142349 5952 142365 6016
rect 142429 5952 142445 6016
rect 142509 5952 142525 6016
rect 142589 5952 142597 6016
rect 142277 4928 142597 5952
rect 142277 4864 142285 4928
rect 142349 4864 142365 4928
rect 142429 4864 142445 4928
rect 142509 4864 142525 4928
rect 142589 4864 142597 4928
rect 142277 3840 142597 4864
rect 142277 3776 142285 3840
rect 142349 3776 142365 3840
rect 142429 3776 142445 3840
rect 142509 3776 142525 3840
rect 142589 3776 142597 3840
rect 142277 2752 142597 3776
rect 142277 2688 142285 2752
rect 142349 2688 142365 2752
rect 142429 2688 142445 2752
rect 142509 2688 142525 2752
rect 142589 2688 142597 2752
rect 71610 2144 71618 2208
rect 71682 2144 71698 2208
rect 71762 2144 71778 2208
rect 71842 2144 71858 2208
rect 71922 2144 71931 2208
rect 71610 2128 71931 2144
rect 127206 101 127266 2262
rect 142277 2128 142597 2688
rect 212944 7648 213264 7664
rect 212944 7584 212952 7648
rect 213016 7584 213032 7648
rect 213096 7584 213112 7648
rect 213176 7584 213192 7648
rect 213256 7584 213264 7648
rect 212944 6560 213264 7584
rect 212944 6496 212952 6560
rect 213016 6496 213032 6560
rect 213096 6496 213112 6560
rect 213176 6496 213192 6560
rect 213256 6496 213264 6560
rect 212944 5472 213264 6496
rect 212944 5408 212952 5472
rect 213016 5408 213032 5472
rect 213096 5408 213112 5472
rect 213176 5408 213192 5472
rect 213256 5408 213264 5472
rect 212944 4384 213264 5408
rect 212944 4320 212952 4384
rect 213016 4320 213032 4384
rect 213096 4320 213112 4384
rect 213176 4320 213192 4384
rect 213256 4320 213264 4384
rect 212944 3296 213264 4320
rect 212944 3232 212952 3296
rect 213016 3232 213032 3296
rect 213096 3232 213112 3296
rect 213176 3232 213192 3296
rect 213256 3232 213264 3296
rect 212944 2208 213264 3232
rect 283610 7104 283930 7664
rect 283610 7040 283618 7104
rect 283682 7040 283698 7104
rect 283762 7040 283778 7104
rect 283842 7040 283858 7104
rect 283922 7040 283930 7104
rect 283610 6016 283930 7040
rect 283610 5952 283618 6016
rect 283682 5952 283698 6016
rect 283762 5952 283778 6016
rect 283842 5952 283858 6016
rect 283922 5952 283930 6016
rect 283610 4928 283930 5952
rect 283610 4864 283618 4928
rect 283682 4864 283698 4928
rect 283762 4864 283778 4928
rect 283842 4864 283858 4928
rect 283922 4864 283930 4928
rect 283610 3840 283930 4864
rect 283610 3776 283618 3840
rect 283682 3776 283698 3840
rect 283762 3776 283778 3840
rect 283842 3776 283858 3840
rect 283922 3776 283930 3840
rect 283610 2752 283930 3776
rect 283610 2688 283618 2752
rect 283682 2688 283698 2752
rect 283762 2688 283778 2752
rect 283842 2688 283858 2752
rect 283922 2688 283930 2752
rect 212944 2144 212952 2208
rect 213016 2144 213032 2208
rect 213096 2144 213112 2208
rect 213176 2144 213192 2208
rect 213256 2144 213264 2208
rect 212944 2128 213264 2144
rect 283610 2128 283930 2688
rect 354277 7648 354597 7664
rect 354277 7584 354285 7648
rect 354349 7584 354365 7648
rect 354429 7584 354445 7648
rect 354509 7584 354525 7648
rect 354589 7584 354597 7648
rect 354277 6560 354597 7584
rect 354277 6496 354285 6560
rect 354349 6496 354365 6560
rect 354429 6496 354445 6560
rect 354509 6496 354525 6560
rect 354589 6496 354597 6560
rect 354277 5472 354597 6496
rect 354277 5408 354285 5472
rect 354349 5408 354365 5472
rect 354429 5408 354445 5472
rect 354509 5408 354525 5472
rect 354589 5408 354597 5472
rect 354277 4384 354597 5408
rect 423446 4589 423506 8606
rect 423627 8604 423628 8606
rect 423692 8604 423693 8668
rect 423627 8603 423693 8604
rect 423443 4588 423509 4589
rect 423443 4524 423444 4588
rect 423508 4524 423509 4588
rect 423443 4523 423509 4524
rect 354277 4320 354285 4384
rect 354349 4320 354365 4384
rect 354429 4320 354445 4384
rect 354509 4320 354525 4384
rect 354589 4320 354597 4384
rect 354277 3296 354597 4320
rect 354277 3232 354285 3296
rect 354349 3232 354365 3296
rect 354429 3232 354445 3296
rect 354509 3232 354525 3296
rect 354589 3232 354597 3296
rect 354277 2208 354597 3232
rect 354277 2144 354285 2208
rect 354349 2144 354365 2208
rect 354429 2144 354445 2208
rect 354509 2144 354525 2208
rect 354589 2144 354597 2208
rect 354277 2128 354597 2144
rect 127203 100 127269 101
rect 127203 36 127204 100
rect 127268 36 127269 100
rect 127203 35 127269 36
<< via4 >>
rect 127118 2262 127354 2498
rect 216542 2412 216778 2498
rect 216542 2348 216628 2412
rect 216628 2348 216692 2412
rect 216692 2348 216778 2412
rect 216542 2262 216778 2348
<< metal5 >>
rect 127076 2498 216820 2540
rect 127076 2262 127118 2498
rect 127354 2262 216542 2498
rect 216778 2262 216820 2498
rect 127076 2220 216820 2262
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_20 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_39
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_51 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_21
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_59 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_87
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_22
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_23
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_118
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_24
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_25
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_26
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_27
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_261
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_28
timestamp 1586364061
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_280
timestamp 1586364061
transform 1 0 26864 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_281
timestamp 1586364061
transform 1 0 26956 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_292
timestamp 1586364061
transform 1 0 27968 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_293
timestamp 1586364061
transform 1 0 28060 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_29
timestamp 1586364061
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_304
timestamp 1586364061
transform 1 0 29072 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_311
timestamp 1586364061
transform 1 0 29716 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_306
timestamp 1586364061
transform 1 0 29256 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_318
timestamp 1586364061
transform 1 0 30360 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_323
timestamp 1586364061
transform 1 0 30820 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_335
timestamp 1586364061
transform 1 0 31924 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_330
timestamp 1586364061
transform 1 0 31464 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_30
timestamp 1586364061
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_342
timestamp 1586364061
transform 1 0 32568 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_354
timestamp 1586364061
transform 1 0 33672 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_342
timestamp 1586364061
transform 1 0 32568 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_354
timestamp 1586364061
transform 1 0 33672 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_31
timestamp 1586364061
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_366
timestamp 1586364061
transform 1 0 34776 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_373
timestamp 1586364061
transform 1 0 35420 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_367
timestamp 1586364061
transform 1 0 34868 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_385
timestamp 1586364061
transform 1 0 36524 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_379
timestamp 1586364061
transform 1 0 35972 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_391
timestamp 1586364061
transform 1 0 37076 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_32
timestamp 1586364061
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_397
timestamp 1586364061
transform 1 0 37628 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_404
timestamp 1586364061
transform 1 0 38272 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_403
timestamp 1586364061
transform 1 0 38180 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 40388 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_416
timestamp 1586364061
transform 1 0 39376 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_428
timestamp 1586364061
transform 1 0 40480 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_415
timestamp 1586364061
transform 1 0 39284 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_428
timestamp 1586364061
transform 1 0 40480 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_33
timestamp 1586364061
transform 1 0 41032 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_435
timestamp 1586364061
transform 1 0 41124 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_440
timestamp 1586364061
transform 1 0 41584 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_447
timestamp 1586364061
transform 1 0 42228 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_459
timestamp 1586364061
transform 1 0 43332 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_452
timestamp 1586364061
transform 1 0 42688 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_34
timestamp 1586364061
transform 1 0 43884 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_466
timestamp 1586364061
transform 1 0 43976 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_478
timestamp 1586364061
transform 1 0 45080 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_464
timestamp 1586364061
transform 1 0 43792 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_476
timestamp 1586364061
transform 1 0 44896 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_35
timestamp 1586364061
transform 1 0 46736 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 46000 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_490
timestamp 1586364061
transform 1 0 46184 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_497
timestamp 1586364061
transform 1 0 46828 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_489
timestamp 1586364061
transform 1 0 46092 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_509
timestamp 1586364061
transform 1 0 47932 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_501
timestamp 1586364061
transform 1 0 47196 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_513
timestamp 1586364061
transform 1 0 48300 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_36
timestamp 1586364061
transform 1 0 49588 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_521
timestamp 1586364061
transform 1 0 49036 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_528
timestamp 1586364061
transform 1 0 49680 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_525
timestamp 1586364061
transform 1 0 49404 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 51612 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_540
timestamp 1586364061
transform 1 0 50784 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_552
timestamp 1586364061
transform 1 0 51888 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_537
timestamp 1586364061
transform 1 0 50508 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_550
timestamp 1586364061
transform 1 0 51704 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_37
timestamp 1586364061
transform 1 0 52440 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_559
timestamp 1586364061
transform 1 0 52532 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_562
timestamp 1586364061
transform 1 0 52808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_571
timestamp 1586364061
transform 1 0 53636 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_583
timestamp 1586364061
transform 1 0 54740 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_574
timestamp 1586364061
transform 1 0 53912 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_586
timestamp 1586364061
transform 1 0 55016 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_38
timestamp 1586364061
transform 1 0 55292 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_590
timestamp 1586364061
transform 1 0 55384 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_602
timestamp 1586364061
transform 1 0 56488 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_598
timestamp 1586364061
transform 1 0 56120 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_39
timestamp 1586364061
transform 1 0 58144 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 57224 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_614
timestamp 1586364061
transform 1 0 57592 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_621
timestamp 1586364061
transform 1 0 58236 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_611
timestamp 1586364061
transform 1 0 57316 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_623
timestamp 1586364061
transform 1 0 58420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_633
timestamp 1586364061
transform 1 0 59340 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_635
timestamp 1586364061
transform 1 0 59524 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_40
timestamp 1586364061
transform 1 0 60996 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_645
timestamp 1586364061
transform 1 0 60444 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_652
timestamp 1586364061
transform 1 0 61088 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_647
timestamp 1586364061
transform 1 0 60628 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_659
timestamp 1586364061
transform 1 0 61732 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 62836 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_664
timestamp 1586364061
transform 1 0 62192 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_676
timestamp 1586364061
transform 1 0 63296 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_672
timestamp 1586364061
transform 1 0 62928 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_41
timestamp 1586364061
transform 1 0 63848 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_683
timestamp 1586364061
transform 1 0 63940 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_695
timestamp 1586364061
transform 1 0 65044 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_684
timestamp 1586364061
transform 1 0 64032 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_42
timestamp 1586364061
transform 1 0 66700 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_707
timestamp 1586364061
transform 1 0 66148 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_696
timestamp 1586364061
transform 1 0 65136 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_708
timestamp 1586364061
transform 1 0 66240 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_714
timestamp 1586364061
transform 1 0 66792 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_726
timestamp 1586364061
transform 1 0 67896 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_720
timestamp 1586364061
transform 1 0 67344 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_43
timestamp 1586364061
transform 1 0 69552 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 68448 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_738
timestamp 1586364061
transform 1 0 69000 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_745
timestamp 1586364061
transform 1 0 69644 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_733
timestamp 1586364061
transform 1 0 68540 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_745
timestamp 1586364061
transform 1 0 69644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_757
timestamp 1586364061
transform 1 0 70748 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_757
timestamp 1586364061
transform 1 0 70748 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_44
timestamp 1586364061
transform 1 0 72404 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_769
timestamp 1586364061
transform 1 0 71852 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_776
timestamp 1586364061
transform 1 0 72496 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_769
timestamp 1586364061
transform 1 0 71852 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_781
timestamp 1586364061
transform 1 0 72956 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 74060 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_788
timestamp 1586364061
transform 1 0 73600 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_800
timestamp 1586364061
transform 1 0 74704 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_794
timestamp 1586364061
transform 1 0 74152 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_45
timestamp 1586364061
transform 1 0 75256 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_807
timestamp 1586364061
transform 1 0 75348 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_819
timestamp 1586364061
transform 1 0 76452 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_806
timestamp 1586364061
transform 1 0 75256 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_818
timestamp 1586364061
transform 1 0 76360 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_46
timestamp 1586364061
transform 1 0 78108 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_831
timestamp 1586364061
transform 1 0 77556 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_838
timestamp 1586364061
transform 1 0 78200 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_830
timestamp 1586364061
transform 1 0 77464 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 79672 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_850
timestamp 1586364061
transform 1 0 79304 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_842
timestamp 1586364061
transform 1 0 78568 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_855
timestamp 1586364061
transform 1 0 79764 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_47
timestamp 1586364061
transform 1 0 80960 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_862
timestamp 1586364061
transform 1 0 80408 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_869
timestamp 1586364061
transform 1 0 81052 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_867
timestamp 1586364061
transform 1 0 80868 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_881
timestamp 1586364061
transform 1 0 82156 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_879
timestamp 1586364061
transform 1 0 81972 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_891
timestamp 1586364061
transform 1 0 83076 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_48
timestamp 1586364061
transform 1 0 83812 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_893
timestamp 1586364061
transform 1 0 83260 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_900
timestamp 1586364061
transform 1 0 83904 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_903
timestamp 1586364061
transform 1 0 84180 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 85284 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_912
timestamp 1586364061
transform 1 0 85008 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_924
timestamp 1586364061
transform 1 0 86112 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_916
timestamp 1586364061
transform 1 0 85376 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_49
timestamp 1586364061
transform 1 0 86664 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_931
timestamp 1586364061
transform 1 0 86756 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_943
timestamp 1586364061
transform 1 0 87860 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_928
timestamp 1586364061
transform 1 0 86480 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_940
timestamp 1586364061
transform 1 0 87584 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_50
timestamp 1586364061
transform 1 0 89516 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_955
timestamp 1586364061
transform 1 0 88964 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_962
timestamp 1586364061
transform 1 0 89608 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_952
timestamp 1586364061
transform 1 0 88688 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 90896 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_974
timestamp 1586364061
transform 1 0 90712 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_964
timestamp 1586364061
transform 1 0 89792 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_977
timestamp 1586364061
transform 1 0 90988 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_51
timestamp 1586364061
transform 1 0 92368 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_986
timestamp 1586364061
transform 1 0 91816 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_993
timestamp 1586364061
transform 1 0 92460 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_989
timestamp 1586364061
transform 1 0 92092 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1005
timestamp 1586364061
transform 1 0 93564 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1001
timestamp 1586364061
transform 1 0 93196 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1013
timestamp 1586364061
transform 1 0 94300 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_52
timestamp 1586364061
transform 1 0 95220 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1017
timestamp 1586364061
transform 1 0 94668 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1024
timestamp 1586364061
transform 1 0 95312 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1025
timestamp 1586364061
transform 1 0 95404 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 96508 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1036
timestamp 1586364061
transform 1 0 96416 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_1048
timestamp 1586364061
transform 1 0 97520 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1038
timestamp 1586364061
transform 1 0 96600 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1050
timestamp 1586364061
transform 1 0 97704 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_53
timestamp 1586364061
transform 1 0 98072 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1055
timestamp 1586364061
transform 1 0 98164 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1067
timestamp 1586364061
transform 1 0 99268 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1062
timestamp 1586364061
transform 1 0 98808 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_54
timestamp 1586364061
transform 1 0 100924 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1079
timestamp 1586364061
transform 1 0 100372 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1086
timestamp 1586364061
transform 1 0 101016 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1074
timestamp 1586364061
transform 1 0 99912 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1086
timestamp 1586364061
transform 1 0 101016 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 102120 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1098
timestamp 1586364061
transform 1 0 102120 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1099
timestamp 1586364061
transform 1 0 102212 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_55
timestamp 1586364061
transform 1 0 103776 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1110
timestamp 1586364061
transform 1 0 103224 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1117
timestamp 1586364061
transform 1 0 103868 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1111
timestamp 1586364061
transform 1 0 103316 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1123
timestamp 1586364061
transform 1 0 104420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1129
timestamp 1586364061
transform 1 0 104972 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_1141
timestamp 1586364061
transform 1 0 106076 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1135
timestamp 1586364061
transform 1 0 105524 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_56
timestamp 1586364061
transform 1 0 106628 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 107732 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1148
timestamp 1586364061
transform 1 0 106720 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1147
timestamp 1586364061
transform 1 0 106628 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1160
timestamp 1586364061
transform 1 0 107824 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_1172
timestamp 1586364061
transform 1 0 108928 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1160
timestamp 1586364061
transform 1 0 107824 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1172
timestamp 1586364061
transform 1 0 108928 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_57
timestamp 1586364061
transform 1 0 109480 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1179
timestamp 1586364061
transform 1 0 109572 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1191
timestamp 1586364061
transform 1 0 110676 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1184
timestamp 1586364061
transform 1 0 110032 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_58
timestamp 1586364061
transform 1 0 112332 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1203
timestamp 1586364061
transform 1 0 111780 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1210
timestamp 1586364061
transform 1 0 112424 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1196
timestamp 1586364061
transform 1 0 111136 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1208
timestamp 1586364061
transform 1 0 112240 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 113344 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1222
timestamp 1586364061
transform 1 0 113528 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1221
timestamp 1586364061
transform 1 0 113436 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_59
timestamp 1586364061
transform 1 0 115184 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1234
timestamp 1586364061
transform 1 0 114632 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1241
timestamp 1586364061
transform 1 0 115276 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1233
timestamp 1586364061
transform 1 0 114540 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1245
timestamp 1586364061
transform 1 0 115644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1253
timestamp 1586364061
transform 1 0 116380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_1265
timestamp 1586364061
transform 1 0 117484 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1257
timestamp 1586364061
transform 1 0 116748 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_60
timestamp 1586364061
transform 1 0 118036 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 118956 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1272
timestamp 1586364061
transform 1 0 118128 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1284
timestamp 1586364061
transform 1 0 119232 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1269
timestamp 1586364061
transform 1 0 117852 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1282
timestamp 1586364061
transform 1 0 119048 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_61
timestamp 1586364061
transform 1 0 120888 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1296
timestamp 1586364061
transform 1 0 120336 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1294
timestamp 1586364061
transform 1 0 120152 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1303
timestamp 1586364061
transform 1 0 120980 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1315
timestamp 1586364061
transform 1 0 122084 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1306
timestamp 1586364061
transform 1 0 121256 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1318
timestamp 1586364061
transform 1 0 122360 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_62
timestamp 1586364061
transform 1 0 123740 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1327
timestamp 1586364061
transform 1 0 123188 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1334
timestamp 1586364061
transform 1 0 123832 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1330
timestamp 1586364061
transform 1 0 123464 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 124568 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1346
timestamp 1586364061
transform 1 0 124936 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1343
timestamp 1586364061
transform 1 0 124660 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1355
timestamp 1586364061
transform 1 0 125764 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_63
timestamp 1586364061
transform 1 0 126592 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1358
timestamp 1586364061
transform 1 0 126040 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1365
timestamp 1586364061
transform 1 0 126684 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1367
timestamp 1586364061
transform 1 0 126868 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1377
timestamp 1586364061
transform 1 0 127788 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_1389
timestamp 1586364061
transform 1 0 128892 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1379
timestamp 1586364061
transform 1 0 127972 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1391
timestamp 1586364061
transform 1 0 129076 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_64
timestamp 1586364061
transform 1 0 129444 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 130180 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1396
timestamp 1586364061
transform 1 0 129536 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1408
timestamp 1586364061
transform 1 0 130640 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1404
timestamp 1586364061
transform 1 0 130272 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_65
timestamp 1586364061
transform 1 0 132296 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1420
timestamp 1586364061
transform 1 0 131744 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1416
timestamp 1586364061
transform 1 0 131376 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1427
timestamp 1586364061
transform 1 0 132388 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1439
timestamp 1586364061
transform 1 0 133492 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1428
timestamp 1586364061
transform 1 0 132480 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1440
timestamp 1586364061
transform 1 0 133584 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_66
timestamp 1586364061
transform 1 0 135148 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1451
timestamp 1586364061
transform 1 0 134596 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1458
timestamp 1586364061
transform 1 0 135240 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1452
timestamp 1586364061
transform 1 0 134688 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 135792 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1470
timestamp 1586364061
transform 1 0 136344 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1465
timestamp 1586364061
transform 1 0 135884 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1477
timestamp 1586364061
transform 1 0 136988 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_67
timestamp 1586364061
transform 1 0 138000 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1482
timestamp 1586364061
transform 1 0 137448 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1489
timestamp 1586364061
transform 1 0 138092 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1489
timestamp 1586364061
transform 1 0 138092 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1501
timestamp 1586364061
transform 1 0 139196 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_1513
timestamp 1586364061
transform 1 0 140300 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1501
timestamp 1586364061
transform 1 0 139196 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1513
timestamp 1586364061
transform 1 0 140300 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_68
timestamp 1586364061
transform 1 0 140852 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 141404 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1520
timestamp 1586364061
transform 1 0 140944 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1532
timestamp 1586364061
transform 1 0 142048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1526
timestamp 1586364061
transform 1 0 141496 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_69
timestamp 1586364061
transform 1 0 143704 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1544
timestamp 1586364061
transform 1 0 143152 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1551
timestamp 1586364061
transform 1 0 143796 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1538
timestamp 1586364061
transform 1 0 142600 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1550
timestamp 1586364061
transform 1 0 143704 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1563
timestamp 1586364061
transform 1 0 144900 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1562
timestamp 1586364061
transform 1 0 144808 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_70
timestamp 1586364061
transform 1 0 146556 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 147016 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1575
timestamp 1586364061
transform 1 0 146004 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1582
timestamp 1586364061
transform 1 0 146648 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1574
timestamp 1586364061
transform 1 0 145912 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1587
timestamp 1586364061
transform 1 0 147108 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1594
timestamp 1586364061
transform 1 0 147752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1599
timestamp 1586364061
transform 1 0 148212 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_71
timestamp 1586364061
transform 1 0 149408 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1606
timestamp 1586364061
transform 1 0 148856 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1613
timestamp 1586364061
transform 1 0 149500 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1611
timestamp 1586364061
transform 1 0 149316 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1623
timestamp 1586364061
transform 1 0 150420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1625
timestamp 1586364061
transform 1 0 150604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_1637
timestamp 1586364061
transform 1 0 151708 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1635
timestamp 1586364061
transform 1 0 151524 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_72
timestamp 1586364061
transform 1 0 152260 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 152628 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1644
timestamp 1586364061
transform 1 0 152352 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1656
timestamp 1586364061
transform 1 0 153456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1648
timestamp 1586364061
transform 1 0 152720 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 155112 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1668
timestamp 1586364061
transform 1 0 154560 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1675
timestamp 1586364061
transform 1 0 155204 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1660
timestamp 1586364061
transform 1 0 153824 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1672
timestamp 1586364061
transform 1 0 154928 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1687
timestamp 1586364061
transform 1 0 156308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1684
timestamp 1586364061
transform 1 0 156032 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 157964 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 158240 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1699
timestamp 1586364061
transform 1 0 157412 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1706
timestamp 1586364061
transform 1 0 158056 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1696
timestamp 1586364061
transform 1 0 157136 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1709
timestamp 1586364061
transform 1 0 158332 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1718
timestamp 1586364061
transform 1 0 159160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_1730
timestamp 1586364061
transform 1 0 160264 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1721
timestamp 1586364061
transform 1 0 159436 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 160816 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1737
timestamp 1586364061
transform 1 0 160908 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1733
timestamp 1586364061
transform 1 0 160540 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1745
timestamp 1586364061
transform 1 0 161644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1749
timestamp 1586364061
transform 1 0 162012 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_1761
timestamp 1586364061
transform 1 0 163116 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1757
timestamp 1586364061
transform 1 0 162748 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 163668 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 163852 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1768
timestamp 1586364061
transform 1 0 163760 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1780
timestamp 1586364061
transform 1 0 164864 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1770
timestamp 1586364061
transform 1 0 163944 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1782
timestamp 1586364061
transform 1 0 165048 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 166520 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1792
timestamp 1586364061
transform 1 0 165968 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1799
timestamp 1586364061
transform 1 0 166612 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1794
timestamp 1586364061
transform 1 0 166152 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1811
timestamp 1586364061
transform 1 0 167716 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1806
timestamp 1586364061
transform 1 0 167256 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1818
timestamp 1586364061
transform 1 0 168360 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 169372 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 169464 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1823
timestamp 1586364061
transform 1 0 168820 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1830
timestamp 1586364061
transform 1 0 169464 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1831
timestamp 1586364061
transform 1 0 169556 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1842
timestamp 1586364061
transform 1 0 170568 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_1854
timestamp 1586364061
transform 1 0 171672 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1843
timestamp 1586364061
transform 1 0 170660 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1855
timestamp 1586364061
transform 1 0 171764 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 172224 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1861
timestamp 1586364061
transform 1 0 172316 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1867
timestamp 1586364061
transform 1 0 172868 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1873
timestamp 1586364061
transform 1 0 173420 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_1885
timestamp 1586364061
transform 1 0 174524 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1879
timestamp 1586364061
transform 1 0 173972 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 175076 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 175076 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1892
timestamp 1586364061
transform 1 0 175168 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1904
timestamp 1586364061
transform 1 0 176272 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1892
timestamp 1586364061
transform 1 0 175168 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1904
timestamp 1586364061
transform 1 0 176272 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 177928 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1916
timestamp 1586364061
transform 1 0 177376 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1923
timestamp 1586364061
transform 1 0 178020 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1916
timestamp 1586364061
transform 1 0 177376 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1935
timestamp 1586364061
transform 1 0 179124 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1928
timestamp 1586364061
transform 1 0 178480 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1940
timestamp 1586364061
transform 1 0 179584 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 180780 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 180688 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_1947
timestamp 1586364061
transform 1 0 180228 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_1954
timestamp 1586364061
transform 1 0 180872 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1953
timestamp 1586364061
transform 1 0 180780 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1966
timestamp 1586364061
transform 1 0 181976 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_1978
timestamp 1586364061
transform 1 0 183080 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_1965
timestamp 1586364061
transform 1 0 181884 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1977
timestamp 1586364061
transform 1 0 182988 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 183632 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_1985
timestamp 1586364061
transform 1 0 183724 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_1997
timestamp 1586364061
transform 1 0 184828 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_1989
timestamp 1586364061
transform 1 0 184092 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 186484 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 186300 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2009
timestamp 1586364061
transform 1 0 185932 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_2001
timestamp 1586364061
transform 1 0 185196 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2014
timestamp 1586364061
transform 1 0 186392 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2016
timestamp 1586364061
transform 1 0 186576 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2028
timestamp 1586364061
transform 1 0 187680 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2026
timestamp 1586364061
transform 1 0 187496 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 189336 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2040
timestamp 1586364061
transform 1 0 188784 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2047
timestamp 1586364061
transform 1 0 189428 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2038
timestamp 1586364061
transform 1 0 188600 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2050
timestamp 1586364061
transform 1 0 189704 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2059
timestamp 1586364061
transform 1 0 190532 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2062
timestamp 1586364061
transform 1 0 190808 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 192188 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 191912 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2071
timestamp 1586364061
transform 1 0 191636 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2078
timestamp 1586364061
transform 1 0 192280 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2075
timestamp 1586364061
transform 1 0 192004 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2090
timestamp 1586364061
transform 1 0 193384 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_2102
timestamp 1586364061
transform 1 0 194488 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_2087
timestamp 1586364061
transform 1 0 193108 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2099
timestamp 1586364061
transform 1 0 194212 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 195040 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2109
timestamp 1586364061
transform 1 0 195132 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2121
timestamp 1586364061
transform 1 0 196236 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2111
timestamp 1586364061
transform 1 0 195316 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 197892 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 197524 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2133
timestamp 1586364061
transform 1 0 197340 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2140
timestamp 1586364061
transform 1 0 197984 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2123
timestamp 1586364061
transform 1 0 196420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2136
timestamp 1586364061
transform 1 0 197616 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2152
timestamp 1586364061
transform 1 0 199088 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2148
timestamp 1586364061
transform 1 0 198720 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 200744 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2164
timestamp 1586364061
transform 1 0 200192 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2171
timestamp 1586364061
transform 1 0 200836 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2160
timestamp 1586364061
transform 1 0 199824 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2172
timestamp 1586364061
transform 1 0 200928 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2183
timestamp 1586364061
transform 1 0 201940 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2184
timestamp 1586364061
transform 1 0 202032 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 203596 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 203136 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2195
timestamp 1586364061
transform 1 0 203044 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2202
timestamp 1586364061
transform 1 0 203688 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2197
timestamp 1586364061
transform 1 0 203228 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2209
timestamp 1586364061
transform 1 0 204332 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2214
timestamp 1586364061
transform 1 0 204792 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_2226
timestamp 1586364061
transform 1 0 205896 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_2221
timestamp 1586364061
transform 1 0 205436 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 206448 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2233
timestamp 1586364061
transform 1 0 206540 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_2245
timestamp 1586364061
transform 1 0 207644 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_2233
timestamp 1586364061
transform 1 0 206540 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2245
timestamp 1586364061
transform 1 0 207644 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _17_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 208012 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 209300 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 208748 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__17__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 208564 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_2253
timestamp 1586364061
transform 1 0 208380 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_2257
timestamp 1586364061
transform 1 0 208748 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2264
timestamp 1586364061
transform 1 0 209392 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2258
timestamp 1586364061
transform 1 0 208840 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2276
timestamp 1586364061
transform 1 0 210496 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2270
timestamp 1586364061
transform 1 0 209944 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2282
timestamp 1586364061
transform 1 0 211048 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 212152 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2288
timestamp 1586364061
transform 1 0 211600 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2295
timestamp 1586364061
transform 1 0 212244 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2294
timestamp 1586364061
transform 1 0 212152 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 214360 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2307
timestamp 1586364061
transform 1 0 213348 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2306
timestamp 1586364061
transform 1 0 213256 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 215004 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2319
timestamp 1586364061
transform 1 0 214452 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2326
timestamp 1586364061
transform 1 0 215096 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2319
timestamp 1586364061
transform 1 0 214452 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2331
timestamp 1586364061
transform 1 0 215556 0 1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_1_2343 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 216660 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__14__B
timestamp 1586364061
transform 1 0 216752 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_2350
timestamp 1586364061
transform 1 0 217304 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_2346
timestamp 1586364061
transform 1 0 216936 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_2350
timestamp 1586364061
transform 1 0 217304 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__13__D
timestamp 1586364061
transform 1 0 217120 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__14__C
timestamp 1586364061
transform 1 0 217672 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__14__D
timestamp 1586364061
transform 1 0 217488 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_2338
timestamp 1586364061
transform 1 0 216200 0 -1 2720
box -38 -48 1142 592
use scs8hd_nor4_4  _14_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 217672 0 1 2720
box -38 -48 1602 592
use scs8hd_inv_8  _08_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 218408 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 217856 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__08__A
timestamp 1586364061
transform 1 0 218224 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_2357
timestamp 1586364061
transform 1 0 217948 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_2371
timestamp 1586364061
transform 1 0 219236 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_2371
timestamp 1586364061
transform 1 0 219236 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_2375
timestamp 1586364061
transform 1 0 219604 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_2379
timestamp 1586364061
transform 1 0 219972 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_2375
timestamp 1586364061
transform 1 0 219604 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__13__B
timestamp 1586364061
transform 1 0 219788 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__13__C
timestamp 1586364061
transform 1 0 219420 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__11__A
timestamp 1586364061
transform 1 0 219788 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__13__A
timestamp 1586364061
transform 1 0 219420 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 219972 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_2389
timestamp 1586364061
transform 1 0 220892 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 220708 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2388
timestamp 1586364061
transform 1 0 220800 0 -1 2720
box -38 -48 1142 592
use scs8hd_inv_8  _11_
timestamp 1586364061
transform 1 0 220064 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 221076 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 221444 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_2400
timestamp 1586364061
transform 1 0 221904 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_2393
timestamp 1586364061
transform 1 0 221260 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_2397
timestamp 1586364061
transform 1 0 221628 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 223560 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__04__A
timestamp 1586364061
transform 1 0 222916 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_2412
timestamp 1586364061
transform 1 0 223008 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2419
timestamp 1586364061
transform 1 0 223652 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_2409
timestamp 1586364061
transform 1 0 222732 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_2413
timestamp 1586364061
transform 1 0 223100 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_1_2425
timestamp 1586364061
transform 1 0 224204 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_2434
timestamp 1586364061
transform 1 0 225032 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_2430
timestamp 1586364061
transform 1 0 224664 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_2431
timestamp 1586364061
transform 1 0 224756 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__05__A
timestamp 1586364061
transform 1 0 224848 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__05__D
timestamp 1586364061
transform 1 0 224480 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__05__C
timestamp 1586364061
transform 1 0 224848 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_2438
timestamp 1586364061
transform 1 0 225400 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__05__B
timestamp 1586364061
transform 1 0 225216 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 225584 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_2441
timestamp 1586364061
transform 1 0 225676 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2434
timestamp 1586364061
transform 1 0 225032 0 -1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 226412 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_0_2446
timestamp 1586364061
transform 1 0 226136 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_2450
timestamp 1586364061
transform 1 0 226504 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2453
timestamp 1586364061
transform 1 0 226780 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2462
timestamp 1586364061
transform 1 0 227608 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_2474
timestamp 1586364061
transform 1 0 228712 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_2465
timestamp 1586364061
transform 1 0 227884 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2477
timestamp 1586364061
transform 1 0 228988 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 229264 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2481
timestamp 1586364061
transform 1 0 229356 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2493
timestamp 1586364061
transform 1 0 230460 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2489
timestamp 1586364061
transform 1 0 230092 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 232116 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 231196 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2505
timestamp 1586364061
transform 1 0 231564 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2512
timestamp 1586364061
transform 1 0 232208 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2502
timestamp 1586364061
transform 1 0 231288 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2514
timestamp 1586364061
transform 1 0 232392 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2524
timestamp 1586364061
transform 1 0 233312 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2526
timestamp 1586364061
transform 1 0 233496 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 234968 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2536
timestamp 1586364061
transform 1 0 234416 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2543
timestamp 1586364061
transform 1 0 235060 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2538
timestamp 1586364061
transform 1 0 234600 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2550
timestamp 1586364061
transform 1 0 235704 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 236808 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2555
timestamp 1586364061
transform 1 0 236164 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_2567
timestamp 1586364061
transform 1 0 237268 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_2563
timestamp 1586364061
transform 1 0 236900 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 237820 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2574
timestamp 1586364061
transform 1 0 237912 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2586
timestamp 1586364061
transform 1 0 239016 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2575
timestamp 1586364061
transform 1 0 238004 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 240672 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2598
timestamp 1586364061
transform 1 0 240120 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_2587
timestamp 1586364061
transform 1 0 239108 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2599
timestamp 1586364061
transform 1 0 240212 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2605
timestamp 1586364061
transform 1 0 240764 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2617
timestamp 1586364061
transform 1 0 241868 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2611
timestamp 1586364061
transform 1 0 241316 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 243524 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 242420 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2629
timestamp 1586364061
transform 1 0 242972 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2636
timestamp 1586364061
transform 1 0 243616 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2624
timestamp 1586364061
transform 1 0 242512 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2636
timestamp 1586364061
transform 1 0 243616 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2648
timestamp 1586364061
transform 1 0 244720 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2648
timestamp 1586364061
transform 1 0 244720 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 246376 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2660
timestamp 1586364061
transform 1 0 245824 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2667
timestamp 1586364061
transform 1 0 246468 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2660
timestamp 1586364061
transform 1 0 245824 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2672
timestamp 1586364061
transform 1 0 246928 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 248032 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2679
timestamp 1586364061
transform 1 0 247572 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_2691
timestamp 1586364061
transform 1 0 248676 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_2685
timestamp 1586364061
transform 1 0 248124 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 249228 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2698
timestamp 1586364061
transform 1 0 249320 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2710
timestamp 1586364061
transform 1 0 250424 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2697
timestamp 1586364061
transform 1 0 249228 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2709
timestamp 1586364061
transform 1 0 250332 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 252080 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2722
timestamp 1586364061
transform 1 0 251528 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2729
timestamp 1586364061
transform 1 0 252172 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2721
timestamp 1586364061
transform 1 0 251436 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 253644 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2741
timestamp 1586364061
transform 1 0 253276 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2733
timestamp 1586364061
transform 1 0 252540 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2746
timestamp 1586364061
transform 1 0 253736 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 254932 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2753
timestamp 1586364061
transform 1 0 254380 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2760
timestamp 1586364061
transform 1 0 255024 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2758
timestamp 1586364061
transform 1 0 254840 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2772
timestamp 1586364061
transform 1 0 256128 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2770
timestamp 1586364061
transform 1 0 255944 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2782
timestamp 1586364061
transform 1 0 257048 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 257784 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2784
timestamp 1586364061
transform 1 0 257232 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2791
timestamp 1586364061
transform 1 0 257876 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2794
timestamp 1586364061
transform 1 0 258152 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 259256 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2803
timestamp 1586364061
transform 1 0 258980 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_2815
timestamp 1586364061
transform 1 0 260084 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_2807
timestamp 1586364061
transform 1 0 259348 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 260636 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2822
timestamp 1586364061
transform 1 0 260728 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2834
timestamp 1586364061
transform 1 0 261832 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2819
timestamp 1586364061
transform 1 0 260452 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2831
timestamp 1586364061
transform 1 0 261556 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 263488 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2846
timestamp 1586364061
transform 1 0 262936 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2853
timestamp 1586364061
transform 1 0 263580 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2843
timestamp 1586364061
transform 1 0 262660 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 264868 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2865
timestamp 1586364061
transform 1 0 264684 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2855
timestamp 1586364061
transform 1 0 263764 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2868
timestamp 1586364061
transform 1 0 264960 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 266340 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2877
timestamp 1586364061
transform 1 0 265788 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2884
timestamp 1586364061
transform 1 0 266432 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2880
timestamp 1586364061
transform 1 0 266064 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2896
timestamp 1586364061
transform 1 0 267536 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2892
timestamp 1586364061
transform 1 0 267168 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2904
timestamp 1586364061
transform 1 0 268272 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 269192 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2908
timestamp 1586364061
transform 1 0 268640 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2915
timestamp 1586364061
transform 1 0 269284 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2916
timestamp 1586364061
transform 1 0 269376 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 270480 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2927
timestamp 1586364061
transform 1 0 270388 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_2939
timestamp 1586364061
transform 1 0 271492 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_2929
timestamp 1586364061
transform 1 0 270572 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2941
timestamp 1586364061
transform 1 0 271676 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 272044 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2946
timestamp 1586364061
transform 1 0 272136 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_2958
timestamp 1586364061
transform 1 0 273240 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2953
timestamp 1586364061
transform 1 0 272780 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 274896 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_2970
timestamp 1586364061
transform 1 0 274344 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_2977
timestamp 1586364061
transform 1 0 274988 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2965
timestamp 1586364061
transform 1 0 273884 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2977
timestamp 1586364061
transform 1 0 274988 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 276092 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_2989
timestamp 1586364061
transform 1 0 276092 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_2990
timestamp 1586364061
transform 1 0 276184 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 277748 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3001
timestamp 1586364061
transform 1 0 277196 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3008
timestamp 1586364061
transform 1 0 277840 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3002
timestamp 1586364061
transform 1 0 277288 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3014
timestamp 1586364061
transform 1 0 278392 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3020
timestamp 1586364061
transform 1 0 278944 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_3032
timestamp 1586364061
transform 1 0 280048 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_3026
timestamp 1586364061
transform 1 0 279496 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 280600 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 281704 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_3039
timestamp 1586364061
transform 1 0 280692 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3038
timestamp 1586364061
transform 1 0 280600 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3051
timestamp 1586364061
transform 1 0 281796 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_3063
timestamp 1586364061
transform 1 0 282900 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_3051
timestamp 1586364061
transform 1 0 281796 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3063
timestamp 1586364061
transform 1 0 282900 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 283452 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_3070
timestamp 1586364061
transform 1 0 283544 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3082
timestamp 1586364061
transform 1 0 284648 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3075
timestamp 1586364061
transform 1 0 284004 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 286304 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3094
timestamp 1586364061
transform 1 0 285752 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3101
timestamp 1586364061
transform 1 0 286396 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3087
timestamp 1586364061
transform 1 0 285108 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3099
timestamp 1586364061
transform 1 0 286212 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 287316 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_3113
timestamp 1586364061
transform 1 0 287500 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3112
timestamp 1586364061
transform 1 0 287408 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 289156 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3125
timestamp 1586364061
transform 1 0 288604 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3132
timestamp 1586364061
transform 1 0 289248 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3124
timestamp 1586364061
transform 1 0 288512 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3136
timestamp 1586364061
transform 1 0 289616 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3144
timestamp 1586364061
transform 1 0 290352 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_3156
timestamp 1586364061
transform 1 0 291456 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_3148
timestamp 1586364061
transform 1 0 290720 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 292008 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 292928 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_3163
timestamp 1586364061
transform 1 0 292100 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3160
timestamp 1586364061
transform 1 0 291824 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3173
timestamp 1586364061
transform 1 0 293020 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3175
timestamp 1586364061
transform 1 0 293204 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_3187
timestamp 1586364061
transform 1 0 294308 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_3185
timestamp 1586364061
transform 1 0 294124 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 294860 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_3194
timestamp 1586364061
transform 1 0 294952 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3206
timestamp 1586364061
transform 1 0 296056 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3197
timestamp 1586364061
transform 1 0 295228 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3209
timestamp 1586364061
transform 1 0 296332 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 297712 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3218
timestamp 1586364061
transform 1 0 297160 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3225
timestamp 1586364061
transform 1 0 297804 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3221
timestamp 1586364061
transform 1 0 297436 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 298540 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_3237
timestamp 1586364061
transform 1 0 298908 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3234
timestamp 1586364061
transform 1 0 298632 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3246
timestamp 1586364061
transform 1 0 299736 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 300564 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3249
timestamp 1586364061
transform 1 0 300012 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3256
timestamp 1586364061
transform 1 0 300656 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3258
timestamp 1586364061
transform 1 0 300840 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3268
timestamp 1586364061
transform 1 0 301760 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_3280
timestamp 1586364061
transform 1 0 302864 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_3270
timestamp 1586364061
transform 1 0 301944 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 303416 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 304152 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_3287
timestamp 1586364061
transform 1 0 303508 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3299
timestamp 1586364061
transform 1 0 304612 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3282
timestamp 1586364061
transform 1 0 303048 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3295
timestamp 1586364061
transform 1 0 304244 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 306268 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3311
timestamp 1586364061
transform 1 0 305716 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_3307
timestamp 1586364061
transform 1 0 305348 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3318
timestamp 1586364061
transform 1 0 306360 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3330
timestamp 1586364061
transform 1 0 307464 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3319
timestamp 1586364061
transform 1 0 306452 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3331
timestamp 1586364061
transform 1 0 307556 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 309120 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3342
timestamp 1586364061
transform 1 0 308568 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3349
timestamp 1586364061
transform 1 0 309212 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3343
timestamp 1586364061
transform 1 0 308660 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 309764 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_3361
timestamp 1586364061
transform 1 0 310316 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3356
timestamp 1586364061
transform 1 0 309856 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3368
timestamp 1586364061
transform 1 0 310960 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 311972 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3373
timestamp 1586364061
transform 1 0 311420 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3380
timestamp 1586364061
transform 1 0 312064 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3380
timestamp 1586364061
transform 1 0 312064 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3392
timestamp 1586364061
transform 1 0 313168 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_3404
timestamp 1586364061
transform 1 0 314272 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_3392
timestamp 1586364061
transform 1 0 313168 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3404
timestamp 1586364061
transform 1 0 314272 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 314824 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 315376 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_3411
timestamp 1586364061
transform 1 0 314916 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3423
timestamp 1586364061
transform 1 0 316020 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3417
timestamp 1586364061
transform 1 0 315468 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 317676 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3435
timestamp 1586364061
transform 1 0 317124 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3442
timestamp 1586364061
transform 1 0 317768 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3429
timestamp 1586364061
transform 1 0 316572 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3441
timestamp 1586364061
transform 1 0 317676 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3454
timestamp 1586364061
transform 1 0 318872 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3453
timestamp 1586364061
transform 1 0 318780 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 320528 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 320988 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3466
timestamp 1586364061
transform 1 0 319976 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3473
timestamp 1586364061
transform 1 0 320620 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3465
timestamp 1586364061
transform 1 0 319884 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3478
timestamp 1586364061
transform 1 0 321080 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3485
timestamp 1586364061
transform 1 0 321724 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3490
timestamp 1586364061
transform 1 0 322184 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 323380 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3497
timestamp 1586364061
transform 1 0 322828 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3504
timestamp 1586364061
transform 1 0 323472 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3502
timestamp 1586364061
transform 1 0 323288 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3516
timestamp 1586364061
transform 1 0 324576 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_3528
timestamp 1586364061
transform 1 0 325680 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_3514
timestamp 1586364061
transform 1 0 324392 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3526
timestamp 1586364061
transform 1 0 325496 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 326232 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 326600 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_3535
timestamp 1586364061
transform 1 0 326324 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3547
timestamp 1586364061
transform 1 0 327428 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3539
timestamp 1586364061
transform 1 0 326692 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 329084 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3559
timestamp 1586364061
transform 1 0 328532 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3566
timestamp 1586364061
transform 1 0 329176 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3551
timestamp 1586364061
transform 1 0 327796 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3563
timestamp 1586364061
transform 1 0 328900 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3578
timestamp 1586364061
transform 1 0 330280 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3575
timestamp 1586364061
transform 1 0 330004 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 331936 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 332212 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3590
timestamp 1586364061
transform 1 0 331384 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3597
timestamp 1586364061
transform 1 0 332028 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3587
timestamp 1586364061
transform 1 0 331108 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3600
timestamp 1586364061
transform 1 0 332304 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3609
timestamp 1586364061
transform 1 0 333132 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3612
timestamp 1586364061
transform 1 0 333408 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 334788 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3621
timestamp 1586364061
transform 1 0 334236 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3628
timestamp 1586364061
transform 1 0 334880 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3624
timestamp 1586364061
transform 1 0 334512 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3636
timestamp 1586364061
transform 1 0 335616 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3640
timestamp 1586364061
transform 1 0 335984 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_3652
timestamp 1586364061
transform 1 0 337088 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_3648
timestamp 1586364061
transform 1 0 336720 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 337640 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 337824 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_3659
timestamp 1586364061
transform 1 0 337732 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3671
timestamp 1586364061
transform 1 0 338836 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3661
timestamp 1586364061
transform 1 0 337916 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3673
timestamp 1586364061
transform 1 0 339020 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 340492 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3683
timestamp 1586364061
transform 1 0 339940 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3690
timestamp 1586364061
transform 1 0 340584 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3685
timestamp 1586364061
transform 1 0 340124 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3702
timestamp 1586364061
transform 1 0 341688 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3697
timestamp 1586364061
transform 1 0 341228 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3709
timestamp 1586364061
transform 1 0 342332 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 343344 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 343436 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3714
timestamp 1586364061
transform 1 0 342792 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3721
timestamp 1586364061
transform 1 0 343436 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3722
timestamp 1586364061
transform 1 0 343528 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3733
timestamp 1586364061
transform 1 0 344540 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_3745
timestamp 1586364061
transform 1 0 345644 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_3734
timestamp 1586364061
transform 1 0 344632 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 346196 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_3752
timestamp 1586364061
transform 1 0 346288 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3746
timestamp 1586364061
transform 1 0 345736 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3758
timestamp 1586364061
transform 1 0 346840 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3764
timestamp 1586364061
transform 1 0 347392 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_3776
timestamp 1586364061
transform 1 0 348496 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_3770
timestamp 1586364061
transform 1 0 347944 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 349048 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 349048 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_3783
timestamp 1586364061
transform 1 0 349140 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3795
timestamp 1586364061
transform 1 0 350244 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3783
timestamp 1586364061
transform 1 0 349140 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3795
timestamp 1586364061
transform 1 0 350244 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 351900 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3807
timestamp 1586364061
transform 1 0 351348 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3814
timestamp 1586364061
transform 1 0 351992 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3807
timestamp 1586364061
transform 1 0 351348 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3826
timestamp 1586364061
transform 1 0 353096 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3819
timestamp 1586364061
transform 1 0 352452 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3831
timestamp 1586364061
transform 1 0 353556 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 354752 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 354660 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3838
timestamp 1586364061
transform 1 0 354200 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3845
timestamp 1586364061
transform 1 0 354844 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3844
timestamp 1586364061
transform 1 0 354752 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3857
timestamp 1586364061
transform 1 0 355948 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_3869
timestamp 1586364061
transform 1 0 357052 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_3856
timestamp 1586364061
transform 1 0 355856 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3868
timestamp 1586364061
transform 1 0 356960 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 357604 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_3876
timestamp 1586364061
transform 1 0 357696 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3888
timestamp 1586364061
transform 1 0 358800 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3880
timestamp 1586364061
transform 1 0 358064 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 360456 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 360272 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3900
timestamp 1586364061
transform 1 0 359904 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_3892
timestamp 1586364061
transform 1 0 359168 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3905
timestamp 1586364061
transform 1 0 360364 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3907
timestamp 1586364061
transform 1 0 360548 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3919
timestamp 1586364061
transform 1 0 361652 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3917
timestamp 1586364061
transform 1 0 361468 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 363308 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3931
timestamp 1586364061
transform 1 0 362756 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3938
timestamp 1586364061
transform 1 0 363400 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3929
timestamp 1586364061
transform 1 0 362572 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3941
timestamp 1586364061
transform 1 0 363676 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3950
timestamp 1586364061
transform 1 0 364504 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3953
timestamp 1586364061
transform 1 0 364780 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 366160 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 365884 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_3962
timestamp 1586364061
transform 1 0 365608 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_3969
timestamp 1586364061
transform 1 0 366252 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3966
timestamp 1586364061
transform 1 0 365976 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3981
timestamp 1586364061
transform 1 0 367356 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_3993
timestamp 1586364061
transform 1 0 368460 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_3978
timestamp 1586364061
transform 1 0 367080 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3990
timestamp 1586364061
transform 1 0 368184 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 369012 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_4000
timestamp 1586364061
transform 1 0 369104 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4012
timestamp 1586364061
transform 1 0 370208 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4002
timestamp 1586364061
transform 1 0 369288 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 371864 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 371496 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_4024
timestamp 1586364061
transform 1 0 371312 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_4031
timestamp 1586364061
transform 1 0 371956 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4014
timestamp 1586364061
transform 1 0 370392 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4027
timestamp 1586364061
transform 1 0 371588 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4043
timestamp 1586364061
transform 1 0 373060 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4039
timestamp 1586364061
transform 1 0 372692 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 374716 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_4055
timestamp 1586364061
transform 1 0 374164 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_4062
timestamp 1586364061
transform 1 0 374808 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4051
timestamp 1586364061
transform 1 0 373796 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4063
timestamp 1586364061
transform 1 0 374900 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4074
timestamp 1586364061
transform 1 0 375912 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4075
timestamp 1586364061
transform 1 0 376004 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 377568 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 377108 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_4086
timestamp 1586364061
transform 1 0 377016 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_4093
timestamp 1586364061
transform 1 0 377660 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4088
timestamp 1586364061
transform 1 0 377200 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4100
timestamp 1586364061
transform 1 0 378304 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4105
timestamp 1586364061
transform 1 0 378764 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_4117
timestamp 1586364061
transform 1 0 379868 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_4112
timestamp 1586364061
transform 1 0 379408 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 380420 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_4124
timestamp 1586364061
transform 1 0 380512 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4136
timestamp 1586364061
transform 1 0 381616 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4124
timestamp 1586364061
transform 1 0 380512 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4136
timestamp 1586364061
transform 1 0 381616 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 383272 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 382720 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_4148
timestamp 1586364061
transform 1 0 382720 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_4155
timestamp 1586364061
transform 1 0 383364 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4149
timestamp 1586364061
transform 1 0 382812 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4167
timestamp 1586364061
transform 1 0 384468 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4161
timestamp 1586364061
transform 1 0 383916 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4173
timestamp 1586364061
transform 1 0 385020 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 386124 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_4179
timestamp 1586364061
transform 1 0 385572 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_4186
timestamp 1586364061
transform 1 0 386216 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4185
timestamp 1586364061
transform 1 0 386124 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 388332 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_4198
timestamp 1586364061
transform 1 0 387320 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4197
timestamp 1586364061
transform 1 0 387228 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 388976 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_4210
timestamp 1586364061
transform 1 0 388424 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_4217
timestamp 1586364061
transform 1 0 389068 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4210
timestamp 1586364061
transform 1 0 388424 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4222
timestamp 1586364061
transform 1 0 389528 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4229
timestamp 1586364061
transform 1 0 390172 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_4241
timestamp 1586364061
transform 1 0 391276 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_4234
timestamp 1586364061
transform 1 0 390632 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 391828 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_4248
timestamp 1586364061
transform 1 0 391920 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4260
timestamp 1586364061
transform 1 0 393024 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4246
timestamp 1586364061
transform 1 0 391736 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4258
timestamp 1586364061
transform 1 0 392840 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 394680 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 393944 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_4272
timestamp 1586364061
transform 1 0 394128 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_4279
timestamp 1586364061
transform 1 0 394772 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4271
timestamp 1586364061
transform 1 0 394036 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4291
timestamp 1586364061
transform 1 0 395876 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4283
timestamp 1586364061
transform 1 0 395140 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4295
timestamp 1586364061
transform 1 0 396244 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 397532 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_4303
timestamp 1586364061
transform 1 0 396980 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_4310
timestamp 1586364061
transform 1 0 397624 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4307
timestamp 1586364061
transform 1 0 397348 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 399556 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_4322
timestamp 1586364061
transform 1 0 398728 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_4334
timestamp 1586364061
transform 1 0 399832 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_4319
timestamp 1586364061
transform 1 0 398452 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4332
timestamp 1586364061
transform 1 0 399648 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 400384 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_4341
timestamp 1586364061
transform 1 0 400476 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4344
timestamp 1586364061
transform 1 0 400752 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4353
timestamp 1586364061
transform 1 0 401580 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_4365
timestamp 1586364061
transform 1 0 402684 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_4356
timestamp 1586364061
transform 1 0 401856 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4368
timestamp 1586364061
transform 1 0 402960 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 403236 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_4372
timestamp 1586364061
transform 1 0 403328 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4384
timestamp 1586364061
transform 1 0 404432 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4380
timestamp 1586364061
transform 1 0 404064 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 406088 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 405168 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_4396
timestamp 1586364061
transform 1 0 405536 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_4403
timestamp 1586364061
transform 1 0 406180 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4393
timestamp 1586364061
transform 1 0 405260 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4405
timestamp 1586364061
transform 1 0 406364 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4415
timestamp 1586364061
transform 1 0 407284 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4417
timestamp 1586364061
transform 1 0 407468 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 408940 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_4427
timestamp 1586364061
transform 1 0 408388 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_4434
timestamp 1586364061
transform 1 0 409032 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4429
timestamp 1586364061
transform 1 0 408572 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4441
timestamp 1586364061
transform 1 0 409676 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 410780 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_4446
timestamp 1586364061
transform 1 0 410136 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_4458
timestamp 1586364061
transform 1 0 411240 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_4454
timestamp 1586364061
transform 1 0 410872 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 411792 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_4465
timestamp 1586364061
transform 1 0 411884 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4477
timestamp 1586364061
transform 1 0 412988 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4466
timestamp 1586364061
transform 1 0 411976 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_4489
timestamp 1586364061
transform 1 0 414092 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_4478
timestamp 1586364061
transform 1 0 413080 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4490
timestamp 1586364061
transform 1 0 414184 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 414644 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_4496
timestamp 1586364061
transform 1 0 414736 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4508
timestamp 1586364061
transform 1 0 415840 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4502
timestamp 1586364061
transform 1 0 415288 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 417496 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 416392 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_4520
timestamp 1586364061
transform 1 0 416944 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_4527
timestamp 1586364061
transform 1 0 417588 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4515
timestamp 1586364061
transform 1 0 416484 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4527
timestamp 1586364061
transform 1 0 417588 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_4539
timestamp 1586364061
transform 1 0 418692 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4539
timestamp 1586364061
transform 1 0 418692 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 420348 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_4551
timestamp 1586364061
transform 1 0 419796 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_4558
timestamp 1586364061
transform 1 0 420440 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4551
timestamp 1586364061
transform 1 0 419796 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_4563
timestamp 1586364061
transform 1 0 420900 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 422832 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 422832 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 422004 0 1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_0_4570
timestamp 1586364061
transform 1 0 421544 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_3  FILLER_0_4578
timestamp 1586364061
transform 1 0 422280 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_4576
timestamp 1586364061
transform 1 0 422096 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_4580
timestamp 1586364061
transform 1 0 422464 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_288
timestamp 1586364061
transform 1 0 27600 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_300
timestamp 1586364061
transform 1 0 28704 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_312
timestamp 1586364061
transform 1 0 29808 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_324
timestamp 1586364061
transform 1 0 30912 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_337
timestamp 1586364061
transform 1 0 32108 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_349
timestamp 1586364061
transform 1 0 33212 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_361
timestamp 1586364061
transform 1 0 34316 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_373
timestamp 1586364061
transform 1 0 35420 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_385
timestamp 1586364061
transform 1 0 36524 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_398
timestamp 1586364061
transform 1 0 37720 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_410
timestamp 1586364061
transform 1 0 38824 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_422
timestamp 1586364061
transform 1 0 39928 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_434
timestamp 1586364061
transform 1 0 41032 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 43240 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_446
timestamp 1586364061
transform 1 0 42136 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_459
timestamp 1586364061
transform 1 0 43332 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_471
timestamp 1586364061
transform 1 0 44436 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_483
timestamp 1586364061
transform 1 0 45540 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_495
timestamp 1586364061
transform 1 0 46644 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_507
timestamp 1586364061
transform 1 0 47748 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 48852 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_520
timestamp 1586364061
transform 1 0 48944 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_532
timestamp 1586364061
transform 1 0 50048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_544
timestamp 1586364061
transform 1 0 51152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_556
timestamp 1586364061
transform 1 0 52256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_568
timestamp 1586364061
transform 1 0 53360 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 54464 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_581
timestamp 1586364061
transform 1 0 54556 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_593
timestamp 1586364061
transform 1 0 55660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_605
timestamp 1586364061
transform 1 0 56764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_617
timestamp 1586364061
transform 1 0 57868 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 60076 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_629
timestamp 1586364061
transform 1 0 58972 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_642
timestamp 1586364061
transform 1 0 60168 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_654
timestamp 1586364061
transform 1 0 61272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_666
timestamp 1586364061
transform 1 0 62376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_678
timestamp 1586364061
transform 1 0 63480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_690
timestamp 1586364061
transform 1 0 64584 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 65688 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_703
timestamp 1586364061
transform 1 0 65780 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_715
timestamp 1586364061
transform 1 0 66884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_727
timestamp 1586364061
transform 1 0 67988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_739
timestamp 1586364061
transform 1 0 69092 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 71300 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_751
timestamp 1586364061
transform 1 0 70196 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_764
timestamp 1586364061
transform 1 0 71392 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_776
timestamp 1586364061
transform 1 0 72496 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_788
timestamp 1586364061
transform 1 0 73600 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_800
timestamp 1586364061
transform 1 0 74704 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_812
timestamp 1586364061
transform 1 0 75808 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 76912 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_825
timestamp 1586364061
transform 1 0 77004 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_837
timestamp 1586364061
transform 1 0 78108 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_849
timestamp 1586364061
transform 1 0 79212 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_861
timestamp 1586364061
transform 1 0 80316 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_873
timestamp 1586364061
transform 1 0 81420 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 82524 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_886
timestamp 1586364061
transform 1 0 82616 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_898
timestamp 1586364061
transform 1 0 83720 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_910
timestamp 1586364061
transform 1 0 84824 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_922
timestamp 1586364061
transform 1 0 85928 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_934
timestamp 1586364061
transform 1 0 87032 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 88136 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_947
timestamp 1586364061
transform 1 0 88228 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_959
timestamp 1586364061
transform 1 0 89332 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_971
timestamp 1586364061
transform 1 0 90436 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_983
timestamp 1586364061
transform 1 0 91540 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_995
timestamp 1586364061
transform 1 0 92644 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 93748 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1008
timestamp 1586364061
transform 1 0 93840 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1020
timestamp 1586364061
transform 1 0 94944 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1032
timestamp 1586364061
transform 1 0 96048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1044
timestamp 1586364061
transform 1 0 97152 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 99360 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1056
timestamp 1586364061
transform 1 0 98256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1069
timestamp 1586364061
transform 1 0 99452 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1081
timestamp 1586364061
transform 1 0 100556 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1093
timestamp 1586364061
transform 1 0 101660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1105
timestamp 1586364061
transform 1 0 102764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1117
timestamp 1586364061
transform 1 0 103868 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 104972 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1130
timestamp 1586364061
transform 1 0 105064 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1142
timestamp 1586364061
transform 1 0 106168 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1154
timestamp 1586364061
transform 1 0 107272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1166
timestamp 1586364061
transform 1 0 108376 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 110584 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1178
timestamp 1586364061
transform 1 0 109480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1191
timestamp 1586364061
transform 1 0 110676 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1203
timestamp 1586364061
transform 1 0 111780 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1215
timestamp 1586364061
transform 1 0 112884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1227
timestamp 1586364061
transform 1 0 113988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1239
timestamp 1586364061
transform 1 0 115092 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 116196 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1252
timestamp 1586364061
transform 1 0 116288 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1264
timestamp 1586364061
transform 1 0 117392 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1276
timestamp 1586364061
transform 1 0 118496 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1288
timestamp 1586364061
transform 1 0 119600 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1300
timestamp 1586364061
transform 1 0 120704 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 121808 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1313
timestamp 1586364061
transform 1 0 121900 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1325
timestamp 1586364061
transform 1 0 123004 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1337
timestamp 1586364061
transform 1 0 124108 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1349
timestamp 1586364061
transform 1 0 125212 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 127420 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1361
timestamp 1586364061
transform 1 0 126316 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1374
timestamp 1586364061
transform 1 0 127512 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1386
timestamp 1586364061
transform 1 0 128616 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1398
timestamp 1586364061
transform 1 0 129720 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1410
timestamp 1586364061
transform 1 0 130824 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1422
timestamp 1586364061
transform 1 0 131928 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 133032 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1435
timestamp 1586364061
transform 1 0 133124 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1447
timestamp 1586364061
transform 1 0 134228 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1459
timestamp 1586364061
transform 1 0 135332 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1471
timestamp 1586364061
transform 1 0 136436 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 138644 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1483
timestamp 1586364061
transform 1 0 137540 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1496
timestamp 1586364061
transform 1 0 138736 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1508
timestamp 1586364061
transform 1 0 139840 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1520
timestamp 1586364061
transform 1 0 140944 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1532
timestamp 1586364061
transform 1 0 142048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1544
timestamp 1586364061
transform 1 0 143152 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 144256 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1557
timestamp 1586364061
transform 1 0 144348 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1569
timestamp 1586364061
transform 1 0 145452 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1581
timestamp 1586364061
transform 1 0 146556 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1593
timestamp 1586364061
transform 1 0 147660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1605
timestamp 1586364061
transform 1 0 148764 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 149868 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1618
timestamp 1586364061
transform 1 0 149960 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1630
timestamp 1586364061
transform 1 0 151064 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1642
timestamp 1586364061
transform 1 0 152168 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1654
timestamp 1586364061
transform 1 0 153272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1666
timestamp 1586364061
transform 1 0 154376 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 155480 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1679
timestamp 1586364061
transform 1 0 155572 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1691
timestamp 1586364061
transform 1 0 156676 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1703
timestamp 1586364061
transform 1 0 157780 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1715
timestamp 1586364061
transform 1 0 158884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1727
timestamp 1586364061
transform 1 0 159988 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 161092 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1740
timestamp 1586364061
transform 1 0 161184 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1752
timestamp 1586364061
transform 1 0 162288 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1764
timestamp 1586364061
transform 1 0 163392 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1776
timestamp 1586364061
transform 1 0 164496 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 166704 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1788
timestamp 1586364061
transform 1 0 165600 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1801
timestamp 1586364061
transform 1 0 166796 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1813
timestamp 1586364061
transform 1 0 167900 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1825
timestamp 1586364061
transform 1 0 169004 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1837
timestamp 1586364061
transform 1 0 170108 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1849
timestamp 1586364061
transform 1 0 171212 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 172316 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1862
timestamp 1586364061
transform 1 0 172408 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1874
timestamp 1586364061
transform 1 0 173512 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1886
timestamp 1586364061
transform 1 0 174616 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1898
timestamp 1586364061
transform 1 0 175720 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 177928 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1910
timestamp 1586364061
transform 1 0 176824 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1923
timestamp 1586364061
transform 1 0 178020 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1935
timestamp 1586364061
transform 1 0 179124 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1947
timestamp 1586364061
transform 1 0 180228 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1959
timestamp 1586364061
transform 1 0 181332 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1971
timestamp 1586364061
transform 1 0 182436 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 183540 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_1984
timestamp 1586364061
transform 1 0 183632 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_1996
timestamp 1586364061
transform 1 0 184736 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2008
timestamp 1586364061
transform 1 0 185840 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2020
timestamp 1586364061
transform 1 0 186944 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2032
timestamp 1586364061
transform 1 0 188048 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 189152 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_2045
timestamp 1586364061
transform 1 0 189244 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2057
timestamp 1586364061
transform 1 0 190348 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2069
timestamp 1586364061
transform 1 0 191452 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2081
timestamp 1586364061
transform 1 0 192556 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2093
timestamp 1586364061
transform 1 0 193660 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 194764 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_2106
timestamp 1586364061
transform 1 0 194856 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2118
timestamp 1586364061
transform 1 0 195960 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2130
timestamp 1586364061
transform 1 0 197064 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2142
timestamp 1586364061
transform 1 0 198168 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2154
timestamp 1586364061
transform 1 0 199272 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 200376 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_2167
timestamp 1586364061
transform 1 0 200468 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2179
timestamp 1586364061
transform 1 0 201572 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2191
timestamp 1586364061
transform 1 0 202676 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2203
timestamp 1586364061
transform 1 0 203780 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 205988 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_2215
timestamp 1586364061
transform 1 0 204884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2228
timestamp 1586364061
transform 1 0 206080 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2240
timestamp 1586364061
transform 1 0 207184 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2252
timestamp 1586364061
transform 1 0 208288 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2264
timestamp 1586364061
transform 1 0 209392 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2276
timestamp 1586364061
transform 1 0 210496 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 211600 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_2289
timestamp 1586364061
transform 1 0 211692 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2301
timestamp 1586364061
transform 1 0 212796 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2313
timestamp 1586364061
transform 1 0 213900 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2325
timestamp 1586364061
transform 1 0 215004 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 217212 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__14__A
timestamp 1586364061
transform 1 0 217672 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_2337
timestamp 1586364061
transform 1 0 216108 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_2_2350
timestamp 1586364061
transform 1 0 217304 0 -1 3808
box -38 -48 406 592
use scs8hd_nor4_4  _13_
timestamp 1586364061
transform 1 0 218592 0 -1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 218224 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_2356
timestamp 1586364061
transform 1 0 217856 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_2362
timestamp 1586364061
transform 1 0 218408 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 220892 0 -1 3808
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__07__A
timestamp 1586364061
transform 1 0 220340 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__12__A
timestamp 1586364061
transform 1 0 220708 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_2381
timestamp 1586364061
transform 1 0 220156 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_2385
timestamp 1586364061
transform 1 0 220524 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_2397
timestamp 1586364061
transform 1 0 221628 0 -1 3808
box -38 -48 1142 592
use scs8hd_buf_1  _04_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 222916 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 222824 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__15__B
timestamp 1586364061
transform 1 0 223376 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_2409
timestamp 1586364061
transform 1 0 222732 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_2414
timestamp 1586364061
transform 1 0 223192 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_2418
timestamp 1586364061
transform 1 0 223560 0 -1 3808
box -38 -48 1142 592
use scs8hd_and4_4  _05_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 224848 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__09__D
timestamp 1586364061
transform 1 0 225860 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_2430
timestamp 1586364061
transform 1 0 224664 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_2441
timestamp 1586364061
transform 1 0 225676 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_2445
timestamp 1586364061
transform 1 0 226044 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2457
timestamp 1586364061
transform 1 0 227148 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 228436 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_2469
timestamp 1586364061
transform 1 0 228252 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_2472
timestamp 1586364061
transform 1 0 228528 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2484
timestamp 1586364061
transform 1 0 229632 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2496
timestamp 1586364061
transform 1 0 230736 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2508
timestamp 1586364061
transform 1 0 231840 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 234048 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_2520
timestamp 1586364061
transform 1 0 232944 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2533
timestamp 1586364061
transform 1 0 234140 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2545
timestamp 1586364061
transform 1 0 235244 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2557
timestamp 1586364061
transform 1 0 236348 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2569
timestamp 1586364061
transform 1 0 237452 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2581
timestamp 1586364061
transform 1 0 238556 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 239660 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_2594
timestamp 1586364061
transform 1 0 239752 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2606
timestamp 1586364061
transform 1 0 240856 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2618
timestamp 1586364061
transform 1 0 241960 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2630
timestamp 1586364061
transform 1 0 243064 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 245272 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_2642
timestamp 1586364061
transform 1 0 244168 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2655
timestamp 1586364061
transform 1 0 245364 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2667
timestamp 1586364061
transform 1 0 246468 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2679
timestamp 1586364061
transform 1 0 247572 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2691
timestamp 1586364061
transform 1 0 248676 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2703
timestamp 1586364061
transform 1 0 249780 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_286
timestamp 1586364061
transform 1 0 250884 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_2716
timestamp 1586364061
transform 1 0 250976 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2728
timestamp 1586364061
transform 1 0 252080 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2740
timestamp 1586364061
transform 1 0 253184 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2752
timestamp 1586364061
transform 1 0 254288 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2764
timestamp 1586364061
transform 1 0 255392 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_287
timestamp 1586364061
transform 1 0 256496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_2777
timestamp 1586364061
transform 1 0 256588 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2789
timestamp 1586364061
transform 1 0 257692 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2801
timestamp 1586364061
transform 1 0 258796 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2813
timestamp 1586364061
transform 1 0 259900 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2825
timestamp 1586364061
transform 1 0 261004 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_288
timestamp 1586364061
transform 1 0 262108 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_2838
timestamp 1586364061
transform 1 0 262200 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2850
timestamp 1586364061
transform 1 0 263304 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2862
timestamp 1586364061
transform 1 0 264408 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2874
timestamp 1586364061
transform 1 0 265512 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2886
timestamp 1586364061
transform 1 0 266616 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_289
timestamp 1586364061
transform 1 0 267720 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_2899
timestamp 1586364061
transform 1 0 267812 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2911
timestamp 1586364061
transform 1 0 268916 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2923
timestamp 1586364061
transform 1 0 270020 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2935
timestamp 1586364061
transform 1 0 271124 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_290
timestamp 1586364061
transform 1 0 273332 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_2947
timestamp 1586364061
transform 1 0 272228 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2960
timestamp 1586364061
transform 1 0 273424 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2972
timestamp 1586364061
transform 1 0 274528 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2984
timestamp 1586364061
transform 1 0 275632 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_2996
timestamp 1586364061
transform 1 0 276736 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3008
timestamp 1586364061
transform 1 0 277840 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_291
timestamp 1586364061
transform 1 0 278944 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3021
timestamp 1586364061
transform 1 0 279036 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3033
timestamp 1586364061
transform 1 0 280140 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3045
timestamp 1586364061
transform 1 0 281244 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3057
timestamp 1586364061
transform 1 0 282348 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_292
timestamp 1586364061
transform 1 0 284556 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3069
timestamp 1586364061
transform 1 0 283452 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3082
timestamp 1586364061
transform 1 0 284648 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3094
timestamp 1586364061
transform 1 0 285752 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3106
timestamp 1586364061
transform 1 0 286856 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3118
timestamp 1586364061
transform 1 0 287960 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3130
timestamp 1586364061
transform 1 0 289064 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_293
timestamp 1586364061
transform 1 0 290168 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3143
timestamp 1586364061
transform 1 0 290260 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3155
timestamp 1586364061
transform 1 0 291364 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3167
timestamp 1586364061
transform 1 0 292468 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3179
timestamp 1586364061
transform 1 0 293572 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3191
timestamp 1586364061
transform 1 0 294676 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_294
timestamp 1586364061
transform 1 0 295780 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3204
timestamp 1586364061
transform 1 0 295872 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3216
timestamp 1586364061
transform 1 0 296976 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3228
timestamp 1586364061
transform 1 0 298080 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3240
timestamp 1586364061
transform 1 0 299184 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_295
timestamp 1586364061
transform 1 0 301392 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3252
timestamp 1586364061
transform 1 0 300288 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3265
timestamp 1586364061
transform 1 0 301484 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3277
timestamp 1586364061
transform 1 0 302588 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3289
timestamp 1586364061
transform 1 0 303692 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3301
timestamp 1586364061
transform 1 0 304796 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3313
timestamp 1586364061
transform 1 0 305900 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_296
timestamp 1586364061
transform 1 0 307004 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3326
timestamp 1586364061
transform 1 0 307096 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3338
timestamp 1586364061
transform 1 0 308200 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3350
timestamp 1586364061
transform 1 0 309304 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3362
timestamp 1586364061
transform 1 0 310408 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_297
timestamp 1586364061
transform 1 0 312616 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3374
timestamp 1586364061
transform 1 0 311512 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3387
timestamp 1586364061
transform 1 0 312708 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3399
timestamp 1586364061
transform 1 0 313812 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3411
timestamp 1586364061
transform 1 0 314916 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3423
timestamp 1586364061
transform 1 0 316020 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3435
timestamp 1586364061
transform 1 0 317124 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_298
timestamp 1586364061
transform 1 0 318228 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3448
timestamp 1586364061
transform 1 0 318320 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3460
timestamp 1586364061
transform 1 0 319424 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3472
timestamp 1586364061
transform 1 0 320528 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3484
timestamp 1586364061
transform 1 0 321632 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3496
timestamp 1586364061
transform 1 0 322736 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_299
timestamp 1586364061
transform 1 0 323840 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3509
timestamp 1586364061
transform 1 0 323932 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3521
timestamp 1586364061
transform 1 0 325036 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3533
timestamp 1586364061
transform 1 0 326140 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3545
timestamp 1586364061
transform 1 0 327244 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3557
timestamp 1586364061
transform 1 0 328348 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_300
timestamp 1586364061
transform 1 0 329452 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3570
timestamp 1586364061
transform 1 0 329544 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3582
timestamp 1586364061
transform 1 0 330648 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3594
timestamp 1586364061
transform 1 0 331752 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3606
timestamp 1586364061
transform 1 0 332856 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3618
timestamp 1586364061
transform 1 0 333960 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_301
timestamp 1586364061
transform 1 0 335064 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3631
timestamp 1586364061
transform 1 0 335156 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3643
timestamp 1586364061
transform 1 0 336260 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3655
timestamp 1586364061
transform 1 0 337364 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3667
timestamp 1586364061
transform 1 0 338468 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_302
timestamp 1586364061
transform 1 0 340676 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3679
timestamp 1586364061
transform 1 0 339572 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3692
timestamp 1586364061
transform 1 0 340768 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3704
timestamp 1586364061
transform 1 0 341872 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3716
timestamp 1586364061
transform 1 0 342976 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3728
timestamp 1586364061
transform 1 0 344080 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3740
timestamp 1586364061
transform 1 0 345184 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_303
timestamp 1586364061
transform 1 0 346288 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3753
timestamp 1586364061
transform 1 0 346380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3765
timestamp 1586364061
transform 1 0 347484 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3777
timestamp 1586364061
transform 1 0 348588 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3789
timestamp 1586364061
transform 1 0 349692 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_304
timestamp 1586364061
transform 1 0 351900 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3801
timestamp 1586364061
transform 1 0 350796 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3814
timestamp 1586364061
transform 1 0 351992 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3826
timestamp 1586364061
transform 1 0 353096 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3838
timestamp 1586364061
transform 1 0 354200 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3850
timestamp 1586364061
transform 1 0 355304 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3862
timestamp 1586364061
transform 1 0 356408 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_305
timestamp 1586364061
transform 1 0 357512 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3875
timestamp 1586364061
transform 1 0 357604 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3887
timestamp 1586364061
transform 1 0 358708 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3899
timestamp 1586364061
transform 1 0 359812 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3911
timestamp 1586364061
transform 1 0 360916 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3923
timestamp 1586364061
transform 1 0 362020 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_306
timestamp 1586364061
transform 1 0 363124 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3936
timestamp 1586364061
transform 1 0 363216 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3948
timestamp 1586364061
transform 1 0 364320 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3960
timestamp 1586364061
transform 1 0 365424 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3972
timestamp 1586364061
transform 1 0 366528 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_3984
timestamp 1586364061
transform 1 0 367632 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_307
timestamp 1586364061
transform 1 0 368736 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_3997
timestamp 1586364061
transform 1 0 368828 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4009
timestamp 1586364061
transform 1 0 369932 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4021
timestamp 1586364061
transform 1 0 371036 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4033
timestamp 1586364061
transform 1 0 372140 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4045
timestamp 1586364061
transform 1 0 373244 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_308
timestamp 1586364061
transform 1 0 374348 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_4058
timestamp 1586364061
transform 1 0 374440 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4070
timestamp 1586364061
transform 1 0 375544 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4082
timestamp 1586364061
transform 1 0 376648 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4094
timestamp 1586364061
transform 1 0 377752 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_309
timestamp 1586364061
transform 1 0 379960 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_4106
timestamp 1586364061
transform 1 0 378856 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4119
timestamp 1586364061
transform 1 0 380052 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4131
timestamp 1586364061
transform 1 0 381156 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4143
timestamp 1586364061
transform 1 0 382260 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4155
timestamp 1586364061
transform 1 0 383364 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4167
timestamp 1586364061
transform 1 0 384468 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_310
timestamp 1586364061
transform 1 0 385572 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_4180
timestamp 1586364061
transform 1 0 385664 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4192
timestamp 1586364061
transform 1 0 386768 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4204
timestamp 1586364061
transform 1 0 387872 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4216
timestamp 1586364061
transform 1 0 388976 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_311
timestamp 1586364061
transform 1 0 391184 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_4228
timestamp 1586364061
transform 1 0 390080 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4241
timestamp 1586364061
transform 1 0 391276 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4253
timestamp 1586364061
transform 1 0 392380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4265
timestamp 1586364061
transform 1 0 393484 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4277
timestamp 1586364061
transform 1 0 394588 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4289
timestamp 1586364061
transform 1 0 395692 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_312
timestamp 1586364061
transform 1 0 396796 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_4302
timestamp 1586364061
transform 1 0 396888 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4314
timestamp 1586364061
transform 1 0 397992 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4326
timestamp 1586364061
transform 1 0 399096 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4338
timestamp 1586364061
transform 1 0 400200 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4350
timestamp 1586364061
transform 1 0 401304 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_313
timestamp 1586364061
transform 1 0 402408 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_4363
timestamp 1586364061
transform 1 0 402500 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4375
timestamp 1586364061
transform 1 0 403604 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4387
timestamp 1586364061
transform 1 0 404708 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4399
timestamp 1586364061
transform 1 0 405812 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_314
timestamp 1586364061
transform 1 0 408020 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_4411
timestamp 1586364061
transform 1 0 406916 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4424
timestamp 1586364061
transform 1 0 408112 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4436
timestamp 1586364061
transform 1 0 409216 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4448
timestamp 1586364061
transform 1 0 410320 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4460
timestamp 1586364061
transform 1 0 411424 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4472
timestamp 1586364061
transform 1 0 412528 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_315
timestamp 1586364061
transform 1 0 413632 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_4485
timestamp 1586364061
transform 1 0 413724 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4497
timestamp 1586364061
transform 1 0 414828 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4509
timestamp 1586364061
transform 1 0 415932 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4521
timestamp 1586364061
transform 1 0 417036 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_316
timestamp 1586364061
transform 1 0 419244 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_4533
timestamp 1586364061
transform 1 0 418140 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4546
timestamp 1586364061
transform 1 0 419336 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_4558
timestamp 1586364061
transform 1 0 420440 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 422832 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_4570
timestamp 1586364061
transform 1 0 421544 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_2_4578
timestamp 1586364061
transform 1 0 422280 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_317
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_318
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_110
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_319
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_320
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_232
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_281
timestamp 1586364061
transform 1 0 26956 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_293
timestamp 1586364061
transform 1 0 28060 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_321
timestamp 1586364061
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_306
timestamp 1586364061
transform 1 0 29256 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_318
timestamp 1586364061
transform 1 0 30360 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_330
timestamp 1586364061
transform 1 0 31464 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_342
timestamp 1586364061
transform 1 0 32568 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_354
timestamp 1586364061
transform 1 0 33672 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_322
timestamp 1586364061
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_367
timestamp 1586364061
transform 1 0 34868 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_379
timestamp 1586364061
transform 1 0 35972 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_391
timestamp 1586364061
transform 1 0 37076 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_403
timestamp 1586364061
transform 1 0 38180 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_323
timestamp 1586364061
transform 1 0 40388 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_415
timestamp 1586364061
transform 1 0 39284 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_428
timestamp 1586364061
transform 1 0 40480 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_440
timestamp 1586364061
transform 1 0 41584 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_452
timestamp 1586364061
transform 1 0 42688 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_464
timestamp 1586364061
transform 1 0 43792 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_476
timestamp 1586364061
transform 1 0 44896 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_324
timestamp 1586364061
transform 1 0 46000 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_489
timestamp 1586364061
transform 1 0 46092 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_501
timestamp 1586364061
transform 1 0 47196 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_513
timestamp 1586364061
transform 1 0 48300 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_525
timestamp 1586364061
transform 1 0 49404 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_325
timestamp 1586364061
transform 1 0 51612 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_537
timestamp 1586364061
transform 1 0 50508 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_550
timestamp 1586364061
transform 1 0 51704 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_562
timestamp 1586364061
transform 1 0 52808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_574
timestamp 1586364061
transform 1 0 53912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_586
timestamp 1586364061
transform 1 0 55016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_598
timestamp 1586364061
transform 1 0 56120 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_326
timestamp 1586364061
transform 1 0 57224 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_611
timestamp 1586364061
transform 1 0 57316 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_623
timestamp 1586364061
transform 1 0 58420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_635
timestamp 1586364061
transform 1 0 59524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_647
timestamp 1586364061
transform 1 0 60628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_659
timestamp 1586364061
transform 1 0 61732 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_327
timestamp 1586364061
transform 1 0 62836 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_672
timestamp 1586364061
transform 1 0 62928 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_684
timestamp 1586364061
transform 1 0 64032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_696
timestamp 1586364061
transform 1 0 65136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_708
timestamp 1586364061
transform 1 0 66240 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_720
timestamp 1586364061
transform 1 0 67344 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_328
timestamp 1586364061
transform 1 0 68448 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_733
timestamp 1586364061
transform 1 0 68540 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_745
timestamp 1586364061
transform 1 0 69644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_757
timestamp 1586364061
transform 1 0 70748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_769
timestamp 1586364061
transform 1 0 71852 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_781
timestamp 1586364061
transform 1 0 72956 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_329
timestamp 1586364061
transform 1 0 74060 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_794
timestamp 1586364061
transform 1 0 74152 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_806
timestamp 1586364061
transform 1 0 75256 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_818
timestamp 1586364061
transform 1 0 76360 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_830
timestamp 1586364061
transform 1 0 77464 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_330
timestamp 1586364061
transform 1 0 79672 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_842
timestamp 1586364061
transform 1 0 78568 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_855
timestamp 1586364061
transform 1 0 79764 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_867
timestamp 1586364061
transform 1 0 80868 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_879
timestamp 1586364061
transform 1 0 81972 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_891
timestamp 1586364061
transform 1 0 83076 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_903
timestamp 1586364061
transform 1 0 84180 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_331
timestamp 1586364061
transform 1 0 85284 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_916
timestamp 1586364061
transform 1 0 85376 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_928
timestamp 1586364061
transform 1 0 86480 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_940
timestamp 1586364061
transform 1 0 87584 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_952
timestamp 1586364061
transform 1 0 88688 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_332
timestamp 1586364061
transform 1 0 90896 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_964
timestamp 1586364061
transform 1 0 89792 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_977
timestamp 1586364061
transform 1 0 90988 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_989
timestamp 1586364061
transform 1 0 92092 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1001
timestamp 1586364061
transform 1 0 93196 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1013
timestamp 1586364061
transform 1 0 94300 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1025
timestamp 1586364061
transform 1 0 95404 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_333
timestamp 1586364061
transform 1 0 96508 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1038
timestamp 1586364061
transform 1 0 96600 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1050
timestamp 1586364061
transform 1 0 97704 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1062
timestamp 1586364061
transform 1 0 98808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1074
timestamp 1586364061
transform 1 0 99912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1086
timestamp 1586364061
transform 1 0 101016 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_334
timestamp 1586364061
transform 1 0 102120 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1099
timestamp 1586364061
transform 1 0 102212 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1111
timestamp 1586364061
transform 1 0 103316 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1123
timestamp 1586364061
transform 1 0 104420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1135
timestamp 1586364061
transform 1 0 105524 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_335
timestamp 1586364061
transform 1 0 107732 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1147
timestamp 1586364061
transform 1 0 106628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1160
timestamp 1586364061
transform 1 0 107824 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1172
timestamp 1586364061
transform 1 0 108928 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1184
timestamp 1586364061
transform 1 0 110032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1196
timestamp 1586364061
transform 1 0 111136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1208
timestamp 1586364061
transform 1 0 112240 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_336
timestamp 1586364061
transform 1 0 113344 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1221
timestamp 1586364061
transform 1 0 113436 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1233
timestamp 1586364061
transform 1 0 114540 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1245
timestamp 1586364061
transform 1 0 115644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1257
timestamp 1586364061
transform 1 0 116748 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_337
timestamp 1586364061
transform 1 0 118956 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1269
timestamp 1586364061
transform 1 0 117852 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1282
timestamp 1586364061
transform 1 0 119048 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1294
timestamp 1586364061
transform 1 0 120152 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1306
timestamp 1586364061
transform 1 0 121256 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1318
timestamp 1586364061
transform 1 0 122360 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1330
timestamp 1586364061
transform 1 0 123464 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_338
timestamp 1586364061
transform 1 0 124568 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1343
timestamp 1586364061
transform 1 0 124660 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1355
timestamp 1586364061
transform 1 0 125764 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1367
timestamp 1586364061
transform 1 0 126868 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1379
timestamp 1586364061
transform 1 0 127972 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1391
timestamp 1586364061
transform 1 0 129076 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_339
timestamp 1586364061
transform 1 0 130180 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1404
timestamp 1586364061
transform 1 0 130272 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1416
timestamp 1586364061
transform 1 0 131376 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1428
timestamp 1586364061
transform 1 0 132480 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1440
timestamp 1586364061
transform 1 0 133584 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1452
timestamp 1586364061
transform 1 0 134688 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_340
timestamp 1586364061
transform 1 0 135792 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1465
timestamp 1586364061
transform 1 0 135884 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1477
timestamp 1586364061
transform 1 0 136988 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1489
timestamp 1586364061
transform 1 0 138092 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1501
timestamp 1586364061
transform 1 0 139196 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1513
timestamp 1586364061
transform 1 0 140300 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_341
timestamp 1586364061
transform 1 0 141404 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1526
timestamp 1586364061
transform 1 0 141496 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1538
timestamp 1586364061
transform 1 0 142600 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1550
timestamp 1586364061
transform 1 0 143704 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1562
timestamp 1586364061
transform 1 0 144808 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_342
timestamp 1586364061
transform 1 0 147016 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1574
timestamp 1586364061
transform 1 0 145912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1587
timestamp 1586364061
transform 1 0 147108 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1599
timestamp 1586364061
transform 1 0 148212 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1611
timestamp 1586364061
transform 1 0 149316 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1623
timestamp 1586364061
transform 1 0 150420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1635
timestamp 1586364061
transform 1 0 151524 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_343
timestamp 1586364061
transform 1 0 152628 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1648
timestamp 1586364061
transform 1 0 152720 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1660
timestamp 1586364061
transform 1 0 153824 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1672
timestamp 1586364061
transform 1 0 154928 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1684
timestamp 1586364061
transform 1 0 156032 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_344
timestamp 1586364061
transform 1 0 158240 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1696
timestamp 1586364061
transform 1 0 157136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1709
timestamp 1586364061
transform 1 0 158332 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1721
timestamp 1586364061
transform 1 0 159436 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1733
timestamp 1586364061
transform 1 0 160540 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1745
timestamp 1586364061
transform 1 0 161644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1757
timestamp 1586364061
transform 1 0 162748 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_345
timestamp 1586364061
transform 1 0 163852 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1770
timestamp 1586364061
transform 1 0 163944 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1782
timestamp 1586364061
transform 1 0 165048 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1794
timestamp 1586364061
transform 1 0 166152 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1806
timestamp 1586364061
transform 1 0 167256 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1818
timestamp 1586364061
transform 1 0 168360 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_346
timestamp 1586364061
transform 1 0 169464 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1831
timestamp 1586364061
transform 1 0 169556 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1843
timestamp 1586364061
transform 1 0 170660 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1855
timestamp 1586364061
transform 1 0 171764 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1867
timestamp 1586364061
transform 1 0 172868 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1879
timestamp 1586364061
transform 1 0 173972 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_347
timestamp 1586364061
transform 1 0 175076 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1892
timestamp 1586364061
transform 1 0 175168 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1904
timestamp 1586364061
transform 1 0 176272 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1916
timestamp 1586364061
transform 1 0 177376 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1928
timestamp 1586364061
transform 1 0 178480 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1940
timestamp 1586364061
transform 1 0 179584 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_348
timestamp 1586364061
transform 1 0 180688 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_1953
timestamp 1586364061
transform 1 0 180780 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1965
timestamp 1586364061
transform 1 0 181884 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1977
timestamp 1586364061
transform 1 0 182988 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_1989
timestamp 1586364061
transform 1 0 184092 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_349
timestamp 1586364061
transform 1 0 186300 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_2001
timestamp 1586364061
transform 1 0 185196 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2014
timestamp 1586364061
transform 1 0 186392 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2026
timestamp 1586364061
transform 1 0 187496 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2038
timestamp 1586364061
transform 1 0 188600 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2050
timestamp 1586364061
transform 1 0 189704 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2062
timestamp 1586364061
transform 1 0 190808 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_350
timestamp 1586364061
transform 1 0 191912 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_2075
timestamp 1586364061
transform 1 0 192004 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2087
timestamp 1586364061
transform 1 0 193108 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2099
timestamp 1586364061
transform 1 0 194212 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2111
timestamp 1586364061
transform 1 0 195316 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_351
timestamp 1586364061
transform 1 0 197524 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_2123
timestamp 1586364061
transform 1 0 196420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2136
timestamp 1586364061
transform 1 0 197616 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2148
timestamp 1586364061
transform 1 0 198720 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2160
timestamp 1586364061
transform 1 0 199824 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2172
timestamp 1586364061
transform 1 0 200928 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2184
timestamp 1586364061
transform 1 0 202032 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_352
timestamp 1586364061
transform 1 0 203136 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_2197
timestamp 1586364061
transform 1 0 203228 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2209
timestamp 1586364061
transform 1 0 204332 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2221
timestamp 1586364061
transform 1 0 205436 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2233
timestamp 1586364061
transform 1 0 206540 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2245
timestamp 1586364061
transform 1 0 207644 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_353
timestamp 1586364061
transform 1 0 208748 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_2258
timestamp 1586364061
transform 1 0 208840 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2270
timestamp 1586364061
transform 1 0 209944 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2282
timestamp 1586364061
transform 1 0 211048 0 1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 212336 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 212704 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_2294
timestamp 1586364061
transform 1 0 212152 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_2298
timestamp 1586364061
transform 1 0 212520 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_354
timestamp 1586364061
transform 1 0 214360 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_2302
timestamp 1586364061
transform 1 0 212888 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_3_2314
timestamp 1586364061
transform 1 0 213992 0 1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_3_2319
timestamp 1586364061
transform 1 0 214452 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_3_2331
timestamp 1586364061
transform 1 0 215556 0 1 3808
box -38 -48 590 592
use scs8hd_inv_8  _06_
timestamp 1586364061
transform 1 0 216292 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__06__A
timestamp 1586364061
transform 1 0 216108 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 217672 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_2348
timestamp 1586364061
transform 1 0 217120 0 1 3808
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 218224 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 218040 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_2356
timestamp 1586364061
transform 1 0 217856 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_2371
timestamp 1586364061
transform 1 0 219236 0 1 3808
box -38 -48 222 592
use scs8hd_and4_4  _07_
timestamp 1586364061
transform 1 0 220064 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_355
timestamp 1586364061
transform 1 0 219972 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__07__B
timestamp 1586364061
transform 1 0 219788 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__07__D
timestamp 1586364061
transform 1 0 219420 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_2375
timestamp 1586364061
transform 1 0 219604 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_2389
timestamp 1586364061
transform 1 0 220892 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__15__C
timestamp 1586364061
transform 1 0 222548 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__12__C
timestamp 1586364061
transform 1 0 221076 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__07__C
timestamp 1586364061
transform 1 0 221444 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__12__D
timestamp 1586364061
transform 1 0 221812 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__12__B
timestamp 1586364061
transform 1 0 222180 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_2393
timestamp 1586364061
transform 1 0 221260 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_2397
timestamp 1586364061
transform 1 0 221628 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_2401
timestamp 1586364061
transform 1 0 221996 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_2405
timestamp 1586364061
transform 1 0 222364 0 1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _15_
timestamp 1586364061
transform 1 0 223100 0 1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__15__A
timestamp 1586364061
transform 1 0 222916 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_2409
timestamp 1586364061
transform 1 0 222732 0 1 3808
box -38 -48 222 592
use scs8hd_and4_4  _09_
timestamp 1586364061
transform 1 0 225676 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_356
timestamp 1586364061
transform 1 0 225584 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__09__A
timestamp 1586364061
transform 1 0 225400 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__09__B
timestamp 1586364061
transform 1 0 225032 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_2430
timestamp 1586364061
transform 1 0 224664 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_2436
timestamp 1586364061
transform 1 0 225216 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_2450
timestamp 1586364061
transform 1 0 226504 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2462
timestamp 1586364061
transform 1 0 227608 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2474
timestamp 1586364061
transform 1 0 228712 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2486
timestamp 1586364061
transform 1 0 229816 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_357
timestamp 1586364061
transform 1 0 231196 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 232300 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_2498
timestamp 1586364061
transform 1 0 230920 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_2502
timestamp 1586364061
transform 1 0 231288 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_3_2510
timestamp 1586364061
transform 1 0 232024 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_2515
timestamp 1586364061
transform 1 0 232484 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 232668 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_2519
timestamp 1586364061
transform 1 0 232852 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2531
timestamp 1586364061
transform 1 0 233956 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2543
timestamp 1586364061
transform 1 0 235060 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_358
timestamp 1586364061
transform 1 0 236808 0 1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_3_2555
timestamp 1586364061
transform 1 0 236164 0 1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_3_2561
timestamp 1586364061
transform 1 0 236716 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_2563
timestamp 1586364061
transform 1 0 236900 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2575
timestamp 1586364061
transform 1 0 238004 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2587
timestamp 1586364061
transform 1 0 239108 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2599
timestamp 1586364061
transform 1 0 240212 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2611
timestamp 1586364061
transform 1 0 241316 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_359
timestamp 1586364061
transform 1 0 242420 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_2624
timestamp 1586364061
transform 1 0 242512 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2636
timestamp 1586364061
transform 1 0 243616 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2648
timestamp 1586364061
transform 1 0 244720 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2660
timestamp 1586364061
transform 1 0 245824 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2672
timestamp 1586364061
transform 1 0 246928 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_360
timestamp 1586364061
transform 1 0 248032 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_2685
timestamp 1586364061
transform 1 0 248124 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2697
timestamp 1586364061
transform 1 0 249228 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2709
timestamp 1586364061
transform 1 0 250332 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2721
timestamp 1586364061
transform 1 0 251436 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_361
timestamp 1586364061
transform 1 0 253644 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_2733
timestamp 1586364061
transform 1 0 252540 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2746
timestamp 1586364061
transform 1 0 253736 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2758
timestamp 1586364061
transform 1 0 254840 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2770
timestamp 1586364061
transform 1 0 255944 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2782
timestamp 1586364061
transform 1 0 257048 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2794
timestamp 1586364061
transform 1 0 258152 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_362
timestamp 1586364061
transform 1 0 259256 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_2807
timestamp 1586364061
transform 1 0 259348 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2819
timestamp 1586364061
transform 1 0 260452 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2831
timestamp 1586364061
transform 1 0 261556 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2843
timestamp 1586364061
transform 1 0 262660 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_363
timestamp 1586364061
transform 1 0 264868 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_2855
timestamp 1586364061
transform 1 0 263764 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2868
timestamp 1586364061
transform 1 0 264960 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2880
timestamp 1586364061
transform 1 0 266064 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2892
timestamp 1586364061
transform 1 0 267168 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2904
timestamp 1586364061
transform 1 0 268272 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2916
timestamp 1586364061
transform 1 0 269376 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_364
timestamp 1586364061
transform 1 0 270480 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_2929
timestamp 1586364061
transform 1 0 270572 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2941
timestamp 1586364061
transform 1 0 271676 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2953
timestamp 1586364061
transform 1 0 272780 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2965
timestamp 1586364061
transform 1 0 273884 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_2977
timestamp 1586364061
transform 1 0 274988 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_365
timestamp 1586364061
transform 1 0 276092 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_2990
timestamp 1586364061
transform 1 0 276184 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3002
timestamp 1586364061
transform 1 0 277288 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3014
timestamp 1586364061
transform 1 0 278392 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3026
timestamp 1586364061
transform 1 0 279496 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_366
timestamp 1586364061
transform 1 0 281704 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3038
timestamp 1586364061
transform 1 0 280600 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3051
timestamp 1586364061
transform 1 0 281796 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3063
timestamp 1586364061
transform 1 0 282900 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3075
timestamp 1586364061
transform 1 0 284004 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3087
timestamp 1586364061
transform 1 0 285108 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3099
timestamp 1586364061
transform 1 0 286212 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_367
timestamp 1586364061
transform 1 0 287316 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3112
timestamp 1586364061
transform 1 0 287408 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3124
timestamp 1586364061
transform 1 0 288512 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3136
timestamp 1586364061
transform 1 0 289616 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3148
timestamp 1586364061
transform 1 0 290720 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_368
timestamp 1586364061
transform 1 0 292928 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3160
timestamp 1586364061
transform 1 0 291824 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3173
timestamp 1586364061
transform 1 0 293020 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3185
timestamp 1586364061
transform 1 0 294124 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3197
timestamp 1586364061
transform 1 0 295228 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3209
timestamp 1586364061
transform 1 0 296332 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3221
timestamp 1586364061
transform 1 0 297436 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_369
timestamp 1586364061
transform 1 0 298540 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3234
timestamp 1586364061
transform 1 0 298632 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3246
timestamp 1586364061
transform 1 0 299736 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3258
timestamp 1586364061
transform 1 0 300840 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3270
timestamp 1586364061
transform 1 0 301944 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_370
timestamp 1586364061
transform 1 0 304152 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3282
timestamp 1586364061
transform 1 0 303048 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3295
timestamp 1586364061
transform 1 0 304244 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3307
timestamp 1586364061
transform 1 0 305348 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3319
timestamp 1586364061
transform 1 0 306452 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3331
timestamp 1586364061
transform 1 0 307556 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3343
timestamp 1586364061
transform 1 0 308660 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_371
timestamp 1586364061
transform 1 0 309764 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3356
timestamp 1586364061
transform 1 0 309856 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3368
timestamp 1586364061
transform 1 0 310960 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3380
timestamp 1586364061
transform 1 0 312064 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3392
timestamp 1586364061
transform 1 0 313168 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3404
timestamp 1586364061
transform 1 0 314272 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_372
timestamp 1586364061
transform 1 0 315376 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3417
timestamp 1586364061
transform 1 0 315468 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3429
timestamp 1586364061
transform 1 0 316572 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3441
timestamp 1586364061
transform 1 0 317676 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3453
timestamp 1586364061
transform 1 0 318780 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_373
timestamp 1586364061
transform 1 0 320988 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3465
timestamp 1586364061
transform 1 0 319884 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3478
timestamp 1586364061
transform 1 0 321080 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3490
timestamp 1586364061
transform 1 0 322184 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3502
timestamp 1586364061
transform 1 0 323288 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3514
timestamp 1586364061
transform 1 0 324392 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3526
timestamp 1586364061
transform 1 0 325496 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_374
timestamp 1586364061
transform 1 0 326600 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3539
timestamp 1586364061
transform 1 0 326692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3551
timestamp 1586364061
transform 1 0 327796 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3563
timestamp 1586364061
transform 1 0 328900 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3575
timestamp 1586364061
transform 1 0 330004 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_375
timestamp 1586364061
transform 1 0 332212 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3587
timestamp 1586364061
transform 1 0 331108 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3600
timestamp 1586364061
transform 1 0 332304 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3612
timestamp 1586364061
transform 1 0 333408 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3624
timestamp 1586364061
transform 1 0 334512 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3636
timestamp 1586364061
transform 1 0 335616 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3648
timestamp 1586364061
transform 1 0 336720 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_376
timestamp 1586364061
transform 1 0 337824 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3661
timestamp 1586364061
transform 1 0 337916 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3673
timestamp 1586364061
transform 1 0 339020 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3685
timestamp 1586364061
transform 1 0 340124 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3697
timestamp 1586364061
transform 1 0 341228 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3709
timestamp 1586364061
transform 1 0 342332 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_377
timestamp 1586364061
transform 1 0 343436 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3722
timestamp 1586364061
transform 1 0 343528 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3734
timestamp 1586364061
transform 1 0 344632 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3746
timestamp 1586364061
transform 1 0 345736 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3758
timestamp 1586364061
transform 1 0 346840 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3770
timestamp 1586364061
transform 1 0 347944 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_378
timestamp 1586364061
transform 1 0 349048 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3783
timestamp 1586364061
transform 1 0 349140 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3795
timestamp 1586364061
transform 1 0 350244 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3807
timestamp 1586364061
transform 1 0 351348 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3819
timestamp 1586364061
transform 1 0 352452 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3831
timestamp 1586364061
transform 1 0 353556 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_379
timestamp 1586364061
transform 1 0 354660 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3844
timestamp 1586364061
transform 1 0 354752 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3856
timestamp 1586364061
transform 1 0 355856 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3868
timestamp 1586364061
transform 1 0 356960 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3880
timestamp 1586364061
transform 1 0 358064 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_380
timestamp 1586364061
transform 1 0 360272 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3892
timestamp 1586364061
transform 1 0 359168 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3905
timestamp 1586364061
transform 1 0 360364 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3917
timestamp 1586364061
transform 1 0 361468 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3929
timestamp 1586364061
transform 1 0 362572 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3941
timestamp 1586364061
transform 1 0 363676 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3953
timestamp 1586364061
transform 1 0 364780 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_381
timestamp 1586364061
transform 1 0 365884 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_3966
timestamp 1586364061
transform 1 0 365976 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3978
timestamp 1586364061
transform 1 0 367080 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_3990
timestamp 1586364061
transform 1 0 368184 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4002
timestamp 1586364061
transform 1 0 369288 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_382
timestamp 1586364061
transform 1 0 371496 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_4014
timestamp 1586364061
transform 1 0 370392 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4027
timestamp 1586364061
transform 1 0 371588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4039
timestamp 1586364061
transform 1 0 372692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4051
timestamp 1586364061
transform 1 0 373796 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4063
timestamp 1586364061
transform 1 0 374900 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4075
timestamp 1586364061
transform 1 0 376004 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_383
timestamp 1586364061
transform 1 0 377108 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_4088
timestamp 1586364061
transform 1 0 377200 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4100
timestamp 1586364061
transform 1 0 378304 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4112
timestamp 1586364061
transform 1 0 379408 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4124
timestamp 1586364061
transform 1 0 380512 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4136
timestamp 1586364061
transform 1 0 381616 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_384
timestamp 1586364061
transform 1 0 382720 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_4149
timestamp 1586364061
transform 1 0 382812 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4161
timestamp 1586364061
transform 1 0 383916 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4173
timestamp 1586364061
transform 1 0 385020 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4185
timestamp 1586364061
transform 1 0 386124 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_385
timestamp 1586364061
transform 1 0 388332 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_4197
timestamp 1586364061
transform 1 0 387228 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4210
timestamp 1586364061
transform 1 0 388424 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4222
timestamp 1586364061
transform 1 0 389528 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4234
timestamp 1586364061
transform 1 0 390632 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4246
timestamp 1586364061
transform 1 0 391736 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4258
timestamp 1586364061
transform 1 0 392840 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_386
timestamp 1586364061
transform 1 0 393944 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_4271
timestamp 1586364061
transform 1 0 394036 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4283
timestamp 1586364061
transform 1 0 395140 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4295
timestamp 1586364061
transform 1 0 396244 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4307
timestamp 1586364061
transform 1 0 397348 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_387
timestamp 1586364061
transform 1 0 399556 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_4319
timestamp 1586364061
transform 1 0 398452 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4332
timestamp 1586364061
transform 1 0 399648 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4344
timestamp 1586364061
transform 1 0 400752 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4356
timestamp 1586364061
transform 1 0 401856 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4368
timestamp 1586364061
transform 1 0 402960 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4380
timestamp 1586364061
transform 1 0 404064 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_388
timestamp 1586364061
transform 1 0 405168 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_4393
timestamp 1586364061
transform 1 0 405260 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4405
timestamp 1586364061
transform 1 0 406364 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4417
timestamp 1586364061
transform 1 0 407468 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4429
timestamp 1586364061
transform 1 0 408572 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4441
timestamp 1586364061
transform 1 0 409676 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_389
timestamp 1586364061
transform 1 0 410780 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_4454
timestamp 1586364061
transform 1 0 410872 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4466
timestamp 1586364061
transform 1 0 411976 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4478
timestamp 1586364061
transform 1 0 413080 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4490
timestamp 1586364061
transform 1 0 414184 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4502
timestamp 1586364061
transform 1 0 415288 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_390
timestamp 1586364061
transform 1 0 416392 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_4515
timestamp 1586364061
transform 1 0 416484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4527
timestamp 1586364061
transform 1 0 417588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4539
timestamp 1586364061
transform 1 0 418692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4551
timestamp 1586364061
transform 1 0 419796 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_4563
timestamp 1586364061
transform 1 0 420900 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 422832 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_391
timestamp 1586364061
transform 1 0 422004 0 1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_3_4576
timestamp 1586364061
transform 1 0 422096 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_4580
timestamp 1586364061
transform 1 0 422464 0 1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_392
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_393
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_394
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_395
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_263
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_396
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_288
timestamp 1586364061
transform 1 0 27600 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_300
timestamp 1586364061
transform 1 0 28704 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_312
timestamp 1586364061
transform 1 0 29808 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_397
timestamp 1586364061
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_324
timestamp 1586364061
transform 1 0 30912 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_337
timestamp 1586364061
transform 1 0 32108 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_349
timestamp 1586364061
transform 1 0 33212 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_361
timestamp 1586364061
transform 1 0 34316 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_373
timestamp 1586364061
transform 1 0 35420 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_385
timestamp 1586364061
transform 1 0 36524 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_398
timestamp 1586364061
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_398
timestamp 1586364061
transform 1 0 37720 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_410
timestamp 1586364061
transform 1 0 38824 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_422
timestamp 1586364061
transform 1 0 39928 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_434
timestamp 1586364061
transform 1 0 41032 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_399
timestamp 1586364061
transform 1 0 43240 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_446
timestamp 1586364061
transform 1 0 42136 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_459
timestamp 1586364061
transform 1 0 43332 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_471
timestamp 1586364061
transform 1 0 44436 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_483
timestamp 1586364061
transform 1 0 45540 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_495
timestamp 1586364061
transform 1 0 46644 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_507
timestamp 1586364061
transform 1 0 47748 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_400
timestamp 1586364061
transform 1 0 48852 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_520
timestamp 1586364061
transform 1 0 48944 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_532
timestamp 1586364061
transform 1 0 50048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_544
timestamp 1586364061
transform 1 0 51152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_556
timestamp 1586364061
transform 1 0 52256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_568
timestamp 1586364061
transform 1 0 53360 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_401
timestamp 1586364061
transform 1 0 54464 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_581
timestamp 1586364061
transform 1 0 54556 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_593
timestamp 1586364061
transform 1 0 55660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_605
timestamp 1586364061
transform 1 0 56764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_617
timestamp 1586364061
transform 1 0 57868 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_402
timestamp 1586364061
transform 1 0 60076 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_629
timestamp 1586364061
transform 1 0 58972 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_642
timestamp 1586364061
transform 1 0 60168 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_654
timestamp 1586364061
transform 1 0 61272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_666
timestamp 1586364061
transform 1 0 62376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_678
timestamp 1586364061
transform 1 0 63480 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_690
timestamp 1586364061
transform 1 0 64584 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_403
timestamp 1586364061
transform 1 0 65688 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_703
timestamp 1586364061
transform 1 0 65780 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_715
timestamp 1586364061
transform 1 0 66884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_727
timestamp 1586364061
transform 1 0 67988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_739
timestamp 1586364061
transform 1 0 69092 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_404
timestamp 1586364061
transform 1 0 71300 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_751
timestamp 1586364061
transform 1 0 70196 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_764
timestamp 1586364061
transform 1 0 71392 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_776
timestamp 1586364061
transform 1 0 72496 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_788
timestamp 1586364061
transform 1 0 73600 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_800
timestamp 1586364061
transform 1 0 74704 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_812
timestamp 1586364061
transform 1 0 75808 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_405
timestamp 1586364061
transform 1 0 76912 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_825
timestamp 1586364061
transform 1 0 77004 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_837
timestamp 1586364061
transform 1 0 78108 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_849
timestamp 1586364061
transform 1 0 79212 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_861
timestamp 1586364061
transform 1 0 80316 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_873
timestamp 1586364061
transform 1 0 81420 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_406
timestamp 1586364061
transform 1 0 82524 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_886
timestamp 1586364061
transform 1 0 82616 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_898
timestamp 1586364061
transform 1 0 83720 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_910
timestamp 1586364061
transform 1 0 84824 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_922
timestamp 1586364061
transform 1 0 85928 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_934
timestamp 1586364061
transform 1 0 87032 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_407
timestamp 1586364061
transform 1 0 88136 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_947
timestamp 1586364061
transform 1 0 88228 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_959
timestamp 1586364061
transform 1 0 89332 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_971
timestamp 1586364061
transform 1 0 90436 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_983
timestamp 1586364061
transform 1 0 91540 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_995
timestamp 1586364061
transform 1 0 92644 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_408
timestamp 1586364061
transform 1 0 93748 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1008
timestamp 1586364061
transform 1 0 93840 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1020
timestamp 1586364061
transform 1 0 94944 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1032
timestamp 1586364061
transform 1 0 96048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1044
timestamp 1586364061
transform 1 0 97152 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_409
timestamp 1586364061
transform 1 0 99360 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1056
timestamp 1586364061
transform 1 0 98256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1069
timestamp 1586364061
transform 1 0 99452 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1081
timestamp 1586364061
transform 1 0 100556 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1093
timestamp 1586364061
transform 1 0 101660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1105
timestamp 1586364061
transform 1 0 102764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1117
timestamp 1586364061
transform 1 0 103868 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_410
timestamp 1586364061
transform 1 0 104972 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1130
timestamp 1586364061
transform 1 0 105064 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1142
timestamp 1586364061
transform 1 0 106168 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1154
timestamp 1586364061
transform 1 0 107272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1166
timestamp 1586364061
transform 1 0 108376 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_411
timestamp 1586364061
transform 1 0 110584 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1178
timestamp 1586364061
transform 1 0 109480 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1191
timestamp 1586364061
transform 1 0 110676 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1203
timestamp 1586364061
transform 1 0 111780 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1215
timestamp 1586364061
transform 1 0 112884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1227
timestamp 1586364061
transform 1 0 113988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1239
timestamp 1586364061
transform 1 0 115092 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_412
timestamp 1586364061
transform 1 0 116196 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1252
timestamp 1586364061
transform 1 0 116288 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1264
timestamp 1586364061
transform 1 0 117392 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1276
timestamp 1586364061
transform 1 0 118496 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1288
timestamp 1586364061
transform 1 0 119600 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1300
timestamp 1586364061
transform 1 0 120704 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_413
timestamp 1586364061
transform 1 0 121808 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1313
timestamp 1586364061
transform 1 0 121900 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1325
timestamp 1586364061
transform 1 0 123004 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1337
timestamp 1586364061
transform 1 0 124108 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1349
timestamp 1586364061
transform 1 0 125212 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_414
timestamp 1586364061
transform 1 0 127420 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1361
timestamp 1586364061
transform 1 0 126316 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1374
timestamp 1586364061
transform 1 0 127512 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1386
timestamp 1586364061
transform 1 0 128616 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1398
timestamp 1586364061
transform 1 0 129720 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1410
timestamp 1586364061
transform 1 0 130824 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1422
timestamp 1586364061
transform 1 0 131928 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_415
timestamp 1586364061
transform 1 0 133032 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1435
timestamp 1586364061
transform 1 0 133124 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1447
timestamp 1586364061
transform 1 0 134228 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1459
timestamp 1586364061
transform 1 0 135332 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1471
timestamp 1586364061
transform 1 0 136436 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_416
timestamp 1586364061
transform 1 0 138644 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1483
timestamp 1586364061
transform 1 0 137540 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1496
timestamp 1586364061
transform 1 0 138736 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1508
timestamp 1586364061
transform 1 0 139840 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1520
timestamp 1586364061
transform 1 0 140944 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1532
timestamp 1586364061
transform 1 0 142048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1544
timestamp 1586364061
transform 1 0 143152 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_417
timestamp 1586364061
transform 1 0 144256 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1557
timestamp 1586364061
transform 1 0 144348 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1569
timestamp 1586364061
transform 1 0 145452 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1581
timestamp 1586364061
transform 1 0 146556 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1593
timestamp 1586364061
transform 1 0 147660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1605
timestamp 1586364061
transform 1 0 148764 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_418
timestamp 1586364061
transform 1 0 149868 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1618
timestamp 1586364061
transform 1 0 149960 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1630
timestamp 1586364061
transform 1 0 151064 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1642
timestamp 1586364061
transform 1 0 152168 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1654
timestamp 1586364061
transform 1 0 153272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1666
timestamp 1586364061
transform 1 0 154376 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_419
timestamp 1586364061
transform 1 0 155480 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1679
timestamp 1586364061
transform 1 0 155572 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1691
timestamp 1586364061
transform 1 0 156676 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1703
timestamp 1586364061
transform 1 0 157780 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1715
timestamp 1586364061
transform 1 0 158884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1727
timestamp 1586364061
transform 1 0 159988 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_420
timestamp 1586364061
transform 1 0 161092 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1740
timestamp 1586364061
transform 1 0 161184 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1752
timestamp 1586364061
transform 1 0 162288 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1764
timestamp 1586364061
transform 1 0 163392 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1776
timestamp 1586364061
transform 1 0 164496 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_421
timestamp 1586364061
transform 1 0 166704 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1788
timestamp 1586364061
transform 1 0 165600 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1801
timestamp 1586364061
transform 1 0 166796 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1813
timestamp 1586364061
transform 1 0 167900 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1825
timestamp 1586364061
transform 1 0 169004 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1837
timestamp 1586364061
transform 1 0 170108 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1849
timestamp 1586364061
transform 1 0 171212 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_422
timestamp 1586364061
transform 1 0 172316 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1862
timestamp 1586364061
transform 1 0 172408 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1874
timestamp 1586364061
transform 1 0 173512 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1886
timestamp 1586364061
transform 1 0 174616 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1898
timestamp 1586364061
transform 1 0 175720 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_423
timestamp 1586364061
transform 1 0 177928 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1910
timestamp 1586364061
transform 1 0 176824 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1923
timestamp 1586364061
transform 1 0 178020 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1935
timestamp 1586364061
transform 1 0 179124 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1947
timestamp 1586364061
transform 1 0 180228 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1959
timestamp 1586364061
transform 1 0 181332 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1971
timestamp 1586364061
transform 1 0 182436 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_424
timestamp 1586364061
transform 1 0 183540 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_1984
timestamp 1586364061
transform 1 0 183632 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_1996
timestamp 1586364061
transform 1 0 184736 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2008
timestamp 1586364061
transform 1 0 185840 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2020
timestamp 1586364061
transform 1 0 186944 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2032
timestamp 1586364061
transform 1 0 188048 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_425
timestamp 1586364061
transform 1 0 189152 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_2045
timestamp 1586364061
transform 1 0 189244 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2057
timestamp 1586364061
transform 1 0 190348 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2069
timestamp 1586364061
transform 1 0 191452 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2081
timestamp 1586364061
transform 1 0 192556 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2093
timestamp 1586364061
transform 1 0 193660 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_426
timestamp 1586364061
transform 1 0 194764 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_2106
timestamp 1586364061
transform 1 0 194856 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2118
timestamp 1586364061
transform 1 0 195960 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2130
timestamp 1586364061
transform 1 0 197064 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2142
timestamp 1586364061
transform 1 0 198168 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2154
timestamp 1586364061
transform 1 0 199272 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_427
timestamp 1586364061
transform 1 0 200376 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_2167
timestamp 1586364061
transform 1 0 200468 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2179
timestamp 1586364061
transform 1 0 201572 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2191
timestamp 1586364061
transform 1 0 202676 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2203
timestamp 1586364061
transform 1 0 203780 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_428
timestamp 1586364061
transform 1 0 205988 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_2215
timestamp 1586364061
transform 1 0 204884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2228
timestamp 1586364061
transform 1 0 206080 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2240
timestamp 1586364061
transform 1 0 207184 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2252
timestamp 1586364061
transform 1 0 208288 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2264
timestamp 1586364061
transform 1 0 209392 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2276
timestamp 1586364061
transform 1 0 210496 0 -1 4896
box -38 -48 1142 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 212336 0 -1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_429
timestamp 1586364061
transform 1 0 211600 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_4_2289
timestamp 1586364061
transform 1 0 211692 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_2295
timestamp 1586364061
transform 1 0 212244 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_2304
timestamp 1586364061
transform 1 0 213072 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2316
timestamp 1586364061
transform 1 0 214176 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2328
timestamp 1586364061
transform 1 0 215280 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_430
timestamp 1586364061
transform 1 0 217212 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 217580 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_2340
timestamp 1586364061
transform 1 0 216384 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_2348
timestamp 1586364061
transform 1 0 217120 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_2350
timestamp 1586364061
transform 1 0 217304 0 -1 4896
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 218408 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 218224 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_2355
timestamp 1586364061
transform 1 0 217764 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_2359
timestamp 1586364061
transform 1 0 218132 0 -1 4896
box -38 -48 130 592
use scs8hd_nor4_4  _12_
timestamp 1586364061
transform 1 0 220524 0 -1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__10__C
timestamp 1586364061
transform 1 0 220340 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_2373
timestamp 1586364061
transform 1 0 219420 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_2381
timestamp 1586364061
transform 1 0 220156 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_2402
timestamp 1586364061
transform 1 0 222088 0 -1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_431
timestamp 1586364061
transform 1 0 222824 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__15__D
timestamp 1586364061
transform 1 0 223100 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_2411
timestamp 1586364061
transform 1 0 222916 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_2415
timestamp 1586364061
transform 1 0 223284 0 -1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__09__C
timestamp 1586364061
transform 1 0 225676 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_2427
timestamp 1586364061
transform 1 0 224388 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_4_2439
timestamp 1586364061
transform 1 0 225492 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_2443
timestamp 1586364061
transform 1 0 225860 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2455
timestamp 1586364061
transform 1 0 226964 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_432
timestamp 1586364061
transform 1 0 228436 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_2467
timestamp 1586364061
transform 1 0 228068 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_2472
timestamp 1586364061
transform 1 0 228528 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2484
timestamp 1586364061
transform 1 0 229632 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2496
timestamp 1586364061
transform 1 0 230736 0 -1 4896
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 232300 0 -1 4896
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_4_2508
timestamp 1586364061
transform 1 0 231840 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_2512
timestamp 1586364061
transform 1 0 232208 0 -1 4896
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_433
timestamp 1586364061
transform 1 0 234048 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_2524
timestamp 1586364061
transform 1 0 233312 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_12  FILLER_4_2533
timestamp 1586364061
transform 1 0 234140 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2545
timestamp 1586364061
transform 1 0 235244 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2557
timestamp 1586364061
transform 1 0 236348 0 -1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 238464 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_2569
timestamp 1586364061
transform 1 0 237452 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_4_2577
timestamp 1586364061
transform 1 0 238188 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_2582
timestamp 1586364061
transform 1 0 238648 0 -1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_434
timestamp 1586364061
transform 1 0 239660 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_2590
timestamp 1586364061
transform 1 0 239384 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_2594
timestamp 1586364061
transform 1 0 239752 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2606
timestamp 1586364061
transform 1 0 240856 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2618
timestamp 1586364061
transform 1 0 241960 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2630
timestamp 1586364061
transform 1 0 243064 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_435
timestamp 1586364061
transform 1 0 245272 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_2642
timestamp 1586364061
transform 1 0 244168 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2655
timestamp 1586364061
transform 1 0 245364 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2667
timestamp 1586364061
transform 1 0 246468 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2679
timestamp 1586364061
transform 1 0 247572 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2691
timestamp 1586364061
transform 1 0 248676 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2703
timestamp 1586364061
transform 1 0 249780 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_436
timestamp 1586364061
transform 1 0 250884 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_2716
timestamp 1586364061
transform 1 0 250976 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2728
timestamp 1586364061
transform 1 0 252080 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2740
timestamp 1586364061
transform 1 0 253184 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2752
timestamp 1586364061
transform 1 0 254288 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2764
timestamp 1586364061
transform 1 0 255392 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_437
timestamp 1586364061
transform 1 0 256496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_2777
timestamp 1586364061
transform 1 0 256588 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2789
timestamp 1586364061
transform 1 0 257692 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2801
timestamp 1586364061
transform 1 0 258796 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2813
timestamp 1586364061
transform 1 0 259900 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2825
timestamp 1586364061
transform 1 0 261004 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_438
timestamp 1586364061
transform 1 0 262108 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_2838
timestamp 1586364061
transform 1 0 262200 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2850
timestamp 1586364061
transform 1 0 263304 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2862
timestamp 1586364061
transform 1 0 264408 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2874
timestamp 1586364061
transform 1 0 265512 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2886
timestamp 1586364061
transform 1 0 266616 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_439
timestamp 1586364061
transform 1 0 267720 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_2899
timestamp 1586364061
transform 1 0 267812 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2911
timestamp 1586364061
transform 1 0 268916 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2923
timestamp 1586364061
transform 1 0 270020 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2935
timestamp 1586364061
transform 1 0 271124 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_440
timestamp 1586364061
transform 1 0 273332 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_2947
timestamp 1586364061
transform 1 0 272228 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2960
timestamp 1586364061
transform 1 0 273424 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2972
timestamp 1586364061
transform 1 0 274528 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2984
timestamp 1586364061
transform 1 0 275632 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_2996
timestamp 1586364061
transform 1 0 276736 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3008
timestamp 1586364061
transform 1 0 277840 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_441
timestamp 1586364061
transform 1 0 278944 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3021
timestamp 1586364061
transform 1 0 279036 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3033
timestamp 1586364061
transform 1 0 280140 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3045
timestamp 1586364061
transform 1 0 281244 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3057
timestamp 1586364061
transform 1 0 282348 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_442
timestamp 1586364061
transform 1 0 284556 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3069
timestamp 1586364061
transform 1 0 283452 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3082
timestamp 1586364061
transform 1 0 284648 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3094
timestamp 1586364061
transform 1 0 285752 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3106
timestamp 1586364061
transform 1 0 286856 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3118
timestamp 1586364061
transform 1 0 287960 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3130
timestamp 1586364061
transform 1 0 289064 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_443
timestamp 1586364061
transform 1 0 290168 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3143
timestamp 1586364061
transform 1 0 290260 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3155
timestamp 1586364061
transform 1 0 291364 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3167
timestamp 1586364061
transform 1 0 292468 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3179
timestamp 1586364061
transform 1 0 293572 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3191
timestamp 1586364061
transform 1 0 294676 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_444
timestamp 1586364061
transform 1 0 295780 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3204
timestamp 1586364061
transform 1 0 295872 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3216
timestamp 1586364061
transform 1 0 296976 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3228
timestamp 1586364061
transform 1 0 298080 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3240
timestamp 1586364061
transform 1 0 299184 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_445
timestamp 1586364061
transform 1 0 301392 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3252
timestamp 1586364061
transform 1 0 300288 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3265
timestamp 1586364061
transform 1 0 301484 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3277
timestamp 1586364061
transform 1 0 302588 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3289
timestamp 1586364061
transform 1 0 303692 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3301
timestamp 1586364061
transform 1 0 304796 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3313
timestamp 1586364061
transform 1 0 305900 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_446
timestamp 1586364061
transform 1 0 307004 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3326
timestamp 1586364061
transform 1 0 307096 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3338
timestamp 1586364061
transform 1 0 308200 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3350
timestamp 1586364061
transform 1 0 309304 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3362
timestamp 1586364061
transform 1 0 310408 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_447
timestamp 1586364061
transform 1 0 312616 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3374
timestamp 1586364061
transform 1 0 311512 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3387
timestamp 1586364061
transform 1 0 312708 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3399
timestamp 1586364061
transform 1 0 313812 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3411
timestamp 1586364061
transform 1 0 314916 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3423
timestamp 1586364061
transform 1 0 316020 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3435
timestamp 1586364061
transform 1 0 317124 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_448
timestamp 1586364061
transform 1 0 318228 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3448
timestamp 1586364061
transform 1 0 318320 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3460
timestamp 1586364061
transform 1 0 319424 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3472
timestamp 1586364061
transform 1 0 320528 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3484
timestamp 1586364061
transform 1 0 321632 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3496
timestamp 1586364061
transform 1 0 322736 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_449
timestamp 1586364061
transform 1 0 323840 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3509
timestamp 1586364061
transform 1 0 323932 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3521
timestamp 1586364061
transform 1 0 325036 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3533
timestamp 1586364061
transform 1 0 326140 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3545
timestamp 1586364061
transform 1 0 327244 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3557
timestamp 1586364061
transform 1 0 328348 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_450
timestamp 1586364061
transform 1 0 329452 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3570
timestamp 1586364061
transform 1 0 329544 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3582
timestamp 1586364061
transform 1 0 330648 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3594
timestamp 1586364061
transform 1 0 331752 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3606
timestamp 1586364061
transform 1 0 332856 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3618
timestamp 1586364061
transform 1 0 333960 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_451
timestamp 1586364061
transform 1 0 335064 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3631
timestamp 1586364061
transform 1 0 335156 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3643
timestamp 1586364061
transform 1 0 336260 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3655
timestamp 1586364061
transform 1 0 337364 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3667
timestamp 1586364061
transform 1 0 338468 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_452
timestamp 1586364061
transform 1 0 340676 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3679
timestamp 1586364061
transform 1 0 339572 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3692
timestamp 1586364061
transform 1 0 340768 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3704
timestamp 1586364061
transform 1 0 341872 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3716
timestamp 1586364061
transform 1 0 342976 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3728
timestamp 1586364061
transform 1 0 344080 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3740
timestamp 1586364061
transform 1 0 345184 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_453
timestamp 1586364061
transform 1 0 346288 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3753
timestamp 1586364061
transform 1 0 346380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3765
timestamp 1586364061
transform 1 0 347484 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3777
timestamp 1586364061
transform 1 0 348588 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3789
timestamp 1586364061
transform 1 0 349692 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_454
timestamp 1586364061
transform 1 0 351900 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3801
timestamp 1586364061
transform 1 0 350796 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3814
timestamp 1586364061
transform 1 0 351992 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3826
timestamp 1586364061
transform 1 0 353096 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3838
timestamp 1586364061
transform 1 0 354200 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3850
timestamp 1586364061
transform 1 0 355304 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3862
timestamp 1586364061
transform 1 0 356408 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_455
timestamp 1586364061
transform 1 0 357512 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3875
timestamp 1586364061
transform 1 0 357604 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3887
timestamp 1586364061
transform 1 0 358708 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3899
timestamp 1586364061
transform 1 0 359812 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3911
timestamp 1586364061
transform 1 0 360916 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3923
timestamp 1586364061
transform 1 0 362020 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_456
timestamp 1586364061
transform 1 0 363124 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3936
timestamp 1586364061
transform 1 0 363216 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3948
timestamp 1586364061
transform 1 0 364320 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3960
timestamp 1586364061
transform 1 0 365424 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3972
timestamp 1586364061
transform 1 0 366528 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_3984
timestamp 1586364061
transform 1 0 367632 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_457
timestamp 1586364061
transform 1 0 368736 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_3997
timestamp 1586364061
transform 1 0 368828 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4009
timestamp 1586364061
transform 1 0 369932 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4021
timestamp 1586364061
transform 1 0 371036 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4033
timestamp 1586364061
transform 1 0 372140 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4045
timestamp 1586364061
transform 1 0 373244 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_458
timestamp 1586364061
transform 1 0 374348 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_4058
timestamp 1586364061
transform 1 0 374440 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4070
timestamp 1586364061
transform 1 0 375544 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4082
timestamp 1586364061
transform 1 0 376648 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4094
timestamp 1586364061
transform 1 0 377752 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_459
timestamp 1586364061
transform 1 0 379960 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_4106
timestamp 1586364061
transform 1 0 378856 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4119
timestamp 1586364061
transform 1 0 380052 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4131
timestamp 1586364061
transform 1 0 381156 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4143
timestamp 1586364061
transform 1 0 382260 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4155
timestamp 1586364061
transform 1 0 383364 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4167
timestamp 1586364061
transform 1 0 384468 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_460
timestamp 1586364061
transform 1 0 385572 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_4180
timestamp 1586364061
transform 1 0 385664 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4192
timestamp 1586364061
transform 1 0 386768 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4204
timestamp 1586364061
transform 1 0 387872 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4216
timestamp 1586364061
transform 1 0 388976 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_461
timestamp 1586364061
transform 1 0 391184 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_4228
timestamp 1586364061
transform 1 0 390080 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4241
timestamp 1586364061
transform 1 0 391276 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4253
timestamp 1586364061
transform 1 0 392380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4265
timestamp 1586364061
transform 1 0 393484 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4277
timestamp 1586364061
transform 1 0 394588 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4289
timestamp 1586364061
transform 1 0 395692 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_462
timestamp 1586364061
transform 1 0 396796 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_4302
timestamp 1586364061
transform 1 0 396888 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4314
timestamp 1586364061
transform 1 0 397992 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4326
timestamp 1586364061
transform 1 0 399096 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4338
timestamp 1586364061
transform 1 0 400200 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4350
timestamp 1586364061
transform 1 0 401304 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_463
timestamp 1586364061
transform 1 0 402408 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_4363
timestamp 1586364061
transform 1 0 402500 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4375
timestamp 1586364061
transform 1 0 403604 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4387
timestamp 1586364061
transform 1 0 404708 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4399
timestamp 1586364061
transform 1 0 405812 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_464
timestamp 1586364061
transform 1 0 408020 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_4411
timestamp 1586364061
transform 1 0 406916 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4424
timestamp 1586364061
transform 1 0 408112 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4436
timestamp 1586364061
transform 1 0 409216 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4448
timestamp 1586364061
transform 1 0 410320 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4460
timestamp 1586364061
transform 1 0 411424 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4472
timestamp 1586364061
transform 1 0 412528 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_465
timestamp 1586364061
transform 1 0 413632 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_4485
timestamp 1586364061
transform 1 0 413724 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4497
timestamp 1586364061
transform 1 0 414828 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4509
timestamp 1586364061
transform 1 0 415932 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4521
timestamp 1586364061
transform 1 0 417036 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_466
timestamp 1586364061
transform 1 0 419244 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_4533
timestamp 1586364061
transform 1 0 418140 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4546
timestamp 1586364061
transform 1 0 419336 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_4558
timestamp 1586364061
transform 1 0 420440 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 422832 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_4570
timestamp 1586364061
transform 1 0 421544 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_4_4578
timestamp 1586364061
transform 1 0 422280 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_467
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_468
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_171
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_469
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_470
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_281
timestamp 1586364061
transform 1 0 26956 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_293
timestamp 1586364061
transform 1 0 28060 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_471
timestamp 1586364061
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_306
timestamp 1586364061
transform 1 0 29256 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_318
timestamp 1586364061
transform 1 0 30360 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_330
timestamp 1586364061
transform 1 0 31464 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_342
timestamp 1586364061
transform 1 0 32568 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_354
timestamp 1586364061
transform 1 0 33672 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_472
timestamp 1586364061
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_367
timestamp 1586364061
transform 1 0 34868 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_379
timestamp 1586364061
transform 1 0 35972 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_391
timestamp 1586364061
transform 1 0 37076 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_403
timestamp 1586364061
transform 1 0 38180 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_473
timestamp 1586364061
transform 1 0 40388 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_415
timestamp 1586364061
transform 1 0 39284 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_428
timestamp 1586364061
transform 1 0 40480 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_440
timestamp 1586364061
transform 1 0 41584 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_452
timestamp 1586364061
transform 1 0 42688 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_464
timestamp 1586364061
transform 1 0 43792 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_476
timestamp 1586364061
transform 1 0 44896 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_474
timestamp 1586364061
transform 1 0 46000 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_489
timestamp 1586364061
transform 1 0 46092 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_501
timestamp 1586364061
transform 1 0 47196 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_513
timestamp 1586364061
transform 1 0 48300 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_525
timestamp 1586364061
transform 1 0 49404 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_475
timestamp 1586364061
transform 1 0 51612 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_537
timestamp 1586364061
transform 1 0 50508 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_550
timestamp 1586364061
transform 1 0 51704 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_562
timestamp 1586364061
transform 1 0 52808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_574
timestamp 1586364061
transform 1 0 53912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_586
timestamp 1586364061
transform 1 0 55016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_598
timestamp 1586364061
transform 1 0 56120 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_476
timestamp 1586364061
transform 1 0 57224 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_611
timestamp 1586364061
transform 1 0 57316 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_623
timestamp 1586364061
transform 1 0 58420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_635
timestamp 1586364061
transform 1 0 59524 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_647
timestamp 1586364061
transform 1 0 60628 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_659
timestamp 1586364061
transform 1 0 61732 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_477
timestamp 1586364061
transform 1 0 62836 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_672
timestamp 1586364061
transform 1 0 62928 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_684
timestamp 1586364061
transform 1 0 64032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_696
timestamp 1586364061
transform 1 0 65136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_708
timestamp 1586364061
transform 1 0 66240 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_720
timestamp 1586364061
transform 1 0 67344 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_478
timestamp 1586364061
transform 1 0 68448 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_733
timestamp 1586364061
transform 1 0 68540 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_745
timestamp 1586364061
transform 1 0 69644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_757
timestamp 1586364061
transform 1 0 70748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_769
timestamp 1586364061
transform 1 0 71852 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_781
timestamp 1586364061
transform 1 0 72956 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_479
timestamp 1586364061
transform 1 0 74060 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_794
timestamp 1586364061
transform 1 0 74152 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_806
timestamp 1586364061
transform 1 0 75256 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_818
timestamp 1586364061
transform 1 0 76360 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_830
timestamp 1586364061
transform 1 0 77464 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_480
timestamp 1586364061
transform 1 0 79672 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_842
timestamp 1586364061
transform 1 0 78568 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_855
timestamp 1586364061
transform 1 0 79764 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_867
timestamp 1586364061
transform 1 0 80868 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_879
timestamp 1586364061
transform 1 0 81972 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_891
timestamp 1586364061
transform 1 0 83076 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_903
timestamp 1586364061
transform 1 0 84180 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_481
timestamp 1586364061
transform 1 0 85284 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_916
timestamp 1586364061
transform 1 0 85376 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_928
timestamp 1586364061
transform 1 0 86480 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_940
timestamp 1586364061
transform 1 0 87584 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_952
timestamp 1586364061
transform 1 0 88688 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_482
timestamp 1586364061
transform 1 0 90896 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_964
timestamp 1586364061
transform 1 0 89792 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_977
timestamp 1586364061
transform 1 0 90988 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_989
timestamp 1586364061
transform 1 0 92092 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1001
timestamp 1586364061
transform 1 0 93196 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1013
timestamp 1586364061
transform 1 0 94300 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1025
timestamp 1586364061
transform 1 0 95404 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_483
timestamp 1586364061
transform 1 0 96508 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1038
timestamp 1586364061
transform 1 0 96600 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1050
timestamp 1586364061
transform 1 0 97704 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1062
timestamp 1586364061
transform 1 0 98808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1074
timestamp 1586364061
transform 1 0 99912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1086
timestamp 1586364061
transform 1 0 101016 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_484
timestamp 1586364061
transform 1 0 102120 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1099
timestamp 1586364061
transform 1 0 102212 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1111
timestamp 1586364061
transform 1 0 103316 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1123
timestamp 1586364061
transform 1 0 104420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1135
timestamp 1586364061
transform 1 0 105524 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_485
timestamp 1586364061
transform 1 0 107732 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1147
timestamp 1586364061
transform 1 0 106628 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1160
timestamp 1586364061
transform 1 0 107824 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1172
timestamp 1586364061
transform 1 0 108928 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1184
timestamp 1586364061
transform 1 0 110032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1196
timestamp 1586364061
transform 1 0 111136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1208
timestamp 1586364061
transform 1 0 112240 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_486
timestamp 1586364061
transform 1 0 113344 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1221
timestamp 1586364061
transform 1 0 113436 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1233
timestamp 1586364061
transform 1 0 114540 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1245
timestamp 1586364061
transform 1 0 115644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1257
timestamp 1586364061
transform 1 0 116748 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_487
timestamp 1586364061
transform 1 0 118956 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1269
timestamp 1586364061
transform 1 0 117852 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1282
timestamp 1586364061
transform 1 0 119048 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1294
timestamp 1586364061
transform 1 0 120152 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1306
timestamp 1586364061
transform 1 0 121256 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1318
timestamp 1586364061
transform 1 0 122360 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1330
timestamp 1586364061
transform 1 0 123464 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_488
timestamp 1586364061
transform 1 0 124568 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1343
timestamp 1586364061
transform 1 0 124660 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1355
timestamp 1586364061
transform 1 0 125764 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1367
timestamp 1586364061
transform 1 0 126868 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1379
timestamp 1586364061
transform 1 0 127972 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1391
timestamp 1586364061
transform 1 0 129076 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_489
timestamp 1586364061
transform 1 0 130180 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1404
timestamp 1586364061
transform 1 0 130272 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1416
timestamp 1586364061
transform 1 0 131376 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1428
timestamp 1586364061
transform 1 0 132480 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1440
timestamp 1586364061
transform 1 0 133584 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1452
timestamp 1586364061
transform 1 0 134688 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_490
timestamp 1586364061
transform 1 0 135792 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1465
timestamp 1586364061
transform 1 0 135884 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1477
timestamp 1586364061
transform 1 0 136988 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1489
timestamp 1586364061
transform 1 0 138092 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1501
timestamp 1586364061
transform 1 0 139196 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1513
timestamp 1586364061
transform 1 0 140300 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_491
timestamp 1586364061
transform 1 0 141404 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1526
timestamp 1586364061
transform 1 0 141496 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1538
timestamp 1586364061
transform 1 0 142600 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1550
timestamp 1586364061
transform 1 0 143704 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1562
timestamp 1586364061
transform 1 0 144808 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_492
timestamp 1586364061
transform 1 0 147016 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1574
timestamp 1586364061
transform 1 0 145912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1587
timestamp 1586364061
transform 1 0 147108 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1599
timestamp 1586364061
transform 1 0 148212 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1611
timestamp 1586364061
transform 1 0 149316 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1623
timestamp 1586364061
transform 1 0 150420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1635
timestamp 1586364061
transform 1 0 151524 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_493
timestamp 1586364061
transform 1 0 152628 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1648
timestamp 1586364061
transform 1 0 152720 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1660
timestamp 1586364061
transform 1 0 153824 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1672
timestamp 1586364061
transform 1 0 154928 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1684
timestamp 1586364061
transform 1 0 156032 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_494
timestamp 1586364061
transform 1 0 158240 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1696
timestamp 1586364061
transform 1 0 157136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1709
timestamp 1586364061
transform 1 0 158332 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1721
timestamp 1586364061
transform 1 0 159436 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1733
timestamp 1586364061
transform 1 0 160540 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1745
timestamp 1586364061
transform 1 0 161644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1757
timestamp 1586364061
transform 1 0 162748 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_495
timestamp 1586364061
transform 1 0 163852 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1770
timestamp 1586364061
transform 1 0 163944 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1782
timestamp 1586364061
transform 1 0 165048 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1794
timestamp 1586364061
transform 1 0 166152 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1806
timestamp 1586364061
transform 1 0 167256 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1818
timestamp 1586364061
transform 1 0 168360 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_496
timestamp 1586364061
transform 1 0 169464 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1831
timestamp 1586364061
transform 1 0 169556 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1843
timestamp 1586364061
transform 1 0 170660 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1855
timestamp 1586364061
transform 1 0 171764 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1867
timestamp 1586364061
transform 1 0 172868 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1879
timestamp 1586364061
transform 1 0 173972 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_497
timestamp 1586364061
transform 1 0 175076 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1892
timestamp 1586364061
transform 1 0 175168 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1904
timestamp 1586364061
transform 1 0 176272 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1916
timestamp 1586364061
transform 1 0 177376 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1928
timestamp 1586364061
transform 1 0 178480 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1940
timestamp 1586364061
transform 1 0 179584 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_498
timestamp 1586364061
transform 1 0 180688 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_1953
timestamp 1586364061
transform 1 0 180780 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1965
timestamp 1586364061
transform 1 0 181884 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1977
timestamp 1586364061
transform 1 0 182988 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_1989
timestamp 1586364061
transform 1 0 184092 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_499
timestamp 1586364061
transform 1 0 186300 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_2001
timestamp 1586364061
transform 1 0 185196 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2014
timestamp 1586364061
transform 1 0 186392 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2026
timestamp 1586364061
transform 1 0 187496 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2038
timestamp 1586364061
transform 1 0 188600 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2050
timestamp 1586364061
transform 1 0 189704 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2062
timestamp 1586364061
transform 1 0 190808 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_500
timestamp 1586364061
transform 1 0 191912 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_2075
timestamp 1586364061
transform 1 0 192004 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2087
timestamp 1586364061
transform 1 0 193108 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2099
timestamp 1586364061
transform 1 0 194212 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2111
timestamp 1586364061
transform 1 0 195316 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_501
timestamp 1586364061
transform 1 0 197524 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_2123
timestamp 1586364061
transform 1 0 196420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2136
timestamp 1586364061
transform 1 0 197616 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2148
timestamp 1586364061
transform 1 0 198720 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2160
timestamp 1586364061
transform 1 0 199824 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2172
timestamp 1586364061
transform 1 0 200928 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2184
timestamp 1586364061
transform 1 0 202032 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_502
timestamp 1586364061
transform 1 0 203136 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_2197
timestamp 1586364061
transform 1 0 203228 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2209
timestamp 1586364061
transform 1 0 204332 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2221
timestamp 1586364061
transform 1 0 205436 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2233
timestamp 1586364061
transform 1 0 206540 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2245
timestamp 1586364061
transform 1 0 207644 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_503
timestamp 1586364061
transform 1 0 208748 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__21__A
timestamp 1586364061
transform 1 0 209300 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_2258
timestamp 1586364061
transform 1 0 208840 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_2262
timestamp 1586364061
transform 1 0 209208 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_2265
timestamp 1586364061
transform 1 0 209484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2277
timestamp 1586364061
transform 1 0 210588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2289
timestamp 1586364061
transform 1 0 211692 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_504
timestamp 1586364061
transform 1 0 214360 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_2301
timestamp 1586364061
transform 1 0 212796 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_5_2313
timestamp 1586364061
transform 1 0 213900 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_2317
timestamp 1586364061
transform 1 0 214268 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 215280 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 215648 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_2319
timestamp 1586364061
transform 1 0 214452 0 1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_5_2327
timestamp 1586364061
transform 1 0 215188 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_2330
timestamp 1586364061
transform 1 0 215464 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_2334
timestamp 1586364061
transform 1 0 215832 0 1 4896
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 217580 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 217396 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_2346
timestamp 1586364061
transform 1 0 216936 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_2350
timestamp 1586364061
transform 1 0 217304 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 219328 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_2364
timestamp 1586364061
transform 1 0 218592 0 1 4896
box -38 -48 774 592
use scs8hd_and4_4  _10_
timestamp 1586364061
transform 1 0 220340 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_505
timestamp 1586364061
transform 1 0 219972 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 219696 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_2374
timestamp 1586364061
transform 1 0 219512 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_2378
timestamp 1586364061
transform 1 0 219880 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_5_2380
timestamp 1586364061
transform 1 0 220064 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__10__B
timestamp 1586364061
transform 1 0 221352 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__10__D
timestamp 1586364061
transform 1 0 221720 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_2392
timestamp 1586364061
transform 1 0 221168 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_2396
timestamp 1586364061
transform 1 0 221536 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_2400
timestamp 1586364061
transform 1 0 221904 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2412
timestamp 1586364061
transform 1 0 223008 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2424
timestamp 1586364061
transform 1 0 224112 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_506
timestamp 1586364061
transform 1 0 225584 0 1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_5_2436
timestamp 1586364061
transform 1 0 225216 0 1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_5_2441
timestamp 1586364061
transform 1 0 225676 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2453
timestamp 1586364061
transform 1 0 226780 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2465
timestamp 1586364061
transform 1 0 227884 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2477
timestamp 1586364061
transform 1 0 228988 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2489
timestamp 1586364061
transform 1 0 230092 0 1 4896
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 232392 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_507
timestamp 1586364061
transform 1 0 231196 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 232208 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_2502
timestamp 1586364061
transform 1 0 231288 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_2510
timestamp 1586364061
transform 1 0 232024 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_2525
timestamp 1586364061
transform 1 0 233404 0 1 4896
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 234140 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 234508 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_2535
timestamp 1586364061
transform 1 0 234324 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_2539
timestamp 1586364061
transform 1 0 234692 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_508
timestamp 1586364061
transform 1 0 236808 0 1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_5_2551
timestamp 1586364061
transform 1 0 235796 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_5_2559
timestamp 1586364061
transform 1 0 236532 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_2563
timestamp 1586364061
transform 1 0 236900 0 1 4896
box -38 -48 1142 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 238464 0 1 4896
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 238280 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_2575
timestamp 1586364061
transform 1 0 238004 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_2588
timestamp 1586364061
transform 1 0 239200 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2600
timestamp 1586364061
transform 1 0 240304 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_2612
timestamp 1586364061
transform 1 0 241408 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_5_2620
timestamp 1586364061
transform 1 0 242144 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_509
timestamp 1586364061
transform 1 0 242420 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_2624
timestamp 1586364061
transform 1 0 242512 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2636
timestamp 1586364061
transform 1 0 243616 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2648
timestamp 1586364061
transform 1 0 244720 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2660
timestamp 1586364061
transform 1 0 245824 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2672
timestamp 1586364061
transform 1 0 246928 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_510
timestamp 1586364061
transform 1 0 248032 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_2685
timestamp 1586364061
transform 1 0 248124 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2697
timestamp 1586364061
transform 1 0 249228 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2709
timestamp 1586364061
transform 1 0 250332 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2721
timestamp 1586364061
transform 1 0 251436 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_511
timestamp 1586364061
transform 1 0 253644 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_2733
timestamp 1586364061
transform 1 0 252540 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2746
timestamp 1586364061
transform 1 0 253736 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2758
timestamp 1586364061
transform 1 0 254840 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2770
timestamp 1586364061
transform 1 0 255944 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2782
timestamp 1586364061
transform 1 0 257048 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2794
timestamp 1586364061
transform 1 0 258152 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_512
timestamp 1586364061
transform 1 0 259256 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_2807
timestamp 1586364061
transform 1 0 259348 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2819
timestamp 1586364061
transform 1 0 260452 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2831
timestamp 1586364061
transform 1 0 261556 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2843
timestamp 1586364061
transform 1 0 262660 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_513
timestamp 1586364061
transform 1 0 264868 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_2855
timestamp 1586364061
transform 1 0 263764 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2868
timestamp 1586364061
transform 1 0 264960 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2880
timestamp 1586364061
transform 1 0 266064 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2892
timestamp 1586364061
transform 1 0 267168 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2904
timestamp 1586364061
transform 1 0 268272 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2916
timestamp 1586364061
transform 1 0 269376 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_514
timestamp 1586364061
transform 1 0 270480 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_2929
timestamp 1586364061
transform 1 0 270572 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2941
timestamp 1586364061
transform 1 0 271676 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2953
timestamp 1586364061
transform 1 0 272780 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2965
timestamp 1586364061
transform 1 0 273884 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_2977
timestamp 1586364061
transform 1 0 274988 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_515
timestamp 1586364061
transform 1 0 276092 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_2990
timestamp 1586364061
transform 1 0 276184 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3002
timestamp 1586364061
transform 1 0 277288 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3014
timestamp 1586364061
transform 1 0 278392 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3026
timestamp 1586364061
transform 1 0 279496 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_516
timestamp 1586364061
transform 1 0 281704 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3038
timestamp 1586364061
transform 1 0 280600 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3051
timestamp 1586364061
transform 1 0 281796 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3063
timestamp 1586364061
transform 1 0 282900 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3075
timestamp 1586364061
transform 1 0 284004 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3087
timestamp 1586364061
transform 1 0 285108 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3099
timestamp 1586364061
transform 1 0 286212 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_517
timestamp 1586364061
transform 1 0 287316 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3112
timestamp 1586364061
transform 1 0 287408 0 1 4896
box -38 -48 1142 592
use scs8hd_buf_2  _20_
timestamp 1586364061
transform 1 0 289432 0 1 4896
box -38 -48 406 592
use scs8hd_decap_8  FILLER_5_3124
timestamp 1586364061
transform 1 0 288512 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_3132
timestamp 1586364061
transform 1 0 289248 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_3138
timestamp 1586364061
transform 1 0 289800 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__20__A
timestamp 1586364061
transform 1 0 289984 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_3142
timestamp 1586364061
transform 1 0 290168 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3154
timestamp 1586364061
transform 1 0 291272 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_518
timestamp 1586364061
transform 1 0 292928 0 1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_5_3166
timestamp 1586364061
transform 1 0 292376 0 1 4896
box -38 -48 590 592
use scs8hd_decap_12  FILLER_5_3173
timestamp 1586364061
transform 1 0 293020 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3185
timestamp 1586364061
transform 1 0 294124 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3197
timestamp 1586364061
transform 1 0 295228 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3209
timestamp 1586364061
transform 1 0 296332 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3221
timestamp 1586364061
transform 1 0 297436 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_519
timestamp 1586364061
transform 1 0 298540 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3234
timestamp 1586364061
transform 1 0 298632 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3246
timestamp 1586364061
transform 1 0 299736 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3258
timestamp 1586364061
transform 1 0 300840 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3270
timestamp 1586364061
transform 1 0 301944 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_520
timestamp 1586364061
transform 1 0 304152 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3282
timestamp 1586364061
transform 1 0 303048 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3295
timestamp 1586364061
transform 1 0 304244 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3307
timestamp 1586364061
transform 1 0 305348 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3319
timestamp 1586364061
transform 1 0 306452 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3331
timestamp 1586364061
transform 1 0 307556 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3343
timestamp 1586364061
transform 1 0 308660 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_521
timestamp 1586364061
transform 1 0 309764 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3356
timestamp 1586364061
transform 1 0 309856 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3368
timestamp 1586364061
transform 1 0 310960 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3380
timestamp 1586364061
transform 1 0 312064 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3392
timestamp 1586364061
transform 1 0 313168 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3404
timestamp 1586364061
transform 1 0 314272 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_522
timestamp 1586364061
transform 1 0 315376 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3417
timestamp 1586364061
transform 1 0 315468 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3429
timestamp 1586364061
transform 1 0 316572 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3441
timestamp 1586364061
transform 1 0 317676 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3453
timestamp 1586364061
transform 1 0 318780 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_523
timestamp 1586364061
transform 1 0 320988 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3465
timestamp 1586364061
transform 1 0 319884 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3478
timestamp 1586364061
transform 1 0 321080 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3490
timestamp 1586364061
transform 1 0 322184 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3502
timestamp 1586364061
transform 1 0 323288 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3514
timestamp 1586364061
transform 1 0 324392 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3526
timestamp 1586364061
transform 1 0 325496 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_524
timestamp 1586364061
transform 1 0 326600 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3539
timestamp 1586364061
transform 1 0 326692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3551
timestamp 1586364061
transform 1 0 327796 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3563
timestamp 1586364061
transform 1 0 328900 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3575
timestamp 1586364061
transform 1 0 330004 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_525
timestamp 1586364061
transform 1 0 332212 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3587
timestamp 1586364061
transform 1 0 331108 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3600
timestamp 1586364061
transform 1 0 332304 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3612
timestamp 1586364061
transform 1 0 333408 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3624
timestamp 1586364061
transform 1 0 334512 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3636
timestamp 1586364061
transform 1 0 335616 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3648
timestamp 1586364061
transform 1 0 336720 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_526
timestamp 1586364061
transform 1 0 337824 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3661
timestamp 1586364061
transform 1 0 337916 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3673
timestamp 1586364061
transform 1 0 339020 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3685
timestamp 1586364061
transform 1 0 340124 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3697
timestamp 1586364061
transform 1 0 341228 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3709
timestamp 1586364061
transform 1 0 342332 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_527
timestamp 1586364061
transform 1 0 343436 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3722
timestamp 1586364061
transform 1 0 343528 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3734
timestamp 1586364061
transform 1 0 344632 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3746
timestamp 1586364061
transform 1 0 345736 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3758
timestamp 1586364061
transform 1 0 346840 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3770
timestamp 1586364061
transform 1 0 347944 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_528
timestamp 1586364061
transform 1 0 349048 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3783
timestamp 1586364061
transform 1 0 349140 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3795
timestamp 1586364061
transform 1 0 350244 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3807
timestamp 1586364061
transform 1 0 351348 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3819
timestamp 1586364061
transform 1 0 352452 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3831
timestamp 1586364061
transform 1 0 353556 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_529
timestamp 1586364061
transform 1 0 354660 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3844
timestamp 1586364061
transform 1 0 354752 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3856
timestamp 1586364061
transform 1 0 355856 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3868
timestamp 1586364061
transform 1 0 356960 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3880
timestamp 1586364061
transform 1 0 358064 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_530
timestamp 1586364061
transform 1 0 360272 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3892
timestamp 1586364061
transform 1 0 359168 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3905
timestamp 1586364061
transform 1 0 360364 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3917
timestamp 1586364061
transform 1 0 361468 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3929
timestamp 1586364061
transform 1 0 362572 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3941
timestamp 1586364061
transform 1 0 363676 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3953
timestamp 1586364061
transform 1 0 364780 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_531
timestamp 1586364061
transform 1 0 365884 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_3966
timestamp 1586364061
transform 1 0 365976 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3978
timestamp 1586364061
transform 1 0 367080 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_3990
timestamp 1586364061
transform 1 0 368184 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4002
timestamp 1586364061
transform 1 0 369288 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_532
timestamp 1586364061
transform 1 0 371496 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_4014
timestamp 1586364061
transform 1 0 370392 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4027
timestamp 1586364061
transform 1 0 371588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4039
timestamp 1586364061
transform 1 0 372692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4051
timestamp 1586364061
transform 1 0 373796 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4063
timestamp 1586364061
transform 1 0 374900 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4075
timestamp 1586364061
transform 1 0 376004 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_533
timestamp 1586364061
transform 1 0 377108 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_4088
timestamp 1586364061
transform 1 0 377200 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4100
timestamp 1586364061
transform 1 0 378304 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4112
timestamp 1586364061
transform 1 0 379408 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4124
timestamp 1586364061
transform 1 0 380512 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4136
timestamp 1586364061
transform 1 0 381616 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_534
timestamp 1586364061
transform 1 0 382720 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_4149
timestamp 1586364061
transform 1 0 382812 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4161
timestamp 1586364061
transform 1 0 383916 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4173
timestamp 1586364061
transform 1 0 385020 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4185
timestamp 1586364061
transform 1 0 386124 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_535
timestamp 1586364061
transform 1 0 388332 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_4197
timestamp 1586364061
transform 1 0 387228 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4210
timestamp 1586364061
transform 1 0 388424 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4222
timestamp 1586364061
transform 1 0 389528 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4234
timestamp 1586364061
transform 1 0 390632 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4246
timestamp 1586364061
transform 1 0 391736 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4258
timestamp 1586364061
transform 1 0 392840 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_536
timestamp 1586364061
transform 1 0 393944 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_4271
timestamp 1586364061
transform 1 0 394036 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4283
timestamp 1586364061
transform 1 0 395140 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4295
timestamp 1586364061
transform 1 0 396244 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4307
timestamp 1586364061
transform 1 0 397348 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_537
timestamp 1586364061
transform 1 0 399556 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_4319
timestamp 1586364061
transform 1 0 398452 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4332
timestamp 1586364061
transform 1 0 399648 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4344
timestamp 1586364061
transform 1 0 400752 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4356
timestamp 1586364061
transform 1 0 401856 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4368
timestamp 1586364061
transform 1 0 402960 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4380
timestamp 1586364061
transform 1 0 404064 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_538
timestamp 1586364061
transform 1 0 405168 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_4393
timestamp 1586364061
transform 1 0 405260 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4405
timestamp 1586364061
transform 1 0 406364 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4417
timestamp 1586364061
transform 1 0 407468 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4429
timestamp 1586364061
transform 1 0 408572 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4441
timestamp 1586364061
transform 1 0 409676 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_539
timestamp 1586364061
transform 1 0 410780 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_4454
timestamp 1586364061
transform 1 0 410872 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4466
timestamp 1586364061
transform 1 0 411976 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4478
timestamp 1586364061
transform 1 0 413080 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4490
timestamp 1586364061
transform 1 0 414184 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4502
timestamp 1586364061
transform 1 0 415288 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_540
timestamp 1586364061
transform 1 0 416392 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_4515
timestamp 1586364061
transform 1 0 416484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4527
timestamp 1586364061
transform 1 0 417588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4539
timestamp 1586364061
transform 1 0 418692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4551
timestamp 1586364061
transform 1 0 419796 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_4563
timestamp 1586364061
transform 1 0 420900 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 422832 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_541
timestamp 1586364061
transform 1 0 422004 0 1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_5_4576
timestamp 1586364061
transform 1 0 422096 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_4580
timestamp 1586364061
transform 1 0 422464 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_542
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_617
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_543
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_618
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_544
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_159
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_171
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_619
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_545
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_220
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_620
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_232
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_263
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_546
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_281
timestamp 1586364061
transform 1 0 26956 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_288
timestamp 1586364061
transform 1 0 27600 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_300
timestamp 1586364061
transform 1 0 28704 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_293
timestamp 1586364061
transform 1 0 28060 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_621
timestamp 1586364061
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_312
timestamp 1586364061
transform 1 0 29808 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_306
timestamp 1586364061
transform 1 0 29256 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_318
timestamp 1586364061
transform 1 0 30360 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_547
timestamp 1586364061
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_324
timestamp 1586364061
transform 1 0 30912 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_337
timestamp 1586364061
transform 1 0 32108 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_330
timestamp 1586364061
transform 1 0 31464 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_349
timestamp 1586364061
transform 1 0 33212 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_342
timestamp 1586364061
transform 1 0 32568 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_354
timestamp 1586364061
transform 1 0 33672 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_622
timestamp 1586364061
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_361
timestamp 1586364061
transform 1 0 34316 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_373
timestamp 1586364061
transform 1 0 35420 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_367
timestamp 1586364061
transform 1 0 34868 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_385
timestamp 1586364061
transform 1 0 36524 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_379
timestamp 1586364061
transform 1 0 35972 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_391
timestamp 1586364061
transform 1 0 37076 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_548
timestamp 1586364061
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_398
timestamp 1586364061
transform 1 0 37720 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_410
timestamp 1586364061
transform 1 0 38824 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_403
timestamp 1586364061
transform 1 0 38180 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_623
timestamp 1586364061
transform 1 0 40388 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_422
timestamp 1586364061
transform 1 0 39928 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_415
timestamp 1586364061
transform 1 0 39284 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_428
timestamp 1586364061
transform 1 0 40480 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_434
timestamp 1586364061
transform 1 0 41032 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_440
timestamp 1586364061
transform 1 0 41584 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_549
timestamp 1586364061
transform 1 0 43240 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_446
timestamp 1586364061
transform 1 0 42136 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_459
timestamp 1586364061
transform 1 0 43332 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_452
timestamp 1586364061
transform 1 0 42688 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_471
timestamp 1586364061
transform 1 0 44436 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_464
timestamp 1586364061
transform 1 0 43792 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_476
timestamp 1586364061
transform 1 0 44896 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_624
timestamp 1586364061
transform 1 0 46000 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_483
timestamp 1586364061
transform 1 0 45540 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_495
timestamp 1586364061
transform 1 0 46644 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_489
timestamp 1586364061
transform 1 0 46092 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_507
timestamp 1586364061
transform 1 0 47748 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_501
timestamp 1586364061
transform 1 0 47196 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_513
timestamp 1586364061
transform 1 0 48300 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_550
timestamp 1586364061
transform 1 0 48852 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_520
timestamp 1586364061
transform 1 0 48944 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_532
timestamp 1586364061
transform 1 0 50048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_525
timestamp 1586364061
transform 1 0 49404 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_625
timestamp 1586364061
transform 1 0 51612 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_544
timestamp 1586364061
transform 1 0 51152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_537
timestamp 1586364061
transform 1 0 50508 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_550
timestamp 1586364061
transform 1 0 51704 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_556
timestamp 1586364061
transform 1 0 52256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_568
timestamp 1586364061
transform 1 0 53360 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_562
timestamp 1586364061
transform 1 0 52808 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_551
timestamp 1586364061
transform 1 0 54464 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_581
timestamp 1586364061
transform 1 0 54556 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_574
timestamp 1586364061
transform 1 0 53912 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_586
timestamp 1586364061
transform 1 0 55016 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_593
timestamp 1586364061
transform 1 0 55660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_605
timestamp 1586364061
transform 1 0 56764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_598
timestamp 1586364061
transform 1 0 56120 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_626
timestamp 1586364061
transform 1 0 57224 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_617
timestamp 1586364061
transform 1 0 57868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_611
timestamp 1586364061
transform 1 0 57316 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_623
timestamp 1586364061
transform 1 0 58420 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_552
timestamp 1586364061
transform 1 0 60076 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_629
timestamp 1586364061
transform 1 0 58972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_642
timestamp 1586364061
transform 1 0 60168 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_635
timestamp 1586364061
transform 1 0 59524 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_654
timestamp 1586364061
transform 1 0 61272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_647
timestamp 1586364061
transform 1 0 60628 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_659
timestamp 1586364061
transform 1 0 61732 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_627
timestamp 1586364061
transform 1 0 62836 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_666
timestamp 1586364061
transform 1 0 62376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_672
timestamp 1586364061
transform 1 0 62928 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_678
timestamp 1586364061
transform 1 0 63480 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_690
timestamp 1586364061
transform 1 0 64584 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_684
timestamp 1586364061
transform 1 0 64032 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_553
timestamp 1586364061
transform 1 0 65688 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_703
timestamp 1586364061
transform 1 0 65780 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_696
timestamp 1586364061
transform 1 0 65136 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_708
timestamp 1586364061
transform 1 0 66240 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_715
timestamp 1586364061
transform 1 0 66884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_727
timestamp 1586364061
transform 1 0 67988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_720
timestamp 1586364061
transform 1 0 67344 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_628
timestamp 1586364061
transform 1 0 68448 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_739
timestamp 1586364061
transform 1 0 69092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_733
timestamp 1586364061
transform 1 0 68540 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_745
timestamp 1586364061
transform 1 0 69644 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_554
timestamp 1586364061
transform 1 0 71300 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_751
timestamp 1586364061
transform 1 0 70196 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_764
timestamp 1586364061
transform 1 0 71392 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_757
timestamp 1586364061
transform 1 0 70748 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_776
timestamp 1586364061
transform 1 0 72496 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_769
timestamp 1586364061
transform 1 0 71852 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_781
timestamp 1586364061
transform 1 0 72956 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_629
timestamp 1586364061
transform 1 0 74060 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_788
timestamp 1586364061
transform 1 0 73600 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_800
timestamp 1586364061
transform 1 0 74704 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_794
timestamp 1586364061
transform 1 0 74152 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_812
timestamp 1586364061
transform 1 0 75808 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_806
timestamp 1586364061
transform 1 0 75256 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_818
timestamp 1586364061
transform 1 0 76360 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_555
timestamp 1586364061
transform 1 0 76912 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_825
timestamp 1586364061
transform 1 0 77004 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_837
timestamp 1586364061
transform 1 0 78108 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_830
timestamp 1586364061
transform 1 0 77464 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_630
timestamp 1586364061
transform 1 0 79672 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_849
timestamp 1586364061
transform 1 0 79212 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_842
timestamp 1586364061
transform 1 0 78568 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_855
timestamp 1586364061
transform 1 0 79764 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_861
timestamp 1586364061
transform 1 0 80316 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_873
timestamp 1586364061
transform 1 0 81420 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_867
timestamp 1586364061
transform 1 0 80868 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_556
timestamp 1586364061
transform 1 0 82524 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_886
timestamp 1586364061
transform 1 0 82616 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_879
timestamp 1586364061
transform 1 0 81972 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_891
timestamp 1586364061
transform 1 0 83076 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_898
timestamp 1586364061
transform 1 0 83720 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_903
timestamp 1586364061
transform 1 0 84180 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_631
timestamp 1586364061
transform 1 0 85284 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_910
timestamp 1586364061
transform 1 0 84824 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_922
timestamp 1586364061
transform 1 0 85928 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_916
timestamp 1586364061
transform 1 0 85376 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_934
timestamp 1586364061
transform 1 0 87032 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_928
timestamp 1586364061
transform 1 0 86480 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_940
timestamp 1586364061
transform 1 0 87584 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_557
timestamp 1586364061
transform 1 0 88136 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_947
timestamp 1586364061
transform 1 0 88228 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_959
timestamp 1586364061
transform 1 0 89332 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_952
timestamp 1586364061
transform 1 0 88688 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_632
timestamp 1586364061
transform 1 0 90896 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_971
timestamp 1586364061
transform 1 0 90436 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_964
timestamp 1586364061
transform 1 0 89792 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_977
timestamp 1586364061
transform 1 0 90988 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_983
timestamp 1586364061
transform 1 0 91540 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_995
timestamp 1586364061
transform 1 0 92644 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_989
timestamp 1586364061
transform 1 0 92092 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_558
timestamp 1586364061
transform 1 0 93748 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1008
timestamp 1586364061
transform 1 0 93840 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1001
timestamp 1586364061
transform 1 0 93196 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1013
timestamp 1586364061
transform 1 0 94300 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1020
timestamp 1586364061
transform 1 0 94944 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1032
timestamp 1586364061
transform 1 0 96048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1025
timestamp 1586364061
transform 1 0 95404 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_633
timestamp 1586364061
transform 1 0 96508 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1044
timestamp 1586364061
transform 1 0 97152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1038
timestamp 1586364061
transform 1 0 96600 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1050
timestamp 1586364061
transform 1 0 97704 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_559
timestamp 1586364061
transform 1 0 99360 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1056
timestamp 1586364061
transform 1 0 98256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1069
timestamp 1586364061
transform 1 0 99452 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1062
timestamp 1586364061
transform 1 0 98808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1081
timestamp 1586364061
transform 1 0 100556 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1074
timestamp 1586364061
transform 1 0 99912 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1086
timestamp 1586364061
transform 1 0 101016 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_634
timestamp 1586364061
transform 1 0 102120 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1093
timestamp 1586364061
transform 1 0 101660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1105
timestamp 1586364061
transform 1 0 102764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1099
timestamp 1586364061
transform 1 0 102212 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1117
timestamp 1586364061
transform 1 0 103868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1111
timestamp 1586364061
transform 1 0 103316 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1123
timestamp 1586364061
transform 1 0 104420 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_560
timestamp 1586364061
transform 1 0 104972 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1130
timestamp 1586364061
transform 1 0 105064 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1135
timestamp 1586364061
transform 1 0 105524 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_635
timestamp 1586364061
transform 1 0 107732 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1142
timestamp 1586364061
transform 1 0 106168 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1154
timestamp 1586364061
transform 1 0 107272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1147
timestamp 1586364061
transform 1 0 106628 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1166
timestamp 1586364061
transform 1 0 108376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1160
timestamp 1586364061
transform 1 0 107824 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1172
timestamp 1586364061
transform 1 0 108928 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_561
timestamp 1586364061
transform 1 0 110584 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1178
timestamp 1586364061
transform 1 0 109480 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1191
timestamp 1586364061
transform 1 0 110676 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1184
timestamp 1586364061
transform 1 0 110032 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1203
timestamp 1586364061
transform 1 0 111780 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1196
timestamp 1586364061
transform 1 0 111136 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1208
timestamp 1586364061
transform 1 0 112240 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_636
timestamp 1586364061
transform 1 0 113344 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1215
timestamp 1586364061
transform 1 0 112884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1227
timestamp 1586364061
transform 1 0 113988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1221
timestamp 1586364061
transform 1 0 113436 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1239
timestamp 1586364061
transform 1 0 115092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1233
timestamp 1586364061
transform 1 0 114540 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1245
timestamp 1586364061
transform 1 0 115644 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_562
timestamp 1586364061
transform 1 0 116196 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1252
timestamp 1586364061
transform 1 0 116288 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1264
timestamp 1586364061
transform 1 0 117392 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1257
timestamp 1586364061
transform 1 0 116748 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_637
timestamp 1586364061
transform 1 0 118956 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1276
timestamp 1586364061
transform 1 0 118496 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1269
timestamp 1586364061
transform 1 0 117852 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1282
timestamp 1586364061
transform 1 0 119048 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1288
timestamp 1586364061
transform 1 0 119600 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1300
timestamp 1586364061
transform 1 0 120704 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1294
timestamp 1586364061
transform 1 0 120152 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_563
timestamp 1586364061
transform 1 0 121808 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1313
timestamp 1586364061
transform 1 0 121900 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1306
timestamp 1586364061
transform 1 0 121256 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1318
timestamp 1586364061
transform 1 0 122360 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1325
timestamp 1586364061
transform 1 0 123004 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1337
timestamp 1586364061
transform 1 0 124108 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1330
timestamp 1586364061
transform 1 0 123464 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_638
timestamp 1586364061
transform 1 0 124568 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1349
timestamp 1586364061
transform 1 0 125212 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1343
timestamp 1586364061
transform 1 0 124660 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1355
timestamp 1586364061
transform 1 0 125764 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_564
timestamp 1586364061
transform 1 0 127420 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1361
timestamp 1586364061
transform 1 0 126316 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1367
timestamp 1586364061
transform 1 0 126868 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1374
timestamp 1586364061
transform 1 0 127512 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1386
timestamp 1586364061
transform 1 0 128616 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1379
timestamp 1586364061
transform 1 0 127972 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1391
timestamp 1586364061
transform 1 0 129076 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_639
timestamp 1586364061
transform 1 0 130180 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1398
timestamp 1586364061
transform 1 0 129720 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1404
timestamp 1586364061
transform 1 0 130272 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1410
timestamp 1586364061
transform 1 0 130824 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1422
timestamp 1586364061
transform 1 0 131928 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1416
timestamp 1586364061
transform 1 0 131376 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_565
timestamp 1586364061
transform 1 0 133032 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1435
timestamp 1586364061
transform 1 0 133124 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1428
timestamp 1586364061
transform 1 0 132480 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1440
timestamp 1586364061
transform 1 0 133584 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1447
timestamp 1586364061
transform 1 0 134228 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1459
timestamp 1586364061
transform 1 0 135332 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1452
timestamp 1586364061
transform 1 0 134688 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_640
timestamp 1586364061
transform 1 0 135792 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1471
timestamp 1586364061
transform 1 0 136436 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1465
timestamp 1586364061
transform 1 0 135884 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1477
timestamp 1586364061
transform 1 0 136988 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_566
timestamp 1586364061
transform 1 0 138644 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1483
timestamp 1586364061
transform 1 0 137540 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1496
timestamp 1586364061
transform 1 0 138736 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1489
timestamp 1586364061
transform 1 0 138092 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1508
timestamp 1586364061
transform 1 0 139840 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1501
timestamp 1586364061
transform 1 0 139196 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1513
timestamp 1586364061
transform 1 0 140300 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_641
timestamp 1586364061
transform 1 0 141404 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1520
timestamp 1586364061
transform 1 0 140944 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1532
timestamp 1586364061
transform 1 0 142048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1526
timestamp 1586364061
transform 1 0 141496 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1544
timestamp 1586364061
transform 1 0 143152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1538
timestamp 1586364061
transform 1 0 142600 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1550
timestamp 1586364061
transform 1 0 143704 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_567
timestamp 1586364061
transform 1 0 144256 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1557
timestamp 1586364061
transform 1 0 144348 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1569
timestamp 1586364061
transform 1 0 145452 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1562
timestamp 1586364061
transform 1 0 144808 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_642
timestamp 1586364061
transform 1 0 147016 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1581
timestamp 1586364061
transform 1 0 146556 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1574
timestamp 1586364061
transform 1 0 145912 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1587
timestamp 1586364061
transform 1 0 147108 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1593
timestamp 1586364061
transform 1 0 147660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1605
timestamp 1586364061
transform 1 0 148764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1599
timestamp 1586364061
transform 1 0 148212 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_568
timestamp 1586364061
transform 1 0 149868 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1618
timestamp 1586364061
transform 1 0 149960 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1611
timestamp 1586364061
transform 1 0 149316 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1623
timestamp 1586364061
transform 1 0 150420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1630
timestamp 1586364061
transform 1 0 151064 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1635
timestamp 1586364061
transform 1 0 151524 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_643
timestamp 1586364061
transform 1 0 152628 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1642
timestamp 1586364061
transform 1 0 152168 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1654
timestamp 1586364061
transform 1 0 153272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1648
timestamp 1586364061
transform 1 0 152720 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1666
timestamp 1586364061
transform 1 0 154376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1660
timestamp 1586364061
transform 1 0 153824 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1672
timestamp 1586364061
transform 1 0 154928 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_569
timestamp 1586364061
transform 1 0 155480 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1679
timestamp 1586364061
transform 1 0 155572 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1691
timestamp 1586364061
transform 1 0 156676 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1684
timestamp 1586364061
transform 1 0 156032 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_644
timestamp 1586364061
transform 1 0 158240 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1703
timestamp 1586364061
transform 1 0 157780 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1696
timestamp 1586364061
transform 1 0 157136 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1709
timestamp 1586364061
transform 1 0 158332 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1715
timestamp 1586364061
transform 1 0 158884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1727
timestamp 1586364061
transform 1 0 159988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1721
timestamp 1586364061
transform 1 0 159436 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_570
timestamp 1586364061
transform 1 0 161092 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1740
timestamp 1586364061
transform 1 0 161184 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1733
timestamp 1586364061
transform 1 0 160540 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1745
timestamp 1586364061
transform 1 0 161644 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1752
timestamp 1586364061
transform 1 0 162288 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1764
timestamp 1586364061
transform 1 0 163392 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1757
timestamp 1586364061
transform 1 0 162748 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_645
timestamp 1586364061
transform 1 0 163852 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1776
timestamp 1586364061
transform 1 0 164496 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1770
timestamp 1586364061
transform 1 0 163944 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1782
timestamp 1586364061
transform 1 0 165048 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_571
timestamp 1586364061
transform 1 0 166704 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1788
timestamp 1586364061
transform 1 0 165600 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1801
timestamp 1586364061
transform 1 0 166796 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1794
timestamp 1586364061
transform 1 0 166152 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1813
timestamp 1586364061
transform 1 0 167900 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1806
timestamp 1586364061
transform 1 0 167256 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1818
timestamp 1586364061
transform 1 0 168360 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_646
timestamp 1586364061
transform 1 0 169464 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1825
timestamp 1586364061
transform 1 0 169004 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1837
timestamp 1586364061
transform 1 0 170108 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1831
timestamp 1586364061
transform 1 0 169556 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1849
timestamp 1586364061
transform 1 0 171212 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1843
timestamp 1586364061
transform 1 0 170660 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1855
timestamp 1586364061
transform 1 0 171764 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_572
timestamp 1586364061
transform 1 0 172316 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1862
timestamp 1586364061
transform 1 0 172408 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1867
timestamp 1586364061
transform 1 0 172868 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1874
timestamp 1586364061
transform 1 0 173512 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1886
timestamp 1586364061
transform 1 0 174616 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1879
timestamp 1586364061
transform 1 0 173972 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_647
timestamp 1586364061
transform 1 0 175076 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1898
timestamp 1586364061
transform 1 0 175720 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1892
timestamp 1586364061
transform 1 0 175168 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1904
timestamp 1586364061
transform 1 0 176272 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_573
timestamp 1586364061
transform 1 0 177928 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1910
timestamp 1586364061
transform 1 0 176824 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1923
timestamp 1586364061
transform 1 0 178020 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1916
timestamp 1586364061
transform 1 0 177376 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1935
timestamp 1586364061
transform 1 0 179124 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1928
timestamp 1586364061
transform 1 0 178480 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1940
timestamp 1586364061
transform 1 0 179584 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_648
timestamp 1586364061
transform 1 0 180688 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1947
timestamp 1586364061
transform 1 0 180228 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1959
timestamp 1586364061
transform 1 0 181332 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1953
timestamp 1586364061
transform 1 0 180780 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1971
timestamp 1586364061
transform 1 0 182436 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1965
timestamp 1586364061
transform 1 0 181884 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1977
timestamp 1586364061
transform 1 0 182988 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_574
timestamp 1586364061
transform 1 0 183540 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_1984
timestamp 1586364061
transform 1 0 183632 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_1996
timestamp 1586364061
transform 1 0 184736 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_1989
timestamp 1586364061
transform 1 0 184092 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_649
timestamp 1586364061
transform 1 0 186300 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2008
timestamp 1586364061
transform 1 0 185840 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2001
timestamp 1586364061
transform 1 0 185196 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2014
timestamp 1586364061
transform 1 0 186392 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2020
timestamp 1586364061
transform 1 0 186944 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2032
timestamp 1586364061
transform 1 0 188048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2026
timestamp 1586364061
transform 1 0 187496 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_575
timestamp 1586364061
transform 1 0 189152 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2045
timestamp 1586364061
transform 1 0 189244 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2038
timestamp 1586364061
transform 1 0 188600 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2050
timestamp 1586364061
transform 1 0 189704 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2057
timestamp 1586364061
transform 1 0 190348 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2069
timestamp 1586364061
transform 1 0 191452 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2062
timestamp 1586364061
transform 1 0 190808 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_650
timestamp 1586364061
transform 1 0 191912 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2081
timestamp 1586364061
transform 1 0 192556 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2075
timestamp 1586364061
transform 1 0 192004 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2093
timestamp 1586364061
transform 1 0 193660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2087
timestamp 1586364061
transform 1 0 193108 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2099
timestamp 1586364061
transform 1 0 194212 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_576
timestamp 1586364061
transform 1 0 194764 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2106
timestamp 1586364061
transform 1 0 194856 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2118
timestamp 1586364061
transform 1 0 195960 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2111
timestamp 1586364061
transform 1 0 195316 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_651
timestamp 1586364061
transform 1 0 197524 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2130
timestamp 1586364061
transform 1 0 197064 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2123
timestamp 1586364061
transform 1 0 196420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2136
timestamp 1586364061
transform 1 0 197616 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2142
timestamp 1586364061
transform 1 0 198168 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2154
timestamp 1586364061
transform 1 0 199272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2148
timestamp 1586364061
transform 1 0 198720 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_577
timestamp 1586364061
transform 1 0 200376 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2167
timestamp 1586364061
transform 1 0 200468 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2160
timestamp 1586364061
transform 1 0 199824 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2172
timestamp 1586364061
transform 1 0 200928 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2179
timestamp 1586364061
transform 1 0 201572 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2191
timestamp 1586364061
transform 1 0 202676 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2184
timestamp 1586364061
transform 1 0 202032 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_652
timestamp 1586364061
transform 1 0 203136 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2203
timestamp 1586364061
transform 1 0 203780 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2197
timestamp 1586364061
transform 1 0 203228 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2209
timestamp 1586364061
transform 1 0 204332 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_578
timestamp 1586364061
transform 1 0 205988 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2215
timestamp 1586364061
transform 1 0 204884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2228
timestamp 1586364061
transform 1 0 206080 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2221
timestamp 1586364061
transform 1 0 205436 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2240
timestamp 1586364061
transform 1 0 207184 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2233
timestamp 1586364061
transform 1 0 206540 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2245
timestamp 1586364061
transform 1 0 207644 0 1 5984
box -38 -48 1142 592
use scs8hd_buf_2  _21_
timestamp 1586364061
transform 1 0 209300 0 -1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_653
timestamp 1586364061
transform 1 0 208748 0 1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_2252
timestamp 1586364061
transform 1 0 208288 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_6_2260
timestamp 1586364061
transform 1 0 209024 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_2258
timestamp 1586364061
transform 1 0 208840 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2267
timestamp 1586364061
transform 1 0 209668 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_6_2279
timestamp 1586364061
transform 1 0 210772 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_7_2270
timestamp 1586364061
transform 1 0 209944 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2282
timestamp 1586364061
transform 1 0 211048 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_579
timestamp 1586364061
transform 1 0 211600 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_2287
timestamp 1586364061
transform 1 0 211508 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2289
timestamp 1586364061
transform 1 0 211692 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_7_2294
timestamp 1586364061
transform 1 0 212152 0 1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_2300
timestamp 1586364061
transform 1 0 212704 0 1 5984
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_654
timestamp 1586364061
transform 1 0 214360 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__23__A
timestamp 1586364061
transform 1 0 212796 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_2301
timestamp 1586364061
transform 1 0 212796 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2313
timestamp 1586364061
transform 1 0 213900 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2303
timestamp 1586364061
transform 1 0 212980 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_7_2315
timestamp 1586364061
transform 1 0 214084 0 1 5984
box -38 -48 314 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 215464 0 1 5984
box -38 -48 774 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 215280 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 215280 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 214912 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_2325
timestamp 1586364061
transform 1 0 215004 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_2336
timestamp 1586364061
transform 1 0 216016 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_2319
timestamp 1586364061
transform 1 0 214452 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_2323
timestamp 1586364061
transform 1 0 214820 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_2326
timestamp 1586364061
transform 1 0 215096 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_580
timestamp 1586364061
transform 1 0 217212 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 216384 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 216200 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_2340
timestamp 1586364061
transform 1 0 216384 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_2348
timestamp 1586364061
transform 1 0 217120 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2350
timestamp 1586364061
transform 1 0 217304 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_2338
timestamp 1586364061
transform 1 0 216200 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_2342
timestamp 1586364061
transform 1 0 216568 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2354
timestamp 1586364061
transform 1 0 217672 0 1 5984
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 219144 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_2362
timestamp 1586364061
transform 1 0 218408 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_2366
timestamp 1586364061
transform 1 0 218776 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_2372
timestamp 1586364061
transform 1 0 219328 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 219696 0 -1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_655
timestamp 1586364061
transform 1 0 219972 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__10__A
timestamp 1586364061
transform 1 0 220892 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 219512 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_2374
timestamp 1586364061
transform 1 0 219512 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_2387
timestamp 1586364061
transform 1 0 220708 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_2376
timestamp 1586364061
transform 1 0 219696 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_2380
timestamp 1586364061
transform 1 0 220064 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2391
timestamp 1586364061
transform 1 0 221076 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_6_2403
timestamp 1586364061
transform 1 0 222180 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_12  FILLER_7_2392
timestamp 1586364061
transform 1 0 221168 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2404
timestamp 1586364061
transform 1 0 222272 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_581
timestamp 1586364061
transform 1 0 222824 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_2409
timestamp 1586364061
transform 1 0 222732 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2411
timestamp 1586364061
transform 1 0 222916 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2423
timestamp 1586364061
transform 1 0 224020 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2416
timestamp 1586364061
transform 1 0 223376 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_656
timestamp 1586364061
transform 1 0 225584 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2435
timestamp 1586364061
transform 1 0 225124 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2428
timestamp 1586364061
transform 1 0 224480 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2441
timestamp 1586364061
transform 1 0 225676 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2447
timestamp 1586364061
transform 1 0 226228 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2459
timestamp 1586364061
transform 1 0 227332 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2453
timestamp 1586364061
transform 1 0 226780 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_582
timestamp 1586364061
transform 1 0 228436 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2472
timestamp 1586364061
transform 1 0 228528 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2465
timestamp 1586364061
transform 1 0 227884 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2477
timestamp 1586364061
transform 1 0 228988 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2484
timestamp 1586364061
transform 1 0 229632 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2496
timestamp 1586364061
transform 1 0 230736 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2489
timestamp 1586364061
transform 1 0 230092 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_657
timestamp 1586364061
transform 1 0 231196 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 232392 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_2508
timestamp 1586364061
transform 1 0 231840 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_12  FILLER_7_2502
timestamp 1586364061
transform 1 0 231288 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2514
timestamp 1586364061
transform 1 0 232392 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_583
timestamp 1586364061
transform 1 0 234048 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2516
timestamp 1586364061
transform 1 0 232576 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_6_2528
timestamp 1586364061
transform 1 0 233680 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_7_2526
timestamp 1586364061
transform 1 0 233496 0 1 5984
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 234140 0 -1 5984
box -38 -48 1050 592
use scs8hd_decap_12  FILLER_6_2544
timestamp 1586364061
transform 1 0 235152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2538
timestamp 1586364061
transform 1 0 234600 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2550
timestamp 1586364061
transform 1 0 235704 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_658
timestamp 1586364061
transform 1 0 236808 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 237268 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_2556
timestamp 1586364061
transform 1 0 236256 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_6_2568
timestamp 1586364061
transform 1 0 237360 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_2563
timestamp 1586364061
transform 1 0 236900 0 1 5984
box -38 -48 406 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 237452 0 1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 237452 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_2571
timestamp 1586364061
transform 1 0 237636 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_6_2583
timestamp 1586364061
transform 1 0 238740 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_7_2577
timestamp 1586364061
transform 1 0 238188 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_584
timestamp 1586364061
transform 1 0 239660 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_2591
timestamp 1586364061
transform 1 0 239476 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_2594
timestamp 1586364061
transform 1 0 239752 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2589
timestamp 1586364061
transform 1 0 239292 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2601
timestamp 1586364061
transform 1 0 240396 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2606
timestamp 1586364061
transform 1 0 240856 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2618
timestamp 1586364061
transform 1 0 241960 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_2613
timestamp 1586364061
transform 1 0 241500 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_2621
timestamp 1586364061
transform 1 0 242236 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_659
timestamp 1586364061
transform 1 0 242420 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2630
timestamp 1586364061
transform 1 0 243064 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2624
timestamp 1586364061
transform 1 0 242512 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2636
timestamp 1586364061
transform 1 0 243616 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_585
timestamp 1586364061
transform 1 0 245272 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2642
timestamp 1586364061
transform 1 0 244168 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2655
timestamp 1586364061
transform 1 0 245364 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2648
timestamp 1586364061
transform 1 0 244720 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2667
timestamp 1586364061
transform 1 0 246468 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2660
timestamp 1586364061
transform 1 0 245824 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2672
timestamp 1586364061
transform 1 0 246928 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_660
timestamp 1586364061
transform 1 0 248032 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2679
timestamp 1586364061
transform 1 0 247572 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2691
timestamp 1586364061
transform 1 0 248676 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2685
timestamp 1586364061
transform 1 0 248124 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2703
timestamp 1586364061
transform 1 0 249780 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2697
timestamp 1586364061
transform 1 0 249228 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2709
timestamp 1586364061
transform 1 0 250332 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_586
timestamp 1586364061
transform 1 0 250884 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2716
timestamp 1586364061
transform 1 0 250976 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2728
timestamp 1586364061
transform 1 0 252080 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2721
timestamp 1586364061
transform 1 0 251436 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_661
timestamp 1586364061
transform 1 0 253644 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2740
timestamp 1586364061
transform 1 0 253184 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2733
timestamp 1586364061
transform 1 0 252540 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2746
timestamp 1586364061
transform 1 0 253736 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2752
timestamp 1586364061
transform 1 0 254288 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2764
timestamp 1586364061
transform 1 0 255392 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2758
timestamp 1586364061
transform 1 0 254840 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_587
timestamp 1586364061
transform 1 0 256496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2777
timestamp 1586364061
transform 1 0 256588 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2770
timestamp 1586364061
transform 1 0 255944 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2782
timestamp 1586364061
transform 1 0 257048 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2789
timestamp 1586364061
transform 1 0 257692 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2794
timestamp 1586364061
transform 1 0 258152 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_662
timestamp 1586364061
transform 1 0 259256 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2801
timestamp 1586364061
transform 1 0 258796 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2813
timestamp 1586364061
transform 1 0 259900 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2807
timestamp 1586364061
transform 1 0 259348 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2825
timestamp 1586364061
transform 1 0 261004 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2819
timestamp 1586364061
transform 1 0 260452 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2831
timestamp 1586364061
transform 1 0 261556 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_588
timestamp 1586364061
transform 1 0 262108 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2838
timestamp 1586364061
transform 1 0 262200 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2850
timestamp 1586364061
transform 1 0 263304 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2843
timestamp 1586364061
transform 1 0 262660 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_663
timestamp 1586364061
transform 1 0 264868 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2862
timestamp 1586364061
transform 1 0 264408 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2855
timestamp 1586364061
transform 1 0 263764 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2868
timestamp 1586364061
transform 1 0 264960 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2874
timestamp 1586364061
transform 1 0 265512 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2886
timestamp 1586364061
transform 1 0 266616 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2880
timestamp 1586364061
transform 1 0 266064 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_589
timestamp 1586364061
transform 1 0 267720 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2899
timestamp 1586364061
transform 1 0 267812 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2892
timestamp 1586364061
transform 1 0 267168 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2904
timestamp 1586364061
transform 1 0 268272 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2911
timestamp 1586364061
transform 1 0 268916 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2923
timestamp 1586364061
transform 1 0 270020 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2916
timestamp 1586364061
transform 1 0 269376 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_664
timestamp 1586364061
transform 1 0 270480 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2935
timestamp 1586364061
transform 1 0 271124 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2929
timestamp 1586364061
transform 1 0 270572 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2941
timestamp 1586364061
transform 1 0 271676 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_590
timestamp 1586364061
transform 1 0 273332 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2947
timestamp 1586364061
transform 1 0 272228 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2960
timestamp 1586364061
transform 1 0 273424 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2953
timestamp 1586364061
transform 1 0 272780 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2972
timestamp 1586364061
transform 1 0 274528 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2965
timestamp 1586364061
transform 1 0 273884 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2977
timestamp 1586364061
transform 1 0 274988 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_665
timestamp 1586364061
transform 1 0 276092 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_2984
timestamp 1586364061
transform 1 0 275632 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_2996
timestamp 1586364061
transform 1 0 276736 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_2990
timestamp 1586364061
transform 1 0 276184 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3008
timestamp 1586364061
transform 1 0 277840 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3002
timestamp 1586364061
transform 1 0 277288 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3014
timestamp 1586364061
transform 1 0 278392 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_591
timestamp 1586364061
transform 1 0 278944 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3021
timestamp 1586364061
transform 1 0 279036 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3026
timestamp 1586364061
transform 1 0 279496 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_666
timestamp 1586364061
transform 1 0 281704 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3033
timestamp 1586364061
transform 1 0 280140 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3045
timestamp 1586364061
transform 1 0 281244 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3038
timestamp 1586364061
transform 1 0 280600 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3057
timestamp 1586364061
transform 1 0 282348 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3051
timestamp 1586364061
transform 1 0 281796 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3063
timestamp 1586364061
transform 1 0 282900 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_592
timestamp 1586364061
transform 1 0 284556 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3069
timestamp 1586364061
transform 1 0 283452 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3082
timestamp 1586364061
transform 1 0 284648 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3075
timestamp 1586364061
transform 1 0 284004 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3094
timestamp 1586364061
transform 1 0 285752 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3087
timestamp 1586364061
transform 1 0 285108 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3099
timestamp 1586364061
transform 1 0 286212 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_667
timestamp 1586364061
transform 1 0 287316 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3106
timestamp 1586364061
transform 1 0 286856 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3118
timestamp 1586364061
transform 1 0 287960 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3112
timestamp 1586364061
transform 1 0 287408 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3130
timestamp 1586364061
transform 1 0 289064 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3124
timestamp 1586364061
transform 1 0 288512 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3136
timestamp 1586364061
transform 1 0 289616 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_593
timestamp 1586364061
transform 1 0 290168 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3143
timestamp 1586364061
transform 1 0 290260 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3155
timestamp 1586364061
transform 1 0 291364 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3148
timestamp 1586364061
transform 1 0 290720 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_668
timestamp 1586364061
transform 1 0 292928 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3167
timestamp 1586364061
transform 1 0 292468 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3160
timestamp 1586364061
transform 1 0 291824 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3173
timestamp 1586364061
transform 1 0 293020 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3179
timestamp 1586364061
transform 1 0 293572 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3191
timestamp 1586364061
transform 1 0 294676 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3185
timestamp 1586364061
transform 1 0 294124 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_594
timestamp 1586364061
transform 1 0 295780 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3204
timestamp 1586364061
transform 1 0 295872 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3197
timestamp 1586364061
transform 1 0 295228 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3209
timestamp 1586364061
transform 1 0 296332 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3216
timestamp 1586364061
transform 1 0 296976 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3228
timestamp 1586364061
transform 1 0 298080 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3221
timestamp 1586364061
transform 1 0 297436 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_669
timestamp 1586364061
transform 1 0 298540 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3240
timestamp 1586364061
transform 1 0 299184 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3234
timestamp 1586364061
transform 1 0 298632 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3246
timestamp 1586364061
transform 1 0 299736 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_595
timestamp 1586364061
transform 1 0 301392 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3252
timestamp 1586364061
transform 1 0 300288 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3258
timestamp 1586364061
transform 1 0 300840 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3265
timestamp 1586364061
transform 1 0 301484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3277
timestamp 1586364061
transform 1 0 302588 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3270
timestamp 1586364061
transform 1 0 301944 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_670
timestamp 1586364061
transform 1 0 304152 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3289
timestamp 1586364061
transform 1 0 303692 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3282
timestamp 1586364061
transform 1 0 303048 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3295
timestamp 1586364061
transform 1 0 304244 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3301
timestamp 1586364061
transform 1 0 304796 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3313
timestamp 1586364061
transform 1 0 305900 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3307
timestamp 1586364061
transform 1 0 305348 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_596
timestamp 1586364061
transform 1 0 307004 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3326
timestamp 1586364061
transform 1 0 307096 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3319
timestamp 1586364061
transform 1 0 306452 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3331
timestamp 1586364061
transform 1 0 307556 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3338
timestamp 1586364061
transform 1 0 308200 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3350
timestamp 1586364061
transform 1 0 309304 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3343
timestamp 1586364061
transform 1 0 308660 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_671
timestamp 1586364061
transform 1 0 309764 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3362
timestamp 1586364061
transform 1 0 310408 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3356
timestamp 1586364061
transform 1 0 309856 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3368
timestamp 1586364061
transform 1 0 310960 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_597
timestamp 1586364061
transform 1 0 312616 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3374
timestamp 1586364061
transform 1 0 311512 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3387
timestamp 1586364061
transform 1 0 312708 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3380
timestamp 1586364061
transform 1 0 312064 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3399
timestamp 1586364061
transform 1 0 313812 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3392
timestamp 1586364061
transform 1 0 313168 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3404
timestamp 1586364061
transform 1 0 314272 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_672
timestamp 1586364061
transform 1 0 315376 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3411
timestamp 1586364061
transform 1 0 314916 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3423
timestamp 1586364061
transform 1 0 316020 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3417
timestamp 1586364061
transform 1 0 315468 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3435
timestamp 1586364061
transform 1 0 317124 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3429
timestamp 1586364061
transform 1 0 316572 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3441
timestamp 1586364061
transform 1 0 317676 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_598
timestamp 1586364061
transform 1 0 318228 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3448
timestamp 1586364061
transform 1 0 318320 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3460
timestamp 1586364061
transform 1 0 319424 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3453
timestamp 1586364061
transform 1 0 318780 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_673
timestamp 1586364061
transform 1 0 320988 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3472
timestamp 1586364061
transform 1 0 320528 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3465
timestamp 1586364061
transform 1 0 319884 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3478
timestamp 1586364061
transform 1 0 321080 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3484
timestamp 1586364061
transform 1 0 321632 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3496
timestamp 1586364061
transform 1 0 322736 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3490
timestamp 1586364061
transform 1 0 322184 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_599
timestamp 1586364061
transform 1 0 323840 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3509
timestamp 1586364061
transform 1 0 323932 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3502
timestamp 1586364061
transform 1 0 323288 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3521
timestamp 1586364061
transform 1 0 325036 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3514
timestamp 1586364061
transform 1 0 324392 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3526
timestamp 1586364061
transform 1 0 325496 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_674
timestamp 1586364061
transform 1 0 326600 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3533
timestamp 1586364061
transform 1 0 326140 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3545
timestamp 1586364061
transform 1 0 327244 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3539
timestamp 1586364061
transform 1 0 326692 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3557
timestamp 1586364061
transform 1 0 328348 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3551
timestamp 1586364061
transform 1 0 327796 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3563
timestamp 1586364061
transform 1 0 328900 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_600
timestamp 1586364061
transform 1 0 329452 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3570
timestamp 1586364061
transform 1 0 329544 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3582
timestamp 1586364061
transform 1 0 330648 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3575
timestamp 1586364061
transform 1 0 330004 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_675
timestamp 1586364061
transform 1 0 332212 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3594
timestamp 1586364061
transform 1 0 331752 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3587
timestamp 1586364061
transform 1 0 331108 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3600
timestamp 1586364061
transform 1 0 332304 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3606
timestamp 1586364061
transform 1 0 332856 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3618
timestamp 1586364061
transform 1 0 333960 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3612
timestamp 1586364061
transform 1 0 333408 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_601
timestamp 1586364061
transform 1 0 335064 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3631
timestamp 1586364061
transform 1 0 335156 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3624
timestamp 1586364061
transform 1 0 334512 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3636
timestamp 1586364061
transform 1 0 335616 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3643
timestamp 1586364061
transform 1 0 336260 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3655
timestamp 1586364061
transform 1 0 337364 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3648
timestamp 1586364061
transform 1 0 336720 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_676
timestamp 1586364061
transform 1 0 337824 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3667
timestamp 1586364061
transform 1 0 338468 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3661
timestamp 1586364061
transform 1 0 337916 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3673
timestamp 1586364061
transform 1 0 339020 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_602
timestamp 1586364061
transform 1 0 340676 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3679
timestamp 1586364061
transform 1 0 339572 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3692
timestamp 1586364061
transform 1 0 340768 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3685
timestamp 1586364061
transform 1 0 340124 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3704
timestamp 1586364061
transform 1 0 341872 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3697
timestamp 1586364061
transform 1 0 341228 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3709
timestamp 1586364061
transform 1 0 342332 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_677
timestamp 1586364061
transform 1 0 343436 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3716
timestamp 1586364061
transform 1 0 342976 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3722
timestamp 1586364061
transform 1 0 343528 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3728
timestamp 1586364061
transform 1 0 344080 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3740
timestamp 1586364061
transform 1 0 345184 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3734
timestamp 1586364061
transform 1 0 344632 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_603
timestamp 1586364061
transform 1 0 346288 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3753
timestamp 1586364061
transform 1 0 346380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3746
timestamp 1586364061
transform 1 0 345736 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3758
timestamp 1586364061
transform 1 0 346840 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3765
timestamp 1586364061
transform 1 0 347484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3777
timestamp 1586364061
transform 1 0 348588 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3770
timestamp 1586364061
transform 1 0 347944 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_678
timestamp 1586364061
transform 1 0 349048 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3789
timestamp 1586364061
transform 1 0 349692 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3783
timestamp 1586364061
transform 1 0 349140 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3795
timestamp 1586364061
transform 1 0 350244 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_604
timestamp 1586364061
transform 1 0 351900 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3801
timestamp 1586364061
transform 1 0 350796 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3814
timestamp 1586364061
transform 1 0 351992 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3807
timestamp 1586364061
transform 1 0 351348 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3826
timestamp 1586364061
transform 1 0 353096 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3819
timestamp 1586364061
transform 1 0 352452 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3831
timestamp 1586364061
transform 1 0 353556 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_679
timestamp 1586364061
transform 1 0 354660 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3838
timestamp 1586364061
transform 1 0 354200 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3850
timestamp 1586364061
transform 1 0 355304 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3844
timestamp 1586364061
transform 1 0 354752 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3862
timestamp 1586364061
transform 1 0 356408 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3856
timestamp 1586364061
transform 1 0 355856 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3868
timestamp 1586364061
transform 1 0 356960 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_605
timestamp 1586364061
transform 1 0 357512 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3875
timestamp 1586364061
transform 1 0 357604 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3887
timestamp 1586364061
transform 1 0 358708 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3880
timestamp 1586364061
transform 1 0 358064 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_680
timestamp 1586364061
transform 1 0 360272 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3899
timestamp 1586364061
transform 1 0 359812 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3892
timestamp 1586364061
transform 1 0 359168 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3905
timestamp 1586364061
transform 1 0 360364 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3911
timestamp 1586364061
transform 1 0 360916 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3923
timestamp 1586364061
transform 1 0 362020 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3917
timestamp 1586364061
transform 1 0 361468 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_606
timestamp 1586364061
transform 1 0 363124 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3936
timestamp 1586364061
transform 1 0 363216 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3929
timestamp 1586364061
transform 1 0 362572 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3941
timestamp 1586364061
transform 1 0 363676 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3948
timestamp 1586364061
transform 1 0 364320 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3953
timestamp 1586364061
transform 1 0 364780 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_681
timestamp 1586364061
transform 1 0 365884 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3960
timestamp 1586364061
transform 1 0 365424 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3972
timestamp 1586364061
transform 1 0 366528 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3966
timestamp 1586364061
transform 1 0 365976 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_3984
timestamp 1586364061
transform 1 0 367632 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3978
timestamp 1586364061
transform 1 0 367080 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3990
timestamp 1586364061
transform 1 0 368184 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_607
timestamp 1586364061
transform 1 0 368736 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_3997
timestamp 1586364061
transform 1 0 368828 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4009
timestamp 1586364061
transform 1 0 369932 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4002
timestamp 1586364061
transform 1 0 369288 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_682
timestamp 1586364061
transform 1 0 371496 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4021
timestamp 1586364061
transform 1 0 371036 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4014
timestamp 1586364061
transform 1 0 370392 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4027
timestamp 1586364061
transform 1 0 371588 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4033
timestamp 1586364061
transform 1 0 372140 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4045
timestamp 1586364061
transform 1 0 373244 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4039
timestamp 1586364061
transform 1 0 372692 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_608
timestamp 1586364061
transform 1 0 374348 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4058
timestamp 1586364061
transform 1 0 374440 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4051
timestamp 1586364061
transform 1 0 373796 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4063
timestamp 1586364061
transform 1 0 374900 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4070
timestamp 1586364061
transform 1 0 375544 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4082
timestamp 1586364061
transform 1 0 376648 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4075
timestamp 1586364061
transform 1 0 376004 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_683
timestamp 1586364061
transform 1 0 377108 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4094
timestamp 1586364061
transform 1 0 377752 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4088
timestamp 1586364061
transform 1 0 377200 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4100
timestamp 1586364061
transform 1 0 378304 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_609
timestamp 1586364061
transform 1 0 379960 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4106
timestamp 1586364061
transform 1 0 378856 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4119
timestamp 1586364061
transform 1 0 380052 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4112
timestamp 1586364061
transform 1 0 379408 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4131
timestamp 1586364061
transform 1 0 381156 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4124
timestamp 1586364061
transform 1 0 380512 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4136
timestamp 1586364061
transform 1 0 381616 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_684
timestamp 1586364061
transform 1 0 382720 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4143
timestamp 1586364061
transform 1 0 382260 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4155
timestamp 1586364061
transform 1 0 383364 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4149
timestamp 1586364061
transform 1 0 382812 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4167
timestamp 1586364061
transform 1 0 384468 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4161
timestamp 1586364061
transform 1 0 383916 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4173
timestamp 1586364061
transform 1 0 385020 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_610
timestamp 1586364061
transform 1 0 385572 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4180
timestamp 1586364061
transform 1 0 385664 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4185
timestamp 1586364061
transform 1 0 386124 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_685
timestamp 1586364061
transform 1 0 388332 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4192
timestamp 1586364061
transform 1 0 386768 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4204
timestamp 1586364061
transform 1 0 387872 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4197
timestamp 1586364061
transform 1 0 387228 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4216
timestamp 1586364061
transform 1 0 388976 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4210
timestamp 1586364061
transform 1 0 388424 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4222
timestamp 1586364061
transform 1 0 389528 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_611
timestamp 1586364061
transform 1 0 391184 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4228
timestamp 1586364061
transform 1 0 390080 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4241
timestamp 1586364061
transform 1 0 391276 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4234
timestamp 1586364061
transform 1 0 390632 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4253
timestamp 1586364061
transform 1 0 392380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4246
timestamp 1586364061
transform 1 0 391736 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4258
timestamp 1586364061
transform 1 0 392840 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_686
timestamp 1586364061
transform 1 0 393944 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4265
timestamp 1586364061
transform 1 0 393484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4277
timestamp 1586364061
transform 1 0 394588 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4271
timestamp 1586364061
transform 1 0 394036 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4289
timestamp 1586364061
transform 1 0 395692 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4283
timestamp 1586364061
transform 1 0 395140 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4295
timestamp 1586364061
transform 1 0 396244 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_612
timestamp 1586364061
transform 1 0 396796 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4302
timestamp 1586364061
transform 1 0 396888 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4314
timestamp 1586364061
transform 1 0 397992 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4307
timestamp 1586364061
transform 1 0 397348 0 1 5984
box -38 -48 1142 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 399648 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_687
timestamp 1586364061
transform 1 0 399556 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
timestamp 1586364061
transform 1 0 399372 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
timestamp 1586364061
transform 1 0 399648 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_4326
timestamp 1586364061
transform 1 0 399096 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_12  FILLER_6_4334
timestamp 1586364061
transform 1 0 399832 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_4319
timestamp 1586364061
transform 1 0 398452 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_4327
timestamp 1586364061
transform 1 0 399188 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_4346
timestamp 1586364061
transform 1 0 400936 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4340
timestamp 1586364061
transform 1 0 400384 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4352
timestamp 1586364061
transform 1 0 401488 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_613
timestamp 1586364061
transform 1 0 402408 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_4358
timestamp 1586364061
transform 1 0 402040 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_4363
timestamp 1586364061
transform 1 0 402500 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4364
timestamp 1586364061
transform 1 0 402592 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4375
timestamp 1586364061
transform 1 0 403604 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4387
timestamp 1586364061
transform 1 0 404708 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4376
timestamp 1586364061
transform 1 0 403696 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_688
timestamp 1586364061
transform 1 0 405168 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4399
timestamp 1586364061
transform 1 0 405812 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_4388
timestamp 1586364061
transform 1 0 404800 0 1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_7_4393
timestamp 1586364061
transform 1 0 405260 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4405
timestamp 1586364061
transform 1 0 406364 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_614
timestamp 1586364061
transform 1 0 408020 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4411
timestamp 1586364061
transform 1 0 406916 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4417
timestamp 1586364061
transform 1 0 407468 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4424
timestamp 1586364061
transform 1 0 408112 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4436
timestamp 1586364061
transform 1 0 409216 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4429
timestamp 1586364061
transform 1 0 408572 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4441
timestamp 1586364061
transform 1 0 409676 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_689
timestamp 1586364061
transform 1 0 410780 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4448
timestamp 1586364061
transform 1 0 410320 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4454
timestamp 1586364061
transform 1 0 410872 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4460
timestamp 1586364061
transform 1 0 411424 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4472
timestamp 1586364061
transform 1 0 412528 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4466
timestamp 1586364061
transform 1 0 411976 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_615
timestamp 1586364061
transform 1 0 413632 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4485
timestamp 1586364061
transform 1 0 413724 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4478
timestamp 1586364061
transform 1 0 413080 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4490
timestamp 1586364061
transform 1 0 414184 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4497
timestamp 1586364061
transform 1 0 414828 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4509
timestamp 1586364061
transform 1 0 415932 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4502
timestamp 1586364061
transform 1 0 415288 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_690
timestamp 1586364061
transform 1 0 416392 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4521
timestamp 1586364061
transform 1 0 417036 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4515
timestamp 1586364061
transform 1 0 416484 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4527
timestamp 1586364061
transform 1 0 417588 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_616
timestamp 1586364061
transform 1 0 419244 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_4533
timestamp 1586364061
transform 1 0 418140 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4546
timestamp 1586364061
transform 1 0 419336 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4539
timestamp 1586364061
transform 1 0 418692 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_4558
timestamp 1586364061
transform 1 0 420440 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4551
timestamp 1586364061
transform 1 0 419796 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_4563
timestamp 1586364061
transform 1 0 420900 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 422832 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 422832 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_691
timestamp 1586364061
transform 1 0 422004 0 1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_4570
timestamp 1586364061
transform 1 0 421544 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_6_4578
timestamp 1586364061
transform 1 0 422280 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_4576
timestamp 1586364061
transform 1 0 422096 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_4580
timestamp 1586364061
transform 1 0 422464 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_692
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_80
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_693
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_141
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_694
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_695
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_263
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_696
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_288
timestamp 1586364061
transform 1 0 27600 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_300
timestamp 1586364061
transform 1 0 28704 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_312
timestamp 1586364061
transform 1 0 29808 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_697
timestamp 1586364061
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_324
timestamp 1586364061
transform 1 0 30912 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_337
timestamp 1586364061
transform 1 0 32108 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_349
timestamp 1586364061
transform 1 0 33212 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_361
timestamp 1586364061
transform 1 0 34316 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_373
timestamp 1586364061
transform 1 0 35420 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_385
timestamp 1586364061
transform 1 0 36524 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_698
timestamp 1586364061
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_398
timestamp 1586364061
transform 1 0 37720 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_410
timestamp 1586364061
transform 1 0 38824 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_422
timestamp 1586364061
transform 1 0 39928 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_434
timestamp 1586364061
transform 1 0 41032 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_699
timestamp 1586364061
transform 1 0 43240 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_446
timestamp 1586364061
transform 1 0 42136 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_459
timestamp 1586364061
transform 1 0 43332 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_471
timestamp 1586364061
transform 1 0 44436 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_483
timestamp 1586364061
transform 1 0 45540 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_495
timestamp 1586364061
transform 1 0 46644 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_507
timestamp 1586364061
transform 1 0 47748 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_700
timestamp 1586364061
transform 1 0 48852 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_520
timestamp 1586364061
transform 1 0 48944 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_532
timestamp 1586364061
transform 1 0 50048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_544
timestamp 1586364061
transform 1 0 51152 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_556
timestamp 1586364061
transform 1 0 52256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_568
timestamp 1586364061
transform 1 0 53360 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_701
timestamp 1586364061
transform 1 0 54464 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_581
timestamp 1586364061
transform 1 0 54556 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_593
timestamp 1586364061
transform 1 0 55660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_605
timestamp 1586364061
transform 1 0 56764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_617
timestamp 1586364061
transform 1 0 57868 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_702
timestamp 1586364061
transform 1 0 60076 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_629
timestamp 1586364061
transform 1 0 58972 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_642
timestamp 1586364061
transform 1 0 60168 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_654
timestamp 1586364061
transform 1 0 61272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_666
timestamp 1586364061
transform 1 0 62376 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_678
timestamp 1586364061
transform 1 0 63480 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_690
timestamp 1586364061
transform 1 0 64584 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_703
timestamp 1586364061
transform 1 0 65688 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_703
timestamp 1586364061
transform 1 0 65780 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_715
timestamp 1586364061
transform 1 0 66884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_727
timestamp 1586364061
transform 1 0 67988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_739
timestamp 1586364061
transform 1 0 69092 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_704
timestamp 1586364061
transform 1 0 71300 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_751
timestamp 1586364061
transform 1 0 70196 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_764
timestamp 1586364061
transform 1 0 71392 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_776
timestamp 1586364061
transform 1 0 72496 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_788
timestamp 1586364061
transform 1 0 73600 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_800
timestamp 1586364061
transform 1 0 74704 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_812
timestamp 1586364061
transform 1 0 75808 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_705
timestamp 1586364061
transform 1 0 76912 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_825
timestamp 1586364061
transform 1 0 77004 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_837
timestamp 1586364061
transform 1 0 78108 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_849
timestamp 1586364061
transform 1 0 79212 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_861
timestamp 1586364061
transform 1 0 80316 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_873
timestamp 1586364061
transform 1 0 81420 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_706
timestamp 1586364061
transform 1 0 82524 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_886
timestamp 1586364061
transform 1 0 82616 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_898
timestamp 1586364061
transform 1 0 83720 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_910
timestamp 1586364061
transform 1 0 84824 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_922
timestamp 1586364061
transform 1 0 85928 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_934
timestamp 1586364061
transform 1 0 87032 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_707
timestamp 1586364061
transform 1 0 88136 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_947
timestamp 1586364061
transform 1 0 88228 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_959
timestamp 1586364061
transform 1 0 89332 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_971
timestamp 1586364061
transform 1 0 90436 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_983
timestamp 1586364061
transform 1 0 91540 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_995
timestamp 1586364061
transform 1 0 92644 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_708
timestamp 1586364061
transform 1 0 93748 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1008
timestamp 1586364061
transform 1 0 93840 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1020
timestamp 1586364061
transform 1 0 94944 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1032
timestamp 1586364061
transform 1 0 96048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1044
timestamp 1586364061
transform 1 0 97152 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_709
timestamp 1586364061
transform 1 0 99360 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1056
timestamp 1586364061
transform 1 0 98256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1069
timestamp 1586364061
transform 1 0 99452 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1081
timestamp 1586364061
transform 1 0 100556 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1093
timestamp 1586364061
transform 1 0 101660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1105
timestamp 1586364061
transform 1 0 102764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1117
timestamp 1586364061
transform 1 0 103868 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_710
timestamp 1586364061
transform 1 0 104972 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1130
timestamp 1586364061
transform 1 0 105064 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1142
timestamp 1586364061
transform 1 0 106168 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1154
timestamp 1586364061
transform 1 0 107272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1166
timestamp 1586364061
transform 1 0 108376 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_711
timestamp 1586364061
transform 1 0 110584 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1178
timestamp 1586364061
transform 1 0 109480 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1191
timestamp 1586364061
transform 1 0 110676 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1203
timestamp 1586364061
transform 1 0 111780 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1215
timestamp 1586364061
transform 1 0 112884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1227
timestamp 1586364061
transform 1 0 113988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1239
timestamp 1586364061
transform 1 0 115092 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_712
timestamp 1586364061
transform 1 0 116196 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1252
timestamp 1586364061
transform 1 0 116288 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1264
timestamp 1586364061
transform 1 0 117392 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1276
timestamp 1586364061
transform 1 0 118496 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1288
timestamp 1586364061
transform 1 0 119600 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1300
timestamp 1586364061
transform 1 0 120704 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_713
timestamp 1586364061
transform 1 0 121808 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1313
timestamp 1586364061
transform 1 0 121900 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1325
timestamp 1586364061
transform 1 0 123004 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1337
timestamp 1586364061
transform 1 0 124108 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1349
timestamp 1586364061
transform 1 0 125212 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_714
timestamp 1586364061
transform 1 0 127420 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1361
timestamp 1586364061
transform 1 0 126316 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1374
timestamp 1586364061
transform 1 0 127512 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1386
timestamp 1586364061
transform 1 0 128616 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1398
timestamp 1586364061
transform 1 0 129720 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1410
timestamp 1586364061
transform 1 0 130824 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1422
timestamp 1586364061
transform 1 0 131928 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_715
timestamp 1586364061
transform 1 0 133032 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1435
timestamp 1586364061
transform 1 0 133124 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1447
timestamp 1586364061
transform 1 0 134228 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1459
timestamp 1586364061
transform 1 0 135332 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1471
timestamp 1586364061
transform 1 0 136436 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_716
timestamp 1586364061
transform 1 0 138644 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1483
timestamp 1586364061
transform 1 0 137540 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1496
timestamp 1586364061
transform 1 0 138736 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1508
timestamp 1586364061
transform 1 0 139840 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1520
timestamp 1586364061
transform 1 0 140944 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1532
timestamp 1586364061
transform 1 0 142048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1544
timestamp 1586364061
transform 1 0 143152 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_717
timestamp 1586364061
transform 1 0 144256 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1557
timestamp 1586364061
transform 1 0 144348 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1569
timestamp 1586364061
transform 1 0 145452 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1581
timestamp 1586364061
transform 1 0 146556 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1593
timestamp 1586364061
transform 1 0 147660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1605
timestamp 1586364061
transform 1 0 148764 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_718
timestamp 1586364061
transform 1 0 149868 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1618
timestamp 1586364061
transform 1 0 149960 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1630
timestamp 1586364061
transform 1 0 151064 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1642
timestamp 1586364061
transform 1 0 152168 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1654
timestamp 1586364061
transform 1 0 153272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1666
timestamp 1586364061
transform 1 0 154376 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_719
timestamp 1586364061
transform 1 0 155480 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1679
timestamp 1586364061
transform 1 0 155572 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1691
timestamp 1586364061
transform 1 0 156676 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1703
timestamp 1586364061
transform 1 0 157780 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1715
timestamp 1586364061
transform 1 0 158884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1727
timestamp 1586364061
transform 1 0 159988 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_720
timestamp 1586364061
transform 1 0 161092 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1740
timestamp 1586364061
transform 1 0 161184 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1752
timestamp 1586364061
transform 1 0 162288 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1764
timestamp 1586364061
transform 1 0 163392 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1776
timestamp 1586364061
transform 1 0 164496 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_721
timestamp 1586364061
transform 1 0 166704 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1788
timestamp 1586364061
transform 1 0 165600 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1801
timestamp 1586364061
transform 1 0 166796 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1813
timestamp 1586364061
transform 1 0 167900 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1825
timestamp 1586364061
transform 1 0 169004 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1837
timestamp 1586364061
transform 1 0 170108 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1849
timestamp 1586364061
transform 1 0 171212 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_722
timestamp 1586364061
transform 1 0 172316 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1862
timestamp 1586364061
transform 1 0 172408 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1874
timestamp 1586364061
transform 1 0 173512 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1886
timestamp 1586364061
transform 1 0 174616 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1898
timestamp 1586364061
transform 1 0 175720 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_723
timestamp 1586364061
transform 1 0 177928 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1910
timestamp 1586364061
transform 1 0 176824 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1923
timestamp 1586364061
transform 1 0 178020 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1935
timestamp 1586364061
transform 1 0 179124 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1947
timestamp 1586364061
transform 1 0 180228 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1959
timestamp 1586364061
transform 1 0 181332 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1971
timestamp 1586364061
transform 1 0 182436 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_724
timestamp 1586364061
transform 1 0 183540 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_1984
timestamp 1586364061
transform 1 0 183632 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_1996
timestamp 1586364061
transform 1 0 184736 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2008
timestamp 1586364061
transform 1 0 185840 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2020
timestamp 1586364061
transform 1 0 186944 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2032
timestamp 1586364061
transform 1 0 188048 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_725
timestamp 1586364061
transform 1 0 189152 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_2045
timestamp 1586364061
transform 1 0 189244 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2057
timestamp 1586364061
transform 1 0 190348 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2069
timestamp 1586364061
transform 1 0 191452 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2081
timestamp 1586364061
transform 1 0 192556 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2093
timestamp 1586364061
transform 1 0 193660 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_726
timestamp 1586364061
transform 1 0 194764 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_2106
timestamp 1586364061
transform 1 0 194856 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2118
timestamp 1586364061
transform 1 0 195960 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2130
timestamp 1586364061
transform 1 0 197064 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2142
timestamp 1586364061
transform 1 0 198168 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2154
timestamp 1586364061
transform 1 0 199272 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_727
timestamp 1586364061
transform 1 0 200376 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_2167
timestamp 1586364061
transform 1 0 200468 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2179
timestamp 1586364061
transform 1 0 201572 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2191
timestamp 1586364061
transform 1 0 202676 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2203
timestamp 1586364061
transform 1 0 203780 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_728
timestamp 1586364061
transform 1 0 205988 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_2215
timestamp 1586364061
transform 1 0 204884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2228
timestamp 1586364061
transform 1 0 206080 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2240
timestamp 1586364061
transform 1 0 207184 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2252
timestamp 1586364061
transform 1 0 208288 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2264
timestamp 1586364061
transform 1 0 209392 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2276
timestamp 1586364061
transform 1 0 210496 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_729
timestamp 1586364061
transform 1 0 211600 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_2289
timestamp 1586364061
transform 1 0 211692 0 -1 7072
box -38 -48 1142 592
use scs8hd_buf_2  _23_
timestamp 1586364061
transform 1 0 212796 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_2305
timestamp 1586364061
transform 1 0 213164 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2317
timestamp 1586364061
transform 1 0 214268 0 -1 7072
box -38 -48 1142 592
use scs8hd_ebufn_1  logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
timestamp 1586364061
transform 1 0 215556 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_2329
timestamp 1586364061
transform 1 0 215372 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_730
timestamp 1586364061
transform 1 0 217212 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_2339
timestamp 1586364061
transform 1 0 216292 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_2347
timestamp 1586364061
transform 1 0 217028 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_2350
timestamp 1586364061
transform 1 0 217304 0 -1 7072
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 219144 0 -1 7072
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_8_2362
timestamp 1586364061
transform 1 0 218408 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_12  FILLER_8_2381
timestamp 1586364061
transform 1 0 220156 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2393
timestamp 1586364061
transform 1 0 221260 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_8_2405
timestamp 1586364061
transform 1 0 222364 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_731
timestamp 1586364061
transform 1 0 222824 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_2409
timestamp 1586364061
transform 1 0 222732 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_2411
timestamp 1586364061
transform 1 0 222916 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2423
timestamp 1586364061
transform 1 0 224020 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2435
timestamp 1586364061
transform 1 0 225124 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2447
timestamp 1586364061
transform 1 0 226228 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2459
timestamp 1586364061
transform 1 0 227332 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_732
timestamp 1586364061
transform 1 0 228436 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_2472
timestamp 1586364061
transform 1 0 228528 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2484
timestamp 1586364061
transform 1 0 229632 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2496
timestamp 1586364061
transform 1 0 230736 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2508
timestamp 1586364061
transform 1 0 231840 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_733
timestamp 1586364061
transform 1 0 234048 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_2520
timestamp 1586364061
transform 1 0 232944 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2533
timestamp 1586364061
transform 1 0 234140 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2545
timestamp 1586364061
transform 1 0 235244 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2557
timestamp 1586364061
transform 1 0 236348 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2569
timestamp 1586364061
transform 1 0 237452 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2581
timestamp 1586364061
transform 1 0 238556 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_734
timestamp 1586364061
transform 1 0 239660 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_2594
timestamp 1586364061
transform 1 0 239752 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2606
timestamp 1586364061
transform 1 0 240856 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2618
timestamp 1586364061
transform 1 0 241960 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2630
timestamp 1586364061
transform 1 0 243064 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_735
timestamp 1586364061
transform 1 0 245272 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_2642
timestamp 1586364061
transform 1 0 244168 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2655
timestamp 1586364061
transform 1 0 245364 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2667
timestamp 1586364061
transform 1 0 246468 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2679
timestamp 1586364061
transform 1 0 247572 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2691
timestamp 1586364061
transform 1 0 248676 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2703
timestamp 1586364061
transform 1 0 249780 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_736
timestamp 1586364061
transform 1 0 250884 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_2716
timestamp 1586364061
transform 1 0 250976 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2728
timestamp 1586364061
transform 1 0 252080 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2740
timestamp 1586364061
transform 1 0 253184 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2752
timestamp 1586364061
transform 1 0 254288 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2764
timestamp 1586364061
transform 1 0 255392 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_737
timestamp 1586364061
transform 1 0 256496 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_2777
timestamp 1586364061
transform 1 0 256588 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2789
timestamp 1586364061
transform 1 0 257692 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2801
timestamp 1586364061
transform 1 0 258796 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2813
timestamp 1586364061
transform 1 0 259900 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2825
timestamp 1586364061
transform 1 0 261004 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_738
timestamp 1586364061
transform 1 0 262108 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_2838
timestamp 1586364061
transform 1 0 262200 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2850
timestamp 1586364061
transform 1 0 263304 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2862
timestamp 1586364061
transform 1 0 264408 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2874
timestamp 1586364061
transform 1 0 265512 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2886
timestamp 1586364061
transform 1 0 266616 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_739
timestamp 1586364061
transform 1 0 267720 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_2899
timestamp 1586364061
transform 1 0 267812 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2911
timestamp 1586364061
transform 1 0 268916 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2923
timestamp 1586364061
transform 1 0 270020 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2935
timestamp 1586364061
transform 1 0 271124 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_740
timestamp 1586364061
transform 1 0 273332 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_2947
timestamp 1586364061
transform 1 0 272228 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2960
timestamp 1586364061
transform 1 0 273424 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2972
timestamp 1586364061
transform 1 0 274528 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2984
timestamp 1586364061
transform 1 0 275632 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_2996
timestamp 1586364061
transform 1 0 276736 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3008
timestamp 1586364061
transform 1 0 277840 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_741
timestamp 1586364061
transform 1 0 278944 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3021
timestamp 1586364061
transform 1 0 279036 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3033
timestamp 1586364061
transform 1 0 280140 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3045
timestamp 1586364061
transform 1 0 281244 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3057
timestamp 1586364061
transform 1 0 282348 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_742
timestamp 1586364061
transform 1 0 284556 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3069
timestamp 1586364061
transform 1 0 283452 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3082
timestamp 1586364061
transform 1 0 284648 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3094
timestamp 1586364061
transform 1 0 285752 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3106
timestamp 1586364061
transform 1 0 286856 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3118
timestamp 1586364061
transform 1 0 287960 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3130
timestamp 1586364061
transform 1 0 289064 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_743
timestamp 1586364061
transform 1 0 290168 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3143
timestamp 1586364061
transform 1 0 290260 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3155
timestamp 1586364061
transform 1 0 291364 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3167
timestamp 1586364061
transform 1 0 292468 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3179
timestamp 1586364061
transform 1 0 293572 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3191
timestamp 1586364061
transform 1 0 294676 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_744
timestamp 1586364061
transform 1 0 295780 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3204
timestamp 1586364061
transform 1 0 295872 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3216
timestamp 1586364061
transform 1 0 296976 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3228
timestamp 1586364061
transform 1 0 298080 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3240
timestamp 1586364061
transform 1 0 299184 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_745
timestamp 1586364061
transform 1 0 301392 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3252
timestamp 1586364061
transform 1 0 300288 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3265
timestamp 1586364061
transform 1 0 301484 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3277
timestamp 1586364061
transform 1 0 302588 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3289
timestamp 1586364061
transform 1 0 303692 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3301
timestamp 1586364061
transform 1 0 304796 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3313
timestamp 1586364061
transform 1 0 305900 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_746
timestamp 1586364061
transform 1 0 307004 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3326
timestamp 1586364061
transform 1 0 307096 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3338
timestamp 1586364061
transform 1 0 308200 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3350
timestamp 1586364061
transform 1 0 309304 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3362
timestamp 1586364061
transform 1 0 310408 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_747
timestamp 1586364061
transform 1 0 312616 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3374
timestamp 1586364061
transform 1 0 311512 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3387
timestamp 1586364061
transform 1 0 312708 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3399
timestamp 1586364061
transform 1 0 313812 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3411
timestamp 1586364061
transform 1 0 314916 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3423
timestamp 1586364061
transform 1 0 316020 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3435
timestamp 1586364061
transform 1 0 317124 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_748
timestamp 1586364061
transform 1 0 318228 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3448
timestamp 1586364061
transform 1 0 318320 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3460
timestamp 1586364061
transform 1 0 319424 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3472
timestamp 1586364061
transform 1 0 320528 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3484
timestamp 1586364061
transform 1 0 321632 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3496
timestamp 1586364061
transform 1 0 322736 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_749
timestamp 1586364061
transform 1 0 323840 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3509
timestamp 1586364061
transform 1 0 323932 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3521
timestamp 1586364061
transform 1 0 325036 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3533
timestamp 1586364061
transform 1 0 326140 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3545
timestamp 1586364061
transform 1 0 327244 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3557
timestamp 1586364061
transform 1 0 328348 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_750
timestamp 1586364061
transform 1 0 329452 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3570
timestamp 1586364061
transform 1 0 329544 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3582
timestamp 1586364061
transform 1 0 330648 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3594
timestamp 1586364061
transform 1 0 331752 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3606
timestamp 1586364061
transform 1 0 332856 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3618
timestamp 1586364061
transform 1 0 333960 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_751
timestamp 1586364061
transform 1 0 335064 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3631
timestamp 1586364061
transform 1 0 335156 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3643
timestamp 1586364061
transform 1 0 336260 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3655
timestamp 1586364061
transform 1 0 337364 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3667
timestamp 1586364061
transform 1 0 338468 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_752
timestamp 1586364061
transform 1 0 340676 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3679
timestamp 1586364061
transform 1 0 339572 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3692
timestamp 1586364061
transform 1 0 340768 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3704
timestamp 1586364061
transform 1 0 341872 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3716
timestamp 1586364061
transform 1 0 342976 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3728
timestamp 1586364061
transform 1 0 344080 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3740
timestamp 1586364061
transform 1 0 345184 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_753
timestamp 1586364061
transform 1 0 346288 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3753
timestamp 1586364061
transform 1 0 346380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3765
timestamp 1586364061
transform 1 0 347484 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3777
timestamp 1586364061
transform 1 0 348588 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3789
timestamp 1586364061
transform 1 0 349692 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_754
timestamp 1586364061
transform 1 0 351900 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3801
timestamp 1586364061
transform 1 0 350796 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3814
timestamp 1586364061
transform 1 0 351992 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3826
timestamp 1586364061
transform 1 0 353096 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3838
timestamp 1586364061
transform 1 0 354200 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3850
timestamp 1586364061
transform 1 0 355304 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3862
timestamp 1586364061
transform 1 0 356408 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_755
timestamp 1586364061
transform 1 0 357512 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3875
timestamp 1586364061
transform 1 0 357604 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3887
timestamp 1586364061
transform 1 0 358708 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3899
timestamp 1586364061
transform 1 0 359812 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3911
timestamp 1586364061
transform 1 0 360916 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3923
timestamp 1586364061
transform 1 0 362020 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_756
timestamp 1586364061
transform 1 0 363124 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3936
timestamp 1586364061
transform 1 0 363216 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3948
timestamp 1586364061
transform 1 0 364320 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3960
timestamp 1586364061
transform 1 0 365424 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3972
timestamp 1586364061
transform 1 0 366528 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_3984
timestamp 1586364061
transform 1 0 367632 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_757
timestamp 1586364061
transform 1 0 368736 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_3997
timestamp 1586364061
transform 1 0 368828 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4009
timestamp 1586364061
transform 1 0 369932 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4021
timestamp 1586364061
transform 1 0 371036 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4033
timestamp 1586364061
transform 1 0 372140 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4045
timestamp 1586364061
transform 1 0 373244 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_758
timestamp 1586364061
transform 1 0 374348 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_4058
timestamp 1586364061
transform 1 0 374440 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4070
timestamp 1586364061
transform 1 0 375544 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4082
timestamp 1586364061
transform 1 0 376648 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4094
timestamp 1586364061
transform 1 0 377752 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_759
timestamp 1586364061
transform 1 0 379960 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_4106
timestamp 1586364061
transform 1 0 378856 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4119
timestamp 1586364061
transform 1 0 380052 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4131
timestamp 1586364061
transform 1 0 381156 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4143
timestamp 1586364061
transform 1 0 382260 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4155
timestamp 1586364061
transform 1 0 383364 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4167
timestamp 1586364061
transform 1 0 384468 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_760
timestamp 1586364061
transform 1 0 385572 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_4180
timestamp 1586364061
transform 1 0 385664 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4192
timestamp 1586364061
transform 1 0 386768 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4204
timestamp 1586364061
transform 1 0 387872 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4216
timestamp 1586364061
transform 1 0 388976 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_761
timestamp 1586364061
transform 1 0 391184 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_4228
timestamp 1586364061
transform 1 0 390080 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4241
timestamp 1586364061
transform 1 0 391276 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4253
timestamp 1586364061
transform 1 0 392380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4265
timestamp 1586364061
transform 1 0 393484 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4277
timestamp 1586364061
transform 1 0 394588 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4289
timestamp 1586364061
transform 1 0 395692 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_762
timestamp 1586364061
transform 1 0 396796 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_4302
timestamp 1586364061
transform 1 0 396888 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4314
timestamp 1586364061
transform 1 0 397992 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4326
timestamp 1586364061
transform 1 0 399096 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4338
timestamp 1586364061
transform 1 0 400200 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4350
timestamp 1586364061
transform 1 0 401304 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_763
timestamp 1586364061
transform 1 0 402408 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_4363
timestamp 1586364061
transform 1 0 402500 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4375
timestamp 1586364061
transform 1 0 403604 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4387
timestamp 1586364061
transform 1 0 404708 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4399
timestamp 1586364061
transform 1 0 405812 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_764
timestamp 1586364061
transform 1 0 408020 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_4411
timestamp 1586364061
transform 1 0 406916 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4424
timestamp 1586364061
transform 1 0 408112 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4436
timestamp 1586364061
transform 1 0 409216 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4448
timestamp 1586364061
transform 1 0 410320 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4460
timestamp 1586364061
transform 1 0 411424 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4472
timestamp 1586364061
transform 1 0 412528 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_765
timestamp 1586364061
transform 1 0 413632 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_4485
timestamp 1586364061
transform 1 0 413724 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4497
timestamp 1586364061
transform 1 0 414828 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4509
timestamp 1586364061
transform 1 0 415932 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4521
timestamp 1586364061
transform 1 0 417036 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_766
timestamp 1586364061
transform 1 0 419244 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_4533
timestamp 1586364061
transform 1 0 418140 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4546
timestamp 1586364061
transform 1 0 419336 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_4558
timestamp 1586364061
transform 1 0 420440 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 422832 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_4570
timestamp 1586364061
transform 1 0 421544 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_4578
timestamp 1586364061
transform 1 0 422280 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_767
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_9_32
timestamp 1586364061
transform 1 0 4048 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_44
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_768
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_56
timestamp 1586364061
transform 1 0 6256 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_63
timestamp 1586364061
transform 1 0 6900 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_75
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_87
timestamp 1586364061
transform 1 0 9108 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_769
timestamp 1586364061
transform 1 0 9660 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_94
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_106
timestamp 1586364061
transform 1 0 10856 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_770
timestamp 1586364061
transform 1 0 12512 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_125
timestamp 1586364061
transform 1 0 12604 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_137
timestamp 1586364061
transform 1 0 13708 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_771
timestamp 1586364061
transform 1 0 15364 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_149
timestamp 1586364061
transform 1 0 14812 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_156
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_168
timestamp 1586364061
transform 1 0 16560 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_772
timestamp 1586364061
transform 1 0 18216 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_180
timestamp 1586364061
transform 1 0 17664 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_187
timestamp 1586364061
transform 1 0 18308 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_199
timestamp 1586364061
transform 1 0 19412 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_211
timestamp 1586364061
transform 1 0 20516 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_773
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_218
timestamp 1586364061
transform 1 0 21160 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_230
timestamp 1586364061
transform 1 0 22264 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_774
timestamp 1586364061
transform 1 0 23920 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_242
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_249
timestamp 1586364061
transform 1 0 24012 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_261
timestamp 1586364061
transform 1 0 25116 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_775
timestamp 1586364061
transform 1 0 26772 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_273
timestamp 1586364061
transform 1 0 26220 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_280
timestamp 1586364061
transform 1 0 26864 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_292
timestamp 1586364061
transform 1 0 27968 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_776
timestamp 1586364061
transform 1 0 29624 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_304
timestamp 1586364061
transform 1 0 29072 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_311
timestamp 1586364061
transform 1 0 29716 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_323
timestamp 1586364061
transform 1 0 30820 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_335
timestamp 1586364061
transform 1 0 31924 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_777
timestamp 1586364061
transform 1 0 32476 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_342
timestamp 1586364061
transform 1 0 32568 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_354
timestamp 1586364061
transform 1 0 33672 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_778
timestamp 1586364061
transform 1 0 35328 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_366
timestamp 1586364061
transform 1 0 34776 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_373
timestamp 1586364061
transform 1 0 35420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_385
timestamp 1586364061
transform 1 0 36524 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_779
timestamp 1586364061
transform 1 0 38180 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_397
timestamp 1586364061
transform 1 0 37628 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_404
timestamp 1586364061
transform 1 0 38272 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_416
timestamp 1586364061
transform 1 0 39376 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_428
timestamp 1586364061
transform 1 0 40480 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_780
timestamp 1586364061
transform 1 0 41032 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_435
timestamp 1586364061
transform 1 0 41124 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_447
timestamp 1586364061
transform 1 0 42228 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_459
timestamp 1586364061
transform 1 0 43332 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_781
timestamp 1586364061
transform 1 0 43884 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_466
timestamp 1586364061
transform 1 0 43976 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_478
timestamp 1586364061
transform 1 0 45080 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_782
timestamp 1586364061
transform 1 0 46736 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_490
timestamp 1586364061
transform 1 0 46184 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_497
timestamp 1586364061
transform 1 0 46828 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_509
timestamp 1586364061
transform 1 0 47932 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_783
timestamp 1586364061
transform 1 0 49588 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_521
timestamp 1586364061
transform 1 0 49036 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_528
timestamp 1586364061
transform 1 0 49680 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_540
timestamp 1586364061
transform 1 0 50784 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_552
timestamp 1586364061
transform 1 0 51888 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_784
timestamp 1586364061
transform 1 0 52440 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_559
timestamp 1586364061
transform 1 0 52532 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_571
timestamp 1586364061
transform 1 0 53636 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_583
timestamp 1586364061
transform 1 0 54740 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_785
timestamp 1586364061
transform 1 0 55292 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_590
timestamp 1586364061
transform 1 0 55384 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_602
timestamp 1586364061
transform 1 0 56488 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_786
timestamp 1586364061
transform 1 0 58144 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_614
timestamp 1586364061
transform 1 0 57592 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_621
timestamp 1586364061
transform 1 0 58236 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_633
timestamp 1586364061
transform 1 0 59340 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_787
timestamp 1586364061
transform 1 0 60996 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_645
timestamp 1586364061
transform 1 0 60444 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_652
timestamp 1586364061
transform 1 0 61088 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_664
timestamp 1586364061
transform 1 0 62192 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_676
timestamp 1586364061
transform 1 0 63296 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_788
timestamp 1586364061
transform 1 0 63848 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_683
timestamp 1586364061
transform 1 0 63940 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_695
timestamp 1586364061
transform 1 0 65044 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_789
timestamp 1586364061
transform 1 0 66700 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_707
timestamp 1586364061
transform 1 0 66148 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_714
timestamp 1586364061
transform 1 0 66792 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_726
timestamp 1586364061
transform 1 0 67896 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_790
timestamp 1586364061
transform 1 0 69552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_738
timestamp 1586364061
transform 1 0 69000 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_745
timestamp 1586364061
transform 1 0 69644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_757
timestamp 1586364061
transform 1 0 70748 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_791
timestamp 1586364061
transform 1 0 72404 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_769
timestamp 1586364061
transform 1 0 71852 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_776
timestamp 1586364061
transform 1 0 72496 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_788
timestamp 1586364061
transform 1 0 73600 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_800
timestamp 1586364061
transform 1 0 74704 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_792
timestamp 1586364061
transform 1 0 75256 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_807
timestamp 1586364061
transform 1 0 75348 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_819
timestamp 1586364061
transform 1 0 76452 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_793
timestamp 1586364061
transform 1 0 78108 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_831
timestamp 1586364061
transform 1 0 77556 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_838
timestamp 1586364061
transform 1 0 78200 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_850
timestamp 1586364061
transform 1 0 79304 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_794
timestamp 1586364061
transform 1 0 80960 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_862
timestamp 1586364061
transform 1 0 80408 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_869
timestamp 1586364061
transform 1 0 81052 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_881
timestamp 1586364061
transform 1 0 82156 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_795
timestamp 1586364061
transform 1 0 83812 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_893
timestamp 1586364061
transform 1 0 83260 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_900
timestamp 1586364061
transform 1 0 83904 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_912
timestamp 1586364061
transform 1 0 85008 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_924
timestamp 1586364061
transform 1 0 86112 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_796
timestamp 1586364061
transform 1 0 86664 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_931
timestamp 1586364061
transform 1 0 86756 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_943
timestamp 1586364061
transform 1 0 87860 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_797
timestamp 1586364061
transform 1 0 89516 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_955
timestamp 1586364061
transform 1 0 88964 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_962
timestamp 1586364061
transform 1 0 89608 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_974
timestamp 1586364061
transform 1 0 90712 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_798
timestamp 1586364061
transform 1 0 92368 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_986
timestamp 1586364061
transform 1 0 91816 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_993
timestamp 1586364061
transform 1 0 92460 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1005
timestamp 1586364061
transform 1 0 93564 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_799
timestamp 1586364061
transform 1 0 95220 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1017
timestamp 1586364061
transform 1 0 94668 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1024
timestamp 1586364061
transform 1 0 95312 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1036
timestamp 1586364061
transform 1 0 96416 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_1048
timestamp 1586364061
transform 1 0 97520 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_800
timestamp 1586364061
transform 1 0 98072 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_1055
timestamp 1586364061
transform 1 0 98164 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1067
timestamp 1586364061
transform 1 0 99268 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_801
timestamp 1586364061
transform 1 0 100924 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1079
timestamp 1586364061
transform 1 0 100372 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1086
timestamp 1586364061
transform 1 0 101016 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1098
timestamp 1586364061
transform 1 0 102120 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_802
timestamp 1586364061
transform 1 0 103776 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1110
timestamp 1586364061
transform 1 0 103224 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1117
timestamp 1586364061
transform 1 0 103868 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1129
timestamp 1586364061
transform 1 0 104972 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_1141
timestamp 1586364061
transform 1 0 106076 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_803
timestamp 1586364061
transform 1 0 106628 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_1148
timestamp 1586364061
transform 1 0 106720 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1160
timestamp 1586364061
transform 1 0 107824 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_1172
timestamp 1586364061
transform 1 0 108928 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_804
timestamp 1586364061
transform 1 0 109480 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_1179
timestamp 1586364061
transform 1 0 109572 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1191
timestamp 1586364061
transform 1 0 110676 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_805
timestamp 1586364061
transform 1 0 112332 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1203
timestamp 1586364061
transform 1 0 111780 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1210
timestamp 1586364061
transform 1 0 112424 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1222
timestamp 1586364061
transform 1 0 113528 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_806
timestamp 1586364061
transform 1 0 115184 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1234
timestamp 1586364061
transform 1 0 114632 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1241
timestamp 1586364061
transform 1 0 115276 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1253
timestamp 1586364061
transform 1 0 116380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_1265
timestamp 1586364061
transform 1 0 117484 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_807
timestamp 1586364061
transform 1 0 118036 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_1272
timestamp 1586364061
transform 1 0 118128 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1284
timestamp 1586364061
transform 1 0 119232 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_808
timestamp 1586364061
transform 1 0 120888 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1296
timestamp 1586364061
transform 1 0 120336 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1303
timestamp 1586364061
transform 1 0 120980 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1315
timestamp 1586364061
transform 1 0 122084 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_809
timestamp 1586364061
transform 1 0 123740 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1327
timestamp 1586364061
transform 1 0 123188 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1334
timestamp 1586364061
transform 1 0 123832 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1346
timestamp 1586364061
transform 1 0 124936 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_810
timestamp 1586364061
transform 1 0 126592 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1358
timestamp 1586364061
transform 1 0 126040 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1365
timestamp 1586364061
transform 1 0 126684 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1377
timestamp 1586364061
transform 1 0 127788 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_1389
timestamp 1586364061
transform 1 0 128892 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_811
timestamp 1586364061
transform 1 0 129444 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_1396
timestamp 1586364061
transform 1 0 129536 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1408
timestamp 1586364061
transform 1 0 130640 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_812
timestamp 1586364061
transform 1 0 132296 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1420
timestamp 1586364061
transform 1 0 131744 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1427
timestamp 1586364061
transform 1 0 132388 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1439
timestamp 1586364061
transform 1 0 133492 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_813
timestamp 1586364061
transform 1 0 135148 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1451
timestamp 1586364061
transform 1 0 134596 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1458
timestamp 1586364061
transform 1 0 135240 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1470
timestamp 1586364061
transform 1 0 136344 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_814
timestamp 1586364061
transform 1 0 138000 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1482
timestamp 1586364061
transform 1 0 137448 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1489
timestamp 1586364061
transform 1 0 138092 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1501
timestamp 1586364061
transform 1 0 139196 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_1513
timestamp 1586364061
transform 1 0 140300 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_815
timestamp 1586364061
transform 1 0 140852 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_1520
timestamp 1586364061
transform 1 0 140944 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1532
timestamp 1586364061
transform 1 0 142048 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_816
timestamp 1586364061
transform 1 0 143704 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1544
timestamp 1586364061
transform 1 0 143152 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1551
timestamp 1586364061
transform 1 0 143796 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1563
timestamp 1586364061
transform 1 0 144900 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_817
timestamp 1586364061
transform 1 0 146556 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1575
timestamp 1586364061
transform 1 0 146004 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1582
timestamp 1586364061
transform 1 0 146648 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1594
timestamp 1586364061
transform 1 0 147752 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_818
timestamp 1586364061
transform 1 0 149408 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1606
timestamp 1586364061
transform 1 0 148856 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1613
timestamp 1586364061
transform 1 0 149500 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1625
timestamp 1586364061
transform 1 0 150604 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_1637
timestamp 1586364061
transform 1 0 151708 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_819
timestamp 1586364061
transform 1 0 152260 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_1644
timestamp 1586364061
transform 1 0 152352 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1656
timestamp 1586364061
transform 1 0 153456 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_820
timestamp 1586364061
transform 1 0 155112 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1668
timestamp 1586364061
transform 1 0 154560 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1675
timestamp 1586364061
transform 1 0 155204 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1687
timestamp 1586364061
transform 1 0 156308 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_821
timestamp 1586364061
transform 1 0 157964 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1699
timestamp 1586364061
transform 1 0 157412 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1706
timestamp 1586364061
transform 1 0 158056 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1718
timestamp 1586364061
transform 1 0 159160 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_1730
timestamp 1586364061
transform 1 0 160264 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_822
timestamp 1586364061
transform 1 0 160816 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_1737
timestamp 1586364061
transform 1 0 160908 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1749
timestamp 1586364061
transform 1 0 162012 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_1761
timestamp 1586364061
transform 1 0 163116 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_823
timestamp 1586364061
transform 1 0 163668 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_1768
timestamp 1586364061
transform 1 0 163760 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1780
timestamp 1586364061
transform 1 0 164864 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_824
timestamp 1586364061
transform 1 0 166520 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1792
timestamp 1586364061
transform 1 0 165968 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1799
timestamp 1586364061
transform 1 0 166612 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1811
timestamp 1586364061
transform 1 0 167716 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_825
timestamp 1586364061
transform 1 0 169372 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1823
timestamp 1586364061
transform 1 0 168820 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1830
timestamp 1586364061
transform 1 0 169464 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1842
timestamp 1586364061
transform 1 0 170568 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_1854
timestamp 1586364061
transform 1 0 171672 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_826
timestamp 1586364061
transform 1 0 172224 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_1861
timestamp 1586364061
transform 1 0 172316 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1873
timestamp 1586364061
transform 1 0 173420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_1885
timestamp 1586364061
transform 1 0 174524 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_827
timestamp 1586364061
transform 1 0 175076 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_1892
timestamp 1586364061
transform 1 0 175168 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1904
timestamp 1586364061
transform 1 0 176272 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_828
timestamp 1586364061
transform 1 0 177928 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1916
timestamp 1586364061
transform 1 0 177376 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1923
timestamp 1586364061
transform 1 0 178020 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1935
timestamp 1586364061
transform 1 0 179124 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_829
timestamp 1586364061
transform 1 0 180780 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_1947
timestamp 1586364061
transform 1 0 180228 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_1954
timestamp 1586364061
transform 1 0 180872 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1966
timestamp 1586364061
transform 1 0 181976 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_1978
timestamp 1586364061
transform 1 0 183080 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_830
timestamp 1586364061
transform 1 0 183632 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_1985
timestamp 1586364061
transform 1 0 183724 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_1997
timestamp 1586364061
transform 1 0 184828 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_831
timestamp 1586364061
transform 1 0 186484 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2009
timestamp 1586364061
transform 1 0 185932 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2016
timestamp 1586364061
transform 1 0 186576 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2028
timestamp 1586364061
transform 1 0 187680 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_832
timestamp 1586364061
transform 1 0 189336 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2040
timestamp 1586364061
transform 1 0 188784 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2047
timestamp 1586364061
transform 1 0 189428 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2059
timestamp 1586364061
transform 1 0 190532 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_833
timestamp 1586364061
transform 1 0 192188 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2071
timestamp 1586364061
transform 1 0 191636 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2078
timestamp 1586364061
transform 1 0 192280 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2090
timestamp 1586364061
transform 1 0 193384 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_2102
timestamp 1586364061
transform 1 0 194488 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_834
timestamp 1586364061
transform 1 0 195040 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_2109
timestamp 1586364061
transform 1 0 195132 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2121
timestamp 1586364061
transform 1 0 196236 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_835
timestamp 1586364061
transform 1 0 197892 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2133
timestamp 1586364061
transform 1 0 197340 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2140
timestamp 1586364061
transform 1 0 197984 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2152
timestamp 1586364061
transform 1 0 199088 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_836
timestamp 1586364061
transform 1 0 200744 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2164
timestamp 1586364061
transform 1 0 200192 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2171
timestamp 1586364061
transform 1 0 200836 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2183
timestamp 1586364061
transform 1 0 201940 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_837
timestamp 1586364061
transform 1 0 203596 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2195
timestamp 1586364061
transform 1 0 203044 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2202
timestamp 1586364061
transform 1 0 203688 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2214
timestamp 1586364061
transform 1 0 204792 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_2226
timestamp 1586364061
transform 1 0 205896 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_838
timestamp 1586364061
transform 1 0 206448 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_2233
timestamp 1586364061
transform 1 0 206540 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2245
timestamp 1586364061
transform 1 0 207644 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_839
timestamp 1586364061
transform 1 0 209300 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2257
timestamp 1586364061
transform 1 0 208748 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2264
timestamp 1586364061
transform 1 0 209392 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2276
timestamp 1586364061
transform 1 0 210496 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_840
timestamp 1586364061
transform 1 0 212152 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2288
timestamp 1586364061
transform 1 0 211600 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2295
timestamp 1586364061
transform 1 0 212244 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2307
timestamp 1586364061
transform 1 0 213348 0 1 7072
box -38 -48 1142 592
use scs8hd_buf_2  _22_
timestamp 1586364061
transform 1 0 215096 0 1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_841
timestamp 1586364061
transform 1 0 215004 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__22__A
timestamp 1586364061
transform 1 0 215648 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_2319
timestamp 1586364061
transform 1 0 214452 0 1 7072
box -38 -48 590 592
use scs8hd_fill_2  FILLER_9_2330
timestamp 1586364061
transform 1 0 215464 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_2334
timestamp 1586364061
transform 1 0 215832 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_2346
timestamp 1586364061
transform 1 0 216936 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_2354
timestamp 1586364061
transform 1 0 217672 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_842
timestamp 1586364061
transform 1 0 217856 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_2357
timestamp 1586364061
transform 1 0 217948 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2369
timestamp 1586364061
transform 1 0 219052 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_843
timestamp 1586364061
transform 1 0 220708 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2381
timestamp 1586364061
transform 1 0 220156 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2388
timestamp 1586364061
transform 1 0 220800 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2400
timestamp 1586364061
transform 1 0 221904 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_844
timestamp 1586364061
transform 1 0 223560 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2412
timestamp 1586364061
transform 1 0 223008 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2419
timestamp 1586364061
transform 1 0 223652 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2431
timestamp 1586364061
transform 1 0 224756 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_2443
timestamp 1586364061
transform 1 0 225860 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_845
timestamp 1586364061
transform 1 0 226412 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_2450
timestamp 1586364061
transform 1 0 226504 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2462
timestamp 1586364061
transform 1 0 227608 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_2474
timestamp 1586364061
transform 1 0 228712 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_846
timestamp 1586364061
transform 1 0 229264 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_2481
timestamp 1586364061
transform 1 0 229356 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2493
timestamp 1586364061
transform 1 0 230460 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_847
timestamp 1586364061
transform 1 0 232116 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2505
timestamp 1586364061
transform 1 0 231564 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2512
timestamp 1586364061
transform 1 0 232208 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2524
timestamp 1586364061
transform 1 0 233312 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_848
timestamp 1586364061
transform 1 0 234968 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2536
timestamp 1586364061
transform 1 0 234416 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2543
timestamp 1586364061
transform 1 0 235060 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2555
timestamp 1586364061
transform 1 0 236164 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_2567
timestamp 1586364061
transform 1 0 237268 0 1 7072
box -38 -48 590 592
use scs8hd_buf_2  _16_
timestamp 1586364061
transform 1 0 237912 0 1 7072
box -38 -48 406 592
use scs8hd_buf_2  _19_
timestamp 1586364061
transform 1 0 239016 0 1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_849
timestamp 1586364061
transform 1 0 237820 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__16__A
timestamp 1586364061
transform 1 0 238464 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_2578
timestamp 1586364061
transform 1 0 238280 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_2582
timestamp 1586364061
transform 1 0 238648 0 1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_850
timestamp 1586364061
transform 1 0 240672 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__19__A
timestamp 1586364061
transform 1 0 239568 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_2590
timestamp 1586364061
transform 1 0 239384 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_2594
timestamp 1586364061
transform 1 0 239752 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_2602
timestamp 1586364061
transform 1 0 240488 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_2605
timestamp 1586364061
transform 1 0 240764 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2617
timestamp 1586364061
transform 1 0 241868 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_851
timestamp 1586364061
transform 1 0 243524 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2629
timestamp 1586364061
transform 1 0 242972 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2636
timestamp 1586364061
transform 1 0 243616 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2648
timestamp 1586364061
transform 1 0 244720 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_852
timestamp 1586364061
transform 1 0 246376 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2660
timestamp 1586364061
transform 1 0 245824 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2667
timestamp 1586364061
transform 1 0 246468 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2679
timestamp 1586364061
transform 1 0 247572 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_2691
timestamp 1586364061
transform 1 0 248676 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_853
timestamp 1586364061
transform 1 0 249228 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_2698
timestamp 1586364061
transform 1 0 249320 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2710
timestamp 1586364061
transform 1 0 250424 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_854
timestamp 1586364061
transform 1 0 252080 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2722
timestamp 1586364061
transform 1 0 251528 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2729
timestamp 1586364061
transform 1 0 252172 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2741
timestamp 1586364061
transform 1 0 253276 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_855
timestamp 1586364061
transform 1 0 254932 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2753
timestamp 1586364061
transform 1 0 254380 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2760
timestamp 1586364061
transform 1 0 255024 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2772
timestamp 1586364061
transform 1 0 256128 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_856
timestamp 1586364061
transform 1 0 257784 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2784
timestamp 1586364061
transform 1 0 257232 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2791
timestamp 1586364061
transform 1 0 257876 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2803
timestamp 1586364061
transform 1 0 258980 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_2815
timestamp 1586364061
transform 1 0 260084 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_857
timestamp 1586364061
transform 1 0 260636 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_2822
timestamp 1586364061
transform 1 0 260728 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2834
timestamp 1586364061
transform 1 0 261832 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_858
timestamp 1586364061
transform 1 0 263488 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2846
timestamp 1586364061
transform 1 0 262936 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2853
timestamp 1586364061
transform 1 0 263580 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2865
timestamp 1586364061
transform 1 0 264684 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_859
timestamp 1586364061
transform 1 0 266340 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2877
timestamp 1586364061
transform 1 0 265788 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2884
timestamp 1586364061
transform 1 0 266432 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2896
timestamp 1586364061
transform 1 0 267536 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_860
timestamp 1586364061
transform 1 0 269192 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2908
timestamp 1586364061
transform 1 0 268640 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2915
timestamp 1586364061
transform 1 0 269284 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2927
timestamp 1586364061
transform 1 0 270388 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_2939
timestamp 1586364061
transform 1 0 271492 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_861
timestamp 1586364061
transform 1 0 272044 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_2946
timestamp 1586364061
transform 1 0 272136 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2958
timestamp 1586364061
transform 1 0 273240 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_862
timestamp 1586364061
transform 1 0 274896 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_2970
timestamp 1586364061
transform 1 0 274344 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_2977
timestamp 1586364061
transform 1 0 274988 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_2989
timestamp 1586364061
transform 1 0 276092 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_863
timestamp 1586364061
transform 1 0 277748 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3001
timestamp 1586364061
transform 1 0 277196 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3008
timestamp 1586364061
transform 1 0 277840 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3020
timestamp 1586364061
transform 1 0 278944 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_3032
timestamp 1586364061
transform 1 0 280048 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_864
timestamp 1586364061
transform 1 0 280600 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_3039
timestamp 1586364061
transform 1 0 280692 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3051
timestamp 1586364061
transform 1 0 281796 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_3063
timestamp 1586364061
transform 1 0 282900 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_865
timestamp 1586364061
transform 1 0 283452 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_3070
timestamp 1586364061
transform 1 0 283544 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3082
timestamp 1586364061
transform 1 0 284648 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_866
timestamp 1586364061
transform 1 0 286304 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3094
timestamp 1586364061
transform 1 0 285752 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3101
timestamp 1586364061
transform 1 0 286396 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3113
timestamp 1586364061
transform 1 0 287500 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_867
timestamp 1586364061
transform 1 0 289156 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3125
timestamp 1586364061
transform 1 0 288604 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3132
timestamp 1586364061
transform 1 0 289248 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3144
timestamp 1586364061
transform 1 0 290352 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_3156
timestamp 1586364061
transform 1 0 291456 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_868
timestamp 1586364061
transform 1 0 292008 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_3163
timestamp 1586364061
transform 1 0 292100 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3175
timestamp 1586364061
transform 1 0 293204 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_3187
timestamp 1586364061
transform 1 0 294308 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_869
timestamp 1586364061
transform 1 0 294860 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_3194
timestamp 1586364061
transform 1 0 294952 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3206
timestamp 1586364061
transform 1 0 296056 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_870
timestamp 1586364061
transform 1 0 297712 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3218
timestamp 1586364061
transform 1 0 297160 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3225
timestamp 1586364061
transform 1 0 297804 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3237
timestamp 1586364061
transform 1 0 298908 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_871
timestamp 1586364061
transform 1 0 300564 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3249
timestamp 1586364061
transform 1 0 300012 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3256
timestamp 1586364061
transform 1 0 300656 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3268
timestamp 1586364061
transform 1 0 301760 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_3280
timestamp 1586364061
transform 1 0 302864 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_872
timestamp 1586364061
transform 1 0 303416 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_3287
timestamp 1586364061
transform 1 0 303508 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3299
timestamp 1586364061
transform 1 0 304612 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_873
timestamp 1586364061
transform 1 0 306268 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3311
timestamp 1586364061
transform 1 0 305716 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3318
timestamp 1586364061
transform 1 0 306360 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3330
timestamp 1586364061
transform 1 0 307464 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_874
timestamp 1586364061
transform 1 0 309120 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3342
timestamp 1586364061
transform 1 0 308568 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3349
timestamp 1586364061
transform 1 0 309212 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3361
timestamp 1586364061
transform 1 0 310316 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_875
timestamp 1586364061
transform 1 0 311972 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3373
timestamp 1586364061
transform 1 0 311420 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3380
timestamp 1586364061
transform 1 0 312064 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3392
timestamp 1586364061
transform 1 0 313168 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_3404
timestamp 1586364061
transform 1 0 314272 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_876
timestamp 1586364061
transform 1 0 314824 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_3411
timestamp 1586364061
transform 1 0 314916 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3423
timestamp 1586364061
transform 1 0 316020 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_877
timestamp 1586364061
transform 1 0 317676 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3435
timestamp 1586364061
transform 1 0 317124 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3442
timestamp 1586364061
transform 1 0 317768 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3454
timestamp 1586364061
transform 1 0 318872 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_878
timestamp 1586364061
transform 1 0 320528 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3466
timestamp 1586364061
transform 1 0 319976 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3473
timestamp 1586364061
transform 1 0 320620 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3485
timestamp 1586364061
transform 1 0 321724 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_879
timestamp 1586364061
transform 1 0 323380 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3497
timestamp 1586364061
transform 1 0 322828 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3504
timestamp 1586364061
transform 1 0 323472 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3516
timestamp 1586364061
transform 1 0 324576 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_3528
timestamp 1586364061
transform 1 0 325680 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_880
timestamp 1586364061
transform 1 0 326232 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_3535
timestamp 1586364061
transform 1 0 326324 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3547
timestamp 1586364061
transform 1 0 327428 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_881
timestamp 1586364061
transform 1 0 329084 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3559
timestamp 1586364061
transform 1 0 328532 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3566
timestamp 1586364061
transform 1 0 329176 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3578
timestamp 1586364061
transform 1 0 330280 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_882
timestamp 1586364061
transform 1 0 331936 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3590
timestamp 1586364061
transform 1 0 331384 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3597
timestamp 1586364061
transform 1 0 332028 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3609
timestamp 1586364061
transform 1 0 333132 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_883
timestamp 1586364061
transform 1 0 334788 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3621
timestamp 1586364061
transform 1 0 334236 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3628
timestamp 1586364061
transform 1 0 334880 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3640
timestamp 1586364061
transform 1 0 335984 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_3652
timestamp 1586364061
transform 1 0 337088 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_884
timestamp 1586364061
transform 1 0 337640 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_3659
timestamp 1586364061
transform 1 0 337732 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3671
timestamp 1586364061
transform 1 0 338836 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_885
timestamp 1586364061
transform 1 0 340492 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3683
timestamp 1586364061
transform 1 0 339940 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3690
timestamp 1586364061
transform 1 0 340584 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3702
timestamp 1586364061
transform 1 0 341688 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_886
timestamp 1586364061
transform 1 0 343344 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3714
timestamp 1586364061
transform 1 0 342792 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3721
timestamp 1586364061
transform 1 0 343436 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3733
timestamp 1586364061
transform 1 0 344540 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_3745
timestamp 1586364061
transform 1 0 345644 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_887
timestamp 1586364061
transform 1 0 346196 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_3752
timestamp 1586364061
transform 1 0 346288 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3764
timestamp 1586364061
transform 1 0 347392 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_3776
timestamp 1586364061
transform 1 0 348496 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_888
timestamp 1586364061
transform 1 0 349048 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_3783
timestamp 1586364061
transform 1 0 349140 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3795
timestamp 1586364061
transform 1 0 350244 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_889
timestamp 1586364061
transform 1 0 351900 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3807
timestamp 1586364061
transform 1 0 351348 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3814
timestamp 1586364061
transform 1 0 351992 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3826
timestamp 1586364061
transform 1 0 353096 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_890
timestamp 1586364061
transform 1 0 354752 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3838
timestamp 1586364061
transform 1 0 354200 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3845
timestamp 1586364061
transform 1 0 354844 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3857
timestamp 1586364061
transform 1 0 355948 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_3869
timestamp 1586364061
transform 1 0 357052 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_891
timestamp 1586364061
transform 1 0 357604 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_3876
timestamp 1586364061
transform 1 0 357696 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3888
timestamp 1586364061
transform 1 0 358800 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_892
timestamp 1586364061
transform 1 0 360456 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3900
timestamp 1586364061
transform 1 0 359904 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3907
timestamp 1586364061
transform 1 0 360548 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3919
timestamp 1586364061
transform 1 0 361652 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_893
timestamp 1586364061
transform 1 0 363308 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3931
timestamp 1586364061
transform 1 0 362756 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3938
timestamp 1586364061
transform 1 0 363400 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3950
timestamp 1586364061
transform 1 0 364504 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_894
timestamp 1586364061
transform 1 0 366160 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_3962
timestamp 1586364061
transform 1 0 365608 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_3969
timestamp 1586364061
transform 1 0 366252 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_3981
timestamp 1586364061
transform 1 0 367356 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_3993
timestamp 1586364061
transform 1 0 368460 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_895
timestamp 1586364061
transform 1 0 369012 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_4000
timestamp 1586364061
transform 1 0 369104 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4012
timestamp 1586364061
transform 1 0 370208 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_896
timestamp 1586364061
transform 1 0 371864 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_4024
timestamp 1586364061
transform 1 0 371312 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_4031
timestamp 1586364061
transform 1 0 371956 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4043
timestamp 1586364061
transform 1 0 373060 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_897
timestamp 1586364061
transform 1 0 374716 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_4055
timestamp 1586364061
transform 1 0 374164 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_4062
timestamp 1586364061
transform 1 0 374808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4074
timestamp 1586364061
transform 1 0 375912 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_898
timestamp 1586364061
transform 1 0 377568 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_4086
timestamp 1586364061
transform 1 0 377016 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_4093
timestamp 1586364061
transform 1 0 377660 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4105
timestamp 1586364061
transform 1 0 378764 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_4117
timestamp 1586364061
transform 1 0 379868 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_899
timestamp 1586364061
transform 1 0 380420 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_4124
timestamp 1586364061
transform 1 0 380512 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4136
timestamp 1586364061
transform 1 0 381616 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_900
timestamp 1586364061
transform 1 0 383272 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_4148
timestamp 1586364061
transform 1 0 382720 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_4155
timestamp 1586364061
transform 1 0 383364 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4167
timestamp 1586364061
transform 1 0 384468 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_901
timestamp 1586364061
transform 1 0 386124 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_4179
timestamp 1586364061
transform 1 0 385572 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_4186
timestamp 1586364061
transform 1 0 386216 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4198
timestamp 1586364061
transform 1 0 387320 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_902
timestamp 1586364061
transform 1 0 388976 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_4210
timestamp 1586364061
transform 1 0 388424 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_4217
timestamp 1586364061
transform 1 0 389068 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4229
timestamp 1586364061
transform 1 0 390172 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_4241
timestamp 1586364061
transform 1 0 391276 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_903
timestamp 1586364061
transform 1 0 391828 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_4248
timestamp 1586364061
transform 1 0 391920 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4260
timestamp 1586364061
transform 1 0 393024 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_904
timestamp 1586364061
transform 1 0 394680 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_4272
timestamp 1586364061
transform 1 0 394128 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_4279
timestamp 1586364061
transform 1 0 394772 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4291
timestamp 1586364061
transform 1 0 395876 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_905
timestamp 1586364061
transform 1 0 397532 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_4303
timestamp 1586364061
transform 1 0 396980 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_4310
timestamp 1586364061
transform 1 0 397624 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4322
timestamp 1586364061
transform 1 0 398728 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_4334
timestamp 1586364061
transform 1 0 399832 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_906
timestamp 1586364061
transform 1 0 400384 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_4341
timestamp 1586364061
transform 1 0 400476 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4353
timestamp 1586364061
transform 1 0 401580 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_4365
timestamp 1586364061
transform 1 0 402684 0 1 7072
box -38 -48 590 592
use scs8hd_buf_2  _18_
timestamp 1586364061
transform 1 0 404156 0 1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_907
timestamp 1586364061
transform 1 0 403236 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__18__A
timestamp 1586364061
transform 1 0 404708 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_4372
timestamp 1586364061
transform 1 0 403328 0 1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_9_4380
timestamp 1586364061
transform 1 0 404064 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_4385
timestamp 1586364061
transform 1 0 404524 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_908
timestamp 1586364061
transform 1 0 406088 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_4389
timestamp 1586364061
transform 1 0 404892 0 1 7072
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_9_4401
timestamp 1586364061
transform 1 0 405996 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_4403
timestamp 1586364061
transform 1 0 406180 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4415
timestamp 1586364061
transform 1 0 407284 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_909
timestamp 1586364061
transform 1 0 408940 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_4427
timestamp 1586364061
transform 1 0 408388 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_4434
timestamp 1586364061
transform 1 0 409032 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4446
timestamp 1586364061
transform 1 0 410136 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_4458
timestamp 1586364061
transform 1 0 411240 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_910
timestamp 1586364061
transform 1 0 411792 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_4465
timestamp 1586364061
transform 1 0 411884 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4477
timestamp 1586364061
transform 1 0 412988 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_4489
timestamp 1586364061
transform 1 0 414092 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_911
timestamp 1586364061
transform 1 0 414644 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_4496
timestamp 1586364061
transform 1 0 414736 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4508
timestamp 1586364061
transform 1 0 415840 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_912
timestamp 1586364061
transform 1 0 417496 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_4520
timestamp 1586364061
transform 1 0 416944 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_4527
timestamp 1586364061
transform 1 0 417588 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_4539
timestamp 1586364061
transform 1 0 418692 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_913
timestamp 1586364061
transform 1 0 420348 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_4551
timestamp 1586364061
transform 1 0 419796 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_4558
timestamp 1586364061
transform 1 0 420440 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 422832 0 1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_9_4570
timestamp 1586364061
transform 1 0 421544 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_9_4578
timestamp 1586364061
transform 1 0 422280 0 1 7072
box -38 -48 314 592
<< labels >>
rlabel metal2 s 26514 9520 26570 10000 6 address[0]
port 0 nsew default input
rlabel metal3 s 0 824 480 944 6 address[1]
port 1 nsew default input
rlabel metal2 s 42338 0 42394 480 6 address[2]
port 2 nsew default input
rlabel metal3 s 423520 2184 424000 2304 6 address[3]
port 3 nsew default input
rlabel metal3 s 423520 3136 424000 3256 6 bottom_width_0_height_0__pin_0_
port 4 nsew default input
rlabel metal3 s 423520 4904 424000 5024 6 bottom_width_0_height_0__pin_10_
port 5 nsew default input
rlabel metal2 s 238482 9520 238538 10000 6 bottom_width_0_height_0__pin_11_
port 6 nsew default tristate
rlabel metal3 s 0 9120 480 9240 6 bottom_width_0_height_0__pin_12_
port 7 nsew default input
rlabel metal2 s 211894 0 211950 480 6 bottom_width_0_height_0__pin_13_
port 8 nsew default tristate
rlabel metal3 s 423520 5856 424000 5976 6 bottom_width_0_height_0__pin_14_
port 9 nsew default input
rlabel metal3 s 423520 6808 424000 6928 6 bottom_width_0_height_0__pin_15_
port 10 nsew default tristate
rlabel metal2 s 79506 9520 79562 10000 6 bottom_width_0_height_0__pin_1_
port 11 nsew default tristate
rlabel metal2 s 127070 0 127126 480 6 bottom_width_0_height_0__pin_2_
port 12 nsew default input
rlabel metal3 s 423520 3952 424000 4072 6 bottom_width_0_height_0__pin_3_
port 13 nsew default tristate
rlabel metal3 s 0 2456 480 2576 6 bottom_width_0_height_0__pin_4_
port 14 nsew default input
rlabel metal3 s 0 4088 480 4208 6 bottom_width_0_height_0__pin_5_
port 15 nsew default tristate
rlabel metal3 s 0 5856 480 5976 6 bottom_width_0_height_0__pin_6_
port 16 nsew default input
rlabel metal3 s 0 7488 480 7608 6 bottom_width_0_height_0__pin_7_
port 17 nsew default tristate
rlabel metal2 s 132498 9520 132554 10000 6 bottom_width_0_height_0__pin_8_
port 18 nsew default input
rlabel metal2 s 185490 9520 185546 10000 6 bottom_width_0_height_0__pin_9_
port 19 nsew default tristate
rlabel metal3 s 423520 1232 424000 1352 6 data_in
port 20 nsew default input
rlabel metal3 s 423520 416 424000 536 6 enable
port 21 nsew default input
rlabel metal3 s 423520 7624 424000 7744 6 gfpga_pad_GPIO_PAD[0]
port 22 nsew default bidirectional
rlabel metal2 s 291474 9520 291530 10000 6 gfpga_pad_GPIO_PAD[1]
port 23 nsew default bidirectional
rlabel metal3 s 423520 8576 424000 8696 6 gfpga_pad_GPIO_PAD[2]
port 24 nsew default bidirectional
rlabel metal2 s 344466 9520 344522 10000 6 gfpga_pad_GPIO_PAD[3]
port 25 nsew default bidirectional
rlabel metal2 s 296718 0 296774 480 6 gfpga_pad_GPIO_PAD[4]
port 26 nsew default bidirectional
rlabel metal3 s 423520 9528 424000 9648 6 gfpga_pad_GPIO_PAD[5]
port 27 nsew default bidirectional
rlabel metal2 s 381542 0 381598 480 6 gfpga_pad_GPIO_PAD[6]
port 28 nsew default bidirectional
rlabel metal2 s 397458 9520 397514 10000 6 gfpga_pad_GPIO_PAD[7]
port 29 nsew default bidirectional
rlabel metal4 s 71611 2128 71931 7664 6 vpwr
port 30 nsew default input
rlabel metal4 s 142277 2128 142597 7664 6 vgnd
port 31 nsew default input
<< end >>
