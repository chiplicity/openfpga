magic
tech sky130A
magscale 1 2
timestamp 1605017285
<< locali >>
rect 22569 22143 22603 22313
rect 24317 14527 24351 14833
<< viali >>
rect 23029 25169 23063 25203
rect 24777 25169 24811 25203
rect 22845 25033 22879 25067
rect 24593 25033 24627 25067
rect 25145 24625 25179 24659
rect 23489 24489 23523 24523
rect 22569 24421 22603 24455
rect 23121 24421 23155 24455
rect 23673 24421 23707 24455
rect 24409 24421 24443 24455
rect 24961 24421 24995 24455
rect 25513 24421 25547 24455
rect 23949 24353 23983 24387
rect 19073 24285 19107 24319
rect 22753 24285 22787 24319
rect 24777 24285 24811 24319
rect 25145 24081 25179 24115
rect 23949 24013 23983 24047
rect 13544 23945 13578 23979
rect 19257 23945 19291 23979
rect 21557 23945 21591 23979
rect 23673 23945 23707 23979
rect 24961 23945 24995 23979
rect 10977 23877 11011 23911
rect 13277 23877 13311 23911
rect 16221 23877 16255 23911
rect 19349 23877 19383 23911
rect 19441 23877 19475 23911
rect 21649 23877 21683 23911
rect 21741 23877 21775 23911
rect 22201 23877 22235 23911
rect 21097 23809 21131 23843
rect 10885 23741 10919 23775
rect 14657 23741 14691 23775
rect 15945 23741 15979 23775
rect 18429 23741 18463 23775
rect 18705 23741 18739 23775
rect 18889 23741 18923 23775
rect 21189 23741 21223 23775
rect 13369 23537 13403 23571
rect 14933 23537 14967 23571
rect 20361 23537 20395 23571
rect 21189 23537 21223 23571
rect 25513 23537 25547 23571
rect 19717 23469 19751 23503
rect 14013 23401 14047 23435
rect 14197 23401 14231 23435
rect 20729 23401 20763 23435
rect 21557 23401 21591 23435
rect 24317 23401 24351 23435
rect 10701 23333 10735 23367
rect 10793 23333 10827 23367
rect 11049 23333 11083 23367
rect 15761 23333 15795 23367
rect 15853 23333 15887 23367
rect 18337 23333 18371 23367
rect 18593 23333 18627 23367
rect 24041 23333 24075 23367
rect 25329 23333 25363 23367
rect 25881 23333 25915 23367
rect 16098 23265 16132 23299
rect 18245 23265 18279 23299
rect 21824 23265 21858 23299
rect 12173 23197 12207 23231
rect 13093 23197 13127 23231
rect 13553 23197 13587 23231
rect 13921 23197 13955 23231
rect 14657 23197 14691 23231
rect 17233 23197 17267 23231
rect 22937 23197 22971 23231
rect 23581 23197 23615 23231
rect 23857 23197 23891 23231
rect 24961 23197 24995 23231
rect 9689 22993 9723 23027
rect 10793 22993 10827 23027
rect 11253 22993 11287 23027
rect 14749 22993 14783 23027
rect 16497 22993 16531 23027
rect 18061 22993 18095 23027
rect 19165 22993 19199 23027
rect 19441 22993 19475 23027
rect 9597 22925 9631 22959
rect 13277 22925 13311 22959
rect 13636 22925 13670 22959
rect 18429 22925 18463 22959
rect 11161 22857 11195 22891
rect 18521 22857 18555 22891
rect 20545 22857 20579 22891
rect 20812 22857 20846 22891
rect 23673 22857 23707 22891
rect 24961 22857 24995 22891
rect 9781 22789 9815 22823
rect 11437 22789 11471 22823
rect 13369 22789 13403 22823
rect 16589 22789 16623 22823
rect 16681 22789 16715 22823
rect 18613 22789 18647 22823
rect 23949 22789 23983 22823
rect 9229 22721 9263 22755
rect 16037 22721 16071 22755
rect 17141 22721 17175 22755
rect 15577 22653 15611 22687
rect 16129 22653 16163 22687
rect 21925 22653 21959 22687
rect 25145 22653 25179 22687
rect 8953 22449 8987 22483
rect 9965 22449 9999 22483
rect 10701 22449 10735 22483
rect 13369 22449 13403 22483
rect 15025 22449 15059 22483
rect 15485 22449 15519 22483
rect 16497 22449 16531 22483
rect 18429 22449 18463 22483
rect 19349 22449 19383 22483
rect 20637 22449 20671 22483
rect 21097 22449 21131 22483
rect 23673 22449 23707 22483
rect 25513 22449 25547 22483
rect 18981 22381 19015 22415
rect 21741 22381 21775 22415
rect 24041 22381 24075 22415
rect 10793 22313 10827 22347
rect 14013 22313 14047 22347
rect 14105 22313 14139 22347
rect 15945 22313 15979 22347
rect 16037 22313 16071 22347
rect 19809 22313 19843 22347
rect 22385 22313 22419 22347
rect 22569 22313 22603 22347
rect 11060 22245 11094 22279
rect 15853 22245 15887 22279
rect 16957 22245 16991 22279
rect 17049 22245 17083 22279
rect 19533 22245 19567 22279
rect 13921 22177 13955 22211
rect 14749 22177 14783 22211
rect 17294 22177 17328 22211
rect 21649 22177 21683 22211
rect 22109 22177 22143 22211
rect 22201 22177 22235 22211
rect 23489 22245 23523 22279
rect 24593 22245 24627 22279
rect 25145 22245 25179 22279
rect 22753 22177 22787 22211
rect 9229 22109 9263 22143
rect 10333 22109 10367 22143
rect 12173 22109 12207 22143
rect 13093 22109 13127 22143
rect 13553 22109 13587 22143
rect 22569 22109 22603 22143
rect 23305 22109 23339 22143
rect 24777 22109 24811 22143
rect 10793 21905 10827 21939
rect 11253 21905 11287 21939
rect 11529 21905 11563 21939
rect 13553 21905 13587 21939
rect 14381 21905 14415 21939
rect 15393 21905 15427 21939
rect 16865 21905 16899 21939
rect 18797 21905 18831 21939
rect 19533 21905 19567 21939
rect 21925 21905 21959 21939
rect 13461 21837 13495 21871
rect 14105 21837 14139 21871
rect 21741 21837 21775 21871
rect 15485 21769 15519 21803
rect 15752 21769 15786 21803
rect 18061 21769 18095 21803
rect 18337 21769 18371 21803
rect 24593 21769 24627 21803
rect 19257 21633 19291 21667
rect 23489 21565 23523 21599
rect 24777 21565 24811 21599
rect 10333 21361 10367 21395
rect 22293 21361 22327 21395
rect 24593 21361 24627 21395
rect 16681 21293 16715 21327
rect 10425 21225 10459 21259
rect 14197 21225 14231 21259
rect 15117 21225 15151 21259
rect 16221 21225 16255 21259
rect 17325 21225 17359 21259
rect 19441 21225 19475 21259
rect 23949 21225 23983 21259
rect 13921 21157 13955 21191
rect 14657 21157 14691 21191
rect 20913 21157 20947 21191
rect 24961 21157 24995 21191
rect 25513 21157 25547 21191
rect 10692 21089 10726 21123
rect 16589 21089 16623 21123
rect 18705 21089 18739 21123
rect 19349 21089 19383 21123
rect 21180 21089 21214 21123
rect 23765 21089 23799 21123
rect 11805 21021 11839 21055
rect 12909 21021 12943 21055
rect 15577 21021 15611 21055
rect 17049 21021 17083 21055
rect 17141 21021 17175 21055
rect 17693 21021 17727 21055
rect 18337 21021 18371 21055
rect 18889 21021 18923 21055
rect 19257 21021 19291 21055
rect 20729 21021 20763 21055
rect 23213 21021 23247 21055
rect 23397 21021 23431 21055
rect 23857 21021 23891 21055
rect 25145 21021 25179 21055
rect 10517 20817 10551 20851
rect 10793 20817 10827 20851
rect 14013 20817 14047 20851
rect 16129 20817 16163 20851
rect 18245 20817 18279 20851
rect 18889 20817 18923 20851
rect 20361 20817 20395 20851
rect 22017 20817 22051 20851
rect 22385 20817 22419 20851
rect 11253 20749 11287 20783
rect 19248 20749 19282 20783
rect 21005 20749 21039 20783
rect 23489 20749 23523 20783
rect 23940 20749 23974 20783
rect 11161 20681 11195 20715
rect 12817 20681 12851 20715
rect 14381 20681 14415 20715
rect 16497 20681 16531 20715
rect 22477 20681 22511 20715
rect 11437 20613 11471 20647
rect 12909 20613 12943 20647
rect 13001 20613 13035 20647
rect 14473 20613 14507 20647
rect 14657 20613 14691 20647
rect 16589 20613 16623 20647
rect 16773 20613 16807 20647
rect 17141 20613 17175 20647
rect 18981 20613 19015 20647
rect 22661 20613 22695 20647
rect 23673 20613 23707 20647
rect 16037 20545 16071 20579
rect 12449 20477 12483 20511
rect 13737 20477 13771 20511
rect 25053 20477 25087 20511
rect 10885 20273 10919 20307
rect 12633 20273 12667 20307
rect 13185 20273 13219 20307
rect 14473 20273 14507 20307
rect 14841 20273 14875 20307
rect 16129 20273 16163 20307
rect 17693 20273 17727 20307
rect 20453 20273 20487 20307
rect 22109 20273 22143 20307
rect 23765 20273 23799 20307
rect 24685 20273 24719 20307
rect 13553 20205 13587 20239
rect 11253 20137 11287 20171
rect 15301 20137 15335 20171
rect 19441 20137 19475 20171
rect 19533 20137 19567 20171
rect 19993 20137 20027 20171
rect 22385 20137 22419 20171
rect 11520 20069 11554 20103
rect 13737 20069 13771 20103
rect 16313 20069 16347 20103
rect 22652 20069 22686 20103
rect 24869 20069 24903 20103
rect 25421 20069 25455 20103
rect 14013 20001 14047 20035
rect 16558 20001 16592 20035
rect 18521 20001 18555 20035
rect 19349 20001 19383 20035
rect 24317 20001 24351 20035
rect 10517 19933 10551 19967
rect 15761 19933 15795 19967
rect 18797 19933 18831 19967
rect 18981 19933 19015 19967
rect 21649 19933 21683 19967
rect 25053 19933 25087 19967
rect 10885 19729 10919 19763
rect 11713 19729 11747 19763
rect 12725 19729 12759 19763
rect 13369 19729 13403 19763
rect 14105 19729 14139 19763
rect 16405 19729 16439 19763
rect 18521 19729 18555 19763
rect 22385 19729 22419 19763
rect 22569 19729 22603 19763
rect 25329 19729 25363 19763
rect 11253 19661 11287 19695
rect 13277 19661 13311 19695
rect 15270 19661 15304 19695
rect 22109 19661 22143 19695
rect 23029 19661 23063 19695
rect 19533 19593 19567 19627
rect 19809 19593 19843 19627
rect 23857 19593 23891 19627
rect 25145 19593 25179 19627
rect 13553 19525 13587 19559
rect 15025 19525 15059 19559
rect 24133 19525 24167 19559
rect 12909 19457 12943 19491
rect 17049 19389 17083 19423
rect 19349 19389 19383 19423
rect 11897 19185 11931 19219
rect 15485 19185 15519 19219
rect 20269 19185 20303 19219
rect 23857 19185 23891 19219
rect 25513 19185 25547 19219
rect 12081 19049 12115 19083
rect 19809 19049 19843 19083
rect 22937 19049 22971 19083
rect 12348 18981 12382 19015
rect 16865 18981 16899 19015
rect 18797 18981 18831 19015
rect 21557 18981 21591 19015
rect 24593 18981 24627 19015
rect 25145 18981 25179 19015
rect 19717 18913 19751 18947
rect 22293 18913 22327 18947
rect 22845 18913 22879 18947
rect 13461 18845 13495 18879
rect 14013 18845 14047 18879
rect 15025 18845 15059 18879
rect 19073 18845 19107 18879
rect 19257 18845 19291 18879
rect 19625 18845 19659 18879
rect 21925 18845 21959 18879
rect 22385 18845 22419 18879
rect 22753 18845 22787 18879
rect 24777 18845 24811 18879
rect 12173 18641 12207 18675
rect 13001 18641 13035 18675
rect 14841 18641 14875 18675
rect 21005 18573 21039 18607
rect 21364 18573 21398 18607
rect 13369 18505 13403 18539
rect 13728 18505 13762 18539
rect 18317 18505 18351 18539
rect 21097 18505 21131 18539
rect 24041 18505 24075 18539
rect 25237 18505 25271 18539
rect 13461 18437 13495 18471
rect 18061 18437 18095 18471
rect 24133 18437 24167 18471
rect 24225 18437 24259 18471
rect 25421 18369 25455 18403
rect 15945 18301 15979 18335
rect 17785 18301 17819 18335
rect 19441 18301 19475 18335
rect 22477 18301 22511 18335
rect 23673 18301 23707 18335
rect 13829 18097 13863 18131
rect 19717 18097 19751 18131
rect 24409 18097 24443 18131
rect 24961 18097 24995 18131
rect 22017 18029 22051 18063
rect 22845 18029 22879 18063
rect 20361 17961 20395 17995
rect 21557 17961 21591 17995
rect 23029 17961 23063 17995
rect 15853 17893 15887 17927
rect 16109 17893 16143 17927
rect 18337 17893 18371 17927
rect 21373 17893 21407 17927
rect 22293 17893 22327 17927
rect 23285 17893 23319 17927
rect 15669 17825 15703 17859
rect 17785 17825 17819 17859
rect 18153 17825 18187 17859
rect 18604 17825 18638 17859
rect 20729 17825 20763 17859
rect 21281 17825 21315 17859
rect 25329 17825 25363 17859
rect 13553 17757 13587 17791
rect 14289 17757 14323 17791
rect 17233 17757 17267 17791
rect 20913 17757 20947 17791
rect 15853 17553 15887 17587
rect 18521 17553 18555 17587
rect 21557 17553 21591 17587
rect 23121 17553 23155 17587
rect 23489 17553 23523 17587
rect 23949 17553 23983 17587
rect 25605 17553 25639 17587
rect 16313 17485 16347 17519
rect 20422 17485 20456 17519
rect 24409 17485 24443 17519
rect 14473 17417 14507 17451
rect 16221 17417 16255 17451
rect 18429 17417 18463 17451
rect 19165 17417 19199 17451
rect 20177 17417 20211 17451
rect 24133 17417 24167 17451
rect 25421 17417 25455 17451
rect 14565 17349 14599 17383
rect 14749 17349 14783 17383
rect 15301 17349 15335 17383
rect 16405 17349 16439 17383
rect 18613 17349 18647 17383
rect 14105 17281 14139 17315
rect 12173 17213 12207 17247
rect 13737 17213 13771 17247
rect 17785 17213 17819 17247
rect 18061 17213 18095 17247
rect 13645 17009 13679 17043
rect 14749 17009 14783 17043
rect 16681 17009 16715 17043
rect 17325 17009 17359 17043
rect 19165 17009 19199 17043
rect 20177 17009 20211 17043
rect 20545 17009 20579 17043
rect 23857 17009 23891 17043
rect 24777 17009 24811 17043
rect 25513 17009 25547 17043
rect 26341 17009 26375 17043
rect 12081 16941 12115 16975
rect 13093 16941 13127 16975
rect 17601 16941 17635 16975
rect 12633 16873 12667 16907
rect 14197 16873 14231 16907
rect 18337 16873 18371 16907
rect 20913 16873 20947 16907
rect 23029 16873 23063 16907
rect 24317 16873 24351 16907
rect 13553 16805 13587 16839
rect 14013 16805 14047 16839
rect 15301 16805 15335 16839
rect 15557 16805 15591 16839
rect 18245 16805 18279 16839
rect 24041 16805 24075 16839
rect 25329 16805 25363 16839
rect 25881 16805 25915 16839
rect 11897 16737 11931 16771
rect 12541 16737 12575 16771
rect 14105 16737 14139 16771
rect 18153 16737 18187 16771
rect 19349 16737 19383 16771
rect 12449 16669 12483 16703
rect 15025 16669 15059 16703
rect 17785 16669 17819 16703
rect 18797 16669 18831 16703
rect 12173 16465 12207 16499
rect 13553 16465 13587 16499
rect 15117 16465 15151 16499
rect 16221 16465 16255 16499
rect 16589 16465 16623 16499
rect 17877 16465 17911 16499
rect 18061 16465 18095 16499
rect 18521 16465 18555 16499
rect 21465 16465 21499 16499
rect 25421 16465 25455 16499
rect 14004 16397 14038 16431
rect 15853 16397 15887 16431
rect 17325 16397 17359 16431
rect 18429 16397 18463 16431
rect 24225 16397 24259 16431
rect 21833 16329 21867 16363
rect 23949 16329 23983 16363
rect 25237 16329 25271 16363
rect 13737 16261 13771 16295
rect 18705 16261 18739 16295
rect 21925 16261 21959 16295
rect 22109 16261 22143 16295
rect 22477 16125 22511 16159
rect 13921 15921 13955 15955
rect 15301 15921 15335 15955
rect 18705 15921 18739 15955
rect 19073 15921 19107 15955
rect 21833 15921 21867 15955
rect 23949 15921 23983 15955
rect 25237 15921 25271 15955
rect 14473 15853 14507 15887
rect 18429 15853 18463 15887
rect 24317 15853 24351 15887
rect 15853 15785 15887 15819
rect 17141 15785 17175 15819
rect 17785 15785 17819 15819
rect 17877 15785 17911 15819
rect 22017 15785 22051 15819
rect 24777 15785 24811 15819
rect 12548 15717 12582 15751
rect 15117 15717 15151 15751
rect 15761 15717 15795 15751
rect 16865 15717 16899 15751
rect 20729 15717 20763 15751
rect 24501 15717 24535 15751
rect 12081 15649 12115 15683
rect 12808 15649 12842 15683
rect 17693 15649 17727 15683
rect 21189 15649 21223 15683
rect 22284 15649 22318 15683
rect 12449 15581 12483 15615
rect 15669 15581 15703 15615
rect 17325 15581 17359 15615
rect 21557 15581 21591 15615
rect 23397 15581 23431 15615
rect 13829 15377 13863 15411
rect 14381 15377 14415 15411
rect 14933 15377 14967 15411
rect 15485 15377 15519 15411
rect 16405 15377 16439 15411
rect 18245 15377 18279 15411
rect 20545 15377 20579 15411
rect 21649 15377 21683 15411
rect 22109 15377 22143 15411
rect 24133 15377 24167 15411
rect 15761 15309 15795 15343
rect 12716 15241 12750 15275
rect 16313 15241 16347 15275
rect 16773 15241 16807 15275
rect 16865 15241 16899 15275
rect 19432 15241 19466 15275
rect 22017 15241 22051 15275
rect 24041 15241 24075 15275
rect 25237 15241 25271 15275
rect 12449 15173 12483 15207
rect 16957 15173 16991 15207
rect 19165 15173 19199 15207
rect 22201 15173 22235 15207
rect 24225 15173 24259 15207
rect 25421 15173 25455 15207
rect 21465 15037 21499 15071
rect 23673 15037 23707 15071
rect 12817 14833 12851 14867
rect 17141 14833 17175 14867
rect 17693 14833 17727 14867
rect 20729 14833 20763 14867
rect 23397 14833 23431 14867
rect 24317 14833 24351 14867
rect 24501 14833 24535 14867
rect 25237 14833 25271 14867
rect 22937 14765 22971 14799
rect 23489 14765 23523 14799
rect 21005 14697 21039 14731
rect 24041 14697 24075 14731
rect 15669 14629 15703 14663
rect 15761 14629 15795 14663
rect 18153 14629 18187 14663
rect 18245 14629 18279 14663
rect 18501 14629 18535 14663
rect 23857 14629 23891 14663
rect 16028 14561 16062 14595
rect 21250 14561 21284 14595
rect 23949 14561 23983 14595
rect 25605 14765 25639 14799
rect 25053 14629 25087 14663
rect 24869 14561 24903 14595
rect 12449 14493 12483 14527
rect 19625 14493 19659 14527
rect 22385 14493 22419 14527
rect 24317 14493 24351 14527
rect 16405 14289 16439 14323
rect 17417 14289 17451 14323
rect 19165 14289 19199 14323
rect 19625 14289 19659 14323
rect 21557 14289 21591 14323
rect 22477 14289 22511 14323
rect 23489 14289 23523 14323
rect 23949 14289 23983 14323
rect 25053 14289 25087 14323
rect 25513 14289 25547 14323
rect 16313 14221 16347 14255
rect 21925 14221 21959 14255
rect 24317 14221 24351 14255
rect 16773 14153 16807 14187
rect 18061 14153 18095 14187
rect 21373 14153 21407 14187
rect 24041 14153 24075 14187
rect 25329 14153 25363 14187
rect 16865 14085 16899 14119
rect 17049 14085 17083 14119
rect 15853 14017 15887 14051
rect 21097 13949 21131 13983
rect 22293 13949 22327 13983
rect 15485 13745 15519 13779
rect 16129 13745 16163 13779
rect 17141 13745 17175 13779
rect 23673 13745 23707 13779
rect 24133 13745 24167 13779
rect 24777 13745 24811 13779
rect 25513 13745 25547 13779
rect 16497 13677 16531 13711
rect 17601 13609 17635 13643
rect 17785 13609 17819 13643
rect 21373 13609 21407 13643
rect 21833 13609 21867 13643
rect 24501 13609 24535 13643
rect 25237 13609 25271 13643
rect 15117 13541 15151 13575
rect 15301 13541 15335 13575
rect 17049 13541 17083 13575
rect 17509 13541 17543 13575
rect 20729 13541 20763 13575
rect 21097 13541 21131 13575
rect 23489 13541 23523 13575
rect 24593 13541 24627 13575
rect 13645 13201 13679 13235
rect 16957 13201 16991 13235
rect 17417 13201 17451 13235
rect 22017 13201 22051 13235
rect 24777 13201 24811 13235
rect 16497 13133 16531 13167
rect 20882 13133 20916 13167
rect 13461 13065 13495 13099
rect 16773 13065 16807 13099
rect 20637 13065 20671 13099
rect 24593 13065 24627 13099
rect 20545 12861 20579 12895
rect 13461 12657 13495 12691
rect 20361 12657 20395 12691
rect 20637 12657 20671 12691
rect 23949 12657 23983 12691
rect 24685 12657 24719 12691
rect 25513 12657 25547 12691
rect 12909 12521 12943 12555
rect 15485 12521 15519 12555
rect 16865 12521 16899 12555
rect 17601 12521 17635 12555
rect 20913 12521 20947 12555
rect 24409 12521 24443 12555
rect 12541 12453 12575 12487
rect 12633 12453 12667 12487
rect 15301 12453 15335 12487
rect 16037 12453 16071 12487
rect 17417 12453 17451 12487
rect 21169 12453 21203 12487
rect 23765 12453 23799 12487
rect 24869 12453 24903 12487
rect 18245 12317 18279 12351
rect 19809 12317 19843 12351
rect 22293 12317 22327 12351
rect 25053 12317 25087 12351
rect 13185 12113 13219 12147
rect 15669 12113 15703 12147
rect 20821 12113 20855 12147
rect 24593 12113 24627 12147
rect 13553 11977 13587 12011
rect 16037 11977 16071 12011
rect 21189 11977 21223 12011
rect 24409 11977 24443 12011
rect 13645 11909 13679 11943
rect 13829 11909 13863 11943
rect 15577 11909 15611 11943
rect 16129 11909 16163 11943
rect 16313 11909 16347 11943
rect 18337 11909 18371 11943
rect 21281 11909 21315 11943
rect 21465 11909 21499 11943
rect 20729 11841 20763 11875
rect 12725 11773 12759 11807
rect 18797 11773 18831 11807
rect 18337 11569 18371 11603
rect 19993 11569 20027 11603
rect 20913 11569 20947 11603
rect 21925 11569 21959 11603
rect 24501 11569 24535 11603
rect 18245 11501 18279 11535
rect 18797 11433 18831 11467
rect 18889 11433 18923 11467
rect 21465 11433 21499 11467
rect 22293 11433 22327 11467
rect 12633 11365 12667 11399
rect 12889 11365 12923 11399
rect 15117 11365 15151 11399
rect 15577 11365 15611 11399
rect 18705 11365 18739 11399
rect 12541 11297 12575 11331
rect 15822 11297 15856 11331
rect 17877 11297 17911 11331
rect 20729 11297 20763 11331
rect 21281 11297 21315 11331
rect 14013 11229 14047 11263
rect 14749 11229 14783 11263
rect 16957 11229 16991 11263
rect 20361 11229 20395 11263
rect 21373 11229 21407 11263
rect 12725 11025 12759 11059
rect 13277 11025 13311 11059
rect 13921 11025 13955 11059
rect 15485 11025 15519 11059
rect 16037 11025 16071 11059
rect 16589 11025 16623 11059
rect 19809 11025 19843 11059
rect 20821 11025 20855 11059
rect 22293 11025 22327 11059
rect 24777 11025 24811 11059
rect 16405 10957 16439 10991
rect 21158 10957 21192 10991
rect 13645 10889 13679 10923
rect 14372 10889 14406 10923
rect 18429 10889 18463 10923
rect 18696 10889 18730 10923
rect 20913 10889 20947 10923
rect 24593 10889 24627 10923
rect 14105 10821 14139 10855
rect 12357 10481 12391 10515
rect 12909 10481 12943 10515
rect 13461 10481 13495 10515
rect 14565 10481 14599 10515
rect 14841 10481 14875 10515
rect 16405 10481 16439 10515
rect 16773 10481 16807 10515
rect 18889 10481 18923 10515
rect 21097 10481 21131 10515
rect 21465 10481 21499 10515
rect 24777 10481 24811 10515
rect 24501 10413 24535 10447
rect 14013 10345 14047 10379
rect 10977 10277 11011 10311
rect 16865 10277 16899 10311
rect 17121 10277 17155 10311
rect 24593 10277 24627 10311
rect 10793 10209 10827 10243
rect 11222 10209 11256 10243
rect 13369 10209 13403 10243
rect 13829 10209 13863 10243
rect 13921 10209 13955 10243
rect 18245 10141 18279 10175
rect 19257 10141 19291 10175
rect 25237 10141 25271 10175
rect 10977 9937 11011 9971
rect 13553 9937 13587 9971
rect 15945 9937 15979 9971
rect 18797 9937 18831 9971
rect 19257 9937 19291 9971
rect 24777 9937 24811 9971
rect 16313 9801 16347 9835
rect 19165 9801 19199 9835
rect 24593 9801 24627 9835
rect 16405 9733 16439 9767
rect 16497 9733 16531 9767
rect 19441 9733 19475 9767
rect 16405 9393 16439 9427
rect 19165 9393 19199 9427
rect 16681 9325 16715 9359
rect 19533 9325 19567 9359
rect 24777 9325 24811 9359
rect 25237 9325 25271 9359
rect 24593 9189 24627 9223
rect 16037 9053 16071 9087
rect 18889 9053 18923 9087
rect 24501 9053 24535 9087
rect 24777 8849 24811 8883
rect 24593 8713 24627 8747
rect 24685 8305 24719 8339
rect 24593 7625 24627 7659
rect 24777 7489 24811 7523
rect 17785 7217 17819 7251
rect 24685 7217 24719 7251
rect 18245 7081 18279 7115
rect 17601 7013 17635 7047
rect 16497 6129 16531 6163
rect 16313 5925 16347 5959
rect 16957 5857 16991 5891
rect 15485 5041 15519 5075
rect 15945 4905 15979 4939
rect 15301 4837 15335 4871
rect 24593 3749 24627 3783
rect 24777 3613 24811 3647
rect 25237 3613 25271 3647
<< metal1 >>
rect 21542 26384 21548 26436
rect 21600 26424 21606 26436
rect 23934 26424 23940 26436
rect 21600 26396 23940 26424
rect 21600 26384 21606 26396
rect 23934 26384 23940 26396
rect 23992 26384 23998 26436
rect 1104 25314 26864 25336
rect 1104 25262 10315 25314
rect 10367 25262 10379 25314
rect 10431 25262 10443 25314
rect 10495 25262 10507 25314
rect 10559 25262 19648 25314
rect 19700 25262 19712 25314
rect 19764 25262 19776 25314
rect 19828 25262 19840 25314
rect 19892 25262 26864 25314
rect 1104 25240 26864 25262
rect 23017 25203 23075 25209
rect 23017 25169 23029 25203
rect 23063 25200 23075 25203
rect 23566 25200 23572 25212
rect 23063 25172 23572 25200
rect 23063 25169 23075 25172
rect 23017 25163 23075 25169
rect 23566 25160 23572 25172
rect 23624 25160 23630 25212
rect 24762 25200 24768 25212
rect 24723 25172 24768 25200
rect 24762 25160 24768 25172
rect 24820 25160 24826 25212
rect 22830 25064 22836 25076
rect 22791 25036 22836 25064
rect 22830 25024 22836 25036
rect 22888 25024 22894 25076
rect 24581 25067 24639 25073
rect 24581 25033 24593 25067
rect 24627 25064 24639 25067
rect 24762 25064 24768 25076
rect 24627 25036 24768 25064
rect 24627 25033 24639 25036
rect 24581 25027 24639 25033
rect 24762 25024 24768 25036
rect 24820 25024 24826 25076
rect 1104 24770 26864 24792
rect 1104 24718 5648 24770
rect 5700 24718 5712 24770
rect 5764 24718 5776 24770
rect 5828 24718 5840 24770
rect 5892 24718 14982 24770
rect 15034 24718 15046 24770
rect 15098 24718 15110 24770
rect 15162 24718 15174 24770
rect 15226 24718 24315 24770
rect 24367 24718 24379 24770
rect 24431 24718 24443 24770
rect 24495 24718 24507 24770
rect 24559 24718 26864 24770
rect 1104 24696 26864 24718
rect 25130 24656 25136 24668
rect 25091 24628 25136 24656
rect 25130 24616 25136 24628
rect 25188 24616 25194 24668
rect 22830 24548 22836 24600
rect 22888 24588 22894 24600
rect 22888 24560 23428 24588
rect 22888 24548 22894 24560
rect 15378 24480 15384 24532
rect 15436 24520 15442 24532
rect 15930 24520 15936 24532
rect 15436 24492 15936 24520
rect 15436 24480 15442 24492
rect 15930 24480 15936 24492
rect 15988 24480 15994 24532
rect 20714 24480 20720 24532
rect 20772 24520 20778 24532
rect 21634 24520 21640 24532
rect 20772 24492 21640 24520
rect 20772 24480 20778 24492
rect 21634 24480 21640 24492
rect 21692 24480 21698 24532
rect 23400 24520 23428 24560
rect 23477 24523 23535 24529
rect 23477 24520 23489 24523
rect 23400 24492 23489 24520
rect 23477 24489 23489 24492
rect 23523 24489 23535 24523
rect 23477 24483 23535 24489
rect 19334 24412 19340 24464
rect 19392 24452 19398 24464
rect 20438 24452 20444 24464
rect 19392 24424 20444 24452
rect 19392 24412 19398 24424
rect 20438 24412 20444 24424
rect 20496 24412 20502 24464
rect 22554 24452 22560 24464
rect 22515 24424 22560 24452
rect 22554 24412 22560 24424
rect 22612 24452 22618 24464
rect 23109 24455 23167 24461
rect 23109 24452 23121 24455
rect 22612 24424 23121 24452
rect 22612 24412 22618 24424
rect 23109 24421 23121 24424
rect 23155 24421 23167 24455
rect 23109 24415 23167 24421
rect 23661 24455 23719 24461
rect 23661 24421 23673 24455
rect 23707 24452 23719 24455
rect 24118 24452 24124 24464
rect 23707 24424 24124 24452
rect 23707 24421 23719 24424
rect 23661 24415 23719 24421
rect 24118 24412 24124 24424
rect 24176 24452 24182 24464
rect 24397 24455 24455 24461
rect 24397 24452 24409 24455
rect 24176 24424 24409 24452
rect 24176 24412 24182 24424
rect 24397 24421 24409 24424
rect 24443 24421 24455 24455
rect 24946 24452 24952 24464
rect 24907 24424 24952 24452
rect 24397 24415 24455 24421
rect 24946 24412 24952 24424
rect 25004 24452 25010 24464
rect 25501 24455 25559 24461
rect 25501 24452 25513 24455
rect 25004 24424 25513 24452
rect 25004 24412 25010 24424
rect 25501 24421 25513 24424
rect 25547 24421 25559 24455
rect 25501 24415 25559 24421
rect 23937 24387 23995 24393
rect 23937 24353 23949 24387
rect 23983 24384 23995 24387
rect 25314 24384 25320 24396
rect 23983 24356 25320 24384
rect 23983 24353 23995 24356
rect 23937 24347 23995 24353
rect 25314 24344 25320 24356
rect 25372 24344 25378 24396
rect 19061 24319 19119 24325
rect 19061 24285 19073 24319
rect 19107 24316 19119 24319
rect 19150 24316 19156 24328
rect 19107 24288 19156 24316
rect 19107 24285 19119 24288
rect 19061 24279 19119 24285
rect 19150 24276 19156 24288
rect 19208 24276 19214 24328
rect 22741 24319 22799 24325
rect 22741 24285 22753 24319
rect 22787 24316 22799 24319
rect 23382 24316 23388 24328
rect 22787 24288 23388 24316
rect 22787 24285 22799 24288
rect 22741 24279 22799 24285
rect 23382 24276 23388 24288
rect 23440 24276 23446 24328
rect 24762 24316 24768 24328
rect 24723 24288 24768 24316
rect 24762 24276 24768 24288
rect 24820 24276 24826 24328
rect 1104 24226 26864 24248
rect 1104 24174 10315 24226
rect 10367 24174 10379 24226
rect 10431 24174 10443 24226
rect 10495 24174 10507 24226
rect 10559 24174 19648 24226
rect 19700 24174 19712 24226
rect 19764 24174 19776 24226
rect 19828 24174 19840 24226
rect 19892 24174 26864 24226
rect 1104 24152 26864 24174
rect 25130 24112 25136 24124
rect 25091 24084 25136 24112
rect 25130 24072 25136 24084
rect 25188 24072 25194 24124
rect 23937 24047 23995 24053
rect 23937 24013 23949 24047
rect 23983 24044 23995 24047
rect 24762 24044 24768 24056
rect 23983 24016 24768 24044
rect 23983 24013 23995 24016
rect 23937 24007 23995 24013
rect 24762 24004 24768 24016
rect 24820 24004 24826 24056
rect 13532 23979 13590 23985
rect 13532 23945 13544 23979
rect 13578 23976 13590 23979
rect 14826 23976 14832 23988
rect 13578 23948 14832 23976
rect 13578 23945 13590 23948
rect 13532 23939 13590 23945
rect 14826 23936 14832 23948
rect 14884 23936 14890 23988
rect 19150 23936 19156 23988
rect 19208 23976 19214 23988
rect 19245 23979 19303 23985
rect 19245 23976 19257 23979
rect 19208 23948 19257 23976
rect 19208 23936 19214 23948
rect 19245 23945 19257 23948
rect 19291 23945 19303 23979
rect 19245 23939 19303 23945
rect 20346 23936 20352 23988
rect 20404 23976 20410 23988
rect 21545 23979 21603 23985
rect 21545 23976 21557 23979
rect 20404 23948 21557 23976
rect 20404 23936 20410 23948
rect 21545 23945 21557 23948
rect 21591 23945 21603 23979
rect 21545 23939 21603 23945
rect 22094 23936 22100 23988
rect 22152 23976 22158 23988
rect 23382 23976 23388 23988
rect 22152 23948 23388 23976
rect 22152 23936 22158 23948
rect 23382 23936 23388 23948
rect 23440 23936 23446 23988
rect 23566 23936 23572 23988
rect 23624 23976 23630 23988
rect 23661 23979 23719 23985
rect 23661 23976 23673 23979
rect 23624 23948 23673 23976
rect 23624 23936 23630 23948
rect 23661 23945 23673 23948
rect 23707 23945 23719 23979
rect 23661 23939 23719 23945
rect 24854 23936 24860 23988
rect 24912 23976 24918 23988
rect 24949 23979 25007 23985
rect 24949 23976 24961 23979
rect 24912 23948 24961 23976
rect 24912 23936 24918 23948
rect 24949 23945 24961 23948
rect 24995 23945 25007 23979
rect 24949 23939 25007 23945
rect 10962 23908 10968 23920
rect 10923 23880 10968 23908
rect 10962 23868 10968 23880
rect 11020 23868 11026 23920
rect 13262 23908 13268 23920
rect 13223 23880 13268 23908
rect 13262 23868 13268 23880
rect 13320 23868 13326 23920
rect 16206 23908 16212 23920
rect 16167 23880 16212 23908
rect 16206 23868 16212 23880
rect 16264 23868 16270 23920
rect 19337 23911 19395 23917
rect 19337 23908 19349 23911
rect 18708 23880 19349 23908
rect 10870 23772 10876 23784
rect 10831 23744 10876 23772
rect 10870 23732 10876 23744
rect 10928 23732 10934 23784
rect 14182 23732 14188 23784
rect 14240 23772 14246 23784
rect 14645 23775 14703 23781
rect 14645 23772 14657 23775
rect 14240 23744 14657 23772
rect 14240 23732 14246 23744
rect 14645 23741 14657 23744
rect 14691 23741 14703 23775
rect 14645 23735 14703 23741
rect 15933 23775 15991 23781
rect 15933 23741 15945 23775
rect 15979 23772 15991 23775
rect 16022 23772 16028 23784
rect 15979 23744 16028 23772
rect 15979 23741 15991 23744
rect 15933 23735 15991 23741
rect 16022 23732 16028 23744
rect 16080 23732 16086 23784
rect 18414 23772 18420 23784
rect 18375 23744 18420 23772
rect 18414 23732 18420 23744
rect 18472 23732 18478 23784
rect 18598 23732 18604 23784
rect 18656 23772 18662 23784
rect 18708 23781 18736 23880
rect 19337 23877 19349 23880
rect 19383 23877 19395 23911
rect 19337 23871 19395 23877
rect 19426 23868 19432 23920
rect 19484 23908 19490 23920
rect 19484 23880 19529 23908
rect 19484 23868 19490 23880
rect 21174 23868 21180 23920
rect 21232 23908 21238 23920
rect 21637 23911 21695 23917
rect 21637 23908 21649 23911
rect 21232 23880 21649 23908
rect 21232 23868 21238 23880
rect 21637 23877 21649 23880
rect 21683 23877 21695 23911
rect 21637 23871 21695 23877
rect 21729 23911 21787 23917
rect 21729 23877 21741 23911
rect 21775 23908 21787 23911
rect 22189 23911 22247 23917
rect 22189 23908 22201 23911
rect 21775 23880 22201 23908
rect 21775 23877 21787 23880
rect 21729 23871 21787 23877
rect 22189 23877 22201 23880
rect 22235 23908 22247 23911
rect 22278 23908 22284 23920
rect 22235 23880 22284 23908
rect 22235 23877 22247 23880
rect 22189 23871 22247 23877
rect 21085 23843 21143 23849
rect 21085 23809 21097 23843
rect 21131 23840 21143 23843
rect 21744 23840 21772 23871
rect 22278 23868 22284 23880
rect 22336 23868 22342 23920
rect 21131 23812 21772 23840
rect 21131 23809 21143 23812
rect 21085 23803 21143 23809
rect 18693 23775 18751 23781
rect 18693 23772 18705 23775
rect 18656 23744 18705 23772
rect 18656 23732 18662 23744
rect 18693 23741 18705 23744
rect 18739 23741 18751 23775
rect 18693 23735 18751 23741
rect 18877 23775 18935 23781
rect 18877 23741 18889 23775
rect 18923 23772 18935 23775
rect 19334 23772 19340 23784
rect 18923 23744 19340 23772
rect 18923 23741 18935 23744
rect 18877 23735 18935 23741
rect 19334 23732 19340 23744
rect 19392 23732 19398 23784
rect 21177 23775 21235 23781
rect 21177 23741 21189 23775
rect 21223 23772 21235 23775
rect 22002 23772 22008 23784
rect 21223 23744 22008 23772
rect 21223 23741 21235 23744
rect 21177 23735 21235 23741
rect 22002 23732 22008 23744
rect 22060 23732 22066 23784
rect 1104 23682 26864 23704
rect 1104 23630 5648 23682
rect 5700 23630 5712 23682
rect 5764 23630 5776 23682
rect 5828 23630 5840 23682
rect 5892 23630 14982 23682
rect 15034 23630 15046 23682
rect 15098 23630 15110 23682
rect 15162 23630 15174 23682
rect 15226 23630 24315 23682
rect 24367 23630 24379 23682
rect 24431 23630 24443 23682
rect 24495 23630 24507 23682
rect 24559 23630 26864 23682
rect 1104 23608 26864 23630
rect 13354 23568 13360 23580
rect 13315 23540 13360 23568
rect 13354 23528 13360 23540
rect 13412 23568 13418 23580
rect 13412 23540 14044 23568
rect 13412 23528 13418 23540
rect 14016 23441 14044 23540
rect 14826 23528 14832 23580
rect 14884 23568 14890 23580
rect 14921 23571 14979 23577
rect 14921 23568 14933 23571
rect 14884 23540 14933 23568
rect 14884 23528 14890 23540
rect 14921 23537 14933 23540
rect 14967 23537 14979 23571
rect 14921 23531 14979 23537
rect 19242 23528 19248 23580
rect 19300 23568 19306 23580
rect 20346 23568 20352 23580
rect 19300 23540 20352 23568
rect 19300 23528 19306 23540
rect 20346 23528 20352 23540
rect 20404 23528 20410 23580
rect 21174 23568 21180 23580
rect 21135 23540 21180 23568
rect 21174 23528 21180 23540
rect 21232 23528 21238 23580
rect 25498 23568 25504 23580
rect 25459 23540 25504 23568
rect 25498 23528 25504 23540
rect 25556 23528 25562 23580
rect 19426 23460 19432 23512
rect 19484 23500 19490 23512
rect 19705 23503 19763 23509
rect 19705 23500 19717 23503
rect 19484 23472 19717 23500
rect 19484 23460 19490 23472
rect 19705 23469 19717 23472
rect 19751 23469 19763 23503
rect 19705 23463 19763 23469
rect 14001 23435 14059 23441
rect 14001 23401 14013 23435
rect 14047 23401 14059 23435
rect 14182 23432 14188 23444
rect 14143 23404 14188 23432
rect 14001 23395 14059 23401
rect 14182 23392 14188 23404
rect 14240 23392 14246 23444
rect 20714 23432 20720 23444
rect 20627 23404 20720 23432
rect 20714 23392 20720 23404
rect 20772 23432 20778 23444
rect 21542 23432 21548 23444
rect 20772 23404 21548 23432
rect 20772 23392 20778 23404
rect 21542 23392 21548 23404
rect 21600 23392 21606 23444
rect 24305 23435 24363 23441
rect 24305 23401 24317 23435
rect 24351 23432 24363 23435
rect 24946 23432 24952 23444
rect 24351 23404 24952 23432
rect 24351 23401 24363 23404
rect 24305 23395 24363 23401
rect 24946 23392 24952 23404
rect 25004 23392 25010 23444
rect 10689 23367 10747 23373
rect 10689 23333 10701 23367
rect 10735 23364 10747 23367
rect 10778 23364 10784 23376
rect 10735 23336 10784 23364
rect 10735 23333 10747 23336
rect 10689 23327 10747 23333
rect 10778 23324 10784 23336
rect 10836 23324 10842 23376
rect 10870 23324 10876 23376
rect 10928 23364 10934 23376
rect 11037 23367 11095 23373
rect 11037 23364 11049 23367
rect 10928 23336 11049 23364
rect 10928 23324 10934 23336
rect 11037 23333 11049 23336
rect 11083 23333 11095 23367
rect 11037 23327 11095 23333
rect 15749 23367 15807 23373
rect 15749 23333 15761 23367
rect 15795 23364 15807 23367
rect 15841 23367 15899 23373
rect 15841 23364 15853 23367
rect 15795 23336 15853 23364
rect 15795 23333 15807 23336
rect 15749 23327 15807 23333
rect 15841 23333 15853 23336
rect 15887 23364 15899 23367
rect 16482 23364 16488 23376
rect 15887 23336 16488 23364
rect 15887 23333 15899 23336
rect 15841 23327 15899 23333
rect 16482 23324 16488 23336
rect 16540 23324 16546 23376
rect 18325 23367 18383 23373
rect 18325 23333 18337 23367
rect 18371 23333 18383 23367
rect 18325 23327 18383 23333
rect 10796 23296 10824 23324
rect 10796 23268 13124 23296
rect 11422 23188 11428 23240
rect 11480 23228 11486 23240
rect 13096 23237 13124 23268
rect 16022 23256 16028 23308
rect 16080 23305 16086 23308
rect 16080 23299 16144 23305
rect 16080 23265 16098 23299
rect 16132 23265 16144 23299
rect 16080 23259 16144 23265
rect 16080 23256 16086 23259
rect 18046 23256 18052 23308
rect 18104 23296 18110 23308
rect 18233 23299 18291 23305
rect 18233 23296 18245 23299
rect 18104 23268 18245 23296
rect 18104 23256 18110 23268
rect 18233 23265 18245 23268
rect 18279 23296 18291 23299
rect 18340 23296 18368 23327
rect 18414 23324 18420 23376
rect 18472 23364 18478 23376
rect 18581 23367 18639 23373
rect 18581 23364 18593 23367
rect 18472 23336 18593 23364
rect 18472 23324 18478 23336
rect 18581 23333 18593 23336
rect 18627 23333 18639 23367
rect 24029 23367 24087 23373
rect 24029 23364 24041 23367
rect 18581 23327 18639 23333
rect 23860 23336 24041 23364
rect 19058 23296 19064 23308
rect 18279 23268 19064 23296
rect 18279 23265 18291 23268
rect 18233 23259 18291 23265
rect 19058 23256 19064 23268
rect 19116 23256 19122 23308
rect 21812 23299 21870 23305
rect 21812 23265 21824 23299
rect 21858 23296 21870 23299
rect 22278 23296 22284 23308
rect 21858 23268 22284 23296
rect 21858 23265 21870 23268
rect 21812 23259 21870 23265
rect 22278 23256 22284 23268
rect 22336 23256 22342 23308
rect 23290 23256 23296 23308
rect 23348 23296 23354 23308
rect 23658 23296 23664 23308
rect 23348 23268 23664 23296
rect 23348 23256 23354 23268
rect 23658 23256 23664 23268
rect 23716 23256 23722 23308
rect 23860 23240 23888 23336
rect 24029 23333 24041 23336
rect 24075 23333 24087 23367
rect 25314 23364 25320 23376
rect 25275 23336 25320 23364
rect 24029 23327 24087 23333
rect 25314 23324 25320 23336
rect 25372 23364 25378 23376
rect 25869 23367 25927 23373
rect 25869 23364 25881 23367
rect 25372 23336 25881 23364
rect 25372 23324 25378 23336
rect 25869 23333 25881 23336
rect 25915 23333 25927 23367
rect 25869 23327 25927 23333
rect 12161 23231 12219 23237
rect 12161 23228 12173 23231
rect 11480 23200 12173 23228
rect 11480 23188 11486 23200
rect 12161 23197 12173 23200
rect 12207 23197 12219 23231
rect 12161 23191 12219 23197
rect 13081 23231 13139 23237
rect 13081 23197 13093 23231
rect 13127 23228 13139 23231
rect 13354 23228 13360 23240
rect 13127 23200 13360 23228
rect 13127 23197 13139 23200
rect 13081 23191 13139 23197
rect 13354 23188 13360 23200
rect 13412 23188 13418 23240
rect 13541 23231 13599 23237
rect 13541 23197 13553 23231
rect 13587 23228 13599 23231
rect 13814 23228 13820 23240
rect 13587 23200 13820 23228
rect 13587 23197 13599 23200
rect 13541 23191 13599 23197
rect 13814 23188 13820 23200
rect 13872 23188 13878 23240
rect 13909 23231 13967 23237
rect 13909 23197 13921 23231
rect 13955 23228 13967 23231
rect 14645 23231 14703 23237
rect 14645 23228 14657 23231
rect 13955 23200 14657 23228
rect 13955 23197 13967 23200
rect 13909 23191 13967 23197
rect 14645 23197 14657 23200
rect 14691 23228 14703 23231
rect 14826 23228 14832 23240
rect 14691 23200 14832 23228
rect 14691 23197 14703 23200
rect 14645 23191 14703 23197
rect 14826 23188 14832 23200
rect 14884 23188 14890 23240
rect 17218 23228 17224 23240
rect 17179 23200 17224 23228
rect 17218 23188 17224 23200
rect 17276 23188 17282 23240
rect 22922 23228 22928 23240
rect 22883 23200 22928 23228
rect 22922 23188 22928 23200
rect 22980 23188 22986 23240
rect 23566 23228 23572 23240
rect 23527 23200 23572 23228
rect 23566 23188 23572 23200
rect 23624 23188 23630 23240
rect 23842 23228 23848 23240
rect 23803 23200 23848 23228
rect 23842 23188 23848 23200
rect 23900 23188 23906 23240
rect 24854 23188 24860 23240
rect 24912 23228 24918 23240
rect 24949 23231 25007 23237
rect 24949 23228 24961 23231
rect 24912 23200 24961 23228
rect 24912 23188 24918 23200
rect 24949 23197 24961 23200
rect 24995 23197 25007 23231
rect 24949 23191 25007 23197
rect 1104 23138 26864 23160
rect 1104 23086 10315 23138
rect 10367 23086 10379 23138
rect 10431 23086 10443 23138
rect 10495 23086 10507 23138
rect 10559 23086 19648 23138
rect 19700 23086 19712 23138
rect 19764 23086 19776 23138
rect 19828 23086 19840 23138
rect 19892 23086 26864 23138
rect 1104 23064 26864 23086
rect 8938 22984 8944 23036
rect 8996 23024 9002 23036
rect 9677 23027 9735 23033
rect 9677 23024 9689 23027
rect 8996 22996 9689 23024
rect 8996 22984 9002 22996
rect 9677 22993 9689 22996
rect 9723 23024 9735 23027
rect 10781 23027 10839 23033
rect 10781 23024 10793 23027
rect 9723 22996 10793 23024
rect 9723 22993 9735 22996
rect 9677 22987 9735 22993
rect 10781 22993 10793 22996
rect 10827 22993 10839 23027
rect 10781 22987 10839 22993
rect 11054 22984 11060 23036
rect 11112 23024 11118 23036
rect 11241 23027 11299 23033
rect 11241 23024 11253 23027
rect 11112 22996 11253 23024
rect 11112 22984 11118 22996
rect 11241 22993 11253 22996
rect 11287 23024 11299 23027
rect 11882 23024 11888 23036
rect 11287 22996 11888 23024
rect 11287 22993 11299 22996
rect 11241 22987 11299 22993
rect 11882 22984 11888 22996
rect 11940 22984 11946 23036
rect 14734 23024 14740 23036
rect 14695 22996 14740 23024
rect 14734 22984 14740 22996
rect 14792 22984 14798 23036
rect 16206 22984 16212 23036
rect 16264 23024 16270 23036
rect 16485 23027 16543 23033
rect 16485 23024 16497 23027
rect 16264 22996 16497 23024
rect 16264 22984 16270 22996
rect 16485 22993 16497 22996
rect 16531 22993 16543 23027
rect 16485 22987 16543 22993
rect 18049 23027 18107 23033
rect 18049 22993 18061 23027
rect 18095 23024 18107 23027
rect 18598 23024 18604 23036
rect 18095 22996 18604 23024
rect 18095 22993 18107 22996
rect 18049 22987 18107 22993
rect 18598 22984 18604 22996
rect 18656 22984 18662 23036
rect 19150 23024 19156 23036
rect 19111 22996 19156 23024
rect 19150 22984 19156 22996
rect 19208 22984 19214 23036
rect 19426 23024 19432 23036
rect 19387 22996 19432 23024
rect 19426 22984 19432 22996
rect 19484 22984 19490 23036
rect 9585 22959 9643 22965
rect 9585 22925 9597 22959
rect 9631 22956 9643 22959
rect 9950 22956 9956 22968
rect 9631 22928 9956 22956
rect 9631 22925 9643 22928
rect 9585 22919 9643 22925
rect 9950 22916 9956 22928
rect 10008 22956 10014 22968
rect 10962 22956 10968 22968
rect 10008 22928 10968 22956
rect 10008 22916 10014 22928
rect 10962 22916 10968 22928
rect 11020 22916 11026 22968
rect 13265 22959 13323 22965
rect 13265 22925 13277 22959
rect 13311 22956 13323 22959
rect 13446 22956 13452 22968
rect 13311 22928 13452 22956
rect 13311 22925 13323 22928
rect 13265 22919 13323 22925
rect 13446 22916 13452 22928
rect 13504 22956 13510 22968
rect 13624 22959 13682 22965
rect 13624 22956 13636 22959
rect 13504 22928 13636 22956
rect 13504 22916 13510 22928
rect 13624 22925 13636 22928
rect 13670 22956 13682 22959
rect 14182 22956 14188 22968
rect 13670 22928 14188 22956
rect 13670 22925 13682 22928
rect 13624 22919 13682 22925
rect 14182 22916 14188 22928
rect 14240 22916 14246 22968
rect 18417 22959 18475 22965
rect 18417 22925 18429 22959
rect 18463 22956 18475 22959
rect 18782 22956 18788 22968
rect 18463 22928 18788 22956
rect 18463 22925 18475 22928
rect 18417 22919 18475 22925
rect 18782 22916 18788 22928
rect 18840 22956 18846 22968
rect 19242 22956 19248 22968
rect 18840 22928 19248 22956
rect 18840 22916 18846 22928
rect 19242 22916 19248 22928
rect 19300 22916 19306 22968
rect 11146 22888 11152 22900
rect 11107 22860 11152 22888
rect 11146 22848 11152 22860
rect 11204 22848 11210 22900
rect 18506 22848 18512 22900
rect 18564 22888 18570 22900
rect 18564 22860 18609 22888
rect 18564 22848 18570 22860
rect 19058 22848 19064 22900
rect 19116 22888 19122 22900
rect 20533 22891 20591 22897
rect 20533 22888 20545 22891
rect 19116 22860 20545 22888
rect 19116 22848 19122 22860
rect 20533 22857 20545 22860
rect 20579 22888 20591 22891
rect 20622 22888 20628 22900
rect 20579 22860 20628 22888
rect 20579 22857 20591 22860
rect 20533 22851 20591 22857
rect 20622 22848 20628 22860
rect 20680 22848 20686 22900
rect 20800 22891 20858 22897
rect 20800 22857 20812 22891
rect 20846 22888 20858 22891
rect 21082 22888 21088 22900
rect 20846 22860 21088 22888
rect 20846 22857 20858 22860
rect 20800 22851 20858 22857
rect 21082 22848 21088 22860
rect 21140 22848 21146 22900
rect 23661 22891 23719 22897
rect 23661 22857 23673 22891
rect 23707 22888 23719 22891
rect 23750 22888 23756 22900
rect 23707 22860 23756 22888
rect 23707 22857 23719 22860
rect 23661 22851 23719 22857
rect 23750 22848 23756 22860
rect 23808 22848 23814 22900
rect 24946 22888 24952 22900
rect 24907 22860 24952 22888
rect 24946 22848 24952 22860
rect 25004 22848 25010 22900
rect 9306 22780 9312 22832
rect 9364 22820 9370 22832
rect 9769 22823 9827 22829
rect 9769 22820 9781 22823
rect 9364 22792 9781 22820
rect 9364 22780 9370 22792
rect 9769 22789 9781 22792
rect 9815 22789 9827 22823
rect 11422 22820 11428 22832
rect 11383 22792 11428 22820
rect 9769 22783 9827 22789
rect 11422 22780 11428 22792
rect 11480 22780 11486 22832
rect 13354 22820 13360 22832
rect 13315 22792 13360 22820
rect 13354 22780 13360 22792
rect 13412 22780 13418 22832
rect 15470 22780 15476 22832
rect 15528 22820 15534 22832
rect 16577 22823 16635 22829
rect 16577 22820 16589 22823
rect 15528 22792 16589 22820
rect 15528 22780 15534 22792
rect 16577 22789 16589 22792
rect 16623 22789 16635 22823
rect 16577 22783 16635 22789
rect 16669 22823 16727 22829
rect 16669 22789 16681 22823
rect 16715 22789 16727 22823
rect 16669 22783 16727 22789
rect 18601 22823 18659 22829
rect 18601 22789 18613 22823
rect 18647 22789 18659 22823
rect 18601 22783 18659 22789
rect 23937 22823 23995 22829
rect 23937 22789 23949 22823
rect 23983 22820 23995 22823
rect 24026 22820 24032 22832
rect 23983 22792 24032 22820
rect 23983 22789 23995 22792
rect 23937 22783 23995 22789
rect 9214 22752 9220 22764
rect 9175 22724 9220 22752
rect 9214 22712 9220 22724
rect 9272 22712 9278 22764
rect 16025 22755 16083 22761
rect 16025 22721 16037 22755
rect 16071 22752 16083 22755
rect 16684 22752 16712 22783
rect 17129 22755 17187 22761
rect 17129 22752 17141 22755
rect 16071 22724 17141 22752
rect 16071 22721 16083 22724
rect 16025 22715 16083 22721
rect 17129 22721 17141 22724
rect 17175 22752 17187 22755
rect 17218 22752 17224 22764
rect 17175 22724 17224 22752
rect 17175 22721 17187 22724
rect 17129 22715 17187 22721
rect 17218 22712 17224 22724
rect 17276 22712 17282 22764
rect 18414 22712 18420 22764
rect 18472 22752 18478 22764
rect 18616 22752 18644 22783
rect 24026 22780 24032 22792
rect 24084 22780 24090 22832
rect 18472 22724 18644 22752
rect 18472 22712 18478 22724
rect 15562 22684 15568 22696
rect 15523 22656 15568 22684
rect 15562 22644 15568 22656
rect 15620 22644 15626 22696
rect 16114 22684 16120 22696
rect 16075 22656 16120 22684
rect 16114 22644 16120 22656
rect 16172 22644 16178 22696
rect 20714 22644 20720 22696
rect 20772 22684 20778 22696
rect 21913 22687 21971 22693
rect 21913 22684 21925 22687
rect 20772 22656 21925 22684
rect 20772 22644 20778 22656
rect 21913 22653 21925 22656
rect 21959 22653 21971 22687
rect 21913 22647 21971 22653
rect 23382 22644 23388 22696
rect 23440 22684 23446 22696
rect 23566 22684 23572 22696
rect 23440 22656 23572 22684
rect 23440 22644 23446 22656
rect 23566 22644 23572 22656
rect 23624 22644 23630 22696
rect 25130 22684 25136 22696
rect 25091 22656 25136 22684
rect 25130 22644 25136 22656
rect 25188 22644 25194 22696
rect 1104 22594 26864 22616
rect 1104 22542 5648 22594
rect 5700 22542 5712 22594
rect 5764 22542 5776 22594
rect 5828 22542 5840 22594
rect 5892 22542 14982 22594
rect 15034 22542 15046 22594
rect 15098 22542 15110 22594
rect 15162 22542 15174 22594
rect 15226 22542 24315 22594
rect 24367 22542 24379 22594
rect 24431 22542 24443 22594
rect 24495 22542 24507 22594
rect 24559 22542 26864 22594
rect 1104 22520 26864 22542
rect 8938 22480 8944 22492
rect 8899 22452 8944 22480
rect 8938 22440 8944 22452
rect 8996 22440 9002 22492
rect 9950 22480 9956 22492
rect 9911 22452 9956 22480
rect 9950 22440 9956 22452
rect 10008 22440 10014 22492
rect 10689 22483 10747 22489
rect 10689 22449 10701 22483
rect 10735 22480 10747 22483
rect 11054 22480 11060 22492
rect 10735 22452 11060 22480
rect 10735 22449 10747 22452
rect 10689 22443 10747 22449
rect 11054 22440 11060 22452
rect 11112 22440 11118 22492
rect 13354 22480 13360 22492
rect 13315 22452 13360 22480
rect 13354 22440 13360 22452
rect 13412 22440 13418 22492
rect 14734 22440 14740 22492
rect 14792 22480 14798 22492
rect 15013 22483 15071 22489
rect 15013 22480 15025 22483
rect 14792 22452 15025 22480
rect 14792 22440 14798 22452
rect 15013 22449 15025 22452
rect 15059 22449 15071 22483
rect 15470 22480 15476 22492
rect 15431 22452 15476 22480
rect 15013 22443 15071 22449
rect 10778 22344 10784 22356
rect 10739 22316 10784 22344
rect 10778 22304 10784 22316
rect 10836 22304 10842 22356
rect 13814 22304 13820 22356
rect 13872 22344 13878 22356
rect 14001 22347 14059 22353
rect 14001 22344 14013 22347
rect 13872 22316 14013 22344
rect 13872 22304 13878 22316
rect 14001 22313 14013 22316
rect 14047 22313 14059 22347
rect 14001 22307 14059 22313
rect 14090 22304 14096 22356
rect 14148 22344 14154 22356
rect 15028 22344 15056 22443
rect 15470 22440 15476 22452
rect 15528 22440 15534 22492
rect 16206 22440 16212 22492
rect 16264 22480 16270 22492
rect 16485 22483 16543 22489
rect 16485 22480 16497 22483
rect 16264 22452 16497 22480
rect 16264 22440 16270 22452
rect 16485 22449 16497 22452
rect 16531 22449 16543 22483
rect 18414 22480 18420 22492
rect 18375 22452 18420 22480
rect 16485 22443 16543 22449
rect 18414 22440 18420 22452
rect 18472 22480 18478 22492
rect 19337 22483 19395 22489
rect 19337 22480 19349 22483
rect 18472 22452 19349 22480
rect 18472 22440 18478 22452
rect 19337 22449 19349 22452
rect 19383 22449 19395 22483
rect 20622 22480 20628 22492
rect 20583 22452 20628 22480
rect 19337 22443 19395 22449
rect 20622 22440 20628 22452
rect 20680 22440 20686 22492
rect 21082 22480 21088 22492
rect 21043 22452 21088 22480
rect 21082 22440 21088 22452
rect 21140 22440 21146 22492
rect 23658 22480 23664 22492
rect 23619 22452 23664 22480
rect 23658 22440 23664 22452
rect 23716 22440 23722 22492
rect 24946 22440 24952 22492
rect 25004 22480 25010 22492
rect 25498 22480 25504 22492
rect 25004 22452 25504 22480
rect 25004 22440 25010 22452
rect 25498 22440 25504 22452
rect 25556 22440 25562 22492
rect 18506 22372 18512 22424
rect 18564 22412 18570 22424
rect 18969 22415 19027 22421
rect 18969 22412 18981 22415
rect 18564 22384 18981 22412
rect 18564 22372 18570 22384
rect 18969 22381 18981 22384
rect 19015 22381 19027 22415
rect 18969 22375 19027 22381
rect 21729 22415 21787 22421
rect 21729 22381 21741 22415
rect 21775 22412 21787 22415
rect 23750 22412 23756 22424
rect 21775 22384 23756 22412
rect 21775 22381 21787 22384
rect 21729 22375 21787 22381
rect 23750 22372 23756 22384
rect 23808 22412 23814 22424
rect 24029 22415 24087 22421
rect 24029 22412 24041 22415
rect 23808 22384 24041 22412
rect 23808 22372 23814 22384
rect 24029 22381 24041 22384
rect 24075 22381 24087 22415
rect 24029 22375 24087 22381
rect 15933 22347 15991 22353
rect 15933 22344 15945 22347
rect 14148 22316 14193 22344
rect 15028 22316 15945 22344
rect 14148 22304 14154 22316
rect 15933 22313 15945 22316
rect 15979 22313 15991 22347
rect 15933 22307 15991 22313
rect 16022 22304 16028 22356
rect 16080 22344 16086 22356
rect 19794 22344 19800 22356
rect 16080 22316 16173 22344
rect 19755 22316 19800 22344
rect 16080 22304 16086 22316
rect 19794 22304 19800 22316
rect 19852 22304 19858 22356
rect 22373 22347 22431 22353
rect 22373 22313 22385 22347
rect 22419 22344 22431 22347
rect 22557 22347 22615 22353
rect 22557 22344 22569 22347
rect 22419 22316 22569 22344
rect 22419 22313 22431 22316
rect 22373 22307 22431 22313
rect 22557 22313 22569 22316
rect 22603 22344 22615 22347
rect 22922 22344 22928 22356
rect 22603 22316 22928 22344
rect 22603 22313 22615 22316
rect 22557 22307 22615 22313
rect 22922 22304 22928 22316
rect 22980 22304 22986 22356
rect 11048 22279 11106 22285
rect 11048 22245 11060 22279
rect 11094 22276 11106 22279
rect 11422 22276 11428 22288
rect 11094 22248 11428 22276
rect 11094 22245 11106 22248
rect 11048 22239 11106 22245
rect 11422 22236 11428 22248
rect 11480 22236 11486 22288
rect 15562 22236 15568 22288
rect 15620 22276 15626 22288
rect 15838 22276 15844 22288
rect 15620 22248 15844 22276
rect 15620 22236 15626 22248
rect 15838 22236 15844 22248
rect 15896 22236 15902 22288
rect 16040 22276 16068 22304
rect 15948 22248 16068 22276
rect 13909 22211 13967 22217
rect 13909 22208 13921 22211
rect 9232 22180 12204 22208
rect 9232 22152 9260 22180
rect 9214 22140 9220 22152
rect 9175 22112 9220 22140
rect 9214 22100 9220 22112
rect 9272 22100 9278 22152
rect 10321 22143 10379 22149
rect 10321 22109 10333 22143
rect 10367 22140 10379 22143
rect 11146 22140 11152 22152
rect 10367 22112 11152 22140
rect 10367 22109 10379 22112
rect 10321 22103 10379 22109
rect 11146 22100 11152 22112
rect 11204 22100 11210 22152
rect 12176 22149 12204 22180
rect 13096 22180 13921 22208
rect 13096 22152 13124 22180
rect 13909 22177 13921 22180
rect 13955 22177 13967 22211
rect 13909 22171 13967 22177
rect 14737 22211 14795 22217
rect 14737 22177 14749 22211
rect 14783 22208 14795 22211
rect 15948 22208 15976 22248
rect 16482 22236 16488 22288
rect 16540 22276 16546 22288
rect 16945 22279 17003 22285
rect 16945 22276 16957 22279
rect 16540 22248 16957 22276
rect 16540 22236 16546 22248
rect 16945 22245 16957 22248
rect 16991 22276 17003 22279
rect 17037 22279 17095 22285
rect 17037 22276 17049 22279
rect 16991 22248 17049 22276
rect 16991 22245 17003 22248
rect 16945 22239 17003 22245
rect 17037 22245 17049 22248
rect 17083 22276 17095 22279
rect 18046 22276 18052 22288
rect 17083 22248 18052 22276
rect 17083 22245 17095 22248
rect 17037 22239 17095 22245
rect 18046 22236 18052 22248
rect 18104 22236 18110 22288
rect 19334 22236 19340 22288
rect 19392 22276 19398 22288
rect 19521 22279 19579 22285
rect 19521 22276 19533 22279
rect 19392 22248 19533 22276
rect 19392 22236 19398 22248
rect 19521 22245 19533 22248
rect 19567 22245 19579 22279
rect 23477 22279 23535 22285
rect 23477 22276 23489 22279
rect 19521 22239 19579 22245
rect 23308 22248 23489 22276
rect 14783 22180 15976 22208
rect 14783 22177 14795 22180
rect 14737 22171 14795 22177
rect 17218 22168 17224 22220
rect 17276 22217 17282 22220
rect 17276 22211 17340 22217
rect 17276 22177 17294 22211
rect 17328 22177 17340 22211
rect 17276 22171 17340 22177
rect 21637 22211 21695 22217
rect 21637 22177 21649 22211
rect 21683 22208 21695 22211
rect 22002 22208 22008 22220
rect 21683 22180 22008 22208
rect 21683 22177 21695 22180
rect 21637 22171 21695 22177
rect 17276 22168 17282 22171
rect 22002 22168 22008 22180
rect 22060 22208 22066 22220
rect 22097 22211 22155 22217
rect 22097 22208 22109 22211
rect 22060 22180 22109 22208
rect 22060 22168 22066 22180
rect 22097 22177 22109 22180
rect 22143 22177 22155 22211
rect 22097 22171 22155 22177
rect 22186 22168 22192 22220
rect 22244 22208 22250 22220
rect 22741 22211 22799 22217
rect 22741 22208 22753 22211
rect 22244 22180 22753 22208
rect 22244 22168 22250 22180
rect 22741 22177 22753 22180
rect 22787 22177 22799 22211
rect 22741 22171 22799 22177
rect 23308 22152 23336 22248
rect 23477 22245 23489 22248
rect 23523 22245 23535 22279
rect 24578 22276 24584 22288
rect 24539 22248 24584 22276
rect 23477 22239 23535 22245
rect 24578 22236 24584 22248
rect 24636 22276 24642 22288
rect 25133 22279 25191 22285
rect 25133 22276 25145 22279
rect 24636 22248 25145 22276
rect 24636 22236 24642 22248
rect 25133 22245 25145 22248
rect 25179 22245 25191 22279
rect 25133 22239 25191 22245
rect 12161 22143 12219 22149
rect 12161 22109 12173 22143
rect 12207 22109 12219 22143
rect 13078 22140 13084 22152
rect 13039 22112 13084 22140
rect 12161 22103 12219 22109
rect 13078 22100 13084 22112
rect 13136 22100 13142 22152
rect 13538 22140 13544 22152
rect 13499 22112 13544 22140
rect 13538 22100 13544 22112
rect 13596 22100 13602 22152
rect 21082 22100 21088 22152
rect 21140 22140 21146 22152
rect 22370 22140 22376 22152
rect 21140 22112 22376 22140
rect 21140 22100 21146 22112
rect 22370 22100 22376 22112
rect 22428 22140 22434 22152
rect 22557 22143 22615 22149
rect 22557 22140 22569 22143
rect 22428 22112 22569 22140
rect 22428 22100 22434 22112
rect 22557 22109 22569 22112
rect 22603 22109 22615 22143
rect 23290 22140 23296 22152
rect 23251 22112 23296 22140
rect 22557 22103 22615 22109
rect 23290 22100 23296 22112
rect 23348 22100 23354 22152
rect 24762 22140 24768 22152
rect 24723 22112 24768 22140
rect 24762 22100 24768 22112
rect 24820 22100 24826 22152
rect 1104 22050 26864 22072
rect 1104 21998 10315 22050
rect 10367 21998 10379 22050
rect 10431 21998 10443 22050
rect 10495 21998 10507 22050
rect 10559 21998 19648 22050
rect 19700 21998 19712 22050
rect 19764 21998 19776 22050
rect 19828 21998 19840 22050
rect 19892 21998 26864 22050
rect 1104 21976 26864 21998
rect 10778 21936 10784 21948
rect 10739 21908 10784 21936
rect 10778 21896 10784 21908
rect 10836 21896 10842 21948
rect 11241 21939 11299 21945
rect 11241 21905 11253 21939
rect 11287 21936 11299 21939
rect 11422 21936 11428 21948
rect 11287 21908 11428 21936
rect 11287 21905 11299 21908
rect 11241 21899 11299 21905
rect 11422 21896 11428 21908
rect 11480 21936 11486 21948
rect 11517 21939 11575 21945
rect 11517 21936 11529 21939
rect 11480 21908 11529 21936
rect 11480 21896 11486 21908
rect 11517 21905 11529 21908
rect 11563 21905 11575 21939
rect 11517 21899 11575 21905
rect 13078 21896 13084 21948
rect 13136 21936 13142 21948
rect 13541 21939 13599 21945
rect 13541 21936 13553 21939
rect 13136 21908 13553 21936
rect 13136 21896 13142 21908
rect 13541 21905 13553 21908
rect 13587 21905 13599 21939
rect 13541 21899 13599 21905
rect 13814 21896 13820 21948
rect 13872 21936 13878 21948
rect 14369 21939 14427 21945
rect 14369 21936 14381 21939
rect 13872 21908 14381 21936
rect 13872 21896 13878 21908
rect 14369 21905 14381 21908
rect 14415 21905 14427 21939
rect 14369 21899 14427 21905
rect 15381 21939 15439 21945
rect 15381 21905 15393 21939
rect 15427 21936 15439 21939
rect 15470 21936 15476 21948
rect 15427 21908 15476 21936
rect 15427 21905 15439 21908
rect 15381 21899 15439 21905
rect 15470 21896 15476 21908
rect 15528 21896 15534 21948
rect 16022 21896 16028 21948
rect 16080 21936 16086 21948
rect 16853 21939 16911 21945
rect 16853 21936 16865 21939
rect 16080 21908 16865 21936
rect 16080 21896 16086 21908
rect 16853 21905 16865 21908
rect 16899 21905 16911 21939
rect 18782 21936 18788 21948
rect 18743 21908 18788 21936
rect 16853 21899 16911 21905
rect 18782 21896 18788 21908
rect 18840 21896 18846 21948
rect 19334 21896 19340 21948
rect 19392 21936 19398 21948
rect 19521 21939 19579 21945
rect 19521 21936 19533 21939
rect 19392 21908 19533 21936
rect 19392 21896 19398 21908
rect 19521 21905 19533 21908
rect 19567 21905 19579 21939
rect 19521 21899 19579 21905
rect 21913 21939 21971 21945
rect 21913 21905 21925 21939
rect 21959 21936 21971 21939
rect 22002 21936 22008 21948
rect 21959 21908 22008 21936
rect 21959 21905 21971 21908
rect 21913 21899 21971 21905
rect 22002 21896 22008 21908
rect 22060 21896 22066 21948
rect 13446 21868 13452 21880
rect 13407 21840 13452 21868
rect 13446 21828 13452 21840
rect 13504 21828 13510 21880
rect 14090 21868 14096 21880
rect 14051 21840 14096 21868
rect 14090 21828 14096 21840
rect 14148 21828 14154 21880
rect 21729 21871 21787 21877
rect 21729 21837 21741 21871
rect 21775 21868 21787 21871
rect 22370 21868 22376 21880
rect 21775 21840 22376 21868
rect 21775 21837 21787 21840
rect 21729 21831 21787 21837
rect 22370 21828 22376 21840
rect 22428 21828 22434 21880
rect 15473 21803 15531 21809
rect 15473 21769 15485 21803
rect 15519 21800 15531 21803
rect 15562 21800 15568 21812
rect 15519 21772 15568 21800
rect 15519 21769 15531 21772
rect 15473 21763 15531 21769
rect 15562 21760 15568 21772
rect 15620 21760 15626 21812
rect 15746 21809 15752 21812
rect 15740 21800 15752 21809
rect 15707 21772 15752 21800
rect 15740 21763 15752 21772
rect 15746 21760 15752 21763
rect 15804 21760 15810 21812
rect 18046 21800 18052 21812
rect 18007 21772 18052 21800
rect 18046 21760 18052 21772
rect 18104 21760 18110 21812
rect 18322 21800 18328 21812
rect 18283 21772 18328 21800
rect 18322 21760 18328 21772
rect 18380 21760 18386 21812
rect 24581 21803 24639 21809
rect 24581 21800 24593 21803
rect 24136 21772 24593 21800
rect 24136 21744 24164 21772
rect 24581 21769 24593 21772
rect 24627 21769 24639 21803
rect 24581 21763 24639 21769
rect 24670 21760 24676 21812
rect 24728 21760 24734 21812
rect 24118 21692 24124 21744
rect 24176 21692 24182 21744
rect 24210 21692 24216 21744
rect 24268 21732 24274 21744
rect 24688 21732 24716 21760
rect 24268 21704 24716 21732
rect 24268 21692 24274 21704
rect 19242 21664 19248 21676
rect 19203 21636 19248 21664
rect 19242 21624 19248 21636
rect 19300 21624 19306 21676
rect 23477 21599 23535 21605
rect 23477 21565 23489 21599
rect 23523 21596 23535 21599
rect 23842 21596 23848 21608
rect 23523 21568 23848 21596
rect 23523 21565 23535 21568
rect 23477 21559 23535 21565
rect 23842 21556 23848 21568
rect 23900 21556 23906 21608
rect 24762 21596 24768 21608
rect 24723 21568 24768 21596
rect 24762 21556 24768 21568
rect 24820 21556 24826 21608
rect 1104 21506 26864 21528
rect 1104 21454 5648 21506
rect 5700 21454 5712 21506
rect 5764 21454 5776 21506
rect 5828 21454 5840 21506
rect 5892 21454 14982 21506
rect 15034 21454 15046 21506
rect 15098 21454 15110 21506
rect 15162 21454 15174 21506
rect 15226 21454 24315 21506
rect 24367 21454 24379 21506
rect 24431 21454 24443 21506
rect 24495 21454 24507 21506
rect 24559 21454 26864 21506
rect 1104 21432 26864 21454
rect 10321 21395 10379 21401
rect 10321 21361 10333 21395
rect 10367 21392 10379 21395
rect 10778 21392 10784 21404
rect 10367 21364 10784 21392
rect 10367 21361 10379 21364
rect 10321 21355 10379 21361
rect 10428 21265 10456 21364
rect 10778 21352 10784 21364
rect 10836 21352 10842 21404
rect 22278 21392 22284 21404
rect 22239 21364 22284 21392
rect 22278 21352 22284 21364
rect 22336 21352 22342 21404
rect 23750 21352 23756 21404
rect 23808 21352 23814 21404
rect 24118 21352 24124 21404
rect 24176 21392 24182 21404
rect 24581 21395 24639 21401
rect 24581 21392 24593 21395
rect 24176 21364 24593 21392
rect 24176 21352 24182 21364
rect 24581 21361 24593 21364
rect 24627 21361 24639 21395
rect 24581 21355 24639 21361
rect 16669 21327 16727 21333
rect 16669 21293 16681 21327
rect 16715 21324 16727 21327
rect 18046 21324 18052 21336
rect 16715 21296 18052 21324
rect 16715 21293 16727 21296
rect 16669 21287 16727 21293
rect 18046 21284 18052 21296
rect 18104 21284 18110 21336
rect 23768 21324 23796 21352
rect 24762 21324 24768 21336
rect 23768 21296 24768 21324
rect 24762 21284 24768 21296
rect 24820 21284 24826 21336
rect 10413 21259 10471 21265
rect 10413 21225 10425 21259
rect 10459 21225 10471 21259
rect 14182 21256 14188 21268
rect 14143 21228 14188 21256
rect 10413 21219 10471 21225
rect 14182 21216 14188 21228
rect 14240 21216 14246 21268
rect 15105 21259 15163 21265
rect 15105 21225 15117 21259
rect 15151 21256 15163 21259
rect 15746 21256 15752 21268
rect 15151 21228 15752 21256
rect 15151 21225 15163 21228
rect 15105 21219 15163 21225
rect 15746 21216 15752 21228
rect 15804 21256 15810 21268
rect 16209 21259 16267 21265
rect 16209 21256 16221 21259
rect 15804 21228 16221 21256
rect 15804 21216 15810 21228
rect 16209 21225 16221 21228
rect 16255 21256 16267 21259
rect 17313 21259 17371 21265
rect 17313 21256 17325 21259
rect 16255 21228 17325 21256
rect 16255 21225 16267 21228
rect 16209 21219 16267 21225
rect 17313 21225 17325 21228
rect 17359 21256 17371 21259
rect 17678 21256 17684 21268
rect 17359 21228 17684 21256
rect 17359 21225 17371 21228
rect 17313 21219 17371 21225
rect 17678 21216 17684 21228
rect 17736 21216 17742 21268
rect 19242 21216 19248 21268
rect 19300 21256 19306 21268
rect 19429 21259 19487 21265
rect 19429 21256 19441 21259
rect 19300 21228 19441 21256
rect 19300 21216 19306 21228
rect 19429 21225 19441 21228
rect 19475 21225 19487 21259
rect 19429 21219 19487 21225
rect 23750 21216 23756 21268
rect 23808 21256 23814 21268
rect 23937 21259 23995 21265
rect 23937 21256 23949 21259
rect 23808 21228 23949 21256
rect 23808 21216 23814 21228
rect 23937 21225 23949 21228
rect 23983 21225 23995 21259
rect 23937 21219 23995 21225
rect 13909 21191 13967 21197
rect 13909 21157 13921 21191
rect 13955 21188 13967 21191
rect 13998 21188 14004 21200
rect 13955 21160 14004 21188
rect 13955 21157 13967 21160
rect 13909 21151 13967 21157
rect 13998 21148 14004 21160
rect 14056 21188 14062 21200
rect 14645 21191 14703 21197
rect 14645 21188 14657 21191
rect 14056 21160 14657 21188
rect 14056 21148 14062 21160
rect 14645 21157 14657 21160
rect 14691 21157 14703 21191
rect 19150 21188 19156 21200
rect 14645 21151 14703 21157
rect 18340 21160 19156 21188
rect 10686 21129 10692 21132
rect 10680 21120 10692 21129
rect 10647 21092 10692 21120
rect 10680 21083 10692 21092
rect 10686 21080 10692 21083
rect 10744 21080 10750 21132
rect 16577 21123 16635 21129
rect 16577 21089 16589 21123
rect 16623 21120 16635 21123
rect 16623 21092 16896 21120
rect 16623 21089 16635 21092
rect 16577 21083 16635 21089
rect 16868 21064 16896 21092
rect 18340 21064 18368 21160
rect 19150 21148 19156 21160
rect 19208 21148 19214 21200
rect 20806 21148 20812 21200
rect 20864 21188 20870 21200
rect 20901 21191 20959 21197
rect 20901 21188 20913 21191
rect 20864 21160 20913 21188
rect 20864 21148 20870 21160
rect 20901 21157 20913 21160
rect 20947 21188 20959 21191
rect 22094 21188 22100 21200
rect 20947 21160 22100 21188
rect 20947 21157 20959 21160
rect 20901 21151 20959 21157
rect 22094 21148 22100 21160
rect 22152 21148 22158 21200
rect 24946 21188 24952 21200
rect 24907 21160 24952 21188
rect 24946 21148 24952 21160
rect 25004 21188 25010 21200
rect 25501 21191 25559 21197
rect 25501 21188 25513 21191
rect 25004 21160 25513 21188
rect 25004 21148 25010 21160
rect 25501 21157 25513 21160
rect 25547 21157 25559 21191
rect 25501 21151 25559 21157
rect 18690 21120 18696 21132
rect 18651 21092 18696 21120
rect 18690 21080 18696 21092
rect 18748 21120 18754 21132
rect 21174 21129 21180 21132
rect 19337 21123 19395 21129
rect 19337 21120 19349 21123
rect 18748 21092 19349 21120
rect 18748 21080 18754 21092
rect 19337 21089 19349 21092
rect 19383 21089 19395 21123
rect 21168 21120 21180 21129
rect 21135 21092 21180 21120
rect 19337 21083 19395 21089
rect 21168 21083 21180 21092
rect 21174 21080 21180 21083
rect 21232 21080 21238 21132
rect 23753 21123 23811 21129
rect 23753 21120 23765 21123
rect 23216 21092 23765 21120
rect 23216 21064 23244 21092
rect 23753 21089 23765 21092
rect 23799 21089 23811 21123
rect 23753 21083 23811 21089
rect 11790 21052 11796 21064
rect 11751 21024 11796 21052
rect 11790 21012 11796 21024
rect 11848 21012 11854 21064
rect 12897 21055 12955 21061
rect 12897 21021 12909 21055
rect 12943 21052 12955 21055
rect 13170 21052 13176 21064
rect 12943 21024 13176 21052
rect 12943 21021 12955 21024
rect 12897 21015 12955 21021
rect 13170 21012 13176 21024
rect 13228 21012 13234 21064
rect 15562 21052 15568 21064
rect 15523 21024 15568 21052
rect 15562 21012 15568 21024
rect 15620 21012 15626 21064
rect 16850 21012 16856 21064
rect 16908 21052 16914 21064
rect 17037 21055 17095 21061
rect 17037 21052 17049 21055
rect 16908 21024 17049 21052
rect 16908 21012 16914 21024
rect 17037 21021 17049 21024
rect 17083 21021 17095 21055
rect 17037 21015 17095 21021
rect 17126 21012 17132 21064
rect 17184 21052 17190 21064
rect 17681 21055 17739 21061
rect 17681 21052 17693 21055
rect 17184 21024 17693 21052
rect 17184 21012 17190 21024
rect 17681 21021 17693 21024
rect 17727 21021 17739 21055
rect 18322 21052 18328 21064
rect 18283 21024 18328 21052
rect 17681 21015 17739 21021
rect 18322 21012 18328 21024
rect 18380 21012 18386 21064
rect 18874 21052 18880 21064
rect 18835 21024 18880 21052
rect 18874 21012 18880 21024
rect 18932 21012 18938 21064
rect 19150 21012 19156 21064
rect 19208 21052 19214 21064
rect 19245 21055 19303 21061
rect 19245 21052 19257 21055
rect 19208 21024 19257 21052
rect 19208 21012 19214 21024
rect 19245 21021 19257 21024
rect 19291 21021 19303 21055
rect 20714 21052 20720 21064
rect 20675 21024 20720 21052
rect 19245 21015 19303 21021
rect 20714 21012 20720 21024
rect 20772 21012 20778 21064
rect 23198 21052 23204 21064
rect 23159 21024 23204 21052
rect 23198 21012 23204 21024
rect 23256 21012 23262 21064
rect 23385 21055 23443 21061
rect 23385 21021 23397 21055
rect 23431 21052 23443 21055
rect 23474 21052 23480 21064
rect 23431 21024 23480 21052
rect 23431 21021 23443 21024
rect 23385 21015 23443 21021
rect 23474 21012 23480 21024
rect 23532 21012 23538 21064
rect 23842 21052 23848 21064
rect 23803 21024 23848 21052
rect 23842 21012 23848 21024
rect 23900 21012 23906 21064
rect 25130 21052 25136 21064
rect 25091 21024 25136 21052
rect 25130 21012 25136 21024
rect 25188 21012 25194 21064
rect 1104 20962 26864 20984
rect 1104 20910 10315 20962
rect 10367 20910 10379 20962
rect 10431 20910 10443 20962
rect 10495 20910 10507 20962
rect 10559 20910 19648 20962
rect 19700 20910 19712 20962
rect 19764 20910 19776 20962
rect 19828 20910 19840 20962
rect 19892 20910 26864 20962
rect 1104 20888 26864 20910
rect 10505 20851 10563 20857
rect 10505 20817 10517 20851
rect 10551 20848 10563 20851
rect 10686 20848 10692 20860
rect 10551 20820 10692 20848
rect 10551 20817 10563 20820
rect 10505 20811 10563 20817
rect 10686 20808 10692 20820
rect 10744 20808 10750 20860
rect 10781 20851 10839 20857
rect 10781 20817 10793 20851
rect 10827 20848 10839 20851
rect 12894 20848 12900 20860
rect 10827 20820 12900 20848
rect 10827 20817 10839 20820
rect 10781 20811 10839 20817
rect 12894 20808 12900 20820
rect 12952 20808 12958 20860
rect 13998 20848 14004 20860
rect 13959 20820 14004 20848
rect 13998 20808 14004 20820
rect 14056 20808 14062 20860
rect 16117 20851 16175 20857
rect 16117 20817 16129 20851
rect 16163 20848 16175 20851
rect 17126 20848 17132 20860
rect 16163 20820 17132 20848
rect 16163 20817 16175 20820
rect 16117 20811 16175 20817
rect 17126 20808 17132 20820
rect 17184 20808 17190 20860
rect 18046 20808 18052 20860
rect 18104 20848 18110 20860
rect 18233 20851 18291 20857
rect 18233 20848 18245 20851
rect 18104 20820 18245 20848
rect 18104 20808 18110 20820
rect 18233 20817 18245 20820
rect 18279 20817 18291 20851
rect 18874 20848 18880 20860
rect 18835 20820 18880 20848
rect 18233 20811 18291 20817
rect 18874 20808 18880 20820
rect 18932 20848 18938 20860
rect 19334 20848 19340 20860
rect 18932 20820 19340 20848
rect 18932 20808 18938 20820
rect 19334 20808 19340 20820
rect 19392 20808 19398 20860
rect 19426 20808 19432 20860
rect 19484 20848 19490 20860
rect 20349 20851 20407 20857
rect 20349 20848 20361 20851
rect 19484 20820 20361 20848
rect 19484 20808 19490 20820
rect 20349 20817 20361 20820
rect 20395 20817 20407 20851
rect 22002 20848 22008 20860
rect 21963 20820 22008 20848
rect 20349 20811 20407 20817
rect 22002 20808 22008 20820
rect 22060 20808 22066 20860
rect 22186 20808 22192 20860
rect 22244 20848 22250 20860
rect 22373 20851 22431 20857
rect 22373 20848 22385 20851
rect 22244 20820 22385 20848
rect 22244 20808 22250 20820
rect 22373 20817 22385 20820
rect 22419 20817 22431 20851
rect 22373 20811 22431 20817
rect 10962 20740 10968 20792
rect 11020 20780 11026 20792
rect 11238 20780 11244 20792
rect 11020 20752 11244 20780
rect 11020 20740 11026 20752
rect 11238 20740 11244 20752
rect 11296 20740 11302 20792
rect 19242 20789 19248 20792
rect 19236 20780 19248 20789
rect 19203 20752 19248 20780
rect 19236 20743 19248 20752
rect 19242 20740 19248 20743
rect 19300 20740 19306 20792
rect 20993 20783 21051 20789
rect 20993 20749 21005 20783
rect 21039 20780 21051 20783
rect 21174 20780 21180 20792
rect 21039 20752 21180 20780
rect 21039 20749 21051 20752
rect 20993 20743 21051 20749
rect 21174 20740 21180 20752
rect 21232 20780 21238 20792
rect 23477 20783 23535 20789
rect 23477 20780 23489 20783
rect 21232 20752 23489 20780
rect 21232 20740 21238 20752
rect 23477 20749 23489 20752
rect 23523 20780 23535 20783
rect 23750 20780 23756 20792
rect 23523 20752 23756 20780
rect 23523 20749 23535 20752
rect 23477 20743 23535 20749
rect 23750 20740 23756 20752
rect 23808 20740 23814 20792
rect 23928 20783 23986 20789
rect 23928 20749 23940 20783
rect 23974 20780 23986 20783
rect 24118 20780 24124 20792
rect 23974 20752 24124 20780
rect 23974 20749 23986 20752
rect 23928 20743 23986 20749
rect 24118 20740 24124 20752
rect 24176 20740 24182 20792
rect 11146 20712 11152 20724
rect 11107 20684 11152 20712
rect 11146 20672 11152 20684
rect 11204 20672 11210 20724
rect 12805 20715 12863 20721
rect 12805 20681 12817 20715
rect 12851 20712 12863 20715
rect 13170 20712 13176 20724
rect 12851 20684 13176 20712
rect 12851 20681 12863 20684
rect 12805 20675 12863 20681
rect 13170 20672 13176 20684
rect 13228 20672 13234 20724
rect 14366 20712 14372 20724
rect 14327 20684 14372 20712
rect 14366 20672 14372 20684
rect 14424 20672 14430 20724
rect 16390 20672 16396 20724
rect 16448 20712 16454 20724
rect 16485 20715 16543 20721
rect 16485 20712 16497 20715
rect 16448 20684 16497 20712
rect 16448 20672 16454 20684
rect 16485 20681 16497 20684
rect 16531 20681 16543 20715
rect 20714 20712 20720 20724
rect 16485 20675 16543 20681
rect 18984 20684 20720 20712
rect 11425 20647 11483 20653
rect 11425 20613 11437 20647
rect 11471 20644 11483 20647
rect 11790 20644 11796 20656
rect 11471 20616 11796 20644
rect 11471 20613 11483 20616
rect 11425 20607 11483 20613
rect 11790 20604 11796 20616
rect 11848 20604 11854 20656
rect 12894 20644 12900 20656
rect 12855 20616 12900 20644
rect 12894 20604 12900 20616
rect 12952 20604 12958 20656
rect 12986 20604 12992 20656
rect 13044 20644 13050 20656
rect 14458 20644 14464 20656
rect 13044 20616 13089 20644
rect 14419 20616 14464 20644
rect 13044 20604 13050 20616
rect 14458 20604 14464 20616
rect 14516 20604 14522 20656
rect 14642 20644 14648 20656
rect 14603 20616 14648 20644
rect 14642 20604 14648 20616
rect 14700 20604 14706 20656
rect 16114 20604 16120 20656
rect 16172 20644 16178 20656
rect 16577 20647 16635 20653
rect 16577 20644 16589 20647
rect 16172 20616 16589 20644
rect 16172 20604 16178 20616
rect 16577 20613 16589 20616
rect 16623 20613 16635 20647
rect 16577 20607 16635 20613
rect 16761 20647 16819 20653
rect 16761 20613 16773 20647
rect 16807 20644 16819 20647
rect 17129 20647 17187 20653
rect 17129 20644 17141 20647
rect 16807 20616 17141 20644
rect 16807 20613 16819 20616
rect 16761 20607 16819 20613
rect 17129 20613 17141 20616
rect 17175 20613 17187 20647
rect 17129 20607 17187 20613
rect 16025 20579 16083 20585
rect 16025 20545 16037 20579
rect 16071 20576 16083 20579
rect 16482 20576 16488 20588
rect 16071 20548 16488 20576
rect 16071 20545 16083 20548
rect 16025 20539 16083 20545
rect 16482 20536 16488 20548
rect 16540 20576 16546 20588
rect 16776 20576 16804 20607
rect 18690 20604 18696 20656
rect 18748 20644 18754 20656
rect 18984 20653 19012 20684
rect 20714 20672 20720 20684
rect 20772 20672 20778 20724
rect 22462 20712 22468 20724
rect 22423 20684 22468 20712
rect 22462 20672 22468 20684
rect 22520 20672 22526 20724
rect 18969 20647 19027 20653
rect 18969 20644 18981 20647
rect 18748 20616 18981 20644
rect 18748 20604 18754 20616
rect 18969 20613 18981 20616
rect 19015 20613 19027 20647
rect 18969 20607 19027 20613
rect 22649 20647 22707 20653
rect 22649 20613 22661 20647
rect 22695 20613 22707 20647
rect 23658 20644 23664 20656
rect 23619 20616 23664 20644
rect 22649 20607 22707 20613
rect 16540 20548 16804 20576
rect 16540 20536 16546 20548
rect 22664 20520 22692 20607
rect 23658 20604 23664 20616
rect 23716 20604 23722 20656
rect 12437 20511 12495 20517
rect 12437 20477 12449 20511
rect 12483 20508 12495 20511
rect 13722 20508 13728 20520
rect 12483 20480 13728 20508
rect 12483 20477 12495 20480
rect 12437 20471 12495 20477
rect 13722 20468 13728 20480
rect 13780 20468 13786 20520
rect 22646 20508 22652 20520
rect 22559 20480 22652 20508
rect 22646 20468 22652 20480
rect 22704 20508 22710 20520
rect 25041 20511 25099 20517
rect 25041 20508 25053 20511
rect 22704 20480 25053 20508
rect 22704 20468 22710 20480
rect 25041 20477 25053 20480
rect 25087 20477 25099 20511
rect 25041 20471 25099 20477
rect 1104 20418 26864 20440
rect 1104 20366 5648 20418
rect 5700 20366 5712 20418
rect 5764 20366 5776 20418
rect 5828 20366 5840 20418
rect 5892 20366 14982 20418
rect 15034 20366 15046 20418
rect 15098 20366 15110 20418
rect 15162 20366 15174 20418
rect 15226 20366 24315 20418
rect 24367 20366 24379 20418
rect 24431 20366 24443 20418
rect 24495 20366 24507 20418
rect 24559 20366 26864 20418
rect 1104 20344 26864 20366
rect 10873 20307 10931 20313
rect 10873 20273 10885 20307
rect 10919 20304 10931 20307
rect 10962 20304 10968 20316
rect 10919 20276 10968 20304
rect 10919 20273 10931 20276
rect 10873 20267 10931 20273
rect 10962 20264 10968 20276
rect 11020 20264 11026 20316
rect 12621 20307 12679 20313
rect 12621 20273 12633 20307
rect 12667 20304 12679 20307
rect 12986 20304 12992 20316
rect 12667 20276 12992 20304
rect 12667 20273 12679 20276
rect 12621 20267 12679 20273
rect 12986 20264 12992 20276
rect 13044 20264 13050 20316
rect 13170 20304 13176 20316
rect 13131 20276 13176 20304
rect 13170 20264 13176 20276
rect 13228 20264 13234 20316
rect 14366 20264 14372 20316
rect 14424 20304 14430 20316
rect 14461 20307 14519 20313
rect 14461 20304 14473 20307
rect 14424 20276 14473 20304
rect 14424 20264 14430 20276
rect 14461 20273 14473 20276
rect 14507 20273 14519 20307
rect 14461 20267 14519 20273
rect 12894 20196 12900 20248
rect 12952 20236 12958 20248
rect 13541 20239 13599 20245
rect 13541 20236 13553 20239
rect 12952 20208 13553 20236
rect 12952 20196 12958 20208
rect 13541 20205 13553 20208
rect 13587 20205 13599 20239
rect 13541 20199 13599 20205
rect 10778 20128 10784 20180
rect 10836 20168 10842 20180
rect 11238 20168 11244 20180
rect 10836 20140 11244 20168
rect 10836 20128 10842 20140
rect 11238 20128 11244 20140
rect 11296 20128 11302 20180
rect 14476 20168 14504 20267
rect 14642 20264 14648 20316
rect 14700 20304 14706 20316
rect 14829 20307 14887 20313
rect 14829 20304 14841 20307
rect 14700 20276 14841 20304
rect 14700 20264 14706 20276
rect 14829 20273 14841 20276
rect 14875 20273 14887 20307
rect 16114 20304 16120 20316
rect 16075 20276 16120 20304
rect 14829 20267 14887 20273
rect 16114 20264 16120 20276
rect 16172 20264 16178 20316
rect 17678 20304 17684 20316
rect 17639 20276 17684 20304
rect 17678 20264 17684 20276
rect 17736 20264 17742 20316
rect 20441 20307 20499 20313
rect 20441 20273 20453 20307
rect 20487 20304 20499 20307
rect 20622 20304 20628 20316
rect 20487 20276 20628 20304
rect 20487 20273 20499 20276
rect 20441 20267 20499 20273
rect 20622 20264 20628 20276
rect 20680 20264 20686 20316
rect 22097 20307 22155 20313
rect 22097 20273 22109 20307
rect 22143 20304 22155 20307
rect 22370 20304 22376 20316
rect 22143 20276 22376 20304
rect 22143 20273 22155 20276
rect 22097 20267 22155 20273
rect 22370 20264 22376 20276
rect 22428 20264 22434 20316
rect 23750 20304 23756 20316
rect 23711 20276 23756 20304
rect 23750 20264 23756 20276
rect 23808 20264 23814 20316
rect 24118 20264 24124 20316
rect 24176 20304 24182 20316
rect 24673 20307 24731 20313
rect 24673 20304 24685 20307
rect 24176 20276 24685 20304
rect 24176 20264 24182 20276
rect 24673 20273 24685 20276
rect 24719 20273 24731 20307
rect 24673 20267 24731 20273
rect 15289 20171 15347 20177
rect 15289 20168 15301 20171
rect 14476 20140 15301 20168
rect 15289 20137 15301 20140
rect 15335 20137 15347 20171
rect 15289 20131 15347 20137
rect 19334 20128 19340 20180
rect 19392 20168 19398 20180
rect 19429 20171 19487 20177
rect 19429 20168 19441 20171
rect 19392 20140 19441 20168
rect 19392 20128 19398 20140
rect 19429 20137 19441 20140
rect 19475 20137 19487 20171
rect 19429 20131 19487 20137
rect 19518 20128 19524 20180
rect 19576 20168 19582 20180
rect 19981 20171 20039 20177
rect 19981 20168 19993 20171
rect 19576 20140 19993 20168
rect 19576 20128 19582 20140
rect 19981 20137 19993 20140
rect 20027 20137 20039 20171
rect 19981 20131 20039 20137
rect 22094 20128 22100 20180
rect 22152 20168 22158 20180
rect 22370 20168 22376 20180
rect 22152 20140 22376 20168
rect 22152 20128 22158 20140
rect 22370 20128 22376 20140
rect 22428 20128 22434 20180
rect 23750 20128 23756 20180
rect 23808 20168 23814 20180
rect 26142 20168 26148 20180
rect 23808 20140 26148 20168
rect 23808 20128 23814 20140
rect 26142 20128 26148 20140
rect 26200 20128 26206 20180
rect 11508 20103 11566 20109
rect 11508 20069 11520 20103
rect 11554 20100 11566 20103
rect 11790 20100 11796 20112
rect 11554 20072 11796 20100
rect 11554 20069 11566 20072
rect 11508 20063 11566 20069
rect 11790 20060 11796 20072
rect 11848 20060 11854 20112
rect 13722 20100 13728 20112
rect 13683 20072 13728 20100
rect 13722 20060 13728 20072
rect 13780 20060 13786 20112
rect 22646 20109 22652 20112
rect 16301 20103 16359 20109
rect 16301 20100 16313 20103
rect 15764 20072 16313 20100
rect 13998 20032 14004 20044
rect 13959 20004 14004 20032
rect 13998 19992 14004 20004
rect 14056 19992 14062 20044
rect 10505 19967 10563 19973
rect 10505 19933 10517 19967
rect 10551 19964 10563 19967
rect 10686 19964 10692 19976
rect 10551 19936 10692 19964
rect 10551 19933 10563 19936
rect 10505 19927 10563 19933
rect 10686 19924 10692 19936
rect 10744 19924 10750 19976
rect 14734 19924 14740 19976
rect 14792 19964 14798 19976
rect 15562 19964 15568 19976
rect 14792 19936 15568 19964
rect 14792 19924 14798 19936
rect 15562 19924 15568 19936
rect 15620 19964 15626 19976
rect 15764 19973 15792 20072
rect 16301 20069 16313 20072
rect 16347 20069 16359 20103
rect 22640 20100 22652 20109
rect 22607 20072 22652 20100
rect 16301 20063 16359 20069
rect 22640 20063 22652 20072
rect 22646 20060 22652 20063
rect 22704 20060 22710 20112
rect 24854 20100 24860 20112
rect 24815 20072 24860 20100
rect 24854 20060 24860 20072
rect 24912 20100 24918 20112
rect 25409 20103 25467 20109
rect 25409 20100 25421 20103
rect 24912 20072 25421 20100
rect 24912 20060 24918 20072
rect 25409 20069 25421 20072
rect 25455 20069 25467 20103
rect 25409 20063 25467 20069
rect 16482 19992 16488 20044
rect 16540 20041 16546 20044
rect 16540 20035 16604 20041
rect 16540 20001 16558 20035
rect 16592 20001 16604 20035
rect 18506 20032 18512 20044
rect 18419 20004 18512 20032
rect 16540 19995 16604 20001
rect 16540 19992 16546 19995
rect 18506 19992 18512 20004
rect 18564 20032 18570 20044
rect 19337 20035 19395 20041
rect 19337 20032 19349 20035
rect 18564 20004 19349 20032
rect 18564 19992 18570 20004
rect 19337 20001 19349 20004
rect 19383 20001 19395 20035
rect 19337 19995 19395 20001
rect 22370 19992 22376 20044
rect 22428 20032 22434 20044
rect 23658 20032 23664 20044
rect 22428 20004 23664 20032
rect 22428 19992 22434 20004
rect 23658 19992 23664 20004
rect 23716 20032 23722 20044
rect 24305 20035 24363 20041
rect 24305 20032 24317 20035
rect 23716 20004 24317 20032
rect 23716 19992 23722 20004
rect 24305 20001 24317 20004
rect 24351 20001 24363 20035
rect 24305 19995 24363 20001
rect 15749 19967 15807 19973
rect 15749 19964 15761 19967
rect 15620 19936 15761 19964
rect 15620 19924 15626 19936
rect 15749 19933 15761 19936
rect 15795 19933 15807 19967
rect 15749 19927 15807 19933
rect 18046 19924 18052 19976
rect 18104 19964 18110 19976
rect 18690 19964 18696 19976
rect 18104 19936 18696 19964
rect 18104 19924 18110 19936
rect 18690 19924 18696 19936
rect 18748 19964 18754 19976
rect 18785 19967 18843 19973
rect 18785 19964 18797 19967
rect 18748 19936 18797 19964
rect 18748 19924 18754 19936
rect 18785 19933 18797 19936
rect 18831 19933 18843 19967
rect 18966 19964 18972 19976
rect 18927 19936 18972 19964
rect 18785 19927 18843 19933
rect 18966 19924 18972 19936
rect 19024 19924 19030 19976
rect 21634 19964 21640 19976
rect 21595 19936 21640 19964
rect 21634 19924 21640 19936
rect 21692 19964 21698 19976
rect 22186 19964 22192 19976
rect 21692 19936 22192 19964
rect 21692 19924 21698 19936
rect 22186 19924 22192 19936
rect 22244 19924 22250 19976
rect 25038 19964 25044 19976
rect 24999 19936 25044 19964
rect 25038 19924 25044 19936
rect 25096 19924 25102 19976
rect 1104 19874 26864 19896
rect 1104 19822 10315 19874
rect 10367 19822 10379 19874
rect 10431 19822 10443 19874
rect 10495 19822 10507 19874
rect 10559 19822 19648 19874
rect 19700 19822 19712 19874
rect 19764 19822 19776 19874
rect 19828 19822 19840 19874
rect 19892 19822 26864 19874
rect 1104 19800 26864 19822
rect 10873 19763 10931 19769
rect 10873 19729 10885 19763
rect 10919 19760 10931 19763
rect 11701 19763 11759 19769
rect 11701 19760 11713 19763
rect 10919 19732 11713 19760
rect 10919 19729 10931 19732
rect 10873 19723 10931 19729
rect 11701 19729 11713 19732
rect 11747 19760 11759 19763
rect 11790 19760 11796 19772
rect 11747 19732 11796 19760
rect 11747 19729 11759 19732
rect 11701 19723 11759 19729
rect 11790 19720 11796 19732
rect 11848 19720 11854 19772
rect 12342 19720 12348 19772
rect 12400 19760 12406 19772
rect 12713 19763 12771 19769
rect 12713 19760 12725 19763
rect 12400 19732 12725 19760
rect 12400 19720 12406 19732
rect 12713 19729 12725 19732
rect 12759 19760 12771 19763
rect 12986 19760 12992 19772
rect 12759 19732 12992 19760
rect 12759 19729 12771 19732
rect 12713 19723 12771 19729
rect 12986 19720 12992 19732
rect 13044 19720 13050 19772
rect 13354 19760 13360 19772
rect 13315 19732 13360 19760
rect 13354 19720 13360 19732
rect 13412 19720 13418 19772
rect 14093 19763 14151 19769
rect 14093 19729 14105 19763
rect 14139 19760 14151 19763
rect 14458 19760 14464 19772
rect 14139 19732 14464 19760
rect 14139 19729 14151 19732
rect 14093 19723 14151 19729
rect 11238 19692 11244 19704
rect 11199 19664 11244 19692
rect 11238 19652 11244 19664
rect 11296 19652 11302 19704
rect 13265 19695 13323 19701
rect 13265 19661 13277 19695
rect 13311 19692 13323 19695
rect 13538 19692 13544 19704
rect 13311 19664 13544 19692
rect 13311 19661 13323 19664
rect 13265 19655 13323 19661
rect 13538 19652 13544 19664
rect 13596 19652 13602 19704
rect 13541 19559 13599 19565
rect 13541 19525 13553 19559
rect 13587 19556 13599 19559
rect 13722 19556 13728 19568
rect 13587 19528 13728 19556
rect 13587 19525 13599 19528
rect 13541 19519 13599 19525
rect 13722 19516 13728 19528
rect 13780 19516 13786 19568
rect 12897 19491 12955 19497
rect 12897 19457 12909 19491
rect 12943 19488 12955 19491
rect 14108 19488 14136 19723
rect 14458 19720 14464 19732
rect 14516 19720 14522 19772
rect 16393 19763 16451 19769
rect 16393 19729 16405 19763
rect 16439 19760 16451 19763
rect 16482 19760 16488 19772
rect 16439 19732 16488 19760
rect 16439 19729 16451 19732
rect 16393 19723 16451 19729
rect 16482 19720 16488 19732
rect 16540 19720 16546 19772
rect 18506 19760 18512 19772
rect 18467 19732 18512 19760
rect 18506 19720 18512 19732
rect 18564 19720 18570 19772
rect 22370 19760 22376 19772
rect 22331 19732 22376 19760
rect 22370 19720 22376 19732
rect 22428 19720 22434 19772
rect 22557 19763 22615 19769
rect 22557 19729 22569 19763
rect 22603 19760 22615 19763
rect 23198 19760 23204 19772
rect 22603 19732 23204 19760
rect 22603 19729 22615 19732
rect 22557 19723 22615 19729
rect 23198 19720 23204 19732
rect 23256 19720 23262 19772
rect 25314 19760 25320 19772
rect 25275 19732 25320 19760
rect 25314 19720 25320 19732
rect 25372 19720 25378 19772
rect 14642 19652 14648 19704
rect 14700 19692 14706 19704
rect 15258 19695 15316 19701
rect 15258 19692 15270 19695
rect 14700 19664 15270 19692
rect 14700 19652 14706 19664
rect 15258 19661 15270 19664
rect 15304 19692 15316 19695
rect 15470 19692 15476 19704
rect 15304 19664 15476 19692
rect 15304 19661 15316 19664
rect 15258 19655 15316 19661
rect 15470 19652 15476 19664
rect 15528 19652 15534 19704
rect 22097 19695 22155 19701
rect 22097 19661 22109 19695
rect 22143 19692 22155 19695
rect 22646 19692 22652 19704
rect 22143 19664 22652 19692
rect 22143 19661 22155 19664
rect 22097 19655 22155 19661
rect 22646 19652 22652 19664
rect 22704 19692 22710 19704
rect 23017 19695 23075 19701
rect 23017 19692 23029 19695
rect 22704 19664 23029 19692
rect 22704 19652 22710 19664
rect 23017 19661 23029 19664
rect 23063 19661 23075 19695
rect 23017 19655 23075 19661
rect 18966 19584 18972 19636
rect 19024 19624 19030 19636
rect 19518 19624 19524 19636
rect 19024 19596 19524 19624
rect 19024 19584 19030 19596
rect 19518 19584 19524 19596
rect 19576 19584 19582 19636
rect 19794 19624 19800 19636
rect 19755 19596 19800 19624
rect 19794 19584 19800 19596
rect 19852 19584 19858 19636
rect 23474 19584 23480 19636
rect 23532 19624 23538 19636
rect 23842 19624 23848 19636
rect 23532 19596 23848 19624
rect 23532 19584 23538 19596
rect 23842 19584 23848 19596
rect 23900 19584 23906 19636
rect 24854 19584 24860 19636
rect 24912 19624 24918 19636
rect 25133 19627 25191 19633
rect 25133 19624 25145 19627
rect 24912 19596 25145 19624
rect 24912 19584 24918 19596
rect 25133 19593 25145 19596
rect 25179 19593 25191 19627
rect 25133 19587 25191 19593
rect 14734 19516 14740 19568
rect 14792 19556 14798 19568
rect 15013 19559 15071 19565
rect 15013 19556 15025 19559
rect 14792 19528 15025 19556
rect 14792 19516 14798 19528
rect 15013 19525 15025 19528
rect 15059 19525 15071 19559
rect 24118 19556 24124 19568
rect 24079 19528 24124 19556
rect 15013 19519 15071 19525
rect 24118 19516 24124 19528
rect 24176 19516 24182 19568
rect 12943 19460 14136 19488
rect 12943 19457 12955 19460
rect 12897 19451 12955 19457
rect 16390 19380 16396 19432
rect 16448 19420 16454 19432
rect 17034 19420 17040 19432
rect 16448 19392 17040 19420
rect 16448 19380 16454 19392
rect 17034 19380 17040 19392
rect 17092 19380 17098 19432
rect 19334 19420 19340 19432
rect 19295 19392 19340 19420
rect 19334 19380 19340 19392
rect 19392 19380 19398 19432
rect 1104 19330 26864 19352
rect 1104 19278 5648 19330
rect 5700 19278 5712 19330
rect 5764 19278 5776 19330
rect 5828 19278 5840 19330
rect 5892 19278 14982 19330
rect 15034 19278 15046 19330
rect 15098 19278 15110 19330
rect 15162 19278 15174 19330
rect 15226 19278 24315 19330
rect 24367 19278 24379 19330
rect 24431 19278 24443 19330
rect 24495 19278 24507 19330
rect 24559 19278 26864 19330
rect 1104 19256 26864 19278
rect 11238 19176 11244 19228
rect 11296 19216 11302 19228
rect 11885 19219 11943 19225
rect 11885 19216 11897 19219
rect 11296 19188 11897 19216
rect 11296 19176 11302 19188
rect 11885 19185 11897 19188
rect 11931 19185 11943 19219
rect 15470 19216 15476 19228
rect 15431 19188 15476 19216
rect 11885 19179 11943 19185
rect 11900 19080 11928 19179
rect 15470 19176 15476 19188
rect 15528 19176 15534 19228
rect 19518 19176 19524 19228
rect 19576 19216 19582 19228
rect 20257 19219 20315 19225
rect 20257 19216 20269 19219
rect 19576 19188 20269 19216
rect 19576 19176 19582 19188
rect 20257 19185 20269 19188
rect 20303 19185 20315 19219
rect 23842 19216 23848 19228
rect 23803 19188 23848 19216
rect 20257 19179 20315 19185
rect 23842 19176 23848 19188
rect 23900 19176 23906 19228
rect 24854 19176 24860 19228
rect 24912 19216 24918 19228
rect 25501 19219 25559 19225
rect 25501 19216 25513 19219
rect 24912 19188 25513 19216
rect 24912 19176 24918 19188
rect 25501 19185 25513 19188
rect 25547 19185 25559 19219
rect 25501 19179 25559 19185
rect 12066 19080 12072 19092
rect 11900 19052 12072 19080
rect 12066 19040 12072 19052
rect 12124 19040 12130 19092
rect 19797 19083 19855 19089
rect 19797 19049 19809 19083
rect 19843 19049 19855 19083
rect 22925 19083 22983 19089
rect 22925 19080 22937 19083
rect 19797 19043 19855 19049
rect 22112 19052 22937 19080
rect 12342 19021 12348 19024
rect 12336 19012 12348 19021
rect 12303 18984 12348 19012
rect 12336 18975 12348 18984
rect 12342 18972 12348 18975
rect 12400 18972 12406 19024
rect 16850 19012 16856 19024
rect 16811 18984 16856 19012
rect 16850 18972 16856 18984
rect 16908 18972 16914 19024
rect 18785 19015 18843 19021
rect 18785 18981 18797 19015
rect 18831 19012 18843 19015
rect 19518 19012 19524 19024
rect 18831 18984 19524 19012
rect 18831 18981 18843 18984
rect 18785 18975 18843 18981
rect 19518 18972 19524 18984
rect 19576 19012 19582 19024
rect 19812 19012 19840 19043
rect 19576 18984 19840 19012
rect 21545 19015 21603 19021
rect 19576 18972 19582 18984
rect 21545 18981 21557 19015
rect 21591 19012 21603 19015
rect 22002 19012 22008 19024
rect 21591 18984 22008 19012
rect 21591 18981 21603 18984
rect 21545 18975 21603 18981
rect 22002 18972 22008 18984
rect 22060 19012 22066 19024
rect 22112 19012 22140 19052
rect 22925 19049 22937 19052
rect 22971 19049 22983 19083
rect 22925 19043 22983 19049
rect 22060 18984 22140 19012
rect 22204 18984 22968 19012
rect 22060 18972 22066 18984
rect 19705 18947 19763 18953
rect 19705 18944 19717 18947
rect 19076 18916 19717 18944
rect 19076 18888 19104 18916
rect 19705 18913 19717 18916
rect 19751 18913 19763 18947
rect 19705 18907 19763 18913
rect 13449 18879 13507 18885
rect 13449 18845 13461 18879
rect 13495 18876 13507 18879
rect 13722 18876 13728 18888
rect 13495 18848 13728 18876
rect 13495 18845 13507 18848
rect 13449 18839 13507 18845
rect 13722 18836 13728 18848
rect 13780 18876 13786 18888
rect 14001 18879 14059 18885
rect 14001 18876 14013 18879
rect 13780 18848 14013 18876
rect 13780 18836 13786 18848
rect 14001 18845 14013 18848
rect 14047 18845 14059 18879
rect 14001 18839 14059 18845
rect 14734 18836 14740 18888
rect 14792 18876 14798 18888
rect 15013 18879 15071 18885
rect 15013 18876 15025 18879
rect 14792 18848 15025 18876
rect 14792 18836 14798 18848
rect 15013 18845 15025 18848
rect 15059 18845 15071 18879
rect 19058 18876 19064 18888
rect 19019 18848 19064 18876
rect 15013 18839 15071 18845
rect 19058 18836 19064 18848
rect 19116 18836 19122 18888
rect 19242 18876 19248 18888
rect 19203 18848 19248 18876
rect 19242 18836 19248 18848
rect 19300 18836 19306 18888
rect 19334 18836 19340 18888
rect 19392 18876 19398 18888
rect 19613 18879 19671 18885
rect 19613 18876 19625 18879
rect 19392 18848 19625 18876
rect 19392 18836 19398 18848
rect 19613 18845 19625 18848
rect 19659 18876 19671 18879
rect 20622 18876 20628 18888
rect 19659 18848 20628 18876
rect 19659 18845 19671 18848
rect 19613 18839 19671 18845
rect 20622 18836 20628 18848
rect 20680 18836 20686 18888
rect 21910 18876 21916 18888
rect 21823 18848 21916 18876
rect 21910 18836 21916 18848
rect 21968 18876 21974 18888
rect 22204 18876 22232 18984
rect 22278 18904 22284 18956
rect 22336 18944 22342 18956
rect 22833 18947 22891 18953
rect 22833 18944 22845 18947
rect 22336 18916 22845 18944
rect 22336 18904 22342 18916
rect 22833 18913 22845 18916
rect 22879 18913 22891 18947
rect 22833 18907 22891 18913
rect 22370 18876 22376 18888
rect 21968 18848 22232 18876
rect 22331 18848 22376 18876
rect 21968 18836 21974 18848
rect 22370 18836 22376 18848
rect 22428 18836 22434 18888
rect 22741 18879 22799 18885
rect 22741 18845 22753 18879
rect 22787 18876 22799 18879
rect 22940 18876 22968 18984
rect 24118 18972 24124 19024
rect 24176 19012 24182 19024
rect 24581 19015 24639 19021
rect 24581 19012 24593 19015
rect 24176 18984 24593 19012
rect 24176 18972 24182 18984
rect 24581 18981 24593 18984
rect 24627 19012 24639 19015
rect 25133 19015 25191 19021
rect 25133 19012 25145 19015
rect 24627 18984 25145 19012
rect 24627 18981 24639 18984
rect 24581 18975 24639 18981
rect 25133 18981 25145 18984
rect 25179 18981 25191 19015
rect 25133 18975 25191 18981
rect 23382 18876 23388 18888
rect 22787 18848 23388 18876
rect 22787 18845 22799 18848
rect 22741 18839 22799 18845
rect 23382 18836 23388 18848
rect 23440 18836 23446 18888
rect 24762 18876 24768 18888
rect 24723 18848 24768 18876
rect 24762 18836 24768 18848
rect 24820 18836 24826 18888
rect 1104 18786 26864 18808
rect 1104 18734 10315 18786
rect 10367 18734 10379 18786
rect 10431 18734 10443 18786
rect 10495 18734 10507 18786
rect 10559 18734 19648 18786
rect 19700 18734 19712 18786
rect 19764 18734 19776 18786
rect 19828 18734 19840 18786
rect 19892 18734 26864 18786
rect 1104 18712 26864 18734
rect 12161 18675 12219 18681
rect 12161 18641 12173 18675
rect 12207 18672 12219 18675
rect 12342 18672 12348 18684
rect 12207 18644 12348 18672
rect 12207 18641 12219 18644
rect 12161 18635 12219 18641
rect 12342 18632 12348 18644
rect 12400 18632 12406 18684
rect 12989 18675 13047 18681
rect 12989 18641 13001 18675
rect 13035 18672 13047 18675
rect 13354 18672 13360 18684
rect 13035 18644 13360 18672
rect 13035 18641 13047 18644
rect 12989 18635 13047 18641
rect 13354 18632 13360 18644
rect 13412 18632 13418 18684
rect 14829 18675 14887 18681
rect 14829 18641 14841 18675
rect 14875 18672 14887 18675
rect 15470 18672 15476 18684
rect 14875 18644 15476 18672
rect 14875 18641 14887 18644
rect 14829 18635 14887 18641
rect 15470 18632 15476 18644
rect 15528 18632 15534 18684
rect 24026 18632 24032 18684
rect 24084 18632 24090 18684
rect 20993 18607 21051 18613
rect 20993 18573 21005 18607
rect 21039 18604 21051 18607
rect 21352 18607 21410 18613
rect 21352 18604 21364 18607
rect 21039 18576 21364 18604
rect 21039 18573 21051 18576
rect 20993 18567 21051 18573
rect 21352 18573 21364 18576
rect 21398 18604 21410 18607
rect 21542 18604 21548 18616
rect 21398 18576 21548 18604
rect 21398 18573 21410 18576
rect 21352 18567 21410 18573
rect 21542 18564 21548 18576
rect 21600 18564 21606 18616
rect 24044 18604 24072 18632
rect 24118 18604 24124 18616
rect 24031 18576 24124 18604
rect 24118 18564 24124 18576
rect 24176 18564 24182 18616
rect 12066 18496 12072 18548
rect 12124 18536 12130 18548
rect 13354 18536 13360 18548
rect 12124 18508 13216 18536
rect 13267 18508 13360 18536
rect 12124 18496 12130 18508
rect 13188 18468 13216 18508
rect 13354 18496 13360 18508
rect 13412 18536 13418 18548
rect 13538 18536 13544 18548
rect 13412 18508 13544 18536
rect 13412 18496 13418 18508
rect 13538 18496 13544 18508
rect 13596 18496 13602 18548
rect 13722 18545 13728 18548
rect 13716 18536 13728 18545
rect 13683 18508 13728 18536
rect 13716 18499 13728 18508
rect 13722 18496 13728 18499
rect 13780 18496 13786 18548
rect 18305 18539 18363 18545
rect 18305 18536 18317 18539
rect 17788 18508 18317 18536
rect 13262 18468 13268 18480
rect 13188 18440 13268 18468
rect 13262 18428 13268 18440
rect 13320 18468 13326 18480
rect 13449 18471 13507 18477
rect 13449 18468 13461 18471
rect 13320 18440 13461 18468
rect 13320 18428 13326 18440
rect 13449 18437 13461 18440
rect 13495 18437 13507 18471
rect 13449 18431 13507 18437
rect 15930 18332 15936 18344
rect 15891 18304 15936 18332
rect 15930 18292 15936 18304
rect 15988 18292 15994 18344
rect 17310 18292 17316 18344
rect 17368 18332 17374 18344
rect 17788 18341 17816 18508
rect 18305 18505 18317 18508
rect 18351 18505 18363 18539
rect 18305 18499 18363 18505
rect 21085 18539 21143 18545
rect 21085 18505 21097 18539
rect 21131 18536 21143 18539
rect 21174 18536 21180 18548
rect 21131 18508 21180 18536
rect 21131 18505 21143 18508
rect 21085 18499 21143 18505
rect 21174 18496 21180 18508
rect 21232 18496 21238 18548
rect 24026 18536 24032 18548
rect 23987 18508 24032 18536
rect 24026 18496 24032 18508
rect 24084 18496 24090 18548
rect 24136 18536 24164 18564
rect 25222 18536 25228 18548
rect 24136 18508 24256 18536
rect 25183 18508 25228 18536
rect 18046 18468 18052 18480
rect 18007 18440 18052 18468
rect 18046 18428 18052 18440
rect 18104 18428 18110 18480
rect 22370 18428 22376 18480
rect 22428 18468 22434 18480
rect 23474 18468 23480 18480
rect 22428 18440 23480 18468
rect 22428 18428 22434 18440
rect 23474 18428 23480 18440
rect 23532 18468 23538 18480
rect 24228 18477 24256 18508
rect 25222 18496 25228 18508
rect 25280 18496 25286 18548
rect 24121 18471 24179 18477
rect 24121 18468 24133 18471
rect 23532 18440 24133 18468
rect 23532 18428 23538 18440
rect 24121 18437 24133 18440
rect 24167 18437 24179 18471
rect 24121 18431 24179 18437
rect 24213 18471 24271 18477
rect 24213 18437 24225 18471
rect 24259 18437 24271 18471
rect 24213 18431 24271 18437
rect 25406 18400 25412 18412
rect 25367 18372 25412 18400
rect 25406 18360 25412 18372
rect 25464 18360 25470 18412
rect 17773 18335 17831 18341
rect 17773 18332 17785 18335
rect 17368 18304 17785 18332
rect 17368 18292 17374 18304
rect 17773 18301 17785 18304
rect 17819 18301 17831 18335
rect 17773 18295 17831 18301
rect 19242 18292 19248 18344
rect 19300 18332 19306 18344
rect 19429 18335 19487 18341
rect 19429 18332 19441 18335
rect 19300 18304 19441 18332
rect 19300 18292 19306 18304
rect 19429 18301 19441 18304
rect 19475 18301 19487 18335
rect 19429 18295 19487 18301
rect 22002 18292 22008 18344
rect 22060 18332 22066 18344
rect 22462 18332 22468 18344
rect 22060 18304 22468 18332
rect 22060 18292 22066 18304
rect 22462 18292 22468 18304
rect 22520 18292 22526 18344
rect 23658 18332 23664 18344
rect 23619 18304 23664 18332
rect 23658 18292 23664 18304
rect 23716 18292 23722 18344
rect 1104 18242 26864 18264
rect 1104 18190 5648 18242
rect 5700 18190 5712 18242
rect 5764 18190 5776 18242
rect 5828 18190 5840 18242
rect 5892 18190 14982 18242
rect 15034 18190 15046 18242
rect 15098 18190 15110 18242
rect 15162 18190 15174 18242
rect 15226 18190 24315 18242
rect 24367 18190 24379 18242
rect 24431 18190 24443 18242
rect 24495 18190 24507 18242
rect 24559 18190 26864 18242
rect 1104 18168 26864 18190
rect 13722 18088 13728 18140
rect 13780 18128 13786 18140
rect 13817 18131 13875 18137
rect 13817 18128 13829 18131
rect 13780 18100 13829 18128
rect 13780 18088 13786 18100
rect 13817 18097 13829 18100
rect 13863 18097 13875 18131
rect 13817 18091 13875 18097
rect 19518 18088 19524 18140
rect 19576 18128 19582 18140
rect 19705 18131 19763 18137
rect 19705 18128 19717 18131
rect 19576 18100 19717 18128
rect 19576 18088 19582 18100
rect 19705 18097 19717 18100
rect 19751 18097 19763 18131
rect 19705 18091 19763 18097
rect 24118 18088 24124 18140
rect 24176 18128 24182 18140
rect 24397 18131 24455 18137
rect 24397 18128 24409 18131
rect 24176 18100 24409 18128
rect 24176 18088 24182 18100
rect 24397 18097 24409 18100
rect 24443 18128 24455 18131
rect 24949 18131 25007 18137
rect 24949 18128 24961 18131
rect 24443 18100 24961 18128
rect 24443 18097 24455 18100
rect 24397 18091 24455 18097
rect 24949 18097 24961 18100
rect 24995 18097 25007 18131
rect 24949 18091 25007 18097
rect 20714 18020 20720 18072
rect 20772 18060 20778 18072
rect 21174 18060 21180 18072
rect 20772 18032 21180 18060
rect 20772 18020 20778 18032
rect 21174 18020 21180 18032
rect 21232 18060 21238 18072
rect 22005 18063 22063 18069
rect 22005 18060 22017 18063
rect 21232 18032 22017 18060
rect 21232 18020 21238 18032
rect 22005 18029 22017 18032
rect 22051 18060 22063 18063
rect 22833 18063 22891 18069
rect 22833 18060 22845 18063
rect 22051 18032 22845 18060
rect 22051 18029 22063 18032
rect 22005 18023 22063 18029
rect 22833 18029 22845 18032
rect 22879 18060 22891 18063
rect 22879 18032 23060 18060
rect 22879 18029 22891 18032
rect 22833 18023 22891 18029
rect 20349 17995 20407 18001
rect 20349 17961 20361 17995
rect 20395 17992 20407 17995
rect 21542 17992 21548 18004
rect 20395 17964 21548 17992
rect 20395 17961 20407 17964
rect 20349 17955 20407 17961
rect 21542 17952 21548 17964
rect 21600 17952 21606 18004
rect 23032 18001 23060 18032
rect 23017 17995 23075 18001
rect 23017 17961 23029 17995
rect 23063 17961 23075 17995
rect 23017 17955 23075 17961
rect 15841 17927 15899 17933
rect 15841 17893 15853 17927
rect 15887 17893 15899 17927
rect 15841 17887 15899 17893
rect 14734 17856 14740 17868
rect 13740 17828 14740 17856
rect 13740 17800 13768 17828
rect 14734 17816 14740 17828
rect 14792 17856 14798 17868
rect 15657 17859 15715 17865
rect 15657 17856 15669 17859
rect 14792 17828 15669 17856
rect 14792 17816 14798 17828
rect 15657 17825 15669 17828
rect 15703 17856 15715 17859
rect 15856 17856 15884 17887
rect 15930 17884 15936 17936
rect 15988 17924 15994 17936
rect 16097 17927 16155 17933
rect 16097 17924 16109 17927
rect 15988 17896 16109 17924
rect 15988 17884 15994 17896
rect 16097 17893 16109 17896
rect 16143 17924 16155 17927
rect 16390 17924 16396 17936
rect 16143 17896 16396 17924
rect 16143 17893 16155 17896
rect 16097 17887 16155 17893
rect 16390 17884 16396 17896
rect 16448 17884 16454 17936
rect 18325 17927 18383 17933
rect 18325 17893 18337 17927
rect 18371 17893 18383 17927
rect 21358 17924 21364 17936
rect 21319 17896 21364 17924
rect 18325 17887 18383 17893
rect 17773 17859 17831 17865
rect 17773 17856 17785 17859
rect 15703 17828 17785 17856
rect 15703 17825 15715 17828
rect 15657 17819 15715 17825
rect 17773 17825 17785 17828
rect 17819 17856 17831 17859
rect 18046 17856 18052 17868
rect 17819 17828 18052 17856
rect 17819 17825 17831 17828
rect 17773 17819 17831 17825
rect 18046 17816 18052 17828
rect 18104 17856 18110 17868
rect 18141 17859 18199 17865
rect 18141 17856 18153 17859
rect 18104 17828 18153 17856
rect 18104 17816 18110 17828
rect 18141 17825 18153 17828
rect 18187 17856 18199 17859
rect 18340 17856 18368 17887
rect 21358 17884 21364 17896
rect 21416 17924 21422 17936
rect 22281 17927 22339 17933
rect 22281 17924 22293 17927
rect 21416 17896 22293 17924
rect 21416 17884 21422 17896
rect 22281 17893 22293 17896
rect 22327 17893 22339 17927
rect 22281 17887 22339 17893
rect 22462 17884 22468 17936
rect 22520 17924 22526 17936
rect 23106 17924 23112 17936
rect 22520 17896 23112 17924
rect 22520 17884 22526 17896
rect 23106 17884 23112 17896
rect 23164 17924 23170 17936
rect 23273 17927 23331 17933
rect 23273 17924 23285 17927
rect 23164 17896 23285 17924
rect 23164 17884 23170 17896
rect 23273 17893 23285 17896
rect 23319 17893 23331 17927
rect 23273 17887 23331 17893
rect 18187 17828 18368 17856
rect 18592 17859 18650 17865
rect 18187 17825 18199 17828
rect 18141 17819 18199 17825
rect 18592 17825 18604 17859
rect 18638 17856 18650 17859
rect 19242 17856 19248 17868
rect 18638 17828 19248 17856
rect 18638 17825 18650 17828
rect 18592 17819 18650 17825
rect 19242 17816 19248 17828
rect 19300 17816 19306 17868
rect 20717 17859 20775 17865
rect 20717 17825 20729 17859
rect 20763 17856 20775 17859
rect 20990 17856 20996 17868
rect 20763 17828 20996 17856
rect 20763 17825 20775 17828
rect 20717 17819 20775 17825
rect 20990 17816 20996 17828
rect 21048 17856 21054 17868
rect 21269 17859 21327 17865
rect 21269 17856 21281 17859
rect 21048 17828 21281 17856
rect 21048 17816 21054 17828
rect 21269 17825 21281 17828
rect 21315 17825 21327 17859
rect 21269 17819 21327 17825
rect 24854 17816 24860 17868
rect 24912 17856 24918 17868
rect 25222 17856 25228 17868
rect 24912 17828 25228 17856
rect 24912 17816 24918 17828
rect 25222 17816 25228 17828
rect 25280 17856 25286 17868
rect 25317 17859 25375 17865
rect 25317 17856 25329 17859
rect 25280 17828 25329 17856
rect 25280 17816 25286 17828
rect 25317 17825 25329 17828
rect 25363 17825 25375 17859
rect 25317 17819 25375 17825
rect 13262 17748 13268 17800
rect 13320 17788 13326 17800
rect 13541 17791 13599 17797
rect 13541 17788 13553 17791
rect 13320 17760 13553 17788
rect 13320 17748 13326 17760
rect 13541 17757 13553 17760
rect 13587 17788 13599 17791
rect 13722 17788 13728 17800
rect 13587 17760 13728 17788
rect 13587 17757 13599 17760
rect 13541 17751 13599 17757
rect 13722 17748 13728 17760
rect 13780 17748 13786 17800
rect 14274 17788 14280 17800
rect 14235 17760 14280 17788
rect 14274 17748 14280 17760
rect 14332 17748 14338 17800
rect 17221 17791 17279 17797
rect 17221 17757 17233 17791
rect 17267 17788 17279 17791
rect 17310 17788 17316 17800
rect 17267 17760 17316 17788
rect 17267 17757 17279 17760
rect 17221 17751 17279 17757
rect 17310 17748 17316 17760
rect 17368 17748 17374 17800
rect 20898 17788 20904 17800
rect 20859 17760 20904 17788
rect 20898 17748 20904 17760
rect 20956 17748 20962 17800
rect 1104 17698 26864 17720
rect 1104 17646 10315 17698
rect 10367 17646 10379 17698
rect 10431 17646 10443 17698
rect 10495 17646 10507 17698
rect 10559 17646 19648 17698
rect 19700 17646 19712 17698
rect 19764 17646 19776 17698
rect 19828 17646 19840 17698
rect 19892 17646 26864 17698
rect 1104 17624 26864 17646
rect 15841 17587 15899 17593
rect 15841 17553 15853 17587
rect 15887 17584 15899 17587
rect 18509 17587 18567 17593
rect 18509 17584 18521 17587
rect 15887 17556 18521 17584
rect 15887 17553 15899 17556
rect 15841 17547 15899 17553
rect 18509 17553 18521 17556
rect 18555 17584 18567 17587
rect 19150 17584 19156 17596
rect 18555 17556 19156 17584
rect 18555 17553 18567 17556
rect 18509 17547 18567 17553
rect 19150 17544 19156 17556
rect 19208 17544 19214 17596
rect 21542 17584 21548 17596
rect 21503 17556 21548 17584
rect 21542 17544 21548 17556
rect 21600 17544 21606 17596
rect 23106 17584 23112 17596
rect 23067 17556 23112 17584
rect 23106 17544 23112 17556
rect 23164 17544 23170 17596
rect 23474 17584 23480 17596
rect 23435 17556 23480 17584
rect 23474 17544 23480 17556
rect 23532 17544 23538 17596
rect 23937 17587 23995 17593
rect 23937 17553 23949 17587
rect 23983 17584 23995 17587
rect 24026 17584 24032 17596
rect 23983 17556 24032 17584
rect 23983 17553 23995 17556
rect 23937 17547 23995 17553
rect 24026 17544 24032 17556
rect 24084 17544 24090 17596
rect 25590 17584 25596 17596
rect 25551 17556 25596 17584
rect 25590 17544 25596 17556
rect 25648 17544 25654 17596
rect 15286 17476 15292 17528
rect 15344 17516 15350 17528
rect 15746 17516 15752 17528
rect 15344 17488 15752 17516
rect 15344 17476 15350 17488
rect 15746 17476 15752 17488
rect 15804 17476 15810 17528
rect 16301 17519 16359 17525
rect 16301 17516 16313 17519
rect 15856 17488 16313 17516
rect 15856 17460 15884 17488
rect 16301 17485 16313 17488
rect 16347 17485 16359 17519
rect 16301 17479 16359 17485
rect 19518 17476 19524 17528
rect 19576 17516 19582 17528
rect 20410 17519 20468 17525
rect 20410 17516 20422 17519
rect 19576 17488 20422 17516
rect 19576 17476 19582 17488
rect 20410 17485 20422 17488
rect 20456 17516 20468 17519
rect 20530 17516 20536 17528
rect 20456 17488 20536 17516
rect 20456 17485 20468 17488
rect 20410 17479 20468 17485
rect 20530 17476 20536 17488
rect 20588 17476 20594 17528
rect 20622 17476 20628 17528
rect 20680 17476 20686 17528
rect 24397 17519 24455 17525
rect 24397 17485 24409 17519
rect 24443 17516 24455 17519
rect 24762 17516 24768 17528
rect 24443 17488 24768 17516
rect 24443 17485 24455 17488
rect 24397 17479 24455 17485
rect 24762 17476 24768 17488
rect 24820 17476 24826 17528
rect 14274 17408 14280 17460
rect 14332 17448 14338 17460
rect 14461 17451 14519 17457
rect 14461 17448 14473 17451
rect 14332 17420 14473 17448
rect 14332 17408 14338 17420
rect 14461 17417 14473 17420
rect 14507 17448 14519 17451
rect 15102 17448 15108 17460
rect 14507 17420 15108 17448
rect 14507 17417 14519 17420
rect 14461 17411 14519 17417
rect 15102 17408 15108 17420
rect 15160 17408 15166 17460
rect 15838 17408 15844 17460
rect 15896 17408 15902 17460
rect 16206 17448 16212 17460
rect 16119 17420 16212 17448
rect 16206 17408 16212 17420
rect 16264 17448 16270 17460
rect 17034 17448 17040 17460
rect 16264 17420 17040 17448
rect 16264 17408 16270 17420
rect 17034 17408 17040 17420
rect 17092 17408 17098 17460
rect 18417 17451 18475 17457
rect 18417 17417 18429 17451
rect 18463 17448 18475 17451
rect 18782 17448 18788 17460
rect 18463 17420 18788 17448
rect 18463 17417 18475 17420
rect 18417 17411 18475 17417
rect 18782 17408 18788 17420
rect 18840 17408 18846 17460
rect 19153 17451 19211 17457
rect 19153 17417 19165 17451
rect 19199 17448 19211 17451
rect 19242 17448 19248 17460
rect 19199 17420 19248 17448
rect 19199 17417 19211 17420
rect 19153 17411 19211 17417
rect 19242 17408 19248 17420
rect 19300 17408 19306 17460
rect 20162 17448 20168 17460
rect 20075 17420 20168 17448
rect 20162 17408 20168 17420
rect 20220 17448 20226 17460
rect 20640 17448 20668 17476
rect 20220 17420 20668 17448
rect 20220 17408 20226 17420
rect 23658 17408 23664 17460
rect 23716 17448 23722 17460
rect 24118 17448 24124 17460
rect 23716 17420 24124 17448
rect 23716 17408 23722 17420
rect 24118 17408 24124 17420
rect 24176 17408 24182 17460
rect 25406 17448 25412 17460
rect 25319 17420 25412 17448
rect 25406 17408 25412 17420
rect 25464 17448 25470 17460
rect 26326 17448 26332 17460
rect 25464 17420 26332 17448
rect 25464 17408 25470 17420
rect 26326 17408 26332 17420
rect 26384 17408 26390 17460
rect 14550 17380 14556 17392
rect 14511 17352 14556 17380
rect 14550 17340 14556 17352
rect 14608 17340 14614 17392
rect 14734 17380 14740 17392
rect 14647 17352 14740 17380
rect 14734 17340 14740 17352
rect 14792 17380 14798 17392
rect 15289 17383 15347 17389
rect 15289 17380 15301 17383
rect 14792 17352 15301 17380
rect 14792 17340 14798 17352
rect 15289 17349 15301 17352
rect 15335 17349 15347 17383
rect 16390 17380 16396 17392
rect 16351 17352 16396 17380
rect 15289 17343 15347 17349
rect 16390 17340 16396 17352
rect 16448 17340 16454 17392
rect 18601 17383 18659 17389
rect 18601 17380 18613 17383
rect 17788 17352 18613 17380
rect 14090 17312 14096 17324
rect 14051 17284 14096 17312
rect 14090 17272 14096 17284
rect 14148 17272 14154 17324
rect 17788 17256 17816 17352
rect 18601 17349 18613 17352
rect 18647 17349 18659 17383
rect 18601 17343 18659 17349
rect 12158 17244 12164 17256
rect 12119 17216 12164 17244
rect 12158 17204 12164 17216
rect 12216 17204 12222 17256
rect 13725 17247 13783 17253
rect 13725 17213 13737 17247
rect 13771 17244 13783 17247
rect 14182 17244 14188 17256
rect 13771 17216 14188 17244
rect 13771 17213 13783 17216
rect 13725 17207 13783 17213
rect 14182 17204 14188 17216
rect 14240 17204 14246 17256
rect 17770 17244 17776 17256
rect 17731 17216 17776 17244
rect 17770 17204 17776 17216
rect 17828 17204 17834 17256
rect 18049 17247 18107 17253
rect 18049 17213 18061 17247
rect 18095 17244 18107 17247
rect 18506 17244 18512 17256
rect 18095 17216 18512 17244
rect 18095 17213 18107 17216
rect 18049 17207 18107 17213
rect 18506 17204 18512 17216
rect 18564 17204 18570 17256
rect 1104 17154 26864 17176
rect 1104 17102 5648 17154
rect 5700 17102 5712 17154
rect 5764 17102 5776 17154
rect 5828 17102 5840 17154
rect 5892 17102 14982 17154
rect 15034 17102 15046 17154
rect 15098 17102 15110 17154
rect 15162 17102 15174 17154
rect 15226 17102 24315 17154
rect 24367 17102 24379 17154
rect 24431 17102 24443 17154
rect 24495 17102 24507 17154
rect 24559 17102 26864 17154
rect 1104 17080 26864 17102
rect 13538 17000 13544 17052
rect 13596 17040 13602 17052
rect 13633 17043 13691 17049
rect 13633 17040 13645 17043
rect 13596 17012 13645 17040
rect 13596 17000 13602 17012
rect 13633 17009 13645 17012
rect 13679 17040 13691 17043
rect 14550 17040 14556 17052
rect 13679 17012 14556 17040
rect 13679 17009 13691 17012
rect 13633 17003 13691 17009
rect 14550 17000 14556 17012
rect 14608 17000 14614 17052
rect 14734 17040 14740 17052
rect 14695 17012 14740 17040
rect 14734 17000 14740 17012
rect 14792 17000 14798 17052
rect 16390 17000 16396 17052
rect 16448 17040 16454 17052
rect 16669 17043 16727 17049
rect 16669 17040 16681 17043
rect 16448 17012 16681 17040
rect 16448 17000 16454 17012
rect 16669 17009 16681 17012
rect 16715 17009 16727 17043
rect 17310 17040 17316 17052
rect 17223 17012 17316 17040
rect 16669 17003 16727 17009
rect 17310 17000 17316 17012
rect 17368 17040 17374 17052
rect 17770 17040 17776 17052
rect 17368 17012 17776 17040
rect 17368 17000 17374 17012
rect 17770 17000 17776 17012
rect 17828 17000 17834 17052
rect 19150 17040 19156 17052
rect 19111 17012 19156 17040
rect 19150 17000 19156 17012
rect 19208 17000 19214 17052
rect 20162 17040 20168 17052
rect 20123 17012 20168 17040
rect 20162 17000 20168 17012
rect 20220 17000 20226 17052
rect 20530 17040 20536 17052
rect 20491 17012 20536 17040
rect 20530 17000 20536 17012
rect 20588 17000 20594 17052
rect 23842 17040 23848 17052
rect 23803 17012 23848 17040
rect 23842 17000 23848 17012
rect 23900 17000 23906 17052
rect 24118 17000 24124 17052
rect 24176 17040 24182 17052
rect 24765 17043 24823 17049
rect 24765 17040 24777 17043
rect 24176 17012 24777 17040
rect 24176 17000 24182 17012
rect 24765 17009 24777 17012
rect 24811 17009 24823 17043
rect 25498 17040 25504 17052
rect 25459 17012 25504 17040
rect 24765 17003 24823 17009
rect 25498 17000 25504 17012
rect 25556 17000 25562 17052
rect 26326 17040 26332 17052
rect 26287 17012 26332 17040
rect 26326 17000 26332 17012
rect 26384 17000 26390 17052
rect 12069 16975 12127 16981
rect 12069 16941 12081 16975
rect 12115 16972 12127 16975
rect 13081 16975 13139 16981
rect 13081 16972 13093 16975
rect 12115 16944 13093 16972
rect 12115 16941 12127 16944
rect 12069 16935 12127 16941
rect 13081 16941 13093 16944
rect 13127 16941 13139 16975
rect 13081 16935 13139 16941
rect 12158 16864 12164 16916
rect 12216 16904 12222 16916
rect 12618 16904 12624 16916
rect 12216 16876 12624 16904
rect 12216 16864 12222 16876
rect 12618 16864 12624 16876
rect 12676 16864 12682 16916
rect 13096 16904 13124 16935
rect 14182 16904 14188 16916
rect 13096 16876 13492 16904
rect 14143 16876 14188 16904
rect 12250 16796 12256 16848
rect 12308 16836 12314 16848
rect 13354 16836 13360 16848
rect 12308 16808 13360 16836
rect 12308 16796 12314 16808
rect 11882 16768 11888 16780
rect 11843 16740 11888 16768
rect 11882 16728 11888 16740
rect 11940 16768 11946 16780
rect 12529 16771 12587 16777
rect 12529 16768 12541 16771
rect 11940 16740 12541 16768
rect 11940 16728 11946 16740
rect 12529 16737 12541 16740
rect 12575 16737 12587 16771
rect 12529 16731 12587 16737
rect 12437 16703 12495 16709
rect 12437 16669 12449 16703
rect 12483 16700 12495 16703
rect 12636 16700 12664 16808
rect 13354 16796 13360 16808
rect 13412 16796 13418 16848
rect 13464 16768 13492 16876
rect 14182 16864 14188 16876
rect 14240 16864 14246 16916
rect 14752 16904 14780 17000
rect 17586 16972 17592 16984
rect 17547 16944 17592 16972
rect 17586 16932 17592 16944
rect 17644 16932 17650 16984
rect 15102 16904 15108 16916
rect 14752 16876 15108 16904
rect 15102 16864 15108 16876
rect 15160 16904 15166 16916
rect 15160 16876 15424 16904
rect 15160 16864 15166 16876
rect 13541 16839 13599 16845
rect 13541 16805 13553 16839
rect 13587 16836 13599 16839
rect 13998 16836 14004 16848
rect 13587 16808 14004 16836
rect 13587 16805 13599 16808
rect 13541 16799 13599 16805
rect 13998 16796 14004 16808
rect 14056 16796 14062 16848
rect 15289 16839 15347 16845
rect 15289 16836 15301 16839
rect 15028 16808 15301 16836
rect 14093 16771 14151 16777
rect 14093 16768 14105 16771
rect 13464 16740 14105 16768
rect 14093 16737 14105 16740
rect 14139 16737 14151 16771
rect 14093 16731 14151 16737
rect 12483 16672 12664 16700
rect 12483 16669 12495 16672
rect 12437 16663 12495 16669
rect 13722 16660 13728 16712
rect 13780 16700 13786 16712
rect 15028 16709 15056 16808
rect 15289 16805 15301 16808
rect 15335 16805 15347 16839
rect 15396 16836 15424 16876
rect 15545 16839 15603 16845
rect 15545 16836 15557 16839
rect 15396 16808 15557 16836
rect 15289 16799 15347 16805
rect 15545 16805 15557 16808
rect 15591 16805 15603 16839
rect 15545 16799 15603 16805
rect 17034 16796 17040 16848
rect 17092 16836 17098 16848
rect 17604 16836 17632 16932
rect 17788 16904 17816 17000
rect 24026 16972 24032 16984
rect 23032 16944 24032 16972
rect 18325 16907 18383 16913
rect 18325 16904 18337 16907
rect 17788 16876 18337 16904
rect 18325 16873 18337 16876
rect 18371 16873 18383 16907
rect 18325 16867 18383 16873
rect 20901 16907 20959 16913
rect 20901 16873 20913 16907
rect 20947 16904 20959 16907
rect 20990 16904 20996 16916
rect 20947 16876 20996 16904
rect 20947 16873 20959 16876
rect 20901 16867 20959 16873
rect 20990 16864 20996 16876
rect 21048 16864 21054 16916
rect 23032 16913 23060 16944
rect 24026 16932 24032 16944
rect 24084 16932 24090 16984
rect 26234 16932 26240 16984
rect 26292 16972 26298 16984
rect 27522 16972 27528 16984
rect 26292 16944 27528 16972
rect 26292 16932 26298 16944
rect 27522 16932 27528 16944
rect 27580 16932 27586 16984
rect 23017 16907 23075 16913
rect 23017 16873 23029 16907
rect 23063 16873 23075 16907
rect 23017 16867 23075 16873
rect 24305 16907 24363 16913
rect 24305 16873 24317 16907
rect 24351 16904 24363 16907
rect 25406 16904 25412 16916
rect 24351 16876 25412 16904
rect 24351 16873 24363 16876
rect 24305 16867 24363 16873
rect 25406 16864 25412 16876
rect 25464 16864 25470 16916
rect 18233 16839 18291 16845
rect 18233 16836 18245 16839
rect 17092 16808 18245 16836
rect 17092 16796 17098 16808
rect 18233 16805 18245 16808
rect 18279 16805 18291 16839
rect 18233 16799 18291 16805
rect 23842 16796 23848 16848
rect 23900 16836 23906 16848
rect 24029 16839 24087 16845
rect 24029 16836 24041 16839
rect 23900 16808 24041 16836
rect 23900 16796 23906 16808
rect 24029 16805 24041 16808
rect 24075 16805 24087 16839
rect 25314 16836 25320 16848
rect 25275 16808 25320 16836
rect 24029 16799 24087 16805
rect 25314 16796 25320 16808
rect 25372 16836 25378 16848
rect 25869 16839 25927 16845
rect 25869 16836 25881 16839
rect 25372 16808 25881 16836
rect 25372 16796 25378 16808
rect 25869 16805 25881 16808
rect 25915 16805 25927 16839
rect 25869 16799 25927 16805
rect 17862 16728 17868 16780
rect 17920 16768 17926 16780
rect 18141 16771 18199 16777
rect 18141 16768 18153 16771
rect 17920 16740 18153 16768
rect 17920 16728 17926 16740
rect 18141 16737 18153 16740
rect 18187 16768 18199 16771
rect 19337 16771 19395 16777
rect 19337 16768 19349 16771
rect 18187 16740 19349 16768
rect 18187 16737 18199 16740
rect 18141 16731 18199 16737
rect 19337 16737 19349 16740
rect 19383 16737 19395 16771
rect 19337 16731 19395 16737
rect 15013 16703 15071 16709
rect 15013 16700 15025 16703
rect 13780 16672 15025 16700
rect 13780 16660 13786 16672
rect 15013 16669 15025 16672
rect 15059 16669 15071 16703
rect 17770 16700 17776 16712
rect 17731 16672 17776 16700
rect 15013 16663 15071 16669
rect 17770 16660 17776 16672
rect 17828 16660 17834 16712
rect 18782 16700 18788 16712
rect 18743 16672 18788 16700
rect 18782 16660 18788 16672
rect 18840 16660 18846 16712
rect 1104 16610 26864 16632
rect 1104 16558 10315 16610
rect 10367 16558 10379 16610
rect 10431 16558 10443 16610
rect 10495 16558 10507 16610
rect 10559 16558 19648 16610
rect 19700 16558 19712 16610
rect 19764 16558 19776 16610
rect 19828 16558 19840 16610
rect 19892 16558 26864 16610
rect 1104 16536 26864 16558
rect 12161 16499 12219 16505
rect 12161 16465 12173 16499
rect 12207 16496 12219 16499
rect 12250 16496 12256 16508
rect 12207 16468 12256 16496
rect 12207 16465 12219 16468
rect 12161 16459 12219 16465
rect 12250 16456 12256 16468
rect 12308 16456 12314 16508
rect 13538 16496 13544 16508
rect 13499 16468 13544 16496
rect 13538 16456 13544 16468
rect 13596 16456 13602 16508
rect 15102 16496 15108 16508
rect 15063 16468 15108 16496
rect 15102 16456 15108 16468
rect 15160 16456 15166 16508
rect 16206 16496 16212 16508
rect 16167 16468 16212 16496
rect 16206 16456 16212 16468
rect 16264 16456 16270 16508
rect 16390 16456 16396 16508
rect 16448 16496 16454 16508
rect 16577 16499 16635 16505
rect 16577 16496 16589 16499
rect 16448 16468 16589 16496
rect 16448 16456 16454 16468
rect 16577 16465 16589 16468
rect 16623 16465 16635 16499
rect 17862 16496 17868 16508
rect 17823 16468 17868 16496
rect 16577 16459 16635 16465
rect 17862 16456 17868 16468
rect 17920 16456 17926 16508
rect 18046 16496 18052 16508
rect 18007 16468 18052 16496
rect 18046 16456 18052 16468
rect 18104 16456 18110 16508
rect 18506 16496 18512 16508
rect 18467 16468 18512 16496
rect 18506 16456 18512 16468
rect 18564 16456 18570 16508
rect 21453 16499 21511 16505
rect 21453 16465 21465 16499
rect 21499 16496 21511 16499
rect 21818 16496 21824 16508
rect 21499 16468 21824 16496
rect 21499 16465 21511 16468
rect 21453 16459 21511 16465
rect 21818 16456 21824 16468
rect 21876 16456 21882 16508
rect 25406 16496 25412 16508
rect 25367 16468 25412 16496
rect 25406 16456 25412 16468
rect 25464 16456 25470 16508
rect 13992 16431 14050 16437
rect 13992 16397 14004 16431
rect 14038 16428 14050 16431
rect 14182 16428 14188 16440
rect 14038 16400 14188 16428
rect 14038 16397 14050 16400
rect 13992 16391 14050 16397
rect 14182 16388 14188 16400
rect 14240 16388 14246 16440
rect 15838 16428 15844 16440
rect 15799 16400 15844 16428
rect 15838 16388 15844 16400
rect 15896 16388 15902 16440
rect 16224 16428 16252 16456
rect 17313 16431 17371 16437
rect 17313 16428 17325 16431
rect 16224 16400 17325 16428
rect 17313 16397 17325 16400
rect 17359 16428 17371 16431
rect 17678 16428 17684 16440
rect 17359 16400 17684 16428
rect 17359 16397 17371 16400
rect 17313 16391 17371 16397
rect 17678 16388 17684 16400
rect 17736 16388 17742 16440
rect 17770 16388 17776 16440
rect 17828 16428 17834 16440
rect 18417 16431 18475 16437
rect 18417 16428 18429 16431
rect 17828 16400 18429 16428
rect 17828 16388 17834 16400
rect 18417 16397 18429 16400
rect 18463 16428 18475 16431
rect 19058 16428 19064 16440
rect 18463 16400 19064 16428
rect 18463 16397 18475 16400
rect 18417 16391 18475 16397
rect 19058 16388 19064 16400
rect 19116 16388 19122 16440
rect 24213 16431 24271 16437
rect 24213 16397 24225 16431
rect 24259 16428 24271 16431
rect 25314 16428 25320 16440
rect 24259 16400 25320 16428
rect 24259 16397 24271 16400
rect 24213 16391 24271 16397
rect 25314 16388 25320 16400
rect 25372 16388 25378 16440
rect 21634 16320 21640 16372
rect 21692 16360 21698 16372
rect 21821 16363 21879 16369
rect 21821 16360 21833 16363
rect 21692 16332 21833 16360
rect 21692 16320 21698 16332
rect 21821 16329 21833 16332
rect 21867 16329 21879 16363
rect 21821 16323 21879 16329
rect 23842 16320 23848 16372
rect 23900 16360 23906 16372
rect 23937 16363 23995 16369
rect 23937 16360 23949 16363
rect 23900 16332 23949 16360
rect 23900 16320 23906 16332
rect 23937 16329 23949 16332
rect 23983 16329 23995 16363
rect 25222 16360 25228 16372
rect 25183 16332 25228 16360
rect 23937 16323 23995 16329
rect 25222 16320 25228 16332
rect 25280 16320 25286 16372
rect 12434 16252 12440 16304
rect 12492 16292 12498 16304
rect 13722 16292 13728 16304
rect 12492 16264 13728 16292
rect 12492 16252 12498 16264
rect 13722 16252 13728 16264
rect 13780 16252 13786 16304
rect 18598 16252 18604 16304
rect 18656 16292 18662 16304
rect 18693 16295 18751 16301
rect 18693 16292 18705 16295
rect 18656 16264 18705 16292
rect 18656 16252 18662 16264
rect 18693 16261 18705 16264
rect 18739 16292 18751 16295
rect 19242 16292 19248 16304
rect 18739 16264 19248 16292
rect 18739 16261 18751 16264
rect 18693 16255 18751 16261
rect 19242 16252 19248 16264
rect 19300 16252 19306 16304
rect 21910 16292 21916 16304
rect 21871 16264 21916 16292
rect 21910 16252 21916 16264
rect 21968 16252 21974 16304
rect 22097 16295 22155 16301
rect 22097 16261 22109 16295
rect 22143 16292 22155 16295
rect 22143 16264 22416 16292
rect 22143 16261 22155 16264
rect 22097 16255 22155 16261
rect 22388 16168 22416 16264
rect 22370 16116 22376 16168
rect 22428 16156 22434 16168
rect 22465 16159 22523 16165
rect 22465 16156 22477 16159
rect 22428 16128 22477 16156
rect 22428 16116 22434 16128
rect 22465 16125 22477 16128
rect 22511 16125 22523 16159
rect 22465 16119 22523 16125
rect 1104 16066 26864 16088
rect 1104 16014 5648 16066
rect 5700 16014 5712 16066
rect 5764 16014 5776 16066
rect 5828 16014 5840 16066
rect 5892 16014 14982 16066
rect 15034 16014 15046 16066
rect 15098 16014 15110 16066
rect 15162 16014 15174 16066
rect 15226 16014 24315 16066
rect 24367 16014 24379 16066
rect 24431 16014 24443 16066
rect 24495 16014 24507 16066
rect 24559 16014 26864 16066
rect 1104 15992 26864 16014
rect 13909 15955 13967 15961
rect 13909 15921 13921 15955
rect 13955 15952 13967 15955
rect 14182 15952 14188 15964
rect 13955 15924 14188 15952
rect 13955 15921 13967 15924
rect 13909 15915 13967 15921
rect 14182 15912 14188 15924
rect 14240 15912 14246 15964
rect 15286 15952 15292 15964
rect 15247 15924 15292 15952
rect 15286 15912 15292 15924
rect 15344 15912 15350 15964
rect 18506 15912 18512 15964
rect 18564 15952 18570 15964
rect 18693 15955 18751 15961
rect 18693 15952 18705 15955
rect 18564 15924 18705 15952
rect 18564 15912 18570 15924
rect 18693 15921 18705 15924
rect 18739 15921 18751 15955
rect 19058 15952 19064 15964
rect 19019 15924 19064 15952
rect 18693 15915 18751 15921
rect 19058 15912 19064 15924
rect 19116 15912 19122 15964
rect 20714 15912 20720 15964
rect 20772 15952 20778 15964
rect 21821 15955 21879 15961
rect 21821 15952 21833 15955
rect 20772 15924 21833 15952
rect 20772 15912 20778 15924
rect 21821 15921 21833 15924
rect 21867 15921 21879 15955
rect 21821 15915 21879 15921
rect 13722 15844 13728 15896
rect 13780 15884 13786 15896
rect 14461 15887 14519 15893
rect 14461 15884 14473 15887
rect 13780 15856 14473 15884
rect 13780 15844 13786 15856
rect 14461 15853 14473 15856
rect 14507 15853 14519 15887
rect 14461 15847 14519 15853
rect 18417 15887 18475 15893
rect 18417 15853 18429 15887
rect 18463 15884 18475 15887
rect 18598 15884 18604 15896
rect 18463 15856 18604 15884
rect 18463 15853 18475 15856
rect 18417 15847 18475 15853
rect 18598 15844 18604 15856
rect 18656 15844 18662 15896
rect 15838 15816 15844 15828
rect 15799 15788 15844 15816
rect 15838 15776 15844 15788
rect 15896 15776 15902 15828
rect 17126 15816 17132 15828
rect 17087 15788 17132 15816
rect 17126 15776 17132 15788
rect 17184 15816 17190 15828
rect 17773 15819 17831 15825
rect 17773 15816 17785 15819
rect 17184 15788 17785 15816
rect 17184 15776 17190 15788
rect 17773 15785 17785 15788
rect 17819 15785 17831 15819
rect 17773 15779 17831 15785
rect 17865 15819 17923 15825
rect 17865 15785 17877 15819
rect 17911 15785 17923 15819
rect 21836 15816 21864 15915
rect 23842 15912 23848 15964
rect 23900 15952 23906 15964
rect 23937 15955 23995 15961
rect 23937 15952 23949 15955
rect 23900 15924 23949 15952
rect 23900 15912 23906 15924
rect 23937 15921 23949 15924
rect 23983 15921 23995 15955
rect 25222 15952 25228 15964
rect 25183 15924 25228 15952
rect 23937 15915 23995 15921
rect 25222 15912 25228 15924
rect 25280 15912 25286 15964
rect 23750 15844 23756 15896
rect 23808 15884 23814 15896
rect 24305 15887 24363 15893
rect 24305 15884 24317 15887
rect 23808 15856 24317 15884
rect 23808 15844 23814 15856
rect 24305 15853 24317 15856
rect 24351 15853 24363 15887
rect 24305 15847 24363 15853
rect 22005 15819 22063 15825
rect 22005 15816 22017 15819
rect 21836 15788 22017 15816
rect 17865 15779 17923 15785
rect 22005 15785 22017 15788
rect 22051 15785 22063 15819
rect 22005 15779 22063 15785
rect 12434 15708 12440 15760
rect 12492 15748 12498 15760
rect 12536 15751 12594 15757
rect 12536 15748 12548 15751
rect 12492 15720 12548 15748
rect 12492 15708 12498 15720
rect 12536 15717 12548 15720
rect 12582 15717 12594 15751
rect 12536 15711 12594 15717
rect 14826 15708 14832 15760
rect 14884 15748 14890 15760
rect 15105 15751 15163 15757
rect 15105 15748 15117 15751
rect 14884 15720 15117 15748
rect 14884 15708 14890 15720
rect 15105 15717 15117 15720
rect 15151 15748 15163 15751
rect 15749 15751 15807 15757
rect 15749 15748 15761 15751
rect 15151 15720 15761 15748
rect 15151 15717 15163 15720
rect 15105 15711 15163 15717
rect 15749 15717 15761 15720
rect 15795 15748 15807 15751
rect 16298 15748 16304 15760
rect 15795 15720 16304 15748
rect 15795 15717 15807 15720
rect 15749 15711 15807 15717
rect 16298 15708 16304 15720
rect 16356 15708 16362 15760
rect 16853 15751 16911 15757
rect 16853 15717 16865 15751
rect 16899 15748 16911 15751
rect 17880 15748 17908 15779
rect 23566 15776 23572 15828
rect 23624 15816 23630 15828
rect 23842 15816 23848 15828
rect 23624 15788 23848 15816
rect 23624 15776 23630 15788
rect 23842 15776 23848 15788
rect 23900 15776 23906 15828
rect 18230 15748 18236 15760
rect 16899 15720 18236 15748
rect 16899 15717 16911 15720
rect 16853 15711 16911 15717
rect 18230 15708 18236 15720
rect 18288 15708 18294 15760
rect 20717 15751 20775 15757
rect 20717 15717 20729 15751
rect 20763 15748 20775 15751
rect 21910 15748 21916 15760
rect 20763 15720 21916 15748
rect 20763 15717 20775 15720
rect 20717 15711 20775 15717
rect 21910 15708 21916 15720
rect 21968 15708 21974 15760
rect 24320 15748 24348 15847
rect 24765 15819 24823 15825
rect 24765 15785 24777 15819
rect 24811 15816 24823 15819
rect 25240 15816 25268 15912
rect 24811 15788 25268 15816
rect 24811 15785 24823 15788
rect 24765 15779 24823 15785
rect 24489 15751 24547 15757
rect 24489 15748 24501 15751
rect 24320 15720 24501 15748
rect 24489 15717 24501 15720
rect 24535 15717 24547 15751
rect 24489 15711 24547 15717
rect 12069 15683 12127 15689
rect 12069 15649 12081 15683
rect 12115 15680 12127 15683
rect 12618 15680 12624 15692
rect 12115 15652 12624 15680
rect 12115 15649 12127 15652
rect 12069 15643 12127 15649
rect 12618 15640 12624 15652
rect 12676 15680 12682 15692
rect 12796 15683 12854 15689
rect 12796 15680 12808 15683
rect 12676 15652 12808 15680
rect 12676 15640 12682 15652
rect 12796 15649 12808 15652
rect 12842 15680 12854 15683
rect 13814 15680 13820 15692
rect 12842 15652 13820 15680
rect 12842 15649 12854 15652
rect 12796 15643 12854 15649
rect 13814 15640 13820 15652
rect 13872 15640 13878 15692
rect 17678 15680 17684 15692
rect 17639 15652 17684 15680
rect 17678 15640 17684 15652
rect 17736 15640 17742 15692
rect 21177 15683 21235 15689
rect 21177 15649 21189 15683
rect 21223 15680 21235 15683
rect 22272 15683 22330 15689
rect 22272 15680 22284 15683
rect 21223 15652 22284 15680
rect 21223 15649 21235 15652
rect 21177 15643 21235 15649
rect 22272 15649 22284 15652
rect 22318 15680 22330 15683
rect 22370 15680 22376 15692
rect 22318 15652 22376 15680
rect 22318 15649 22330 15652
rect 22272 15643 22330 15649
rect 22370 15640 22376 15652
rect 22428 15640 22434 15692
rect 12434 15572 12440 15624
rect 12492 15612 12498 15624
rect 15654 15612 15660 15624
rect 12492 15584 12537 15612
rect 15615 15584 15660 15612
rect 12492 15572 12498 15584
rect 15654 15572 15660 15584
rect 15712 15572 15718 15624
rect 17310 15612 17316 15624
rect 17271 15584 17316 15612
rect 17310 15572 17316 15584
rect 17368 15572 17374 15624
rect 21545 15615 21603 15621
rect 21545 15581 21557 15615
rect 21591 15612 21603 15615
rect 21634 15612 21640 15624
rect 21591 15584 21640 15612
rect 21591 15581 21603 15584
rect 21545 15575 21603 15581
rect 21634 15572 21640 15584
rect 21692 15572 21698 15624
rect 22922 15572 22928 15624
rect 22980 15612 22986 15624
rect 23385 15615 23443 15621
rect 23385 15612 23397 15615
rect 22980 15584 23397 15612
rect 22980 15572 22986 15584
rect 23385 15581 23397 15584
rect 23431 15581 23443 15615
rect 23385 15575 23443 15581
rect 23474 15572 23480 15624
rect 23532 15612 23538 15624
rect 23750 15612 23756 15624
rect 23532 15584 23756 15612
rect 23532 15572 23538 15584
rect 23750 15572 23756 15584
rect 23808 15572 23814 15624
rect 1104 15522 26864 15544
rect 1104 15470 10315 15522
rect 10367 15470 10379 15522
rect 10431 15470 10443 15522
rect 10495 15470 10507 15522
rect 10559 15470 19648 15522
rect 19700 15470 19712 15522
rect 19764 15470 19776 15522
rect 19828 15470 19840 15522
rect 19892 15470 26864 15522
rect 1104 15448 26864 15470
rect 13814 15408 13820 15420
rect 13775 15380 13820 15408
rect 13814 15368 13820 15380
rect 13872 15368 13878 15420
rect 14182 15368 14188 15420
rect 14240 15408 14246 15420
rect 14369 15411 14427 15417
rect 14369 15408 14381 15411
rect 14240 15380 14381 15408
rect 14240 15368 14246 15380
rect 14369 15377 14381 15380
rect 14415 15377 14427 15411
rect 14369 15371 14427 15377
rect 14921 15411 14979 15417
rect 14921 15377 14933 15411
rect 14967 15408 14979 15411
rect 15473 15411 15531 15417
rect 15473 15408 15485 15411
rect 14967 15380 15485 15408
rect 14967 15377 14979 15380
rect 14921 15371 14979 15377
rect 15473 15377 15485 15380
rect 15519 15408 15531 15411
rect 15654 15408 15660 15420
rect 15519 15380 15660 15408
rect 15519 15377 15531 15380
rect 15473 15371 15531 15377
rect 14384 15340 14412 15371
rect 15654 15368 15660 15380
rect 15712 15368 15718 15420
rect 16390 15408 16396 15420
rect 16351 15380 16396 15408
rect 16390 15368 16396 15380
rect 16448 15368 16454 15420
rect 18230 15408 18236 15420
rect 18191 15380 18236 15408
rect 18230 15368 18236 15380
rect 18288 15408 18294 15420
rect 20533 15411 20591 15417
rect 20533 15408 20545 15411
rect 18288 15380 20545 15408
rect 18288 15368 18294 15380
rect 20533 15377 20545 15380
rect 20579 15377 20591 15411
rect 20533 15371 20591 15377
rect 21637 15411 21695 15417
rect 21637 15377 21649 15411
rect 21683 15408 21695 15411
rect 21910 15408 21916 15420
rect 21683 15380 21916 15408
rect 21683 15377 21695 15380
rect 21637 15371 21695 15377
rect 21910 15368 21916 15380
rect 21968 15368 21974 15420
rect 22097 15411 22155 15417
rect 22097 15408 22109 15411
rect 22020 15380 22109 15408
rect 15749 15343 15807 15349
rect 15749 15340 15761 15343
rect 14384 15312 15761 15340
rect 15749 15309 15761 15312
rect 15795 15340 15807 15343
rect 15838 15340 15844 15352
rect 15795 15312 15844 15340
rect 15795 15309 15807 15312
rect 15749 15303 15807 15309
rect 15838 15300 15844 15312
rect 15896 15300 15902 15352
rect 21266 15300 21272 15352
rect 21324 15340 21330 15352
rect 22020 15340 22048 15380
rect 22097 15377 22109 15380
rect 22143 15377 22155 15411
rect 24118 15408 24124 15420
rect 24079 15380 24124 15408
rect 22097 15371 22155 15377
rect 24118 15368 24124 15380
rect 24176 15368 24182 15420
rect 21324 15312 22048 15340
rect 21324 15300 21330 15312
rect 12710 15281 12716 15284
rect 12704 15235 12716 15281
rect 12768 15272 12774 15284
rect 16301 15275 16359 15281
rect 12768 15244 12804 15272
rect 12710 15232 12716 15235
rect 12768 15232 12774 15244
rect 16301 15241 16313 15275
rect 16347 15272 16359 15275
rect 16390 15272 16396 15284
rect 16347 15244 16396 15272
rect 16347 15241 16359 15244
rect 16301 15235 16359 15241
rect 16390 15232 16396 15244
rect 16448 15272 16454 15284
rect 16761 15275 16819 15281
rect 16761 15272 16773 15275
rect 16448 15244 16773 15272
rect 16448 15232 16454 15244
rect 16761 15241 16773 15244
rect 16807 15241 16819 15275
rect 16761 15235 16819 15241
rect 16850 15232 16856 15284
rect 16908 15272 16914 15284
rect 19420 15275 19478 15281
rect 16908 15244 16953 15272
rect 16908 15232 16914 15244
rect 19420 15241 19432 15275
rect 19466 15272 19478 15275
rect 20162 15272 20168 15284
rect 19466 15244 20168 15272
rect 19466 15241 19478 15244
rect 19420 15235 19478 15241
rect 20162 15232 20168 15244
rect 20220 15232 20226 15284
rect 20806 15232 20812 15284
rect 20864 15272 20870 15284
rect 22002 15272 22008 15284
rect 20864 15244 22008 15272
rect 20864 15232 20870 15244
rect 22002 15232 22008 15244
rect 22060 15232 22066 15284
rect 23474 15232 23480 15284
rect 23532 15272 23538 15284
rect 24029 15275 24087 15281
rect 24029 15272 24041 15275
rect 23532 15244 24041 15272
rect 23532 15232 23538 15244
rect 24029 15241 24041 15244
rect 24075 15241 24087 15275
rect 24029 15235 24087 15241
rect 25130 15232 25136 15284
rect 25188 15272 25194 15284
rect 25225 15275 25283 15281
rect 25225 15272 25237 15275
rect 25188 15244 25237 15272
rect 25188 15232 25194 15244
rect 25225 15241 25237 15244
rect 25271 15241 25283 15275
rect 25225 15235 25283 15241
rect 12434 15164 12440 15216
rect 12492 15204 12498 15216
rect 16942 15204 16948 15216
rect 12492 15176 12537 15204
rect 16903 15176 16948 15204
rect 12492 15164 12498 15176
rect 16942 15164 16948 15176
rect 17000 15164 17006 15216
rect 19150 15204 19156 15216
rect 19111 15176 19156 15204
rect 19150 15164 19156 15176
rect 19208 15164 19214 15216
rect 22189 15207 22247 15213
rect 22189 15204 22201 15207
rect 21468 15176 22201 15204
rect 21174 15028 21180 15080
rect 21232 15068 21238 15080
rect 21468 15077 21496 15176
rect 22189 15173 22201 15176
rect 22235 15173 22247 15207
rect 22189 15167 22247 15173
rect 24213 15207 24271 15213
rect 24213 15173 24225 15207
rect 24259 15173 24271 15207
rect 25406 15204 25412 15216
rect 25367 15176 25412 15204
rect 24213 15167 24271 15173
rect 24026 15096 24032 15148
rect 24084 15136 24090 15148
rect 24228 15136 24256 15167
rect 25406 15164 25412 15176
rect 25464 15164 25470 15216
rect 24084 15108 24256 15136
rect 24084 15096 24090 15108
rect 21453 15071 21511 15077
rect 21453 15068 21465 15071
rect 21232 15040 21465 15068
rect 21232 15028 21238 15040
rect 21453 15037 21465 15040
rect 21499 15037 21511 15071
rect 23658 15068 23664 15080
rect 23619 15040 23664 15068
rect 21453 15031 21511 15037
rect 23658 15028 23664 15040
rect 23716 15028 23722 15080
rect 1104 14978 26864 15000
rect 1104 14926 5648 14978
rect 5700 14926 5712 14978
rect 5764 14926 5776 14978
rect 5828 14926 5840 14978
rect 5892 14926 14982 14978
rect 15034 14926 15046 14978
rect 15098 14926 15110 14978
rect 15162 14926 15174 14978
rect 15226 14926 24315 14978
rect 24367 14926 24379 14978
rect 24431 14926 24443 14978
rect 24495 14926 24507 14978
rect 24559 14926 26864 14978
rect 1104 14904 26864 14926
rect 12710 14824 12716 14876
rect 12768 14864 12774 14876
rect 12805 14867 12863 14873
rect 12805 14864 12817 14867
rect 12768 14836 12817 14864
rect 12768 14824 12774 14836
rect 12805 14833 12817 14836
rect 12851 14833 12863 14867
rect 12805 14827 12863 14833
rect 16942 14824 16948 14876
rect 17000 14864 17006 14876
rect 17129 14867 17187 14873
rect 17129 14864 17141 14867
rect 17000 14836 17141 14864
rect 17000 14824 17006 14836
rect 17129 14833 17141 14836
rect 17175 14864 17187 14867
rect 17681 14867 17739 14873
rect 17681 14864 17693 14867
rect 17175 14836 17693 14864
rect 17175 14833 17187 14836
rect 17129 14827 17187 14833
rect 17681 14833 17693 14836
rect 17727 14833 17739 14867
rect 20714 14864 20720 14876
rect 20675 14836 20720 14864
rect 17681 14827 17739 14833
rect 20714 14824 20720 14836
rect 20772 14824 20778 14876
rect 23382 14864 23388 14876
rect 23343 14836 23388 14864
rect 23382 14824 23388 14836
rect 23440 14824 23446 14876
rect 24118 14824 24124 14876
rect 24176 14864 24182 14876
rect 24305 14867 24363 14873
rect 24305 14864 24317 14867
rect 24176 14836 24317 14864
rect 24176 14824 24182 14836
rect 24305 14833 24317 14836
rect 24351 14864 24363 14867
rect 24489 14867 24547 14873
rect 24489 14864 24501 14867
rect 24351 14836 24501 14864
rect 24351 14833 24363 14836
rect 24305 14827 24363 14833
rect 24489 14833 24501 14836
rect 24535 14833 24547 14867
rect 24489 14827 24547 14833
rect 25225 14867 25283 14873
rect 25225 14833 25237 14867
rect 25271 14864 25283 14867
rect 25314 14864 25320 14876
rect 25271 14836 25320 14864
rect 25271 14833 25283 14836
rect 25225 14827 25283 14833
rect 25314 14824 25320 14836
rect 25372 14824 25378 14876
rect 20732 14728 20760 14824
rect 22922 14796 22928 14808
rect 22883 14768 22928 14796
rect 22922 14756 22928 14768
rect 22980 14756 22986 14808
rect 23477 14799 23535 14805
rect 23477 14765 23489 14799
rect 23523 14796 23535 14799
rect 25130 14796 25136 14808
rect 23523 14768 25136 14796
rect 23523 14765 23535 14768
rect 23477 14759 23535 14765
rect 25130 14756 25136 14768
rect 25188 14796 25194 14808
rect 25593 14799 25651 14805
rect 25593 14796 25605 14799
rect 25188 14768 25605 14796
rect 25188 14756 25194 14768
rect 25593 14765 25605 14768
rect 25639 14765 25651 14799
rect 25593 14759 25651 14765
rect 20993 14731 21051 14737
rect 20993 14728 21005 14731
rect 20732 14700 21005 14728
rect 20993 14697 21005 14700
rect 21039 14697 21051 14731
rect 22940 14728 22968 14756
rect 24029 14731 24087 14737
rect 24029 14728 24041 14731
rect 22940 14700 24041 14728
rect 20993 14691 21051 14697
rect 24029 14697 24041 14700
rect 24075 14697 24087 14731
rect 24029 14691 24087 14697
rect 15657 14663 15715 14669
rect 15657 14629 15669 14663
rect 15703 14660 15715 14663
rect 15749 14663 15807 14669
rect 15749 14660 15761 14663
rect 15703 14632 15761 14660
rect 15703 14629 15715 14632
rect 15657 14623 15715 14629
rect 15749 14629 15761 14632
rect 15795 14660 15807 14663
rect 18141 14663 18199 14669
rect 18141 14660 18153 14663
rect 15795 14632 18153 14660
rect 15795 14629 15807 14632
rect 15749 14623 15807 14629
rect 18141 14629 18153 14632
rect 18187 14660 18199 14663
rect 18233 14663 18291 14669
rect 18233 14660 18245 14663
rect 18187 14632 18245 14660
rect 18187 14629 18199 14632
rect 18141 14623 18199 14629
rect 18233 14629 18245 14632
rect 18279 14629 18291 14663
rect 18233 14623 18291 14629
rect 16022 14601 16028 14604
rect 16016 14592 16028 14601
rect 15983 14564 16028 14592
rect 16016 14555 16028 14564
rect 16022 14552 16028 14555
rect 16080 14552 16086 14604
rect 18248 14592 18276 14623
rect 18322 14620 18328 14672
rect 18380 14660 18386 14672
rect 18489 14663 18547 14669
rect 18489 14660 18501 14663
rect 18380 14632 18501 14660
rect 18380 14620 18386 14632
rect 18489 14629 18501 14632
rect 18535 14629 18547 14663
rect 18489 14623 18547 14629
rect 23658 14620 23664 14672
rect 23716 14660 23722 14672
rect 23845 14663 23903 14669
rect 23845 14660 23857 14663
rect 23716 14632 23857 14660
rect 23716 14620 23722 14632
rect 23845 14629 23857 14632
rect 23891 14629 23903 14663
rect 25038 14660 25044 14672
rect 24999 14632 25044 14660
rect 23845 14623 23903 14629
rect 25038 14620 25044 14632
rect 25096 14620 25102 14672
rect 19150 14592 19156 14604
rect 18248 14564 19156 14592
rect 19150 14552 19156 14564
rect 19208 14552 19214 14604
rect 21174 14552 21180 14604
rect 21232 14601 21238 14604
rect 21232 14595 21296 14601
rect 21232 14561 21250 14595
rect 21284 14561 21296 14595
rect 21232 14555 21296 14561
rect 21232 14552 21238 14555
rect 23474 14552 23480 14604
rect 23532 14592 23538 14604
rect 23937 14595 23995 14601
rect 23937 14592 23949 14595
rect 23532 14564 23949 14592
rect 23532 14552 23538 14564
rect 23937 14561 23949 14564
rect 23983 14592 23995 14595
rect 24857 14595 24915 14601
rect 24857 14592 24869 14595
rect 23983 14564 24869 14592
rect 23983 14561 23995 14564
rect 23937 14555 23995 14561
rect 24857 14561 24869 14564
rect 24903 14561 24915 14595
rect 24857 14555 24915 14561
rect 12434 14484 12440 14536
rect 12492 14524 12498 14536
rect 12492 14496 12537 14524
rect 12492 14484 12498 14496
rect 19334 14484 19340 14536
rect 19392 14524 19398 14536
rect 19613 14527 19671 14533
rect 19613 14524 19625 14527
rect 19392 14496 19625 14524
rect 19392 14484 19398 14496
rect 19613 14493 19625 14496
rect 19659 14493 19671 14527
rect 22370 14524 22376 14536
rect 22283 14496 22376 14524
rect 19613 14487 19671 14493
rect 22370 14484 22376 14496
rect 22428 14524 22434 14536
rect 24026 14524 24032 14536
rect 22428 14496 24032 14524
rect 22428 14484 22434 14496
rect 24026 14484 24032 14496
rect 24084 14484 24090 14536
rect 24302 14524 24308 14536
rect 24263 14496 24308 14524
rect 24302 14484 24308 14496
rect 24360 14484 24366 14536
rect 1104 14434 26864 14456
rect 1104 14382 10315 14434
rect 10367 14382 10379 14434
rect 10431 14382 10443 14434
rect 10495 14382 10507 14434
rect 10559 14382 19648 14434
rect 19700 14382 19712 14434
rect 19764 14382 19776 14434
rect 19828 14382 19840 14434
rect 19892 14382 26864 14434
rect 1104 14360 26864 14382
rect 16390 14320 16396 14332
rect 16351 14292 16396 14320
rect 16390 14280 16396 14292
rect 16448 14280 16454 14332
rect 17310 14280 17316 14332
rect 17368 14320 17374 14332
rect 17405 14323 17463 14329
rect 17405 14320 17417 14323
rect 17368 14292 17417 14320
rect 17368 14280 17374 14292
rect 17405 14289 17417 14292
rect 17451 14289 17463 14323
rect 19150 14320 19156 14332
rect 19111 14292 19156 14320
rect 17405 14283 17463 14289
rect 19150 14280 19156 14292
rect 19208 14280 19214 14332
rect 19613 14323 19671 14329
rect 19613 14289 19625 14323
rect 19659 14320 19671 14323
rect 20162 14320 20168 14332
rect 19659 14292 20168 14320
rect 19659 14289 19671 14292
rect 19613 14283 19671 14289
rect 20162 14280 20168 14292
rect 20220 14280 20226 14332
rect 21082 14280 21088 14332
rect 21140 14320 21146 14332
rect 21545 14323 21603 14329
rect 21545 14320 21557 14323
rect 21140 14292 21557 14320
rect 21140 14280 21146 14292
rect 21545 14289 21557 14292
rect 21591 14289 21603 14323
rect 21545 14283 21603 14289
rect 22465 14323 22523 14329
rect 22465 14289 22477 14323
rect 22511 14320 22523 14323
rect 23382 14320 23388 14332
rect 22511 14292 23388 14320
rect 22511 14289 22523 14292
rect 22465 14283 22523 14289
rect 23382 14280 23388 14292
rect 23440 14280 23446 14332
rect 23477 14323 23535 14329
rect 23477 14289 23489 14323
rect 23523 14320 23535 14323
rect 23658 14320 23664 14332
rect 23523 14292 23664 14320
rect 23523 14289 23535 14292
rect 23477 14283 23535 14289
rect 23658 14280 23664 14292
rect 23716 14280 23722 14332
rect 23937 14323 23995 14329
rect 23937 14289 23949 14323
rect 23983 14320 23995 14323
rect 24026 14320 24032 14332
rect 23983 14292 24032 14320
rect 23983 14289 23995 14292
rect 23937 14283 23995 14289
rect 24026 14280 24032 14292
rect 24084 14280 24090 14332
rect 25038 14320 25044 14332
rect 24320 14292 25044 14320
rect 16301 14255 16359 14261
rect 16301 14221 16313 14255
rect 16347 14252 16359 14255
rect 16850 14252 16856 14264
rect 16347 14224 16856 14252
rect 16347 14221 16359 14224
rect 16301 14215 16359 14221
rect 16850 14212 16856 14224
rect 16908 14212 16914 14264
rect 21266 14212 21272 14264
rect 21324 14252 21330 14264
rect 24320 14261 24348 14292
rect 25038 14280 25044 14292
rect 25096 14280 25102 14332
rect 25498 14320 25504 14332
rect 25459 14292 25504 14320
rect 25498 14280 25504 14292
rect 25556 14280 25562 14332
rect 21913 14255 21971 14261
rect 21913 14252 21925 14255
rect 21324 14224 21925 14252
rect 21324 14212 21330 14224
rect 21913 14221 21925 14224
rect 21959 14221 21971 14255
rect 21913 14215 21971 14221
rect 24305 14255 24363 14261
rect 24305 14221 24317 14255
rect 24351 14221 24363 14255
rect 24305 14215 24363 14221
rect 16114 14144 16120 14196
rect 16172 14184 16178 14196
rect 16761 14187 16819 14193
rect 16761 14184 16773 14187
rect 16172 14156 16773 14184
rect 16172 14144 16178 14156
rect 16761 14153 16773 14156
rect 16807 14184 16819 14187
rect 18049 14187 18107 14193
rect 18049 14184 18061 14187
rect 16807 14156 18061 14184
rect 16807 14153 16819 14156
rect 16761 14147 16819 14153
rect 18049 14153 18061 14156
rect 18095 14153 18107 14187
rect 21358 14184 21364 14196
rect 21319 14156 21364 14184
rect 18049 14147 18107 14153
rect 21358 14144 21364 14156
rect 21416 14144 21422 14196
rect 24029 14187 24087 14193
rect 24029 14153 24041 14187
rect 24075 14184 24087 14187
rect 24762 14184 24768 14196
rect 24075 14156 24768 14184
rect 24075 14153 24087 14156
rect 24029 14147 24087 14153
rect 24762 14144 24768 14156
rect 24820 14144 24826 14196
rect 25317 14187 25375 14193
rect 25317 14153 25329 14187
rect 25363 14184 25375 14187
rect 25406 14184 25412 14196
rect 25363 14156 25412 14184
rect 25363 14153 25375 14156
rect 25317 14147 25375 14153
rect 25406 14144 25412 14156
rect 25464 14144 25470 14196
rect 16853 14119 16911 14125
rect 16853 14085 16865 14119
rect 16899 14116 16911 14119
rect 16942 14116 16948 14128
rect 16899 14088 16948 14116
rect 16899 14085 16911 14088
rect 16853 14079 16911 14085
rect 16942 14076 16948 14088
rect 17000 14076 17006 14128
rect 17037 14119 17095 14125
rect 17037 14085 17049 14119
rect 17083 14116 17095 14119
rect 17770 14116 17776 14128
rect 17083 14088 17776 14116
rect 17083 14085 17095 14088
rect 17037 14079 17095 14085
rect 15841 14051 15899 14057
rect 15841 14017 15853 14051
rect 15887 14048 15899 14051
rect 16022 14048 16028 14060
rect 15887 14020 16028 14048
rect 15887 14017 15899 14020
rect 15841 14011 15899 14017
rect 16022 14008 16028 14020
rect 16080 14048 16086 14060
rect 17052 14048 17080 14079
rect 17770 14076 17776 14088
rect 17828 14076 17834 14128
rect 16080 14020 17080 14048
rect 16080 14008 16086 14020
rect 24026 14008 24032 14060
rect 24084 14048 24090 14060
rect 24302 14048 24308 14060
rect 24084 14020 24308 14048
rect 24084 14008 24090 14020
rect 24302 14008 24308 14020
rect 24360 14008 24366 14060
rect 21085 13983 21143 13989
rect 21085 13949 21097 13983
rect 21131 13980 21143 13983
rect 21174 13980 21180 13992
rect 21131 13952 21180 13980
rect 21131 13949 21143 13952
rect 21085 13943 21143 13949
rect 21174 13940 21180 13952
rect 21232 13980 21238 13992
rect 22002 13980 22008 13992
rect 21232 13952 22008 13980
rect 21232 13940 21238 13952
rect 22002 13940 22008 13952
rect 22060 13940 22066 13992
rect 22278 13980 22284 13992
rect 22239 13952 22284 13980
rect 22278 13940 22284 13952
rect 22336 13940 22342 13992
rect 1104 13890 26864 13912
rect 1104 13838 5648 13890
rect 5700 13838 5712 13890
rect 5764 13838 5776 13890
rect 5828 13838 5840 13890
rect 5892 13838 14982 13890
rect 15034 13838 15046 13890
rect 15098 13838 15110 13890
rect 15162 13838 15174 13890
rect 15226 13838 24315 13890
rect 24367 13838 24379 13890
rect 24431 13838 24443 13890
rect 24495 13838 24507 13890
rect 24559 13838 26864 13890
rect 1104 13816 26864 13838
rect 15378 13736 15384 13788
rect 15436 13776 15442 13788
rect 15473 13779 15531 13785
rect 15473 13776 15485 13779
rect 15436 13748 15485 13776
rect 15436 13736 15442 13748
rect 15473 13745 15485 13748
rect 15519 13745 15531 13779
rect 16114 13776 16120 13788
rect 16075 13748 16120 13776
rect 15473 13739 15531 13745
rect 16114 13736 16120 13748
rect 16172 13736 16178 13788
rect 16850 13736 16856 13788
rect 16908 13776 16914 13788
rect 17129 13779 17187 13785
rect 17129 13776 17141 13779
rect 16908 13748 17141 13776
rect 16908 13736 16914 13748
rect 17129 13745 17141 13748
rect 17175 13745 17187 13779
rect 23658 13776 23664 13788
rect 23619 13748 23664 13776
rect 17129 13739 17187 13745
rect 23658 13736 23664 13748
rect 23716 13736 23722 13788
rect 24118 13776 24124 13788
rect 24079 13748 24124 13776
rect 24118 13736 24124 13748
rect 24176 13736 24182 13788
rect 24670 13736 24676 13788
rect 24728 13776 24734 13788
rect 24765 13779 24823 13785
rect 24765 13776 24777 13779
rect 24728 13748 24777 13776
rect 24728 13736 24734 13748
rect 24765 13745 24777 13748
rect 24811 13745 24823 13779
rect 24765 13739 24823 13745
rect 25406 13736 25412 13788
rect 25464 13776 25470 13788
rect 25501 13779 25559 13785
rect 25501 13776 25513 13779
rect 25464 13748 25513 13776
rect 25464 13736 25470 13748
rect 25501 13745 25513 13748
rect 25547 13745 25559 13779
rect 25501 13739 25559 13745
rect 16485 13711 16543 13717
rect 16485 13677 16497 13711
rect 16531 13708 16543 13711
rect 16942 13708 16948 13720
rect 16531 13680 16948 13708
rect 16531 13677 16543 13680
rect 16485 13671 16543 13677
rect 16942 13668 16948 13680
rect 17000 13668 17006 13720
rect 17310 13600 17316 13652
rect 17368 13640 17374 13652
rect 17589 13643 17647 13649
rect 17589 13640 17601 13643
rect 17368 13612 17601 13640
rect 17368 13600 17374 13612
rect 17589 13609 17601 13612
rect 17635 13609 17647 13643
rect 17770 13640 17776 13652
rect 17731 13612 17776 13640
rect 17589 13603 17647 13609
rect 17770 13600 17776 13612
rect 17828 13600 17834 13652
rect 21358 13640 21364 13652
rect 21271 13612 21364 13640
rect 21358 13600 21364 13612
rect 21416 13640 21422 13652
rect 21821 13643 21879 13649
rect 21821 13640 21833 13643
rect 21416 13612 21833 13640
rect 21416 13600 21422 13612
rect 21821 13609 21833 13612
rect 21867 13609 21879 13643
rect 21821 13603 21879 13609
rect 24489 13643 24547 13649
rect 24489 13609 24501 13643
rect 24535 13640 24547 13643
rect 24762 13640 24768 13652
rect 24535 13612 24768 13640
rect 24535 13609 24547 13612
rect 24489 13603 24547 13609
rect 24762 13600 24768 13612
rect 24820 13600 24826 13652
rect 25222 13640 25228 13652
rect 25183 13612 25228 13640
rect 25222 13600 25228 13612
rect 25280 13600 25286 13652
rect 15105 13575 15163 13581
rect 15105 13541 15117 13575
rect 15151 13572 15163 13575
rect 15289 13575 15347 13581
rect 15289 13572 15301 13575
rect 15151 13544 15301 13572
rect 15151 13541 15163 13544
rect 15105 13535 15163 13541
rect 15289 13541 15301 13544
rect 15335 13572 15347 13575
rect 15470 13572 15476 13584
rect 15335 13544 15476 13572
rect 15335 13541 15347 13544
rect 15289 13535 15347 13541
rect 15470 13532 15476 13544
rect 15528 13532 15534 13584
rect 17037 13575 17095 13581
rect 17037 13541 17049 13575
rect 17083 13572 17095 13575
rect 17494 13572 17500 13584
rect 17083 13544 17500 13572
rect 17083 13541 17095 13544
rect 17037 13535 17095 13541
rect 17494 13532 17500 13544
rect 17552 13532 17558 13584
rect 20714 13572 20720 13584
rect 20675 13544 20720 13572
rect 20714 13532 20720 13544
rect 20772 13572 20778 13584
rect 21085 13575 21143 13581
rect 21085 13572 21097 13575
rect 20772 13544 21097 13572
rect 20772 13532 20778 13544
rect 21085 13541 21097 13544
rect 21131 13541 21143 13575
rect 21085 13535 21143 13541
rect 23477 13575 23535 13581
rect 23477 13541 23489 13575
rect 23523 13572 23535 13575
rect 24118 13572 24124 13584
rect 23523 13544 24124 13572
rect 23523 13541 23535 13544
rect 23477 13535 23535 13541
rect 24118 13532 24124 13544
rect 24176 13532 24182 13584
rect 24581 13575 24639 13581
rect 24581 13541 24593 13575
rect 24627 13572 24639 13575
rect 25240 13572 25268 13600
rect 24627 13544 25268 13572
rect 24627 13541 24639 13544
rect 24581 13535 24639 13541
rect 1104 13346 26864 13368
rect 1104 13294 10315 13346
rect 10367 13294 10379 13346
rect 10431 13294 10443 13346
rect 10495 13294 10507 13346
rect 10559 13294 19648 13346
rect 19700 13294 19712 13346
rect 19764 13294 19776 13346
rect 19828 13294 19840 13346
rect 19892 13294 26864 13346
rect 1104 13272 26864 13294
rect 13630 13232 13636 13244
rect 13591 13204 13636 13232
rect 13630 13192 13636 13204
rect 13688 13192 13694 13244
rect 16945 13235 17003 13241
rect 16945 13201 16957 13235
rect 16991 13232 17003 13235
rect 17218 13232 17224 13244
rect 16991 13204 17224 13232
rect 16991 13201 17003 13204
rect 16945 13195 17003 13201
rect 17218 13192 17224 13204
rect 17276 13192 17282 13244
rect 17405 13235 17463 13241
rect 17405 13201 17417 13235
rect 17451 13232 17463 13235
rect 17770 13232 17776 13244
rect 17451 13204 17776 13232
rect 17451 13201 17463 13204
rect 17405 13195 17463 13201
rect 16485 13167 16543 13173
rect 16485 13133 16497 13167
rect 16531 13164 16543 13167
rect 17420 13164 17448 13195
rect 17770 13192 17776 13204
rect 17828 13192 17834 13244
rect 22002 13232 22008 13244
rect 21963 13204 22008 13232
rect 22002 13192 22008 13204
rect 22060 13192 22066 13244
rect 24210 13192 24216 13244
rect 24268 13232 24274 13244
rect 24765 13235 24823 13241
rect 24765 13232 24777 13235
rect 24268 13204 24777 13232
rect 24268 13192 24274 13204
rect 24765 13201 24777 13204
rect 24811 13201 24823 13235
rect 24765 13195 24823 13201
rect 16531 13136 17448 13164
rect 16531 13133 16543 13136
rect 16485 13127 16543 13133
rect 20806 13124 20812 13176
rect 20864 13173 20870 13176
rect 20864 13167 20928 13173
rect 20864 13133 20882 13167
rect 20916 13133 20928 13167
rect 20864 13127 20928 13133
rect 20864 13124 20870 13127
rect 13446 13096 13452 13108
rect 13407 13068 13452 13096
rect 13446 13056 13452 13068
rect 13504 13056 13510 13108
rect 16758 13096 16764 13108
rect 16719 13068 16764 13096
rect 16758 13056 16764 13068
rect 16816 13056 16822 13108
rect 20622 13096 20628 13108
rect 20583 13068 20628 13096
rect 20622 13056 20628 13068
rect 20680 13056 20686 13108
rect 24578 13096 24584 13108
rect 24539 13068 24584 13096
rect 24578 13056 24584 13068
rect 24636 13056 24642 13108
rect 20533 12895 20591 12901
rect 20533 12861 20545 12895
rect 20579 12892 20591 12895
rect 20990 12892 20996 12904
rect 20579 12864 20996 12892
rect 20579 12861 20591 12864
rect 20533 12855 20591 12861
rect 20990 12852 20996 12864
rect 21048 12852 21054 12904
rect 1104 12802 26864 12824
rect 1104 12750 5648 12802
rect 5700 12750 5712 12802
rect 5764 12750 5776 12802
rect 5828 12750 5840 12802
rect 5892 12750 14982 12802
rect 15034 12750 15046 12802
rect 15098 12750 15110 12802
rect 15162 12750 15174 12802
rect 15226 12750 24315 12802
rect 24367 12750 24379 12802
rect 24431 12750 24443 12802
rect 24495 12750 24507 12802
rect 24559 12750 26864 12802
rect 1104 12728 26864 12750
rect 13446 12688 13452 12700
rect 13407 12660 13452 12688
rect 13446 12648 13452 12660
rect 13504 12648 13510 12700
rect 20254 12648 20260 12700
rect 20312 12688 20318 12700
rect 20349 12691 20407 12697
rect 20349 12688 20361 12691
rect 20312 12660 20361 12688
rect 20312 12648 20318 12660
rect 20349 12657 20361 12660
rect 20395 12688 20407 12691
rect 20622 12688 20628 12700
rect 20395 12660 20628 12688
rect 20395 12657 20407 12660
rect 20349 12651 20407 12657
rect 20622 12648 20628 12660
rect 20680 12648 20686 12700
rect 23934 12688 23940 12700
rect 23895 12660 23940 12688
rect 23934 12648 23940 12660
rect 23992 12648 23998 12700
rect 24670 12688 24676 12700
rect 24631 12660 24676 12688
rect 24670 12648 24676 12660
rect 24728 12648 24734 12700
rect 25501 12691 25559 12697
rect 25501 12657 25513 12691
rect 25547 12688 25559 12691
rect 25590 12688 25596 12700
rect 25547 12660 25596 12688
rect 25547 12657 25559 12660
rect 25501 12651 25559 12657
rect 12897 12555 12955 12561
rect 12897 12521 12909 12555
rect 12943 12552 12955 12555
rect 13464 12552 13492 12648
rect 15470 12552 15476 12564
rect 12943 12524 13492 12552
rect 15431 12524 15476 12552
rect 12943 12521 12955 12524
rect 12897 12515 12955 12521
rect 15470 12512 15476 12524
rect 15528 12512 15534 12564
rect 16758 12512 16764 12564
rect 16816 12552 16822 12564
rect 16853 12555 16911 12561
rect 16853 12552 16865 12555
rect 16816 12524 16865 12552
rect 16816 12512 16822 12524
rect 16853 12521 16865 12524
rect 16899 12552 16911 12555
rect 17589 12555 17647 12561
rect 17589 12552 17601 12555
rect 16899 12524 17601 12552
rect 16899 12521 16911 12524
rect 16853 12515 16911 12521
rect 17589 12521 17601 12524
rect 17635 12521 17647 12555
rect 20640 12552 20668 12648
rect 20901 12555 20959 12561
rect 20901 12552 20913 12555
rect 20640 12524 20913 12552
rect 17589 12515 17647 12521
rect 20901 12521 20913 12524
rect 20947 12521 20959 12555
rect 24394 12552 24400 12564
rect 24355 12524 24400 12552
rect 20901 12515 20959 12521
rect 24394 12512 24400 12524
rect 24452 12512 24458 12564
rect 12526 12484 12532 12496
rect 12439 12456 12532 12484
rect 12526 12444 12532 12456
rect 12584 12484 12590 12496
rect 12621 12487 12679 12493
rect 12621 12484 12633 12487
rect 12584 12456 12633 12484
rect 12584 12444 12590 12456
rect 12621 12453 12633 12456
rect 12667 12453 12679 12487
rect 12621 12447 12679 12453
rect 15289 12487 15347 12493
rect 15289 12453 15301 12487
rect 15335 12484 15347 12487
rect 15654 12484 15660 12496
rect 15335 12456 15660 12484
rect 15335 12453 15347 12456
rect 15289 12447 15347 12453
rect 15654 12444 15660 12456
rect 15712 12484 15718 12496
rect 16025 12487 16083 12493
rect 16025 12484 16037 12487
rect 15712 12456 16037 12484
rect 15712 12444 15718 12456
rect 16025 12453 16037 12456
rect 16071 12453 16083 12487
rect 16025 12447 16083 12453
rect 17405 12487 17463 12493
rect 17405 12453 17417 12487
rect 17451 12484 17463 12487
rect 17451 12456 18276 12484
rect 17451 12453 17463 12456
rect 17405 12447 17463 12453
rect 18248 12357 18276 12456
rect 20990 12444 20996 12496
rect 21048 12484 21054 12496
rect 21157 12487 21215 12493
rect 21157 12484 21169 12487
rect 21048 12456 21169 12484
rect 21048 12444 21054 12456
rect 21157 12453 21169 12456
rect 21203 12453 21215 12487
rect 21157 12447 21215 12453
rect 23753 12487 23811 12493
rect 23753 12453 23765 12487
rect 23799 12484 23811 12487
rect 24412 12484 24440 12512
rect 23799 12456 24440 12484
rect 24857 12487 24915 12493
rect 23799 12453 23811 12456
rect 23753 12447 23811 12453
rect 24857 12453 24869 12487
rect 24903 12484 24915 12487
rect 25516 12484 25544 12651
rect 25590 12648 25596 12660
rect 25648 12648 25654 12700
rect 24903 12456 25544 12484
rect 24903 12453 24915 12456
rect 24857 12447 24915 12453
rect 23842 12376 23848 12428
rect 23900 12416 23906 12428
rect 24118 12416 24124 12428
rect 23900 12388 24124 12416
rect 23900 12376 23906 12388
rect 24118 12376 24124 12388
rect 24176 12376 24182 12428
rect 18233 12351 18291 12357
rect 18233 12317 18245 12351
rect 18279 12348 18291 12351
rect 18322 12348 18328 12360
rect 18279 12320 18328 12348
rect 18279 12317 18291 12320
rect 18233 12311 18291 12317
rect 18322 12308 18328 12320
rect 18380 12308 18386 12360
rect 19797 12351 19855 12357
rect 19797 12317 19809 12351
rect 19843 12348 19855 12351
rect 19978 12348 19984 12360
rect 19843 12320 19984 12348
rect 19843 12317 19855 12320
rect 19797 12311 19855 12317
rect 19978 12308 19984 12320
rect 20036 12308 20042 12360
rect 21910 12308 21916 12360
rect 21968 12348 21974 12360
rect 22281 12351 22339 12357
rect 22281 12348 22293 12351
rect 21968 12320 22293 12348
rect 21968 12308 21974 12320
rect 22281 12317 22293 12320
rect 22327 12317 22339 12351
rect 22281 12311 22339 12317
rect 25041 12351 25099 12357
rect 25041 12317 25053 12351
rect 25087 12348 25099 12351
rect 25682 12348 25688 12360
rect 25087 12320 25688 12348
rect 25087 12317 25099 12320
rect 25041 12311 25099 12317
rect 25682 12308 25688 12320
rect 25740 12308 25746 12360
rect 1104 12258 26864 12280
rect 1104 12206 10315 12258
rect 10367 12206 10379 12258
rect 10431 12206 10443 12258
rect 10495 12206 10507 12258
rect 10559 12206 19648 12258
rect 19700 12206 19712 12258
rect 19764 12206 19776 12258
rect 19828 12206 19840 12258
rect 19892 12206 26864 12258
rect 1104 12184 26864 12206
rect 12526 12104 12532 12156
rect 12584 12144 12590 12156
rect 13173 12147 13231 12153
rect 13173 12144 13185 12147
rect 12584 12116 13185 12144
rect 12584 12104 12590 12116
rect 13173 12113 13185 12116
rect 13219 12113 13231 12147
rect 15654 12144 15660 12156
rect 15615 12116 15660 12144
rect 13173 12107 13231 12113
rect 15654 12104 15660 12116
rect 15712 12104 15718 12156
rect 20714 12104 20720 12156
rect 20772 12144 20778 12156
rect 20809 12147 20867 12153
rect 20809 12144 20821 12147
rect 20772 12116 20821 12144
rect 20772 12104 20778 12116
rect 20809 12113 20821 12116
rect 20855 12113 20867 12147
rect 20809 12107 20867 12113
rect 24026 12104 24032 12156
rect 24084 12144 24090 12156
rect 24581 12147 24639 12153
rect 24581 12144 24593 12147
rect 24084 12116 24593 12144
rect 24084 12104 24090 12116
rect 24581 12113 24593 12116
rect 24627 12113 24639 12147
rect 24581 12107 24639 12113
rect 13262 11968 13268 12020
rect 13320 12008 13326 12020
rect 13541 12011 13599 12017
rect 13541 12008 13553 12011
rect 13320 11980 13553 12008
rect 13320 11968 13326 11980
rect 13541 11977 13553 11980
rect 13587 11977 13599 12011
rect 16022 12008 16028 12020
rect 15983 11980 16028 12008
rect 13541 11971 13599 11977
rect 16022 11968 16028 11980
rect 16080 11968 16086 12020
rect 19978 11968 19984 12020
rect 20036 12008 20042 12020
rect 21177 12011 21235 12017
rect 21177 12008 21189 12011
rect 20036 11980 21189 12008
rect 20036 11968 20042 11980
rect 21177 11977 21189 11980
rect 21223 11977 21235 12011
rect 24394 12008 24400 12020
rect 24355 11980 24400 12008
rect 21177 11971 21235 11977
rect 24394 11968 24400 11980
rect 24452 11968 24458 12020
rect 13630 11940 13636 11952
rect 13591 11912 13636 11940
rect 13630 11900 13636 11912
rect 13688 11900 13694 11952
rect 13817 11943 13875 11949
rect 13817 11909 13829 11943
rect 13863 11940 13875 11943
rect 13998 11940 14004 11952
rect 13863 11912 14004 11940
rect 13863 11909 13875 11912
rect 13817 11903 13875 11909
rect 13998 11900 14004 11912
rect 14056 11900 14062 11952
rect 15565 11943 15623 11949
rect 15565 11909 15577 11943
rect 15611 11940 15623 11943
rect 15930 11940 15936 11952
rect 15611 11912 15936 11940
rect 15611 11909 15623 11912
rect 15565 11903 15623 11909
rect 15930 11900 15936 11912
rect 15988 11940 15994 11952
rect 16117 11943 16175 11949
rect 16117 11940 16129 11943
rect 15988 11912 16129 11940
rect 15988 11900 15994 11912
rect 16117 11909 16129 11912
rect 16163 11909 16175 11943
rect 16117 11903 16175 11909
rect 16301 11943 16359 11949
rect 16301 11909 16313 11943
rect 16347 11940 16359 11943
rect 16390 11940 16396 11952
rect 16347 11912 16396 11940
rect 16347 11909 16359 11912
rect 16301 11903 16359 11909
rect 16390 11900 16396 11912
rect 16448 11900 16454 11952
rect 18230 11900 18236 11952
rect 18288 11940 18294 11952
rect 18325 11943 18383 11949
rect 18325 11940 18337 11943
rect 18288 11912 18337 11940
rect 18288 11900 18294 11912
rect 18325 11909 18337 11912
rect 18371 11909 18383 11943
rect 18325 11903 18383 11909
rect 20898 11900 20904 11952
rect 20956 11940 20962 11952
rect 21269 11943 21327 11949
rect 21269 11940 21281 11943
rect 20956 11912 21281 11940
rect 20956 11900 20962 11912
rect 21269 11909 21281 11912
rect 21315 11909 21327 11943
rect 21269 11903 21327 11909
rect 21453 11943 21511 11949
rect 21453 11909 21465 11943
rect 21499 11940 21511 11943
rect 21910 11940 21916 11952
rect 21499 11912 21916 11940
rect 21499 11909 21511 11912
rect 21453 11903 21511 11909
rect 20717 11875 20775 11881
rect 20717 11841 20729 11875
rect 20763 11872 20775 11875
rect 20806 11872 20812 11884
rect 20763 11844 20812 11872
rect 20763 11841 20775 11844
rect 20717 11835 20775 11841
rect 20806 11832 20812 11844
rect 20864 11872 20870 11884
rect 21468 11872 21496 11903
rect 21910 11900 21916 11912
rect 21968 11900 21974 11952
rect 20864 11844 21496 11872
rect 20864 11832 20870 11844
rect 12710 11804 12716 11816
rect 12671 11776 12716 11804
rect 12710 11764 12716 11776
rect 12768 11764 12774 11816
rect 18782 11804 18788 11816
rect 18743 11776 18788 11804
rect 18782 11764 18788 11776
rect 18840 11764 18846 11816
rect 1104 11714 26864 11736
rect 1104 11662 5648 11714
rect 5700 11662 5712 11714
rect 5764 11662 5776 11714
rect 5828 11662 5840 11714
rect 5892 11662 14982 11714
rect 15034 11662 15046 11714
rect 15098 11662 15110 11714
rect 15162 11662 15174 11714
rect 15226 11662 24315 11714
rect 24367 11662 24379 11714
rect 24431 11662 24443 11714
rect 24495 11662 24507 11714
rect 24559 11662 26864 11714
rect 1104 11640 26864 11662
rect 18322 11600 18328 11612
rect 18283 11572 18328 11600
rect 18322 11560 18328 11572
rect 18380 11560 18386 11612
rect 19978 11600 19984 11612
rect 19939 11572 19984 11600
rect 19978 11560 19984 11572
rect 20036 11560 20042 11612
rect 20898 11600 20904 11612
rect 20859 11572 20904 11600
rect 20898 11560 20904 11572
rect 20956 11560 20962 11612
rect 21910 11600 21916 11612
rect 21871 11572 21916 11600
rect 21910 11560 21916 11572
rect 21968 11560 21974 11612
rect 24489 11603 24547 11609
rect 24489 11569 24501 11603
rect 24535 11600 24547 11603
rect 24670 11600 24676 11612
rect 24535 11572 24676 11600
rect 24535 11569 24547 11572
rect 24489 11563 24547 11569
rect 24670 11560 24676 11572
rect 24728 11560 24734 11612
rect 18230 11532 18236 11544
rect 18191 11504 18236 11532
rect 18230 11492 18236 11504
rect 18288 11492 18294 11544
rect 12621 11399 12679 11405
rect 12621 11365 12633 11399
rect 12667 11365 12679 11399
rect 12621 11359 12679 11365
rect 12434 11288 12440 11340
rect 12492 11328 12498 11340
rect 12529 11331 12587 11337
rect 12529 11328 12541 11331
rect 12492 11300 12541 11328
rect 12492 11288 12498 11300
rect 12529 11297 12541 11300
rect 12575 11328 12587 11331
rect 12636 11328 12664 11359
rect 12710 11356 12716 11408
rect 12768 11396 12774 11408
rect 12877 11399 12935 11405
rect 12877 11396 12889 11399
rect 12768 11368 12889 11396
rect 12768 11356 12774 11368
rect 12877 11365 12889 11368
rect 12923 11365 12935 11399
rect 12877 11359 12935 11365
rect 14550 11356 14556 11408
rect 14608 11396 14614 11408
rect 15105 11399 15163 11405
rect 15105 11396 15117 11399
rect 14608 11368 15117 11396
rect 14608 11356 14614 11368
rect 15105 11365 15117 11368
rect 15151 11396 15163 11399
rect 15565 11399 15623 11405
rect 15565 11396 15577 11399
rect 15151 11368 15577 11396
rect 15151 11365 15163 11368
rect 15105 11359 15163 11365
rect 15565 11365 15577 11368
rect 15611 11396 15623 11399
rect 16298 11396 16304 11408
rect 15611 11368 16304 11396
rect 15611 11365 15623 11368
rect 15565 11359 15623 11365
rect 16298 11356 16304 11368
rect 16356 11356 16362 11408
rect 18248 11396 18276 11492
rect 18782 11464 18788 11476
rect 18743 11436 18788 11464
rect 18782 11424 18788 11436
rect 18840 11424 18846 11476
rect 18877 11467 18935 11473
rect 18877 11433 18889 11467
rect 18923 11433 18935 11467
rect 18877 11427 18935 11433
rect 18693 11399 18751 11405
rect 18693 11396 18705 11399
rect 18248 11368 18705 11396
rect 18693 11365 18705 11368
rect 18739 11365 18751 11399
rect 18693 11359 18751 11365
rect 14568 11328 14596 11356
rect 18892 11340 18920 11427
rect 20990 11424 20996 11476
rect 21048 11464 21054 11476
rect 21453 11467 21511 11473
rect 21453 11464 21465 11467
rect 21048 11436 21465 11464
rect 21048 11424 21054 11436
rect 21453 11433 21465 11436
rect 21499 11464 21511 11467
rect 22186 11464 22192 11476
rect 21499 11436 22192 11464
rect 21499 11433 21511 11436
rect 21453 11427 21511 11433
rect 22186 11424 22192 11436
rect 22244 11464 22250 11476
rect 22281 11467 22339 11473
rect 22281 11464 22293 11467
rect 22244 11436 22293 11464
rect 22244 11424 22250 11436
rect 22281 11433 22293 11436
rect 22327 11433 22339 11467
rect 22281 11427 22339 11433
rect 15810 11331 15868 11337
rect 15810 11328 15822 11331
rect 12575 11300 14596 11328
rect 14752 11300 15822 11328
rect 12575 11297 12587 11300
rect 12529 11291 12587 11297
rect 14752 11272 14780 11300
rect 15810 11297 15822 11300
rect 15856 11328 15868 11331
rect 16482 11328 16488 11340
rect 15856 11300 16488 11328
rect 15856 11297 15868 11300
rect 15810 11291 15868 11297
rect 16482 11288 16488 11300
rect 16540 11288 16546 11340
rect 17865 11331 17923 11337
rect 17865 11297 17877 11331
rect 17911 11328 17923 11331
rect 18874 11328 18880 11340
rect 17911 11300 18880 11328
rect 17911 11297 17923 11300
rect 17865 11291 17923 11297
rect 18874 11288 18880 11300
rect 18932 11288 18938 11340
rect 20717 11331 20775 11337
rect 20717 11297 20729 11331
rect 20763 11328 20775 11331
rect 21266 11328 21272 11340
rect 20763 11300 21272 11328
rect 20763 11297 20775 11300
rect 20717 11291 20775 11297
rect 21266 11288 21272 11300
rect 21324 11288 21330 11340
rect 13998 11260 14004 11272
rect 13959 11232 14004 11260
rect 13998 11220 14004 11232
rect 14056 11220 14062 11272
rect 14734 11260 14740 11272
rect 14695 11232 14740 11260
rect 14734 11220 14740 11232
rect 14792 11220 14798 11272
rect 16390 11220 16396 11272
rect 16448 11260 16454 11272
rect 16945 11263 17003 11269
rect 16945 11260 16957 11263
rect 16448 11232 16957 11260
rect 16448 11220 16454 11232
rect 16945 11229 16957 11232
rect 16991 11229 17003 11263
rect 16945 11223 17003 11229
rect 19518 11220 19524 11272
rect 19576 11260 19582 11272
rect 20349 11263 20407 11269
rect 20349 11260 20361 11263
rect 19576 11232 20361 11260
rect 19576 11220 19582 11232
rect 20349 11229 20361 11232
rect 20395 11260 20407 11263
rect 21361 11263 21419 11269
rect 21361 11260 21373 11263
rect 20395 11232 21373 11260
rect 20395 11229 20407 11232
rect 20349 11223 20407 11229
rect 21361 11229 21373 11232
rect 21407 11229 21419 11263
rect 21361 11223 21419 11229
rect 1104 11170 26864 11192
rect 1104 11118 10315 11170
rect 10367 11118 10379 11170
rect 10431 11118 10443 11170
rect 10495 11118 10507 11170
rect 10559 11118 19648 11170
rect 19700 11118 19712 11170
rect 19764 11118 19776 11170
rect 19828 11118 19840 11170
rect 19892 11118 26864 11170
rect 1104 11096 26864 11118
rect 12713 11059 12771 11065
rect 12713 11025 12725 11059
rect 12759 11056 12771 11059
rect 13262 11056 13268 11068
rect 12759 11028 13268 11056
rect 12759 11025 12771 11028
rect 12713 11019 12771 11025
rect 13262 11016 13268 11028
rect 13320 11016 13326 11068
rect 13630 11016 13636 11068
rect 13688 11056 13694 11068
rect 13909 11059 13967 11065
rect 13909 11056 13921 11059
rect 13688 11028 13921 11056
rect 13688 11016 13694 11028
rect 13909 11025 13921 11028
rect 13955 11025 13967 11059
rect 13909 11019 13967 11025
rect 14734 11016 14740 11068
rect 14792 11056 14798 11068
rect 15473 11059 15531 11065
rect 15473 11056 15485 11059
rect 14792 11028 15485 11056
rect 14792 11016 14798 11028
rect 15473 11025 15485 11028
rect 15519 11025 15531 11059
rect 16022 11056 16028 11068
rect 15983 11028 16028 11056
rect 15473 11019 15531 11025
rect 16022 11016 16028 11028
rect 16080 11056 16086 11068
rect 16577 11059 16635 11065
rect 16577 11056 16589 11059
rect 16080 11028 16589 11056
rect 16080 11016 16086 11028
rect 16577 11025 16589 11028
rect 16623 11025 16635 11059
rect 16577 11019 16635 11025
rect 18874 11016 18880 11068
rect 18932 11056 18938 11068
rect 19797 11059 19855 11065
rect 19797 11056 19809 11059
rect 18932 11028 19809 11056
rect 18932 11016 18938 11028
rect 19797 11025 19809 11028
rect 19843 11025 19855 11059
rect 19797 11019 19855 11025
rect 20809 11059 20867 11065
rect 20809 11025 20821 11059
rect 20855 11056 20867 11059
rect 20898 11056 20904 11068
rect 20855 11028 20904 11056
rect 20855 11025 20867 11028
rect 20809 11019 20867 11025
rect 16390 10988 16396 11000
rect 16351 10960 16396 10988
rect 16390 10948 16396 10960
rect 16448 10948 16454 11000
rect 19812 10988 19840 11019
rect 20898 11016 20904 11028
rect 20956 11016 20962 11068
rect 22186 11016 22192 11068
rect 22244 11056 22250 11068
rect 22281 11059 22339 11065
rect 22281 11056 22293 11059
rect 22244 11028 22293 11056
rect 22244 11016 22250 11028
rect 22281 11025 22293 11028
rect 22327 11025 22339 11059
rect 24762 11056 24768 11068
rect 24723 11028 24768 11056
rect 22281 11019 22339 11025
rect 24762 11016 24768 11028
rect 24820 11016 24826 11068
rect 21146 10991 21204 10997
rect 21146 10988 21158 10991
rect 19812 10960 21158 10988
rect 21146 10957 21158 10960
rect 21192 10988 21204 10991
rect 21358 10988 21364 11000
rect 21192 10960 21364 10988
rect 21192 10957 21204 10960
rect 21146 10951 21204 10957
rect 21358 10948 21364 10960
rect 21416 10948 21422 11000
rect 13633 10923 13691 10929
rect 13633 10889 13645 10923
rect 13679 10920 13691 10923
rect 13998 10920 14004 10932
rect 13679 10892 14004 10920
rect 13679 10889 13691 10892
rect 13633 10883 13691 10889
rect 13998 10880 14004 10892
rect 14056 10920 14062 10932
rect 14360 10923 14418 10929
rect 14360 10920 14372 10923
rect 14056 10892 14372 10920
rect 14056 10880 14062 10892
rect 14360 10889 14372 10892
rect 14406 10920 14418 10923
rect 14826 10920 14832 10932
rect 14406 10892 14832 10920
rect 14406 10889 14418 10892
rect 14360 10883 14418 10889
rect 14826 10880 14832 10892
rect 14884 10880 14890 10932
rect 18417 10923 18475 10929
rect 18417 10889 18429 10923
rect 18463 10920 18475 10923
rect 18506 10920 18512 10932
rect 18463 10892 18512 10920
rect 18463 10889 18475 10892
rect 18417 10883 18475 10889
rect 18506 10880 18512 10892
rect 18564 10880 18570 10932
rect 18690 10929 18696 10932
rect 18684 10920 18696 10929
rect 18651 10892 18696 10920
rect 18684 10883 18696 10892
rect 18690 10880 18696 10883
rect 18748 10880 18754 10932
rect 20254 10880 20260 10932
rect 20312 10920 20318 10932
rect 20901 10923 20959 10929
rect 20901 10920 20913 10923
rect 20312 10892 20913 10920
rect 20312 10880 20318 10892
rect 20901 10889 20913 10892
rect 20947 10920 20959 10923
rect 20990 10920 20996 10932
rect 20947 10892 20996 10920
rect 20947 10889 20959 10892
rect 20901 10883 20959 10889
rect 20990 10880 20996 10892
rect 21048 10880 21054 10932
rect 24581 10923 24639 10929
rect 24581 10889 24593 10923
rect 24627 10920 24639 10923
rect 24670 10920 24676 10932
rect 24627 10892 24676 10920
rect 24627 10889 24639 10892
rect 24581 10883 24639 10889
rect 24670 10880 24676 10892
rect 24728 10880 24734 10932
rect 14093 10855 14151 10861
rect 14093 10821 14105 10855
rect 14139 10821 14151 10855
rect 14093 10815 14151 10821
rect 14108 10716 14136 10815
rect 14458 10716 14464 10728
rect 14108 10688 14464 10716
rect 14458 10676 14464 10688
rect 14516 10676 14522 10728
rect 1104 10626 26864 10648
rect 1104 10574 5648 10626
rect 5700 10574 5712 10626
rect 5764 10574 5776 10626
rect 5828 10574 5840 10626
rect 5892 10574 14982 10626
rect 15034 10574 15046 10626
rect 15098 10574 15110 10626
rect 15162 10574 15174 10626
rect 15226 10574 24315 10626
rect 24367 10574 24379 10626
rect 24431 10574 24443 10626
rect 24495 10574 24507 10626
rect 24559 10574 26864 10626
rect 1104 10552 26864 10574
rect 12345 10515 12403 10521
rect 12345 10481 12357 10515
rect 12391 10512 12403 10515
rect 12710 10512 12716 10524
rect 12391 10484 12716 10512
rect 12391 10481 12403 10484
rect 12345 10475 12403 10481
rect 12710 10472 12716 10484
rect 12768 10512 12774 10524
rect 12897 10515 12955 10521
rect 12897 10512 12909 10515
rect 12768 10484 12909 10512
rect 12768 10472 12774 10484
rect 12897 10481 12909 10484
rect 12943 10481 12955 10515
rect 12897 10475 12955 10481
rect 13449 10515 13507 10521
rect 13449 10481 13461 10515
rect 13495 10512 13507 10515
rect 13630 10512 13636 10524
rect 13495 10484 13636 10512
rect 13495 10481 13507 10484
rect 13449 10475 13507 10481
rect 12912 10376 12940 10475
rect 13630 10472 13636 10484
rect 13688 10472 13694 10524
rect 14550 10512 14556 10524
rect 14511 10484 14556 10512
rect 14550 10472 14556 10484
rect 14608 10472 14614 10524
rect 14826 10512 14832 10524
rect 14787 10484 14832 10512
rect 14826 10472 14832 10484
rect 14884 10472 14890 10524
rect 16390 10512 16396 10524
rect 16351 10484 16396 10512
rect 16390 10472 16396 10484
rect 16448 10472 16454 10524
rect 16761 10515 16819 10521
rect 16761 10481 16773 10515
rect 16807 10512 16819 10515
rect 16850 10512 16856 10524
rect 16807 10484 16856 10512
rect 16807 10481 16819 10484
rect 16761 10475 16819 10481
rect 16850 10472 16856 10484
rect 16908 10512 16914 10524
rect 18874 10512 18880 10524
rect 16908 10484 18880 10512
rect 16908 10472 16914 10484
rect 18874 10472 18880 10484
rect 18932 10472 18938 10524
rect 20990 10472 20996 10524
rect 21048 10512 21054 10524
rect 21085 10515 21143 10521
rect 21085 10512 21097 10515
rect 21048 10484 21097 10512
rect 21048 10472 21054 10484
rect 21085 10481 21097 10484
rect 21131 10481 21143 10515
rect 21085 10475 21143 10481
rect 21358 10472 21364 10524
rect 21416 10512 21422 10524
rect 21453 10515 21511 10521
rect 21453 10512 21465 10515
rect 21416 10484 21465 10512
rect 21416 10472 21422 10484
rect 21453 10481 21465 10484
rect 21499 10481 21511 10515
rect 21453 10475 21511 10481
rect 23474 10472 23480 10524
rect 23532 10512 23538 10524
rect 24765 10515 24823 10521
rect 24765 10512 24777 10515
rect 23532 10484 24777 10512
rect 23532 10472 23538 10484
rect 24765 10481 24777 10484
rect 24811 10481 24823 10515
rect 24765 10475 24823 10481
rect 14001 10379 14059 10385
rect 14001 10376 14013 10379
rect 12912 10348 14013 10376
rect 14001 10345 14013 10348
rect 14047 10345 14059 10379
rect 16408 10376 16436 10472
rect 24489 10447 24547 10453
rect 24489 10413 24501 10447
rect 24535 10444 24547 10447
rect 24670 10444 24676 10456
rect 24535 10416 24676 10444
rect 24535 10413 24547 10416
rect 24489 10407 24547 10413
rect 24670 10404 24676 10416
rect 24728 10404 24734 10456
rect 16408 10348 16988 10376
rect 14001 10339 14059 10345
rect 10962 10308 10968 10320
rect 10923 10280 10968 10308
rect 10962 10268 10968 10280
rect 11020 10308 11026 10320
rect 12434 10308 12440 10320
rect 11020 10280 12440 10308
rect 11020 10268 11026 10280
rect 12434 10268 12440 10280
rect 12492 10268 12498 10320
rect 16298 10268 16304 10320
rect 16356 10308 16362 10320
rect 16850 10308 16856 10320
rect 16356 10280 16856 10308
rect 16356 10268 16362 10280
rect 16850 10268 16856 10280
rect 16908 10268 16914 10320
rect 16960 10308 16988 10348
rect 17109 10311 17167 10317
rect 17109 10308 17121 10311
rect 16960 10280 17121 10308
rect 17109 10277 17121 10280
rect 17155 10277 17167 10311
rect 17109 10271 17167 10277
rect 24581 10311 24639 10317
rect 24581 10277 24593 10311
rect 24627 10308 24639 10311
rect 24627 10280 25268 10308
rect 24627 10277 24639 10280
rect 24581 10271 24639 10277
rect 10778 10240 10784 10252
rect 10739 10212 10784 10240
rect 10778 10200 10784 10212
rect 10836 10240 10842 10252
rect 11210 10243 11268 10249
rect 11210 10240 11222 10243
rect 10836 10212 11222 10240
rect 10836 10200 10842 10212
rect 11210 10209 11222 10212
rect 11256 10209 11268 10243
rect 11210 10203 11268 10209
rect 13357 10243 13415 10249
rect 13357 10209 13369 10243
rect 13403 10240 13415 10243
rect 13814 10240 13820 10252
rect 13403 10212 13820 10240
rect 13403 10209 13415 10212
rect 13357 10203 13415 10209
rect 13814 10200 13820 10212
rect 13872 10200 13878 10252
rect 13906 10200 13912 10252
rect 13964 10240 13970 10252
rect 16390 10240 16396 10252
rect 13964 10212 16396 10240
rect 13964 10200 13970 10212
rect 16390 10200 16396 10212
rect 16448 10200 16454 10252
rect 18690 10240 18696 10252
rect 18248 10212 18696 10240
rect 18248 10181 18276 10212
rect 18690 10200 18696 10212
rect 18748 10240 18754 10252
rect 18748 10212 19288 10240
rect 18748 10200 18754 10212
rect 19260 10184 19288 10212
rect 25240 10184 25268 10280
rect 18233 10175 18291 10181
rect 18233 10141 18245 10175
rect 18279 10141 18291 10175
rect 19242 10172 19248 10184
rect 19203 10144 19248 10172
rect 18233 10135 18291 10141
rect 19242 10132 19248 10144
rect 19300 10132 19306 10184
rect 25222 10172 25228 10184
rect 25183 10144 25228 10172
rect 25222 10132 25228 10144
rect 25280 10132 25286 10184
rect 1104 10082 26864 10104
rect 1104 10030 10315 10082
rect 10367 10030 10379 10082
rect 10431 10030 10443 10082
rect 10495 10030 10507 10082
rect 10559 10030 19648 10082
rect 19700 10030 19712 10082
rect 19764 10030 19776 10082
rect 19828 10030 19840 10082
rect 19892 10030 26864 10082
rect 1104 10008 26864 10030
rect 10962 9968 10968 9980
rect 10923 9940 10968 9968
rect 10962 9928 10968 9940
rect 11020 9928 11026 9980
rect 13541 9971 13599 9977
rect 13541 9937 13553 9971
rect 13587 9968 13599 9971
rect 13906 9968 13912 9980
rect 13587 9940 13912 9968
rect 13587 9937 13599 9940
rect 13541 9931 13599 9937
rect 13906 9928 13912 9940
rect 13964 9928 13970 9980
rect 15930 9968 15936 9980
rect 15891 9940 15936 9968
rect 15930 9928 15936 9940
rect 15988 9928 15994 9980
rect 18782 9968 18788 9980
rect 18743 9940 18788 9968
rect 18782 9928 18788 9940
rect 18840 9928 18846 9980
rect 19150 9928 19156 9980
rect 19208 9968 19214 9980
rect 19245 9971 19303 9977
rect 19245 9968 19257 9971
rect 19208 9940 19257 9968
rect 19208 9928 19214 9940
rect 19245 9937 19257 9940
rect 19291 9968 19303 9971
rect 19518 9968 19524 9980
rect 19291 9940 19524 9968
rect 19291 9937 19303 9940
rect 19245 9931 19303 9937
rect 19518 9928 19524 9940
rect 19576 9928 19582 9980
rect 24762 9968 24768 9980
rect 24723 9940 24768 9968
rect 24762 9928 24768 9940
rect 24820 9928 24826 9980
rect 16022 9792 16028 9844
rect 16080 9832 16086 9844
rect 16301 9835 16359 9841
rect 16301 9832 16313 9835
rect 16080 9804 16313 9832
rect 16080 9792 16086 9804
rect 16301 9801 16313 9804
rect 16347 9801 16359 9835
rect 16301 9795 16359 9801
rect 18874 9792 18880 9844
rect 18932 9832 18938 9844
rect 19153 9835 19211 9841
rect 19153 9832 19165 9835
rect 18932 9804 19165 9832
rect 18932 9792 18938 9804
rect 19153 9801 19165 9804
rect 19199 9801 19211 9835
rect 19153 9795 19211 9801
rect 24581 9835 24639 9841
rect 24581 9801 24593 9835
rect 24627 9832 24639 9835
rect 24670 9832 24676 9844
rect 24627 9804 24676 9832
rect 24627 9801 24639 9804
rect 24581 9795 24639 9801
rect 24670 9792 24676 9804
rect 24728 9792 24734 9844
rect 16390 9764 16396 9776
rect 16351 9736 16396 9764
rect 16390 9724 16396 9736
rect 16448 9724 16454 9776
rect 16482 9724 16488 9776
rect 16540 9764 16546 9776
rect 19426 9764 19432 9776
rect 16540 9736 16585 9764
rect 19387 9736 19432 9764
rect 16540 9724 16546 9736
rect 19426 9724 19432 9736
rect 19484 9724 19490 9776
rect 1104 9538 26864 9560
rect 1104 9486 5648 9538
rect 5700 9486 5712 9538
rect 5764 9486 5776 9538
rect 5828 9486 5840 9538
rect 5892 9486 14982 9538
rect 15034 9486 15046 9538
rect 15098 9486 15110 9538
rect 15162 9486 15174 9538
rect 15226 9486 24315 9538
rect 24367 9486 24379 9538
rect 24431 9486 24443 9538
rect 24495 9486 24507 9538
rect 24559 9486 26864 9538
rect 1104 9464 26864 9486
rect 16390 9424 16396 9436
rect 16351 9396 16396 9424
rect 16390 9384 16396 9396
rect 16448 9384 16454 9436
rect 16482 9384 16488 9436
rect 16540 9384 16546 9436
rect 19150 9424 19156 9436
rect 19111 9396 19156 9424
rect 19150 9384 19156 9396
rect 19208 9384 19214 9436
rect 16500 9356 16528 9384
rect 16669 9359 16727 9365
rect 16669 9356 16681 9359
rect 16500 9328 16681 9356
rect 16669 9325 16681 9328
rect 16715 9325 16727 9359
rect 16669 9319 16727 9325
rect 19426 9316 19432 9368
rect 19484 9356 19490 9368
rect 19521 9359 19579 9365
rect 19521 9356 19533 9359
rect 19484 9328 19533 9356
rect 19484 9316 19490 9328
rect 19521 9325 19533 9328
rect 19567 9325 19579 9359
rect 24762 9356 24768 9368
rect 24723 9328 24768 9356
rect 19521 9319 19579 9325
rect 24762 9316 24768 9328
rect 24820 9316 24826 9368
rect 25222 9356 25228 9368
rect 25183 9328 25228 9356
rect 25222 9316 25228 9328
rect 25280 9316 25286 9368
rect 24581 9223 24639 9229
rect 24581 9220 24593 9223
rect 24504 9192 24593 9220
rect 24504 9096 24532 9192
rect 24581 9189 24593 9192
rect 24627 9189 24639 9223
rect 24581 9183 24639 9189
rect 16022 9084 16028 9096
rect 15983 9056 16028 9084
rect 16022 9044 16028 9056
rect 16080 9044 16086 9096
rect 18874 9084 18880 9096
rect 18835 9056 18880 9084
rect 18874 9044 18880 9056
rect 18932 9044 18938 9096
rect 24486 9084 24492 9096
rect 24447 9056 24492 9084
rect 24486 9044 24492 9056
rect 24544 9044 24550 9096
rect 1104 8994 26864 9016
rect 1104 8942 10315 8994
rect 10367 8942 10379 8994
rect 10431 8942 10443 8994
rect 10495 8942 10507 8994
rect 10559 8942 19648 8994
rect 19700 8942 19712 8994
rect 19764 8942 19776 8994
rect 19828 8942 19840 8994
rect 19892 8942 26864 8994
rect 1104 8920 26864 8942
rect 24762 8880 24768 8892
rect 24723 8852 24768 8880
rect 24762 8840 24768 8852
rect 24820 8840 24826 8892
rect 24581 8747 24639 8753
rect 24581 8713 24593 8747
rect 24627 8744 24639 8747
rect 24670 8744 24676 8756
rect 24627 8716 24676 8744
rect 24627 8713 24639 8716
rect 24581 8707 24639 8713
rect 24670 8704 24676 8716
rect 24728 8704 24734 8756
rect 1104 8450 26864 8472
rect 1104 8398 5648 8450
rect 5700 8398 5712 8450
rect 5764 8398 5776 8450
rect 5828 8398 5840 8450
rect 5892 8398 14982 8450
rect 15034 8398 15046 8450
rect 15098 8398 15110 8450
rect 15162 8398 15174 8450
rect 15226 8398 24315 8450
rect 24367 8398 24379 8450
rect 24431 8398 24443 8450
rect 24495 8398 24507 8450
rect 24559 8398 26864 8450
rect 1104 8376 26864 8398
rect 24670 8336 24676 8348
rect 24631 8308 24676 8336
rect 24670 8296 24676 8308
rect 24728 8296 24734 8348
rect 1104 7906 26864 7928
rect 1104 7854 10315 7906
rect 10367 7854 10379 7906
rect 10431 7854 10443 7906
rect 10495 7854 10507 7906
rect 10559 7854 19648 7906
rect 19700 7854 19712 7906
rect 19764 7854 19776 7906
rect 19828 7854 19840 7906
rect 19892 7854 26864 7906
rect 1104 7832 26864 7854
rect 24578 7656 24584 7668
rect 24539 7628 24584 7656
rect 24578 7616 24584 7628
rect 24636 7616 24642 7668
rect 24762 7520 24768 7532
rect 24723 7492 24768 7520
rect 24762 7480 24768 7492
rect 24820 7480 24826 7532
rect 1104 7362 26864 7384
rect 1104 7310 5648 7362
rect 5700 7310 5712 7362
rect 5764 7310 5776 7362
rect 5828 7310 5840 7362
rect 5892 7310 14982 7362
rect 15034 7310 15046 7362
rect 15098 7310 15110 7362
rect 15162 7310 15174 7362
rect 15226 7310 24315 7362
rect 24367 7310 24379 7362
rect 24431 7310 24443 7362
rect 24495 7310 24507 7362
rect 24559 7310 26864 7362
rect 1104 7288 26864 7310
rect 17773 7251 17831 7257
rect 17773 7217 17785 7251
rect 17819 7248 17831 7251
rect 17862 7248 17868 7260
rect 17819 7220 17868 7248
rect 17819 7217 17831 7220
rect 17773 7211 17831 7217
rect 17862 7208 17868 7220
rect 17920 7208 17926 7260
rect 23750 7208 23756 7260
rect 23808 7248 23814 7260
rect 23934 7248 23940 7260
rect 23808 7220 23940 7248
rect 23808 7208 23814 7220
rect 23934 7208 23940 7220
rect 23992 7208 23998 7260
rect 24670 7248 24676 7260
rect 24631 7220 24676 7248
rect 24670 7208 24676 7220
rect 24728 7208 24734 7260
rect 18230 7112 18236 7124
rect 17604 7084 18236 7112
rect 17604 7053 17632 7084
rect 18230 7072 18236 7084
rect 18288 7072 18294 7124
rect 17589 7047 17647 7053
rect 17589 7013 17601 7047
rect 17635 7013 17647 7047
rect 17589 7007 17647 7013
rect 1104 6818 26864 6840
rect 1104 6766 10315 6818
rect 10367 6766 10379 6818
rect 10431 6766 10443 6818
rect 10495 6766 10507 6818
rect 10559 6766 19648 6818
rect 19700 6766 19712 6818
rect 19764 6766 19776 6818
rect 19828 6766 19840 6818
rect 19892 6766 26864 6818
rect 1104 6744 26864 6766
rect 1104 6274 26864 6296
rect 1104 6222 5648 6274
rect 5700 6222 5712 6274
rect 5764 6222 5776 6274
rect 5828 6222 5840 6274
rect 5892 6222 14982 6274
rect 15034 6222 15046 6274
rect 15098 6222 15110 6274
rect 15162 6222 15174 6274
rect 15226 6222 24315 6274
rect 24367 6222 24379 6274
rect 24431 6222 24443 6274
rect 24495 6222 24507 6274
rect 24559 6222 26864 6274
rect 1104 6200 26864 6222
rect 16482 6160 16488 6172
rect 16443 6132 16488 6160
rect 16482 6120 16488 6132
rect 16540 6120 16546 6172
rect 16301 5959 16359 5965
rect 16301 5925 16313 5959
rect 16347 5925 16359 5959
rect 16301 5919 16359 5925
rect 16316 5888 16344 5919
rect 16942 5888 16948 5900
rect 16316 5860 16948 5888
rect 16942 5848 16948 5860
rect 17000 5848 17006 5900
rect 1104 5730 26864 5752
rect 1104 5678 10315 5730
rect 10367 5678 10379 5730
rect 10431 5678 10443 5730
rect 10495 5678 10507 5730
rect 10559 5678 19648 5730
rect 19700 5678 19712 5730
rect 19764 5678 19776 5730
rect 19828 5678 19840 5730
rect 19892 5678 26864 5730
rect 1104 5656 26864 5678
rect 1104 5186 26864 5208
rect 1104 5134 5648 5186
rect 5700 5134 5712 5186
rect 5764 5134 5776 5186
rect 5828 5134 5840 5186
rect 5892 5134 14982 5186
rect 15034 5134 15046 5186
rect 15098 5134 15110 5186
rect 15162 5134 15174 5186
rect 15226 5134 24315 5186
rect 24367 5134 24379 5186
rect 24431 5134 24443 5186
rect 24495 5134 24507 5186
rect 24559 5134 26864 5186
rect 1104 5112 26864 5134
rect 15473 5075 15531 5081
rect 15473 5041 15485 5075
rect 15519 5072 15531 5075
rect 15746 5072 15752 5084
rect 15519 5044 15752 5072
rect 15519 5041 15531 5044
rect 15473 5035 15531 5041
rect 15746 5032 15752 5044
rect 15804 5032 15810 5084
rect 15930 4936 15936 4948
rect 15304 4908 15936 4936
rect 15304 4877 15332 4908
rect 15930 4896 15936 4908
rect 15988 4896 15994 4948
rect 15289 4871 15347 4877
rect 15289 4837 15301 4871
rect 15335 4837 15347 4871
rect 15289 4831 15347 4837
rect 1104 4642 26864 4664
rect 1104 4590 10315 4642
rect 10367 4590 10379 4642
rect 10431 4590 10443 4642
rect 10495 4590 10507 4642
rect 10559 4590 19648 4642
rect 19700 4590 19712 4642
rect 19764 4590 19776 4642
rect 19828 4590 19840 4642
rect 19892 4590 26864 4642
rect 1104 4568 26864 4590
rect 1104 4098 26864 4120
rect 1104 4046 5648 4098
rect 5700 4046 5712 4098
rect 5764 4046 5776 4098
rect 5828 4046 5840 4098
rect 5892 4046 14982 4098
rect 15034 4046 15046 4098
rect 15098 4046 15110 4098
rect 15162 4046 15174 4098
rect 15226 4046 24315 4098
rect 24367 4046 24379 4098
rect 24431 4046 24443 4098
rect 24495 4046 24507 4098
rect 24559 4046 26864 4098
rect 1104 4024 26864 4046
rect 24581 3783 24639 3789
rect 24581 3749 24593 3783
rect 24627 3780 24639 3783
rect 24627 3752 25268 3780
rect 24627 3749 24639 3752
rect 24581 3743 24639 3749
rect 25240 3656 25268 3752
rect 24762 3644 24768 3656
rect 24723 3616 24768 3644
rect 24762 3604 24768 3616
rect 24820 3604 24826 3656
rect 25222 3644 25228 3656
rect 25183 3616 25228 3644
rect 25222 3604 25228 3616
rect 25280 3604 25286 3656
rect 1104 3554 26864 3576
rect 1104 3502 10315 3554
rect 10367 3502 10379 3554
rect 10431 3502 10443 3554
rect 10495 3502 10507 3554
rect 10559 3502 19648 3554
rect 19700 3502 19712 3554
rect 19764 3502 19776 3554
rect 19828 3502 19840 3554
rect 19892 3502 26864 3554
rect 1104 3480 26864 3502
rect 1104 3010 26864 3032
rect 1104 2958 5648 3010
rect 5700 2958 5712 3010
rect 5764 2958 5776 3010
rect 5828 2958 5840 3010
rect 5892 2958 14982 3010
rect 15034 2958 15046 3010
rect 15098 2958 15110 3010
rect 15162 2958 15174 3010
rect 15226 2958 24315 3010
rect 24367 2958 24379 3010
rect 24431 2958 24443 3010
rect 24495 2958 24507 3010
rect 24559 2958 26864 3010
rect 1104 2936 26864 2958
rect 1104 2466 26864 2488
rect 1104 2414 10315 2466
rect 10367 2414 10379 2466
rect 10431 2414 10443 2466
rect 10495 2414 10507 2466
rect 10559 2414 19648 2466
rect 19700 2414 19712 2466
rect 19764 2414 19776 2466
rect 19828 2414 19840 2466
rect 19892 2414 26864 2466
rect 1104 2392 26864 2414
rect 1104 1922 26864 1944
rect 1104 1870 5648 1922
rect 5700 1870 5712 1922
rect 5764 1870 5776 1922
rect 5828 1870 5840 1922
rect 5892 1870 14982 1922
rect 15034 1870 15046 1922
rect 15098 1870 15110 1922
rect 15162 1870 15174 1922
rect 15226 1870 24315 1922
rect 24367 1870 24379 1922
rect 24431 1870 24443 1922
rect 24495 1870 24507 1922
rect 24559 1870 26864 1922
rect 1104 1848 26864 1870
<< via1 >>
rect 21548 26384 21600 26436
rect 23940 26384 23992 26436
rect 10315 25262 10367 25314
rect 10379 25262 10431 25314
rect 10443 25262 10495 25314
rect 10507 25262 10559 25314
rect 19648 25262 19700 25314
rect 19712 25262 19764 25314
rect 19776 25262 19828 25314
rect 19840 25262 19892 25314
rect 23572 25160 23624 25212
rect 24768 25203 24820 25212
rect 24768 25169 24777 25203
rect 24777 25169 24811 25203
rect 24811 25169 24820 25203
rect 24768 25160 24820 25169
rect 22836 25067 22888 25076
rect 22836 25033 22845 25067
rect 22845 25033 22879 25067
rect 22879 25033 22888 25067
rect 22836 25024 22888 25033
rect 24768 25024 24820 25076
rect 5648 24718 5700 24770
rect 5712 24718 5764 24770
rect 5776 24718 5828 24770
rect 5840 24718 5892 24770
rect 14982 24718 15034 24770
rect 15046 24718 15098 24770
rect 15110 24718 15162 24770
rect 15174 24718 15226 24770
rect 24315 24718 24367 24770
rect 24379 24718 24431 24770
rect 24443 24718 24495 24770
rect 24507 24718 24559 24770
rect 25136 24659 25188 24668
rect 25136 24625 25145 24659
rect 25145 24625 25179 24659
rect 25179 24625 25188 24659
rect 25136 24616 25188 24625
rect 22836 24548 22888 24600
rect 15384 24480 15436 24532
rect 15936 24480 15988 24532
rect 20720 24480 20772 24532
rect 21640 24480 21692 24532
rect 19340 24412 19392 24464
rect 20444 24412 20496 24464
rect 22560 24455 22612 24464
rect 22560 24421 22569 24455
rect 22569 24421 22603 24455
rect 22603 24421 22612 24455
rect 22560 24412 22612 24421
rect 24124 24412 24176 24464
rect 24952 24455 25004 24464
rect 24952 24421 24961 24455
rect 24961 24421 24995 24455
rect 24995 24421 25004 24455
rect 24952 24412 25004 24421
rect 25320 24344 25372 24396
rect 19156 24276 19208 24328
rect 23388 24276 23440 24328
rect 24768 24319 24820 24328
rect 24768 24285 24777 24319
rect 24777 24285 24811 24319
rect 24811 24285 24820 24319
rect 24768 24276 24820 24285
rect 10315 24174 10367 24226
rect 10379 24174 10431 24226
rect 10443 24174 10495 24226
rect 10507 24174 10559 24226
rect 19648 24174 19700 24226
rect 19712 24174 19764 24226
rect 19776 24174 19828 24226
rect 19840 24174 19892 24226
rect 25136 24115 25188 24124
rect 25136 24081 25145 24115
rect 25145 24081 25179 24115
rect 25179 24081 25188 24115
rect 25136 24072 25188 24081
rect 24768 24004 24820 24056
rect 14832 23936 14884 23988
rect 19156 23936 19208 23988
rect 20352 23936 20404 23988
rect 22100 23936 22152 23988
rect 23388 23936 23440 23988
rect 23572 23936 23624 23988
rect 24860 23936 24912 23988
rect 10968 23911 11020 23920
rect 10968 23877 10977 23911
rect 10977 23877 11011 23911
rect 11011 23877 11020 23911
rect 10968 23868 11020 23877
rect 13268 23911 13320 23920
rect 13268 23877 13277 23911
rect 13277 23877 13311 23911
rect 13311 23877 13320 23911
rect 13268 23868 13320 23877
rect 16212 23911 16264 23920
rect 16212 23877 16221 23911
rect 16221 23877 16255 23911
rect 16255 23877 16264 23911
rect 16212 23868 16264 23877
rect 10876 23775 10928 23784
rect 10876 23741 10885 23775
rect 10885 23741 10919 23775
rect 10919 23741 10928 23775
rect 10876 23732 10928 23741
rect 14188 23732 14240 23784
rect 16028 23732 16080 23784
rect 18420 23775 18472 23784
rect 18420 23741 18429 23775
rect 18429 23741 18463 23775
rect 18463 23741 18472 23775
rect 18420 23732 18472 23741
rect 18604 23732 18656 23784
rect 19432 23911 19484 23920
rect 19432 23877 19441 23911
rect 19441 23877 19475 23911
rect 19475 23877 19484 23911
rect 19432 23868 19484 23877
rect 21180 23868 21232 23920
rect 22284 23868 22336 23920
rect 19340 23732 19392 23784
rect 22008 23732 22060 23784
rect 5648 23630 5700 23682
rect 5712 23630 5764 23682
rect 5776 23630 5828 23682
rect 5840 23630 5892 23682
rect 14982 23630 15034 23682
rect 15046 23630 15098 23682
rect 15110 23630 15162 23682
rect 15174 23630 15226 23682
rect 24315 23630 24367 23682
rect 24379 23630 24431 23682
rect 24443 23630 24495 23682
rect 24507 23630 24559 23682
rect 13360 23571 13412 23580
rect 13360 23537 13369 23571
rect 13369 23537 13403 23571
rect 13403 23537 13412 23571
rect 13360 23528 13412 23537
rect 14832 23528 14884 23580
rect 19248 23528 19300 23580
rect 20352 23571 20404 23580
rect 20352 23537 20361 23571
rect 20361 23537 20395 23571
rect 20395 23537 20404 23571
rect 20352 23528 20404 23537
rect 21180 23571 21232 23580
rect 21180 23537 21189 23571
rect 21189 23537 21223 23571
rect 21223 23537 21232 23571
rect 21180 23528 21232 23537
rect 25504 23571 25556 23580
rect 25504 23537 25513 23571
rect 25513 23537 25547 23571
rect 25547 23537 25556 23571
rect 25504 23528 25556 23537
rect 19432 23460 19484 23512
rect 14188 23435 14240 23444
rect 14188 23401 14197 23435
rect 14197 23401 14231 23435
rect 14231 23401 14240 23435
rect 14188 23392 14240 23401
rect 20720 23435 20772 23444
rect 20720 23401 20729 23435
rect 20729 23401 20763 23435
rect 20763 23401 20772 23435
rect 21548 23435 21600 23444
rect 20720 23392 20772 23401
rect 21548 23401 21557 23435
rect 21557 23401 21591 23435
rect 21591 23401 21600 23435
rect 21548 23392 21600 23401
rect 24952 23392 25004 23444
rect 10784 23367 10836 23376
rect 10784 23333 10793 23367
rect 10793 23333 10827 23367
rect 10827 23333 10836 23367
rect 10784 23324 10836 23333
rect 10876 23324 10928 23376
rect 16488 23324 16540 23376
rect 11428 23188 11480 23240
rect 16028 23256 16080 23308
rect 18052 23256 18104 23308
rect 18420 23324 18472 23376
rect 19064 23256 19116 23308
rect 22284 23256 22336 23308
rect 23296 23256 23348 23308
rect 23664 23256 23716 23308
rect 25320 23367 25372 23376
rect 25320 23333 25329 23367
rect 25329 23333 25363 23367
rect 25363 23333 25372 23367
rect 25320 23324 25372 23333
rect 13360 23188 13412 23240
rect 13820 23188 13872 23240
rect 14832 23188 14884 23240
rect 17224 23231 17276 23240
rect 17224 23197 17233 23231
rect 17233 23197 17267 23231
rect 17267 23197 17276 23231
rect 17224 23188 17276 23197
rect 22928 23231 22980 23240
rect 22928 23197 22937 23231
rect 22937 23197 22971 23231
rect 22971 23197 22980 23231
rect 22928 23188 22980 23197
rect 23572 23231 23624 23240
rect 23572 23197 23581 23231
rect 23581 23197 23615 23231
rect 23615 23197 23624 23231
rect 23572 23188 23624 23197
rect 23848 23231 23900 23240
rect 23848 23197 23857 23231
rect 23857 23197 23891 23231
rect 23891 23197 23900 23231
rect 23848 23188 23900 23197
rect 24860 23188 24912 23240
rect 10315 23086 10367 23138
rect 10379 23086 10431 23138
rect 10443 23086 10495 23138
rect 10507 23086 10559 23138
rect 19648 23086 19700 23138
rect 19712 23086 19764 23138
rect 19776 23086 19828 23138
rect 19840 23086 19892 23138
rect 8944 22984 8996 23036
rect 11060 22984 11112 23036
rect 11888 22984 11940 23036
rect 14740 23027 14792 23036
rect 14740 22993 14749 23027
rect 14749 22993 14783 23027
rect 14783 22993 14792 23027
rect 14740 22984 14792 22993
rect 16212 22984 16264 23036
rect 18604 22984 18656 23036
rect 19156 23027 19208 23036
rect 19156 22993 19165 23027
rect 19165 22993 19199 23027
rect 19199 22993 19208 23027
rect 19156 22984 19208 22993
rect 19432 23027 19484 23036
rect 19432 22993 19441 23027
rect 19441 22993 19475 23027
rect 19475 22993 19484 23027
rect 19432 22984 19484 22993
rect 9956 22916 10008 22968
rect 10968 22916 11020 22968
rect 13452 22916 13504 22968
rect 14188 22916 14240 22968
rect 18788 22916 18840 22968
rect 19248 22916 19300 22968
rect 11152 22891 11204 22900
rect 11152 22857 11161 22891
rect 11161 22857 11195 22891
rect 11195 22857 11204 22891
rect 11152 22848 11204 22857
rect 18512 22891 18564 22900
rect 18512 22857 18521 22891
rect 18521 22857 18555 22891
rect 18555 22857 18564 22891
rect 18512 22848 18564 22857
rect 19064 22848 19116 22900
rect 20628 22848 20680 22900
rect 21088 22848 21140 22900
rect 23756 22848 23808 22900
rect 24952 22891 25004 22900
rect 24952 22857 24961 22891
rect 24961 22857 24995 22891
rect 24995 22857 25004 22891
rect 24952 22848 25004 22857
rect 9312 22780 9364 22832
rect 11428 22823 11480 22832
rect 11428 22789 11437 22823
rect 11437 22789 11471 22823
rect 11471 22789 11480 22823
rect 11428 22780 11480 22789
rect 13360 22823 13412 22832
rect 13360 22789 13369 22823
rect 13369 22789 13403 22823
rect 13403 22789 13412 22823
rect 13360 22780 13412 22789
rect 15476 22780 15528 22832
rect 9220 22755 9272 22764
rect 9220 22721 9229 22755
rect 9229 22721 9263 22755
rect 9263 22721 9272 22755
rect 9220 22712 9272 22721
rect 17224 22712 17276 22764
rect 18420 22712 18472 22764
rect 24032 22780 24084 22832
rect 15568 22687 15620 22696
rect 15568 22653 15577 22687
rect 15577 22653 15611 22687
rect 15611 22653 15620 22687
rect 15568 22644 15620 22653
rect 16120 22687 16172 22696
rect 16120 22653 16129 22687
rect 16129 22653 16163 22687
rect 16163 22653 16172 22687
rect 16120 22644 16172 22653
rect 20720 22644 20772 22696
rect 23388 22644 23440 22696
rect 23572 22644 23624 22696
rect 25136 22687 25188 22696
rect 25136 22653 25145 22687
rect 25145 22653 25179 22687
rect 25179 22653 25188 22687
rect 25136 22644 25188 22653
rect 5648 22542 5700 22594
rect 5712 22542 5764 22594
rect 5776 22542 5828 22594
rect 5840 22542 5892 22594
rect 14982 22542 15034 22594
rect 15046 22542 15098 22594
rect 15110 22542 15162 22594
rect 15174 22542 15226 22594
rect 24315 22542 24367 22594
rect 24379 22542 24431 22594
rect 24443 22542 24495 22594
rect 24507 22542 24559 22594
rect 8944 22483 8996 22492
rect 8944 22449 8953 22483
rect 8953 22449 8987 22483
rect 8987 22449 8996 22483
rect 8944 22440 8996 22449
rect 9956 22483 10008 22492
rect 9956 22449 9965 22483
rect 9965 22449 9999 22483
rect 9999 22449 10008 22483
rect 9956 22440 10008 22449
rect 11060 22440 11112 22492
rect 13360 22483 13412 22492
rect 13360 22449 13369 22483
rect 13369 22449 13403 22483
rect 13403 22449 13412 22483
rect 13360 22440 13412 22449
rect 14740 22440 14792 22492
rect 15476 22483 15528 22492
rect 10784 22347 10836 22356
rect 10784 22313 10793 22347
rect 10793 22313 10827 22347
rect 10827 22313 10836 22347
rect 10784 22304 10836 22313
rect 13820 22304 13872 22356
rect 14096 22347 14148 22356
rect 14096 22313 14105 22347
rect 14105 22313 14139 22347
rect 14139 22313 14148 22347
rect 15476 22449 15485 22483
rect 15485 22449 15519 22483
rect 15519 22449 15528 22483
rect 15476 22440 15528 22449
rect 16212 22440 16264 22492
rect 18420 22483 18472 22492
rect 18420 22449 18429 22483
rect 18429 22449 18463 22483
rect 18463 22449 18472 22483
rect 18420 22440 18472 22449
rect 20628 22483 20680 22492
rect 20628 22449 20637 22483
rect 20637 22449 20671 22483
rect 20671 22449 20680 22483
rect 20628 22440 20680 22449
rect 21088 22483 21140 22492
rect 21088 22449 21097 22483
rect 21097 22449 21131 22483
rect 21131 22449 21140 22483
rect 21088 22440 21140 22449
rect 23664 22483 23716 22492
rect 23664 22449 23673 22483
rect 23673 22449 23707 22483
rect 23707 22449 23716 22483
rect 23664 22440 23716 22449
rect 24952 22440 25004 22492
rect 25504 22483 25556 22492
rect 25504 22449 25513 22483
rect 25513 22449 25547 22483
rect 25547 22449 25556 22483
rect 25504 22440 25556 22449
rect 18512 22372 18564 22424
rect 23756 22372 23808 22424
rect 14096 22304 14148 22313
rect 16028 22347 16080 22356
rect 16028 22313 16037 22347
rect 16037 22313 16071 22347
rect 16071 22313 16080 22347
rect 19800 22347 19852 22356
rect 16028 22304 16080 22313
rect 19800 22313 19809 22347
rect 19809 22313 19843 22347
rect 19843 22313 19852 22347
rect 19800 22304 19852 22313
rect 22928 22304 22980 22356
rect 11428 22236 11480 22288
rect 15568 22236 15620 22288
rect 15844 22279 15896 22288
rect 15844 22245 15853 22279
rect 15853 22245 15887 22279
rect 15887 22245 15896 22279
rect 15844 22236 15896 22245
rect 9220 22143 9272 22152
rect 9220 22109 9229 22143
rect 9229 22109 9263 22143
rect 9263 22109 9272 22143
rect 9220 22100 9272 22109
rect 11152 22100 11204 22152
rect 16488 22236 16540 22288
rect 18052 22236 18104 22288
rect 19340 22236 19392 22288
rect 17224 22168 17276 22220
rect 22008 22168 22060 22220
rect 22192 22211 22244 22220
rect 22192 22177 22201 22211
rect 22201 22177 22235 22211
rect 22235 22177 22244 22211
rect 22192 22168 22244 22177
rect 24584 22279 24636 22288
rect 24584 22245 24593 22279
rect 24593 22245 24627 22279
rect 24627 22245 24636 22279
rect 24584 22236 24636 22245
rect 13084 22143 13136 22152
rect 13084 22109 13093 22143
rect 13093 22109 13127 22143
rect 13127 22109 13136 22143
rect 13084 22100 13136 22109
rect 13544 22143 13596 22152
rect 13544 22109 13553 22143
rect 13553 22109 13587 22143
rect 13587 22109 13596 22143
rect 13544 22100 13596 22109
rect 21088 22100 21140 22152
rect 22376 22100 22428 22152
rect 23296 22143 23348 22152
rect 23296 22109 23305 22143
rect 23305 22109 23339 22143
rect 23339 22109 23348 22143
rect 23296 22100 23348 22109
rect 24768 22143 24820 22152
rect 24768 22109 24777 22143
rect 24777 22109 24811 22143
rect 24811 22109 24820 22143
rect 24768 22100 24820 22109
rect 10315 21998 10367 22050
rect 10379 21998 10431 22050
rect 10443 21998 10495 22050
rect 10507 21998 10559 22050
rect 19648 21998 19700 22050
rect 19712 21998 19764 22050
rect 19776 21998 19828 22050
rect 19840 21998 19892 22050
rect 10784 21939 10836 21948
rect 10784 21905 10793 21939
rect 10793 21905 10827 21939
rect 10827 21905 10836 21939
rect 10784 21896 10836 21905
rect 11428 21896 11480 21948
rect 13084 21896 13136 21948
rect 13820 21896 13872 21948
rect 15476 21896 15528 21948
rect 16028 21896 16080 21948
rect 18788 21939 18840 21948
rect 18788 21905 18797 21939
rect 18797 21905 18831 21939
rect 18831 21905 18840 21939
rect 18788 21896 18840 21905
rect 19340 21896 19392 21948
rect 22008 21896 22060 21948
rect 13452 21871 13504 21880
rect 13452 21837 13461 21871
rect 13461 21837 13495 21871
rect 13495 21837 13504 21871
rect 13452 21828 13504 21837
rect 14096 21871 14148 21880
rect 14096 21837 14105 21871
rect 14105 21837 14139 21871
rect 14139 21837 14148 21871
rect 14096 21828 14148 21837
rect 22376 21828 22428 21880
rect 15568 21760 15620 21812
rect 15752 21803 15804 21812
rect 15752 21769 15786 21803
rect 15786 21769 15804 21803
rect 15752 21760 15804 21769
rect 18052 21803 18104 21812
rect 18052 21769 18061 21803
rect 18061 21769 18095 21803
rect 18095 21769 18104 21803
rect 18052 21760 18104 21769
rect 18328 21803 18380 21812
rect 18328 21769 18337 21803
rect 18337 21769 18371 21803
rect 18371 21769 18380 21803
rect 18328 21760 18380 21769
rect 24676 21760 24728 21812
rect 24124 21692 24176 21744
rect 24216 21692 24268 21744
rect 19248 21667 19300 21676
rect 19248 21633 19257 21667
rect 19257 21633 19291 21667
rect 19291 21633 19300 21667
rect 19248 21624 19300 21633
rect 23848 21556 23900 21608
rect 24768 21599 24820 21608
rect 24768 21565 24777 21599
rect 24777 21565 24811 21599
rect 24811 21565 24820 21599
rect 24768 21556 24820 21565
rect 5648 21454 5700 21506
rect 5712 21454 5764 21506
rect 5776 21454 5828 21506
rect 5840 21454 5892 21506
rect 14982 21454 15034 21506
rect 15046 21454 15098 21506
rect 15110 21454 15162 21506
rect 15174 21454 15226 21506
rect 24315 21454 24367 21506
rect 24379 21454 24431 21506
rect 24443 21454 24495 21506
rect 24507 21454 24559 21506
rect 10784 21352 10836 21404
rect 22284 21395 22336 21404
rect 22284 21361 22293 21395
rect 22293 21361 22327 21395
rect 22327 21361 22336 21395
rect 22284 21352 22336 21361
rect 23756 21352 23808 21404
rect 24124 21352 24176 21404
rect 18052 21284 18104 21336
rect 24768 21284 24820 21336
rect 14188 21259 14240 21268
rect 14188 21225 14197 21259
rect 14197 21225 14231 21259
rect 14231 21225 14240 21259
rect 14188 21216 14240 21225
rect 15752 21216 15804 21268
rect 17684 21216 17736 21268
rect 19248 21216 19300 21268
rect 23756 21216 23808 21268
rect 14004 21148 14056 21200
rect 10692 21123 10744 21132
rect 10692 21089 10726 21123
rect 10726 21089 10744 21123
rect 10692 21080 10744 21089
rect 19156 21148 19208 21200
rect 20812 21148 20864 21200
rect 22100 21148 22152 21200
rect 24952 21191 25004 21200
rect 24952 21157 24961 21191
rect 24961 21157 24995 21191
rect 24995 21157 25004 21191
rect 24952 21148 25004 21157
rect 18696 21123 18748 21132
rect 18696 21089 18705 21123
rect 18705 21089 18739 21123
rect 18739 21089 18748 21123
rect 18696 21080 18748 21089
rect 21180 21123 21232 21132
rect 21180 21089 21214 21123
rect 21214 21089 21232 21123
rect 21180 21080 21232 21089
rect 11796 21055 11848 21064
rect 11796 21021 11805 21055
rect 11805 21021 11839 21055
rect 11839 21021 11848 21055
rect 11796 21012 11848 21021
rect 13176 21012 13228 21064
rect 15568 21055 15620 21064
rect 15568 21021 15577 21055
rect 15577 21021 15611 21055
rect 15611 21021 15620 21055
rect 15568 21012 15620 21021
rect 16856 21012 16908 21064
rect 17132 21055 17184 21064
rect 17132 21021 17141 21055
rect 17141 21021 17175 21055
rect 17175 21021 17184 21055
rect 17132 21012 17184 21021
rect 18328 21055 18380 21064
rect 18328 21021 18337 21055
rect 18337 21021 18371 21055
rect 18371 21021 18380 21055
rect 18328 21012 18380 21021
rect 18880 21055 18932 21064
rect 18880 21021 18889 21055
rect 18889 21021 18923 21055
rect 18923 21021 18932 21055
rect 18880 21012 18932 21021
rect 19156 21012 19208 21064
rect 20720 21055 20772 21064
rect 20720 21021 20729 21055
rect 20729 21021 20763 21055
rect 20763 21021 20772 21055
rect 20720 21012 20772 21021
rect 23204 21055 23256 21064
rect 23204 21021 23213 21055
rect 23213 21021 23247 21055
rect 23247 21021 23256 21055
rect 23204 21012 23256 21021
rect 23480 21012 23532 21064
rect 23848 21055 23900 21064
rect 23848 21021 23857 21055
rect 23857 21021 23891 21055
rect 23891 21021 23900 21055
rect 23848 21012 23900 21021
rect 25136 21055 25188 21064
rect 25136 21021 25145 21055
rect 25145 21021 25179 21055
rect 25179 21021 25188 21055
rect 25136 21012 25188 21021
rect 10315 20910 10367 20962
rect 10379 20910 10431 20962
rect 10443 20910 10495 20962
rect 10507 20910 10559 20962
rect 19648 20910 19700 20962
rect 19712 20910 19764 20962
rect 19776 20910 19828 20962
rect 19840 20910 19892 20962
rect 10692 20808 10744 20860
rect 12900 20808 12952 20860
rect 14004 20851 14056 20860
rect 14004 20817 14013 20851
rect 14013 20817 14047 20851
rect 14047 20817 14056 20851
rect 14004 20808 14056 20817
rect 17132 20808 17184 20860
rect 18052 20808 18104 20860
rect 18880 20851 18932 20860
rect 18880 20817 18889 20851
rect 18889 20817 18923 20851
rect 18923 20817 18932 20851
rect 18880 20808 18932 20817
rect 19340 20808 19392 20860
rect 19432 20808 19484 20860
rect 22008 20851 22060 20860
rect 22008 20817 22017 20851
rect 22017 20817 22051 20851
rect 22051 20817 22060 20851
rect 22008 20808 22060 20817
rect 22192 20808 22244 20860
rect 10968 20740 11020 20792
rect 11244 20783 11296 20792
rect 11244 20749 11253 20783
rect 11253 20749 11287 20783
rect 11287 20749 11296 20783
rect 11244 20740 11296 20749
rect 19248 20783 19300 20792
rect 19248 20749 19282 20783
rect 19282 20749 19300 20783
rect 19248 20740 19300 20749
rect 21180 20740 21232 20792
rect 23756 20740 23808 20792
rect 24124 20740 24176 20792
rect 11152 20715 11204 20724
rect 11152 20681 11161 20715
rect 11161 20681 11195 20715
rect 11195 20681 11204 20715
rect 11152 20672 11204 20681
rect 13176 20672 13228 20724
rect 14372 20715 14424 20724
rect 14372 20681 14381 20715
rect 14381 20681 14415 20715
rect 14415 20681 14424 20715
rect 14372 20672 14424 20681
rect 16396 20672 16448 20724
rect 11796 20604 11848 20656
rect 12900 20647 12952 20656
rect 12900 20613 12909 20647
rect 12909 20613 12943 20647
rect 12943 20613 12952 20647
rect 12900 20604 12952 20613
rect 12992 20647 13044 20656
rect 12992 20613 13001 20647
rect 13001 20613 13035 20647
rect 13035 20613 13044 20647
rect 14464 20647 14516 20656
rect 12992 20604 13044 20613
rect 14464 20613 14473 20647
rect 14473 20613 14507 20647
rect 14507 20613 14516 20647
rect 14464 20604 14516 20613
rect 14648 20647 14700 20656
rect 14648 20613 14657 20647
rect 14657 20613 14691 20647
rect 14691 20613 14700 20647
rect 14648 20604 14700 20613
rect 16120 20604 16172 20656
rect 16488 20536 16540 20588
rect 18696 20604 18748 20656
rect 20720 20672 20772 20724
rect 22468 20715 22520 20724
rect 22468 20681 22477 20715
rect 22477 20681 22511 20715
rect 22511 20681 22520 20715
rect 22468 20672 22520 20681
rect 23664 20647 23716 20656
rect 23664 20613 23673 20647
rect 23673 20613 23707 20647
rect 23707 20613 23716 20647
rect 23664 20604 23716 20613
rect 13728 20511 13780 20520
rect 13728 20477 13737 20511
rect 13737 20477 13771 20511
rect 13771 20477 13780 20511
rect 13728 20468 13780 20477
rect 22652 20468 22704 20520
rect 5648 20366 5700 20418
rect 5712 20366 5764 20418
rect 5776 20366 5828 20418
rect 5840 20366 5892 20418
rect 14982 20366 15034 20418
rect 15046 20366 15098 20418
rect 15110 20366 15162 20418
rect 15174 20366 15226 20418
rect 24315 20366 24367 20418
rect 24379 20366 24431 20418
rect 24443 20366 24495 20418
rect 24507 20366 24559 20418
rect 10968 20264 11020 20316
rect 12992 20264 13044 20316
rect 13176 20307 13228 20316
rect 13176 20273 13185 20307
rect 13185 20273 13219 20307
rect 13219 20273 13228 20307
rect 13176 20264 13228 20273
rect 14372 20264 14424 20316
rect 12900 20196 12952 20248
rect 10784 20128 10836 20180
rect 11244 20171 11296 20180
rect 11244 20137 11253 20171
rect 11253 20137 11287 20171
rect 11287 20137 11296 20171
rect 11244 20128 11296 20137
rect 14648 20264 14700 20316
rect 16120 20307 16172 20316
rect 16120 20273 16129 20307
rect 16129 20273 16163 20307
rect 16163 20273 16172 20307
rect 16120 20264 16172 20273
rect 17684 20307 17736 20316
rect 17684 20273 17693 20307
rect 17693 20273 17727 20307
rect 17727 20273 17736 20307
rect 17684 20264 17736 20273
rect 20628 20264 20680 20316
rect 22376 20264 22428 20316
rect 23756 20307 23808 20316
rect 23756 20273 23765 20307
rect 23765 20273 23799 20307
rect 23799 20273 23808 20307
rect 23756 20264 23808 20273
rect 24124 20264 24176 20316
rect 19340 20128 19392 20180
rect 19524 20171 19576 20180
rect 19524 20137 19533 20171
rect 19533 20137 19567 20171
rect 19567 20137 19576 20171
rect 19524 20128 19576 20137
rect 22100 20128 22152 20180
rect 22376 20171 22428 20180
rect 22376 20137 22385 20171
rect 22385 20137 22419 20171
rect 22419 20137 22428 20171
rect 22376 20128 22428 20137
rect 23756 20128 23808 20180
rect 26148 20128 26200 20180
rect 11796 20060 11848 20112
rect 13728 20103 13780 20112
rect 13728 20069 13737 20103
rect 13737 20069 13771 20103
rect 13771 20069 13780 20103
rect 13728 20060 13780 20069
rect 14004 20035 14056 20044
rect 14004 20001 14013 20035
rect 14013 20001 14047 20035
rect 14047 20001 14056 20035
rect 14004 19992 14056 20001
rect 10692 19924 10744 19976
rect 14740 19924 14792 19976
rect 15568 19924 15620 19976
rect 22652 20103 22704 20112
rect 22652 20069 22686 20103
rect 22686 20069 22704 20103
rect 22652 20060 22704 20069
rect 24860 20103 24912 20112
rect 24860 20069 24869 20103
rect 24869 20069 24903 20103
rect 24903 20069 24912 20103
rect 24860 20060 24912 20069
rect 16488 19992 16540 20044
rect 18512 20035 18564 20044
rect 18512 20001 18521 20035
rect 18521 20001 18555 20035
rect 18555 20001 18564 20035
rect 18512 19992 18564 20001
rect 22376 19992 22428 20044
rect 23664 19992 23716 20044
rect 18052 19924 18104 19976
rect 18696 19924 18748 19976
rect 18972 19967 19024 19976
rect 18972 19933 18981 19967
rect 18981 19933 19015 19967
rect 19015 19933 19024 19967
rect 18972 19924 19024 19933
rect 21640 19967 21692 19976
rect 21640 19933 21649 19967
rect 21649 19933 21683 19967
rect 21683 19933 21692 19967
rect 21640 19924 21692 19933
rect 22192 19924 22244 19976
rect 25044 19967 25096 19976
rect 25044 19933 25053 19967
rect 25053 19933 25087 19967
rect 25087 19933 25096 19967
rect 25044 19924 25096 19933
rect 10315 19822 10367 19874
rect 10379 19822 10431 19874
rect 10443 19822 10495 19874
rect 10507 19822 10559 19874
rect 19648 19822 19700 19874
rect 19712 19822 19764 19874
rect 19776 19822 19828 19874
rect 19840 19822 19892 19874
rect 11796 19720 11848 19772
rect 12348 19720 12400 19772
rect 12992 19720 13044 19772
rect 13360 19763 13412 19772
rect 13360 19729 13369 19763
rect 13369 19729 13403 19763
rect 13403 19729 13412 19763
rect 13360 19720 13412 19729
rect 11244 19695 11296 19704
rect 11244 19661 11253 19695
rect 11253 19661 11287 19695
rect 11287 19661 11296 19695
rect 11244 19652 11296 19661
rect 13544 19652 13596 19704
rect 13728 19516 13780 19568
rect 14464 19720 14516 19772
rect 16488 19720 16540 19772
rect 18512 19763 18564 19772
rect 18512 19729 18521 19763
rect 18521 19729 18555 19763
rect 18555 19729 18564 19763
rect 18512 19720 18564 19729
rect 22376 19763 22428 19772
rect 22376 19729 22385 19763
rect 22385 19729 22419 19763
rect 22419 19729 22428 19763
rect 22376 19720 22428 19729
rect 23204 19720 23256 19772
rect 25320 19763 25372 19772
rect 25320 19729 25329 19763
rect 25329 19729 25363 19763
rect 25363 19729 25372 19763
rect 25320 19720 25372 19729
rect 14648 19652 14700 19704
rect 15476 19652 15528 19704
rect 22652 19652 22704 19704
rect 18972 19584 19024 19636
rect 19524 19627 19576 19636
rect 19524 19593 19533 19627
rect 19533 19593 19567 19627
rect 19567 19593 19576 19627
rect 19524 19584 19576 19593
rect 19800 19627 19852 19636
rect 19800 19593 19809 19627
rect 19809 19593 19843 19627
rect 19843 19593 19852 19627
rect 19800 19584 19852 19593
rect 23480 19584 23532 19636
rect 23848 19627 23900 19636
rect 23848 19593 23857 19627
rect 23857 19593 23891 19627
rect 23891 19593 23900 19627
rect 23848 19584 23900 19593
rect 24860 19584 24912 19636
rect 14740 19516 14792 19568
rect 24124 19559 24176 19568
rect 24124 19525 24133 19559
rect 24133 19525 24167 19559
rect 24167 19525 24176 19559
rect 24124 19516 24176 19525
rect 16396 19380 16448 19432
rect 17040 19423 17092 19432
rect 17040 19389 17049 19423
rect 17049 19389 17083 19423
rect 17083 19389 17092 19423
rect 17040 19380 17092 19389
rect 19340 19423 19392 19432
rect 19340 19389 19349 19423
rect 19349 19389 19383 19423
rect 19383 19389 19392 19423
rect 19340 19380 19392 19389
rect 5648 19278 5700 19330
rect 5712 19278 5764 19330
rect 5776 19278 5828 19330
rect 5840 19278 5892 19330
rect 14982 19278 15034 19330
rect 15046 19278 15098 19330
rect 15110 19278 15162 19330
rect 15174 19278 15226 19330
rect 24315 19278 24367 19330
rect 24379 19278 24431 19330
rect 24443 19278 24495 19330
rect 24507 19278 24559 19330
rect 11244 19176 11296 19228
rect 15476 19219 15528 19228
rect 15476 19185 15485 19219
rect 15485 19185 15519 19219
rect 15519 19185 15528 19219
rect 15476 19176 15528 19185
rect 19524 19176 19576 19228
rect 23848 19219 23900 19228
rect 23848 19185 23857 19219
rect 23857 19185 23891 19219
rect 23891 19185 23900 19219
rect 23848 19176 23900 19185
rect 24860 19176 24912 19228
rect 12072 19083 12124 19092
rect 12072 19049 12081 19083
rect 12081 19049 12115 19083
rect 12115 19049 12124 19083
rect 12072 19040 12124 19049
rect 12348 19015 12400 19024
rect 12348 18981 12382 19015
rect 12382 18981 12400 19015
rect 12348 18972 12400 18981
rect 16856 19015 16908 19024
rect 16856 18981 16865 19015
rect 16865 18981 16899 19015
rect 16899 18981 16908 19015
rect 16856 18972 16908 18981
rect 19524 18972 19576 19024
rect 22008 18972 22060 19024
rect 13728 18836 13780 18888
rect 14740 18836 14792 18888
rect 19064 18879 19116 18888
rect 19064 18845 19073 18879
rect 19073 18845 19107 18879
rect 19107 18845 19116 18879
rect 19064 18836 19116 18845
rect 19248 18879 19300 18888
rect 19248 18845 19257 18879
rect 19257 18845 19291 18879
rect 19291 18845 19300 18879
rect 19248 18836 19300 18845
rect 19340 18836 19392 18888
rect 20628 18836 20680 18888
rect 21916 18879 21968 18888
rect 21916 18845 21925 18879
rect 21925 18845 21959 18879
rect 21959 18845 21968 18879
rect 22284 18947 22336 18956
rect 22284 18913 22293 18947
rect 22293 18913 22327 18947
rect 22327 18913 22336 18947
rect 22284 18904 22336 18913
rect 22376 18879 22428 18888
rect 21916 18836 21968 18845
rect 22376 18845 22385 18879
rect 22385 18845 22419 18879
rect 22419 18845 22428 18879
rect 22376 18836 22428 18845
rect 24124 18972 24176 19024
rect 23388 18836 23440 18888
rect 24768 18879 24820 18888
rect 24768 18845 24777 18879
rect 24777 18845 24811 18879
rect 24811 18845 24820 18879
rect 24768 18836 24820 18845
rect 10315 18734 10367 18786
rect 10379 18734 10431 18786
rect 10443 18734 10495 18786
rect 10507 18734 10559 18786
rect 19648 18734 19700 18786
rect 19712 18734 19764 18786
rect 19776 18734 19828 18786
rect 19840 18734 19892 18786
rect 12348 18632 12400 18684
rect 13360 18632 13412 18684
rect 15476 18632 15528 18684
rect 24032 18632 24084 18684
rect 21548 18564 21600 18616
rect 24124 18564 24176 18616
rect 12072 18496 12124 18548
rect 13360 18539 13412 18548
rect 13360 18505 13369 18539
rect 13369 18505 13403 18539
rect 13403 18505 13412 18539
rect 13360 18496 13412 18505
rect 13544 18496 13596 18548
rect 13728 18539 13780 18548
rect 13728 18505 13762 18539
rect 13762 18505 13780 18539
rect 13728 18496 13780 18505
rect 13268 18428 13320 18480
rect 15936 18335 15988 18344
rect 15936 18301 15945 18335
rect 15945 18301 15979 18335
rect 15979 18301 15988 18335
rect 15936 18292 15988 18301
rect 17316 18292 17368 18344
rect 21180 18496 21232 18548
rect 24032 18539 24084 18548
rect 24032 18505 24041 18539
rect 24041 18505 24075 18539
rect 24075 18505 24084 18539
rect 24032 18496 24084 18505
rect 25228 18539 25280 18548
rect 18052 18471 18104 18480
rect 18052 18437 18061 18471
rect 18061 18437 18095 18471
rect 18095 18437 18104 18471
rect 18052 18428 18104 18437
rect 22376 18428 22428 18480
rect 23480 18428 23532 18480
rect 25228 18505 25237 18539
rect 25237 18505 25271 18539
rect 25271 18505 25280 18539
rect 25228 18496 25280 18505
rect 25412 18403 25464 18412
rect 25412 18369 25421 18403
rect 25421 18369 25455 18403
rect 25455 18369 25464 18403
rect 25412 18360 25464 18369
rect 19248 18292 19300 18344
rect 22008 18292 22060 18344
rect 22468 18335 22520 18344
rect 22468 18301 22477 18335
rect 22477 18301 22511 18335
rect 22511 18301 22520 18335
rect 22468 18292 22520 18301
rect 23664 18335 23716 18344
rect 23664 18301 23673 18335
rect 23673 18301 23707 18335
rect 23707 18301 23716 18335
rect 23664 18292 23716 18301
rect 5648 18190 5700 18242
rect 5712 18190 5764 18242
rect 5776 18190 5828 18242
rect 5840 18190 5892 18242
rect 14982 18190 15034 18242
rect 15046 18190 15098 18242
rect 15110 18190 15162 18242
rect 15174 18190 15226 18242
rect 24315 18190 24367 18242
rect 24379 18190 24431 18242
rect 24443 18190 24495 18242
rect 24507 18190 24559 18242
rect 13728 18088 13780 18140
rect 19524 18088 19576 18140
rect 24124 18088 24176 18140
rect 20720 18020 20772 18072
rect 21180 18020 21232 18072
rect 21548 17995 21600 18004
rect 21548 17961 21557 17995
rect 21557 17961 21591 17995
rect 21591 17961 21600 17995
rect 21548 17952 21600 17961
rect 14740 17816 14792 17868
rect 15936 17884 15988 17936
rect 16396 17884 16448 17936
rect 21364 17927 21416 17936
rect 18052 17816 18104 17868
rect 21364 17893 21373 17927
rect 21373 17893 21407 17927
rect 21407 17893 21416 17927
rect 21364 17884 21416 17893
rect 22468 17884 22520 17936
rect 23112 17884 23164 17936
rect 19248 17816 19300 17868
rect 20996 17816 21048 17868
rect 24860 17816 24912 17868
rect 25228 17816 25280 17868
rect 13268 17748 13320 17800
rect 13728 17748 13780 17800
rect 14280 17791 14332 17800
rect 14280 17757 14289 17791
rect 14289 17757 14323 17791
rect 14323 17757 14332 17791
rect 14280 17748 14332 17757
rect 17316 17748 17368 17800
rect 20904 17791 20956 17800
rect 20904 17757 20913 17791
rect 20913 17757 20947 17791
rect 20947 17757 20956 17791
rect 20904 17748 20956 17757
rect 10315 17646 10367 17698
rect 10379 17646 10431 17698
rect 10443 17646 10495 17698
rect 10507 17646 10559 17698
rect 19648 17646 19700 17698
rect 19712 17646 19764 17698
rect 19776 17646 19828 17698
rect 19840 17646 19892 17698
rect 19156 17544 19208 17596
rect 21548 17587 21600 17596
rect 21548 17553 21557 17587
rect 21557 17553 21591 17587
rect 21591 17553 21600 17587
rect 21548 17544 21600 17553
rect 23112 17587 23164 17596
rect 23112 17553 23121 17587
rect 23121 17553 23155 17587
rect 23155 17553 23164 17587
rect 23112 17544 23164 17553
rect 23480 17587 23532 17596
rect 23480 17553 23489 17587
rect 23489 17553 23523 17587
rect 23523 17553 23532 17587
rect 23480 17544 23532 17553
rect 24032 17544 24084 17596
rect 25596 17587 25648 17596
rect 25596 17553 25605 17587
rect 25605 17553 25639 17587
rect 25639 17553 25648 17587
rect 25596 17544 25648 17553
rect 15292 17476 15344 17528
rect 15752 17476 15804 17528
rect 19524 17476 19576 17528
rect 20536 17476 20588 17528
rect 20628 17476 20680 17528
rect 24768 17476 24820 17528
rect 14280 17408 14332 17460
rect 15108 17408 15160 17460
rect 15844 17408 15896 17460
rect 16212 17451 16264 17460
rect 16212 17417 16221 17451
rect 16221 17417 16255 17451
rect 16255 17417 16264 17451
rect 16212 17408 16264 17417
rect 17040 17408 17092 17460
rect 18788 17408 18840 17460
rect 19248 17408 19300 17460
rect 20168 17451 20220 17460
rect 20168 17417 20177 17451
rect 20177 17417 20211 17451
rect 20211 17417 20220 17451
rect 20168 17408 20220 17417
rect 23664 17408 23716 17460
rect 24124 17451 24176 17460
rect 24124 17417 24133 17451
rect 24133 17417 24167 17451
rect 24167 17417 24176 17451
rect 24124 17408 24176 17417
rect 25412 17451 25464 17460
rect 25412 17417 25421 17451
rect 25421 17417 25455 17451
rect 25455 17417 25464 17451
rect 25412 17408 25464 17417
rect 26332 17408 26384 17460
rect 14556 17383 14608 17392
rect 14556 17349 14565 17383
rect 14565 17349 14599 17383
rect 14599 17349 14608 17383
rect 14556 17340 14608 17349
rect 14740 17383 14792 17392
rect 14740 17349 14749 17383
rect 14749 17349 14783 17383
rect 14783 17349 14792 17383
rect 14740 17340 14792 17349
rect 16396 17383 16448 17392
rect 16396 17349 16405 17383
rect 16405 17349 16439 17383
rect 16439 17349 16448 17383
rect 16396 17340 16448 17349
rect 14096 17315 14148 17324
rect 14096 17281 14105 17315
rect 14105 17281 14139 17315
rect 14139 17281 14148 17315
rect 14096 17272 14148 17281
rect 12164 17247 12216 17256
rect 12164 17213 12173 17247
rect 12173 17213 12207 17247
rect 12207 17213 12216 17247
rect 12164 17204 12216 17213
rect 14188 17204 14240 17256
rect 17776 17247 17828 17256
rect 17776 17213 17785 17247
rect 17785 17213 17819 17247
rect 17819 17213 17828 17247
rect 17776 17204 17828 17213
rect 18512 17204 18564 17256
rect 5648 17102 5700 17154
rect 5712 17102 5764 17154
rect 5776 17102 5828 17154
rect 5840 17102 5892 17154
rect 14982 17102 15034 17154
rect 15046 17102 15098 17154
rect 15110 17102 15162 17154
rect 15174 17102 15226 17154
rect 24315 17102 24367 17154
rect 24379 17102 24431 17154
rect 24443 17102 24495 17154
rect 24507 17102 24559 17154
rect 13544 17000 13596 17052
rect 14556 17000 14608 17052
rect 14740 17043 14792 17052
rect 14740 17009 14749 17043
rect 14749 17009 14783 17043
rect 14783 17009 14792 17043
rect 14740 17000 14792 17009
rect 16396 17000 16448 17052
rect 17316 17043 17368 17052
rect 17316 17009 17325 17043
rect 17325 17009 17359 17043
rect 17359 17009 17368 17043
rect 17316 17000 17368 17009
rect 17776 17000 17828 17052
rect 19156 17043 19208 17052
rect 19156 17009 19165 17043
rect 19165 17009 19199 17043
rect 19199 17009 19208 17043
rect 19156 17000 19208 17009
rect 20168 17043 20220 17052
rect 20168 17009 20177 17043
rect 20177 17009 20211 17043
rect 20211 17009 20220 17043
rect 20168 17000 20220 17009
rect 20536 17043 20588 17052
rect 20536 17009 20545 17043
rect 20545 17009 20579 17043
rect 20579 17009 20588 17043
rect 20536 17000 20588 17009
rect 23848 17043 23900 17052
rect 23848 17009 23857 17043
rect 23857 17009 23891 17043
rect 23891 17009 23900 17043
rect 23848 17000 23900 17009
rect 24124 17000 24176 17052
rect 25504 17043 25556 17052
rect 25504 17009 25513 17043
rect 25513 17009 25547 17043
rect 25547 17009 25556 17043
rect 25504 17000 25556 17009
rect 26332 17043 26384 17052
rect 26332 17009 26341 17043
rect 26341 17009 26375 17043
rect 26375 17009 26384 17043
rect 26332 17000 26384 17009
rect 12164 16864 12216 16916
rect 12624 16907 12676 16916
rect 12624 16873 12633 16907
rect 12633 16873 12667 16907
rect 12667 16873 12676 16907
rect 12624 16864 12676 16873
rect 14188 16907 14240 16916
rect 12256 16796 12308 16848
rect 11888 16771 11940 16780
rect 11888 16737 11897 16771
rect 11897 16737 11931 16771
rect 11931 16737 11940 16771
rect 11888 16728 11940 16737
rect 13360 16796 13412 16848
rect 14188 16873 14197 16907
rect 14197 16873 14231 16907
rect 14231 16873 14240 16907
rect 14188 16864 14240 16873
rect 17592 16975 17644 16984
rect 17592 16941 17601 16975
rect 17601 16941 17635 16975
rect 17635 16941 17644 16975
rect 17592 16932 17644 16941
rect 15108 16864 15160 16916
rect 14004 16839 14056 16848
rect 14004 16805 14013 16839
rect 14013 16805 14047 16839
rect 14047 16805 14056 16839
rect 14004 16796 14056 16805
rect 13728 16660 13780 16712
rect 17040 16796 17092 16848
rect 20996 16864 21048 16916
rect 24032 16932 24084 16984
rect 26240 16932 26292 16984
rect 27528 16932 27580 16984
rect 25412 16864 25464 16916
rect 23848 16796 23900 16848
rect 25320 16839 25372 16848
rect 25320 16805 25329 16839
rect 25329 16805 25363 16839
rect 25363 16805 25372 16839
rect 25320 16796 25372 16805
rect 17868 16728 17920 16780
rect 17776 16703 17828 16712
rect 17776 16669 17785 16703
rect 17785 16669 17819 16703
rect 17819 16669 17828 16703
rect 17776 16660 17828 16669
rect 18788 16703 18840 16712
rect 18788 16669 18797 16703
rect 18797 16669 18831 16703
rect 18831 16669 18840 16703
rect 18788 16660 18840 16669
rect 10315 16558 10367 16610
rect 10379 16558 10431 16610
rect 10443 16558 10495 16610
rect 10507 16558 10559 16610
rect 19648 16558 19700 16610
rect 19712 16558 19764 16610
rect 19776 16558 19828 16610
rect 19840 16558 19892 16610
rect 12256 16456 12308 16508
rect 13544 16499 13596 16508
rect 13544 16465 13553 16499
rect 13553 16465 13587 16499
rect 13587 16465 13596 16499
rect 13544 16456 13596 16465
rect 15108 16499 15160 16508
rect 15108 16465 15117 16499
rect 15117 16465 15151 16499
rect 15151 16465 15160 16499
rect 15108 16456 15160 16465
rect 16212 16499 16264 16508
rect 16212 16465 16221 16499
rect 16221 16465 16255 16499
rect 16255 16465 16264 16499
rect 16212 16456 16264 16465
rect 16396 16456 16448 16508
rect 17868 16499 17920 16508
rect 17868 16465 17877 16499
rect 17877 16465 17911 16499
rect 17911 16465 17920 16499
rect 17868 16456 17920 16465
rect 18052 16499 18104 16508
rect 18052 16465 18061 16499
rect 18061 16465 18095 16499
rect 18095 16465 18104 16499
rect 18052 16456 18104 16465
rect 18512 16499 18564 16508
rect 18512 16465 18521 16499
rect 18521 16465 18555 16499
rect 18555 16465 18564 16499
rect 18512 16456 18564 16465
rect 21824 16456 21876 16508
rect 25412 16499 25464 16508
rect 25412 16465 25421 16499
rect 25421 16465 25455 16499
rect 25455 16465 25464 16499
rect 25412 16456 25464 16465
rect 14188 16388 14240 16440
rect 15844 16431 15896 16440
rect 15844 16397 15853 16431
rect 15853 16397 15887 16431
rect 15887 16397 15896 16431
rect 15844 16388 15896 16397
rect 17684 16388 17736 16440
rect 17776 16388 17828 16440
rect 19064 16388 19116 16440
rect 25320 16388 25372 16440
rect 21640 16320 21692 16372
rect 23848 16320 23900 16372
rect 25228 16363 25280 16372
rect 25228 16329 25237 16363
rect 25237 16329 25271 16363
rect 25271 16329 25280 16363
rect 25228 16320 25280 16329
rect 12440 16252 12492 16304
rect 13728 16295 13780 16304
rect 13728 16261 13737 16295
rect 13737 16261 13771 16295
rect 13771 16261 13780 16295
rect 13728 16252 13780 16261
rect 18604 16252 18656 16304
rect 19248 16252 19300 16304
rect 21916 16295 21968 16304
rect 21916 16261 21925 16295
rect 21925 16261 21959 16295
rect 21959 16261 21968 16295
rect 21916 16252 21968 16261
rect 22376 16116 22428 16168
rect 5648 16014 5700 16066
rect 5712 16014 5764 16066
rect 5776 16014 5828 16066
rect 5840 16014 5892 16066
rect 14982 16014 15034 16066
rect 15046 16014 15098 16066
rect 15110 16014 15162 16066
rect 15174 16014 15226 16066
rect 24315 16014 24367 16066
rect 24379 16014 24431 16066
rect 24443 16014 24495 16066
rect 24507 16014 24559 16066
rect 14188 15912 14240 15964
rect 15292 15955 15344 15964
rect 15292 15921 15301 15955
rect 15301 15921 15335 15955
rect 15335 15921 15344 15955
rect 15292 15912 15344 15921
rect 18512 15912 18564 15964
rect 19064 15955 19116 15964
rect 19064 15921 19073 15955
rect 19073 15921 19107 15955
rect 19107 15921 19116 15955
rect 19064 15912 19116 15921
rect 20720 15912 20772 15964
rect 13728 15844 13780 15896
rect 18604 15844 18656 15896
rect 15844 15819 15896 15828
rect 15844 15785 15853 15819
rect 15853 15785 15887 15819
rect 15887 15785 15896 15819
rect 15844 15776 15896 15785
rect 17132 15819 17184 15828
rect 17132 15785 17141 15819
rect 17141 15785 17175 15819
rect 17175 15785 17184 15819
rect 17132 15776 17184 15785
rect 23848 15912 23900 15964
rect 25228 15955 25280 15964
rect 25228 15921 25237 15955
rect 25237 15921 25271 15955
rect 25271 15921 25280 15955
rect 25228 15912 25280 15921
rect 23756 15844 23808 15896
rect 12440 15708 12492 15760
rect 14832 15708 14884 15760
rect 16304 15708 16356 15760
rect 23572 15776 23624 15828
rect 23848 15776 23900 15828
rect 18236 15708 18288 15760
rect 21916 15708 21968 15760
rect 12624 15640 12676 15692
rect 13820 15640 13872 15692
rect 17684 15683 17736 15692
rect 17684 15649 17693 15683
rect 17693 15649 17727 15683
rect 17727 15649 17736 15683
rect 17684 15640 17736 15649
rect 22376 15640 22428 15692
rect 12440 15615 12492 15624
rect 12440 15581 12449 15615
rect 12449 15581 12483 15615
rect 12483 15581 12492 15615
rect 15660 15615 15712 15624
rect 12440 15572 12492 15581
rect 15660 15581 15669 15615
rect 15669 15581 15703 15615
rect 15703 15581 15712 15615
rect 15660 15572 15712 15581
rect 17316 15615 17368 15624
rect 17316 15581 17325 15615
rect 17325 15581 17359 15615
rect 17359 15581 17368 15615
rect 17316 15572 17368 15581
rect 21640 15572 21692 15624
rect 22928 15572 22980 15624
rect 23480 15572 23532 15624
rect 23756 15572 23808 15624
rect 10315 15470 10367 15522
rect 10379 15470 10431 15522
rect 10443 15470 10495 15522
rect 10507 15470 10559 15522
rect 19648 15470 19700 15522
rect 19712 15470 19764 15522
rect 19776 15470 19828 15522
rect 19840 15470 19892 15522
rect 13820 15411 13872 15420
rect 13820 15377 13829 15411
rect 13829 15377 13863 15411
rect 13863 15377 13872 15411
rect 13820 15368 13872 15377
rect 14188 15368 14240 15420
rect 15660 15368 15712 15420
rect 16396 15411 16448 15420
rect 16396 15377 16405 15411
rect 16405 15377 16439 15411
rect 16439 15377 16448 15411
rect 16396 15368 16448 15377
rect 18236 15411 18288 15420
rect 18236 15377 18245 15411
rect 18245 15377 18279 15411
rect 18279 15377 18288 15411
rect 18236 15368 18288 15377
rect 21916 15368 21968 15420
rect 15844 15300 15896 15352
rect 21272 15300 21324 15352
rect 24124 15411 24176 15420
rect 24124 15377 24133 15411
rect 24133 15377 24167 15411
rect 24167 15377 24176 15411
rect 24124 15368 24176 15377
rect 12716 15275 12768 15284
rect 12716 15241 12750 15275
rect 12750 15241 12768 15275
rect 12716 15232 12768 15241
rect 16396 15232 16448 15284
rect 16856 15275 16908 15284
rect 16856 15241 16865 15275
rect 16865 15241 16899 15275
rect 16899 15241 16908 15275
rect 16856 15232 16908 15241
rect 20168 15232 20220 15284
rect 20812 15232 20864 15284
rect 22008 15275 22060 15284
rect 22008 15241 22017 15275
rect 22017 15241 22051 15275
rect 22051 15241 22060 15275
rect 22008 15232 22060 15241
rect 23480 15232 23532 15284
rect 25136 15232 25188 15284
rect 12440 15207 12492 15216
rect 12440 15173 12449 15207
rect 12449 15173 12483 15207
rect 12483 15173 12492 15207
rect 16948 15207 17000 15216
rect 12440 15164 12492 15173
rect 16948 15173 16957 15207
rect 16957 15173 16991 15207
rect 16991 15173 17000 15207
rect 16948 15164 17000 15173
rect 19156 15207 19208 15216
rect 19156 15173 19165 15207
rect 19165 15173 19199 15207
rect 19199 15173 19208 15207
rect 19156 15164 19208 15173
rect 21180 15028 21232 15080
rect 25412 15207 25464 15216
rect 24032 15096 24084 15148
rect 25412 15173 25421 15207
rect 25421 15173 25455 15207
rect 25455 15173 25464 15207
rect 25412 15164 25464 15173
rect 23664 15071 23716 15080
rect 23664 15037 23673 15071
rect 23673 15037 23707 15071
rect 23707 15037 23716 15071
rect 23664 15028 23716 15037
rect 5648 14926 5700 14978
rect 5712 14926 5764 14978
rect 5776 14926 5828 14978
rect 5840 14926 5892 14978
rect 14982 14926 15034 14978
rect 15046 14926 15098 14978
rect 15110 14926 15162 14978
rect 15174 14926 15226 14978
rect 24315 14926 24367 14978
rect 24379 14926 24431 14978
rect 24443 14926 24495 14978
rect 24507 14926 24559 14978
rect 12716 14824 12768 14876
rect 16948 14824 17000 14876
rect 20720 14867 20772 14876
rect 20720 14833 20729 14867
rect 20729 14833 20763 14867
rect 20763 14833 20772 14867
rect 20720 14824 20772 14833
rect 23388 14867 23440 14876
rect 23388 14833 23397 14867
rect 23397 14833 23431 14867
rect 23431 14833 23440 14867
rect 23388 14824 23440 14833
rect 24124 14824 24176 14876
rect 25320 14824 25372 14876
rect 22928 14799 22980 14808
rect 22928 14765 22937 14799
rect 22937 14765 22971 14799
rect 22971 14765 22980 14799
rect 22928 14756 22980 14765
rect 25136 14756 25188 14808
rect 16028 14595 16080 14604
rect 16028 14561 16062 14595
rect 16062 14561 16080 14595
rect 16028 14552 16080 14561
rect 18328 14620 18380 14672
rect 23664 14620 23716 14672
rect 25044 14663 25096 14672
rect 25044 14629 25053 14663
rect 25053 14629 25087 14663
rect 25087 14629 25096 14663
rect 25044 14620 25096 14629
rect 19156 14552 19208 14604
rect 21180 14552 21232 14604
rect 23480 14552 23532 14604
rect 12440 14527 12492 14536
rect 12440 14493 12449 14527
rect 12449 14493 12483 14527
rect 12483 14493 12492 14527
rect 12440 14484 12492 14493
rect 19340 14484 19392 14536
rect 22376 14527 22428 14536
rect 22376 14493 22385 14527
rect 22385 14493 22419 14527
rect 22419 14493 22428 14527
rect 22376 14484 22428 14493
rect 24032 14484 24084 14536
rect 24308 14527 24360 14536
rect 24308 14493 24317 14527
rect 24317 14493 24351 14527
rect 24351 14493 24360 14527
rect 24308 14484 24360 14493
rect 10315 14382 10367 14434
rect 10379 14382 10431 14434
rect 10443 14382 10495 14434
rect 10507 14382 10559 14434
rect 19648 14382 19700 14434
rect 19712 14382 19764 14434
rect 19776 14382 19828 14434
rect 19840 14382 19892 14434
rect 16396 14323 16448 14332
rect 16396 14289 16405 14323
rect 16405 14289 16439 14323
rect 16439 14289 16448 14323
rect 16396 14280 16448 14289
rect 17316 14280 17368 14332
rect 19156 14323 19208 14332
rect 19156 14289 19165 14323
rect 19165 14289 19199 14323
rect 19199 14289 19208 14323
rect 19156 14280 19208 14289
rect 20168 14280 20220 14332
rect 21088 14280 21140 14332
rect 23388 14280 23440 14332
rect 23664 14280 23716 14332
rect 24032 14280 24084 14332
rect 25044 14323 25096 14332
rect 16856 14212 16908 14264
rect 21272 14212 21324 14264
rect 25044 14289 25053 14323
rect 25053 14289 25087 14323
rect 25087 14289 25096 14323
rect 25044 14280 25096 14289
rect 25504 14323 25556 14332
rect 25504 14289 25513 14323
rect 25513 14289 25547 14323
rect 25547 14289 25556 14323
rect 25504 14280 25556 14289
rect 16120 14144 16172 14196
rect 21364 14187 21416 14196
rect 21364 14153 21373 14187
rect 21373 14153 21407 14187
rect 21407 14153 21416 14187
rect 21364 14144 21416 14153
rect 24768 14144 24820 14196
rect 25412 14144 25464 14196
rect 16948 14076 17000 14128
rect 16028 14008 16080 14060
rect 17776 14076 17828 14128
rect 24032 14008 24084 14060
rect 24308 14008 24360 14060
rect 21180 13940 21232 13992
rect 22008 13940 22060 13992
rect 22284 13983 22336 13992
rect 22284 13949 22293 13983
rect 22293 13949 22327 13983
rect 22327 13949 22336 13983
rect 22284 13940 22336 13949
rect 5648 13838 5700 13890
rect 5712 13838 5764 13890
rect 5776 13838 5828 13890
rect 5840 13838 5892 13890
rect 14982 13838 15034 13890
rect 15046 13838 15098 13890
rect 15110 13838 15162 13890
rect 15174 13838 15226 13890
rect 24315 13838 24367 13890
rect 24379 13838 24431 13890
rect 24443 13838 24495 13890
rect 24507 13838 24559 13890
rect 15384 13736 15436 13788
rect 16120 13779 16172 13788
rect 16120 13745 16129 13779
rect 16129 13745 16163 13779
rect 16163 13745 16172 13779
rect 16120 13736 16172 13745
rect 16856 13736 16908 13788
rect 23664 13779 23716 13788
rect 23664 13745 23673 13779
rect 23673 13745 23707 13779
rect 23707 13745 23716 13779
rect 23664 13736 23716 13745
rect 24124 13779 24176 13788
rect 24124 13745 24133 13779
rect 24133 13745 24167 13779
rect 24167 13745 24176 13779
rect 24124 13736 24176 13745
rect 24676 13736 24728 13788
rect 25412 13736 25464 13788
rect 16948 13668 17000 13720
rect 17316 13600 17368 13652
rect 17776 13643 17828 13652
rect 17776 13609 17785 13643
rect 17785 13609 17819 13643
rect 17819 13609 17828 13643
rect 17776 13600 17828 13609
rect 21364 13643 21416 13652
rect 21364 13609 21373 13643
rect 21373 13609 21407 13643
rect 21407 13609 21416 13643
rect 21364 13600 21416 13609
rect 24768 13600 24820 13652
rect 25228 13643 25280 13652
rect 25228 13609 25237 13643
rect 25237 13609 25271 13643
rect 25271 13609 25280 13643
rect 25228 13600 25280 13609
rect 15476 13532 15528 13584
rect 17500 13575 17552 13584
rect 17500 13541 17509 13575
rect 17509 13541 17543 13575
rect 17543 13541 17552 13575
rect 17500 13532 17552 13541
rect 20720 13575 20772 13584
rect 20720 13541 20729 13575
rect 20729 13541 20763 13575
rect 20763 13541 20772 13575
rect 20720 13532 20772 13541
rect 24124 13532 24176 13584
rect 10315 13294 10367 13346
rect 10379 13294 10431 13346
rect 10443 13294 10495 13346
rect 10507 13294 10559 13346
rect 19648 13294 19700 13346
rect 19712 13294 19764 13346
rect 19776 13294 19828 13346
rect 19840 13294 19892 13346
rect 13636 13235 13688 13244
rect 13636 13201 13645 13235
rect 13645 13201 13679 13235
rect 13679 13201 13688 13235
rect 13636 13192 13688 13201
rect 17224 13192 17276 13244
rect 17776 13192 17828 13244
rect 22008 13235 22060 13244
rect 22008 13201 22017 13235
rect 22017 13201 22051 13235
rect 22051 13201 22060 13235
rect 22008 13192 22060 13201
rect 24216 13192 24268 13244
rect 20812 13124 20864 13176
rect 13452 13099 13504 13108
rect 13452 13065 13461 13099
rect 13461 13065 13495 13099
rect 13495 13065 13504 13099
rect 13452 13056 13504 13065
rect 16764 13099 16816 13108
rect 16764 13065 16773 13099
rect 16773 13065 16807 13099
rect 16807 13065 16816 13099
rect 16764 13056 16816 13065
rect 20628 13099 20680 13108
rect 20628 13065 20637 13099
rect 20637 13065 20671 13099
rect 20671 13065 20680 13099
rect 20628 13056 20680 13065
rect 24584 13099 24636 13108
rect 24584 13065 24593 13099
rect 24593 13065 24627 13099
rect 24627 13065 24636 13099
rect 24584 13056 24636 13065
rect 20996 12852 21048 12904
rect 5648 12750 5700 12802
rect 5712 12750 5764 12802
rect 5776 12750 5828 12802
rect 5840 12750 5892 12802
rect 14982 12750 15034 12802
rect 15046 12750 15098 12802
rect 15110 12750 15162 12802
rect 15174 12750 15226 12802
rect 24315 12750 24367 12802
rect 24379 12750 24431 12802
rect 24443 12750 24495 12802
rect 24507 12750 24559 12802
rect 13452 12691 13504 12700
rect 13452 12657 13461 12691
rect 13461 12657 13495 12691
rect 13495 12657 13504 12691
rect 13452 12648 13504 12657
rect 20260 12648 20312 12700
rect 20628 12691 20680 12700
rect 20628 12657 20637 12691
rect 20637 12657 20671 12691
rect 20671 12657 20680 12691
rect 20628 12648 20680 12657
rect 23940 12691 23992 12700
rect 23940 12657 23949 12691
rect 23949 12657 23983 12691
rect 23983 12657 23992 12691
rect 23940 12648 23992 12657
rect 24676 12691 24728 12700
rect 24676 12657 24685 12691
rect 24685 12657 24719 12691
rect 24719 12657 24728 12691
rect 24676 12648 24728 12657
rect 15476 12555 15528 12564
rect 15476 12521 15485 12555
rect 15485 12521 15519 12555
rect 15519 12521 15528 12555
rect 15476 12512 15528 12521
rect 16764 12512 16816 12564
rect 24400 12555 24452 12564
rect 24400 12521 24409 12555
rect 24409 12521 24443 12555
rect 24443 12521 24452 12555
rect 24400 12512 24452 12521
rect 12532 12487 12584 12496
rect 12532 12453 12541 12487
rect 12541 12453 12575 12487
rect 12575 12453 12584 12487
rect 12532 12444 12584 12453
rect 15660 12444 15712 12496
rect 20996 12444 21048 12496
rect 25596 12648 25648 12700
rect 23848 12376 23900 12428
rect 24124 12376 24176 12428
rect 18328 12308 18380 12360
rect 19984 12308 20036 12360
rect 21916 12308 21968 12360
rect 25688 12308 25740 12360
rect 10315 12206 10367 12258
rect 10379 12206 10431 12258
rect 10443 12206 10495 12258
rect 10507 12206 10559 12258
rect 19648 12206 19700 12258
rect 19712 12206 19764 12258
rect 19776 12206 19828 12258
rect 19840 12206 19892 12258
rect 12532 12104 12584 12156
rect 15660 12147 15712 12156
rect 15660 12113 15669 12147
rect 15669 12113 15703 12147
rect 15703 12113 15712 12147
rect 15660 12104 15712 12113
rect 20720 12104 20772 12156
rect 24032 12104 24084 12156
rect 13268 11968 13320 12020
rect 16028 12011 16080 12020
rect 16028 11977 16037 12011
rect 16037 11977 16071 12011
rect 16071 11977 16080 12011
rect 16028 11968 16080 11977
rect 19984 11968 20036 12020
rect 24400 12011 24452 12020
rect 24400 11977 24409 12011
rect 24409 11977 24443 12011
rect 24443 11977 24452 12011
rect 24400 11968 24452 11977
rect 13636 11943 13688 11952
rect 13636 11909 13645 11943
rect 13645 11909 13679 11943
rect 13679 11909 13688 11943
rect 13636 11900 13688 11909
rect 14004 11900 14056 11952
rect 15936 11900 15988 11952
rect 16396 11900 16448 11952
rect 18236 11900 18288 11952
rect 20904 11900 20956 11952
rect 20812 11832 20864 11884
rect 21916 11900 21968 11952
rect 12716 11807 12768 11816
rect 12716 11773 12725 11807
rect 12725 11773 12759 11807
rect 12759 11773 12768 11807
rect 12716 11764 12768 11773
rect 18788 11807 18840 11816
rect 18788 11773 18797 11807
rect 18797 11773 18831 11807
rect 18831 11773 18840 11807
rect 18788 11764 18840 11773
rect 5648 11662 5700 11714
rect 5712 11662 5764 11714
rect 5776 11662 5828 11714
rect 5840 11662 5892 11714
rect 14982 11662 15034 11714
rect 15046 11662 15098 11714
rect 15110 11662 15162 11714
rect 15174 11662 15226 11714
rect 24315 11662 24367 11714
rect 24379 11662 24431 11714
rect 24443 11662 24495 11714
rect 24507 11662 24559 11714
rect 18328 11603 18380 11612
rect 18328 11569 18337 11603
rect 18337 11569 18371 11603
rect 18371 11569 18380 11603
rect 18328 11560 18380 11569
rect 19984 11603 20036 11612
rect 19984 11569 19993 11603
rect 19993 11569 20027 11603
rect 20027 11569 20036 11603
rect 19984 11560 20036 11569
rect 20904 11603 20956 11612
rect 20904 11569 20913 11603
rect 20913 11569 20947 11603
rect 20947 11569 20956 11603
rect 20904 11560 20956 11569
rect 21916 11603 21968 11612
rect 21916 11569 21925 11603
rect 21925 11569 21959 11603
rect 21959 11569 21968 11603
rect 21916 11560 21968 11569
rect 24676 11560 24728 11612
rect 18236 11535 18288 11544
rect 18236 11501 18245 11535
rect 18245 11501 18279 11535
rect 18279 11501 18288 11535
rect 18236 11492 18288 11501
rect 12440 11288 12492 11340
rect 12716 11356 12768 11408
rect 14556 11356 14608 11408
rect 16304 11356 16356 11408
rect 18788 11467 18840 11476
rect 18788 11433 18797 11467
rect 18797 11433 18831 11467
rect 18831 11433 18840 11467
rect 18788 11424 18840 11433
rect 20996 11424 21048 11476
rect 22192 11424 22244 11476
rect 16488 11288 16540 11340
rect 18880 11288 18932 11340
rect 21272 11331 21324 11340
rect 21272 11297 21281 11331
rect 21281 11297 21315 11331
rect 21315 11297 21324 11331
rect 21272 11288 21324 11297
rect 14004 11263 14056 11272
rect 14004 11229 14013 11263
rect 14013 11229 14047 11263
rect 14047 11229 14056 11263
rect 14004 11220 14056 11229
rect 14740 11263 14792 11272
rect 14740 11229 14749 11263
rect 14749 11229 14783 11263
rect 14783 11229 14792 11263
rect 14740 11220 14792 11229
rect 16396 11220 16448 11272
rect 19524 11220 19576 11272
rect 10315 11118 10367 11170
rect 10379 11118 10431 11170
rect 10443 11118 10495 11170
rect 10507 11118 10559 11170
rect 19648 11118 19700 11170
rect 19712 11118 19764 11170
rect 19776 11118 19828 11170
rect 19840 11118 19892 11170
rect 13268 11059 13320 11068
rect 13268 11025 13277 11059
rect 13277 11025 13311 11059
rect 13311 11025 13320 11059
rect 13268 11016 13320 11025
rect 13636 11016 13688 11068
rect 14740 11016 14792 11068
rect 16028 11059 16080 11068
rect 16028 11025 16037 11059
rect 16037 11025 16071 11059
rect 16071 11025 16080 11059
rect 16028 11016 16080 11025
rect 18880 11016 18932 11068
rect 16396 10991 16448 11000
rect 16396 10957 16405 10991
rect 16405 10957 16439 10991
rect 16439 10957 16448 10991
rect 16396 10948 16448 10957
rect 20904 11016 20956 11068
rect 22192 11016 22244 11068
rect 24768 11059 24820 11068
rect 24768 11025 24777 11059
rect 24777 11025 24811 11059
rect 24811 11025 24820 11059
rect 24768 11016 24820 11025
rect 21364 10948 21416 11000
rect 14004 10880 14056 10932
rect 14832 10880 14884 10932
rect 18512 10880 18564 10932
rect 18696 10923 18748 10932
rect 18696 10889 18730 10923
rect 18730 10889 18748 10923
rect 18696 10880 18748 10889
rect 20260 10880 20312 10932
rect 20996 10880 21048 10932
rect 24676 10880 24728 10932
rect 14464 10676 14516 10728
rect 5648 10574 5700 10626
rect 5712 10574 5764 10626
rect 5776 10574 5828 10626
rect 5840 10574 5892 10626
rect 14982 10574 15034 10626
rect 15046 10574 15098 10626
rect 15110 10574 15162 10626
rect 15174 10574 15226 10626
rect 24315 10574 24367 10626
rect 24379 10574 24431 10626
rect 24443 10574 24495 10626
rect 24507 10574 24559 10626
rect 12716 10472 12768 10524
rect 13636 10472 13688 10524
rect 14556 10515 14608 10524
rect 14556 10481 14565 10515
rect 14565 10481 14599 10515
rect 14599 10481 14608 10515
rect 14556 10472 14608 10481
rect 14832 10515 14884 10524
rect 14832 10481 14841 10515
rect 14841 10481 14875 10515
rect 14875 10481 14884 10515
rect 14832 10472 14884 10481
rect 16396 10515 16448 10524
rect 16396 10481 16405 10515
rect 16405 10481 16439 10515
rect 16439 10481 16448 10515
rect 16396 10472 16448 10481
rect 16856 10472 16908 10524
rect 18880 10515 18932 10524
rect 18880 10481 18889 10515
rect 18889 10481 18923 10515
rect 18923 10481 18932 10515
rect 18880 10472 18932 10481
rect 20996 10472 21048 10524
rect 21364 10472 21416 10524
rect 23480 10472 23532 10524
rect 24676 10404 24728 10456
rect 10968 10311 11020 10320
rect 10968 10277 10977 10311
rect 10977 10277 11011 10311
rect 11011 10277 11020 10311
rect 10968 10268 11020 10277
rect 12440 10268 12492 10320
rect 16304 10268 16356 10320
rect 16856 10311 16908 10320
rect 16856 10277 16865 10311
rect 16865 10277 16899 10311
rect 16899 10277 16908 10311
rect 16856 10268 16908 10277
rect 10784 10243 10836 10252
rect 10784 10209 10793 10243
rect 10793 10209 10827 10243
rect 10827 10209 10836 10243
rect 10784 10200 10836 10209
rect 13820 10243 13872 10252
rect 13820 10209 13829 10243
rect 13829 10209 13863 10243
rect 13863 10209 13872 10243
rect 13820 10200 13872 10209
rect 13912 10243 13964 10252
rect 13912 10209 13921 10243
rect 13921 10209 13955 10243
rect 13955 10209 13964 10243
rect 13912 10200 13964 10209
rect 16396 10200 16448 10252
rect 18696 10200 18748 10252
rect 19248 10175 19300 10184
rect 19248 10141 19257 10175
rect 19257 10141 19291 10175
rect 19291 10141 19300 10175
rect 19248 10132 19300 10141
rect 25228 10175 25280 10184
rect 25228 10141 25237 10175
rect 25237 10141 25271 10175
rect 25271 10141 25280 10175
rect 25228 10132 25280 10141
rect 10315 10030 10367 10082
rect 10379 10030 10431 10082
rect 10443 10030 10495 10082
rect 10507 10030 10559 10082
rect 19648 10030 19700 10082
rect 19712 10030 19764 10082
rect 19776 10030 19828 10082
rect 19840 10030 19892 10082
rect 10968 9971 11020 9980
rect 10968 9937 10977 9971
rect 10977 9937 11011 9971
rect 11011 9937 11020 9971
rect 10968 9928 11020 9937
rect 13912 9928 13964 9980
rect 15936 9971 15988 9980
rect 15936 9937 15945 9971
rect 15945 9937 15979 9971
rect 15979 9937 15988 9971
rect 15936 9928 15988 9937
rect 18788 9971 18840 9980
rect 18788 9937 18797 9971
rect 18797 9937 18831 9971
rect 18831 9937 18840 9971
rect 18788 9928 18840 9937
rect 19156 9928 19208 9980
rect 19524 9928 19576 9980
rect 24768 9971 24820 9980
rect 24768 9937 24777 9971
rect 24777 9937 24811 9971
rect 24811 9937 24820 9971
rect 24768 9928 24820 9937
rect 16028 9792 16080 9844
rect 18880 9792 18932 9844
rect 24676 9792 24728 9844
rect 16396 9767 16448 9776
rect 16396 9733 16405 9767
rect 16405 9733 16439 9767
rect 16439 9733 16448 9767
rect 16396 9724 16448 9733
rect 16488 9767 16540 9776
rect 16488 9733 16497 9767
rect 16497 9733 16531 9767
rect 16531 9733 16540 9767
rect 19432 9767 19484 9776
rect 16488 9724 16540 9733
rect 19432 9733 19441 9767
rect 19441 9733 19475 9767
rect 19475 9733 19484 9767
rect 19432 9724 19484 9733
rect 5648 9486 5700 9538
rect 5712 9486 5764 9538
rect 5776 9486 5828 9538
rect 5840 9486 5892 9538
rect 14982 9486 15034 9538
rect 15046 9486 15098 9538
rect 15110 9486 15162 9538
rect 15174 9486 15226 9538
rect 24315 9486 24367 9538
rect 24379 9486 24431 9538
rect 24443 9486 24495 9538
rect 24507 9486 24559 9538
rect 16396 9427 16448 9436
rect 16396 9393 16405 9427
rect 16405 9393 16439 9427
rect 16439 9393 16448 9427
rect 16396 9384 16448 9393
rect 16488 9384 16540 9436
rect 19156 9427 19208 9436
rect 19156 9393 19165 9427
rect 19165 9393 19199 9427
rect 19199 9393 19208 9427
rect 19156 9384 19208 9393
rect 19432 9316 19484 9368
rect 24768 9359 24820 9368
rect 24768 9325 24777 9359
rect 24777 9325 24811 9359
rect 24811 9325 24820 9359
rect 24768 9316 24820 9325
rect 25228 9359 25280 9368
rect 25228 9325 25237 9359
rect 25237 9325 25271 9359
rect 25271 9325 25280 9359
rect 25228 9316 25280 9325
rect 16028 9087 16080 9096
rect 16028 9053 16037 9087
rect 16037 9053 16071 9087
rect 16071 9053 16080 9087
rect 16028 9044 16080 9053
rect 18880 9087 18932 9096
rect 18880 9053 18889 9087
rect 18889 9053 18923 9087
rect 18923 9053 18932 9087
rect 18880 9044 18932 9053
rect 24492 9087 24544 9096
rect 24492 9053 24501 9087
rect 24501 9053 24535 9087
rect 24535 9053 24544 9087
rect 24492 9044 24544 9053
rect 10315 8942 10367 8994
rect 10379 8942 10431 8994
rect 10443 8942 10495 8994
rect 10507 8942 10559 8994
rect 19648 8942 19700 8994
rect 19712 8942 19764 8994
rect 19776 8942 19828 8994
rect 19840 8942 19892 8994
rect 24768 8883 24820 8892
rect 24768 8849 24777 8883
rect 24777 8849 24811 8883
rect 24811 8849 24820 8883
rect 24768 8840 24820 8849
rect 24676 8704 24728 8756
rect 5648 8398 5700 8450
rect 5712 8398 5764 8450
rect 5776 8398 5828 8450
rect 5840 8398 5892 8450
rect 14982 8398 15034 8450
rect 15046 8398 15098 8450
rect 15110 8398 15162 8450
rect 15174 8398 15226 8450
rect 24315 8398 24367 8450
rect 24379 8398 24431 8450
rect 24443 8398 24495 8450
rect 24507 8398 24559 8450
rect 24676 8339 24728 8348
rect 24676 8305 24685 8339
rect 24685 8305 24719 8339
rect 24719 8305 24728 8339
rect 24676 8296 24728 8305
rect 10315 7854 10367 7906
rect 10379 7854 10431 7906
rect 10443 7854 10495 7906
rect 10507 7854 10559 7906
rect 19648 7854 19700 7906
rect 19712 7854 19764 7906
rect 19776 7854 19828 7906
rect 19840 7854 19892 7906
rect 24584 7659 24636 7668
rect 24584 7625 24593 7659
rect 24593 7625 24627 7659
rect 24627 7625 24636 7659
rect 24584 7616 24636 7625
rect 24768 7523 24820 7532
rect 24768 7489 24777 7523
rect 24777 7489 24811 7523
rect 24811 7489 24820 7523
rect 24768 7480 24820 7489
rect 5648 7310 5700 7362
rect 5712 7310 5764 7362
rect 5776 7310 5828 7362
rect 5840 7310 5892 7362
rect 14982 7310 15034 7362
rect 15046 7310 15098 7362
rect 15110 7310 15162 7362
rect 15174 7310 15226 7362
rect 24315 7310 24367 7362
rect 24379 7310 24431 7362
rect 24443 7310 24495 7362
rect 24507 7310 24559 7362
rect 17868 7208 17920 7260
rect 23756 7208 23808 7260
rect 23940 7208 23992 7260
rect 24676 7251 24728 7260
rect 24676 7217 24685 7251
rect 24685 7217 24719 7251
rect 24719 7217 24728 7251
rect 24676 7208 24728 7217
rect 18236 7115 18288 7124
rect 18236 7081 18245 7115
rect 18245 7081 18279 7115
rect 18279 7081 18288 7115
rect 18236 7072 18288 7081
rect 10315 6766 10367 6818
rect 10379 6766 10431 6818
rect 10443 6766 10495 6818
rect 10507 6766 10559 6818
rect 19648 6766 19700 6818
rect 19712 6766 19764 6818
rect 19776 6766 19828 6818
rect 19840 6766 19892 6818
rect 5648 6222 5700 6274
rect 5712 6222 5764 6274
rect 5776 6222 5828 6274
rect 5840 6222 5892 6274
rect 14982 6222 15034 6274
rect 15046 6222 15098 6274
rect 15110 6222 15162 6274
rect 15174 6222 15226 6274
rect 24315 6222 24367 6274
rect 24379 6222 24431 6274
rect 24443 6222 24495 6274
rect 24507 6222 24559 6274
rect 16488 6163 16540 6172
rect 16488 6129 16497 6163
rect 16497 6129 16531 6163
rect 16531 6129 16540 6163
rect 16488 6120 16540 6129
rect 16948 5891 17000 5900
rect 16948 5857 16957 5891
rect 16957 5857 16991 5891
rect 16991 5857 17000 5891
rect 16948 5848 17000 5857
rect 10315 5678 10367 5730
rect 10379 5678 10431 5730
rect 10443 5678 10495 5730
rect 10507 5678 10559 5730
rect 19648 5678 19700 5730
rect 19712 5678 19764 5730
rect 19776 5678 19828 5730
rect 19840 5678 19892 5730
rect 5648 5134 5700 5186
rect 5712 5134 5764 5186
rect 5776 5134 5828 5186
rect 5840 5134 5892 5186
rect 14982 5134 15034 5186
rect 15046 5134 15098 5186
rect 15110 5134 15162 5186
rect 15174 5134 15226 5186
rect 24315 5134 24367 5186
rect 24379 5134 24431 5186
rect 24443 5134 24495 5186
rect 24507 5134 24559 5186
rect 15752 5032 15804 5084
rect 15936 4939 15988 4948
rect 15936 4905 15945 4939
rect 15945 4905 15979 4939
rect 15979 4905 15988 4939
rect 15936 4896 15988 4905
rect 10315 4590 10367 4642
rect 10379 4590 10431 4642
rect 10443 4590 10495 4642
rect 10507 4590 10559 4642
rect 19648 4590 19700 4642
rect 19712 4590 19764 4642
rect 19776 4590 19828 4642
rect 19840 4590 19892 4642
rect 5648 4046 5700 4098
rect 5712 4046 5764 4098
rect 5776 4046 5828 4098
rect 5840 4046 5892 4098
rect 14982 4046 15034 4098
rect 15046 4046 15098 4098
rect 15110 4046 15162 4098
rect 15174 4046 15226 4098
rect 24315 4046 24367 4098
rect 24379 4046 24431 4098
rect 24443 4046 24495 4098
rect 24507 4046 24559 4098
rect 24768 3647 24820 3656
rect 24768 3613 24777 3647
rect 24777 3613 24811 3647
rect 24811 3613 24820 3647
rect 24768 3604 24820 3613
rect 25228 3647 25280 3656
rect 25228 3613 25237 3647
rect 25237 3613 25271 3647
rect 25271 3613 25280 3647
rect 25228 3604 25280 3613
rect 10315 3502 10367 3554
rect 10379 3502 10431 3554
rect 10443 3502 10495 3554
rect 10507 3502 10559 3554
rect 19648 3502 19700 3554
rect 19712 3502 19764 3554
rect 19776 3502 19828 3554
rect 19840 3502 19892 3554
rect 5648 2958 5700 3010
rect 5712 2958 5764 3010
rect 5776 2958 5828 3010
rect 5840 2958 5892 3010
rect 14982 2958 15034 3010
rect 15046 2958 15098 3010
rect 15110 2958 15162 3010
rect 15174 2958 15226 3010
rect 24315 2958 24367 3010
rect 24379 2958 24431 3010
rect 24443 2958 24495 3010
rect 24507 2958 24559 3010
rect 10315 2414 10367 2466
rect 10379 2414 10431 2466
rect 10443 2414 10495 2466
rect 10507 2414 10559 2466
rect 19648 2414 19700 2466
rect 19712 2414 19764 2466
rect 19776 2414 19828 2466
rect 19840 2414 19892 2466
rect 5648 1870 5700 1922
rect 5712 1870 5764 1922
rect 5776 1870 5828 1922
rect 5840 1870 5892 1922
rect 14982 1870 15034 1922
rect 15046 1870 15098 1922
rect 15110 1870 15162 1922
rect 15174 1870 15226 1922
rect 24315 1870 24367 1922
rect 24379 1870 24431 1922
rect 24443 1870 24495 1922
rect 24507 1870 24559 1922
<< metal2 >>
rect 294 27240 350 27720
rect 938 27240 994 27720
rect 1582 27240 1638 27720
rect 2318 27240 2374 27720
rect 2962 27240 3018 27720
rect 3698 27240 3754 27720
rect 4342 27240 4398 27720
rect 4986 27240 5042 27720
rect 5722 27240 5778 27720
rect 6366 27240 6422 27720
rect 7102 27240 7158 27720
rect 7746 27240 7802 27720
rect 8390 27240 8446 27720
rect 9126 27240 9182 27720
rect 9770 27240 9826 27720
rect 10506 27240 10562 27720
rect 11150 27240 11206 27720
rect 11886 27240 11942 27720
rect 12530 27240 12586 27720
rect 13174 27240 13230 27720
rect 13910 27240 13966 27720
rect 14554 27240 14610 27720
rect 15290 27240 15346 27720
rect 15934 27240 15990 27720
rect 16578 27240 16634 27720
rect 17314 27240 17370 27720
rect 17958 27240 18014 27720
rect 18694 27240 18750 27720
rect 19338 27240 19394 27720
rect 20074 27240 20130 27720
rect 20718 27240 20774 27720
rect 21362 27240 21418 27720
rect 22098 27240 22154 27720
rect 22742 27240 22798 27720
rect 23478 27240 23534 27720
rect 23938 27424 23994 27433
rect 23938 27359 23994 27368
rect 308 16394 336 27240
rect 952 27138 980 27240
rect 952 27110 1348 27138
rect 216 16366 336 16394
rect 216 9753 244 16366
rect 1320 16281 1348 27110
rect 1596 16825 1624 27240
rect 1582 16816 1638 16825
rect 1582 16751 1638 16760
rect 2332 16417 2360 27240
rect 2976 18593 3004 27240
rect 3712 19001 3740 27240
rect 4356 20905 4384 27240
rect 5000 24033 5028 27240
rect 5736 24962 5764 27240
rect 5736 24934 6040 24962
rect 5622 24772 5918 24792
rect 5678 24770 5702 24772
rect 5758 24770 5782 24772
rect 5838 24770 5862 24772
rect 5700 24718 5702 24770
rect 5764 24718 5776 24770
rect 5838 24718 5840 24770
rect 5678 24716 5702 24718
rect 5758 24716 5782 24718
rect 5838 24716 5862 24718
rect 5622 24696 5918 24716
rect 4986 24024 5042 24033
rect 4986 23959 5042 23968
rect 5622 23684 5918 23704
rect 5678 23682 5702 23684
rect 5758 23682 5782 23684
rect 5838 23682 5862 23684
rect 5700 23630 5702 23682
rect 5764 23630 5776 23682
rect 5838 23630 5840 23682
rect 5678 23628 5702 23630
rect 5758 23628 5782 23630
rect 5838 23628 5862 23630
rect 5622 23608 5918 23628
rect 5622 22596 5918 22616
rect 5678 22594 5702 22596
rect 5758 22594 5782 22596
rect 5838 22594 5862 22596
rect 5700 22542 5702 22594
rect 5764 22542 5776 22594
rect 5838 22542 5840 22594
rect 5678 22540 5702 22542
rect 5758 22540 5782 22542
rect 5838 22540 5862 22542
rect 5622 22520 5918 22540
rect 5622 21508 5918 21528
rect 5678 21506 5702 21508
rect 5758 21506 5782 21508
rect 5838 21506 5862 21508
rect 5700 21454 5702 21506
rect 5764 21454 5776 21506
rect 5838 21454 5840 21506
rect 5678 21452 5702 21454
rect 5758 21452 5782 21454
rect 5838 21452 5862 21454
rect 5622 21432 5918 21452
rect 6012 21177 6040 24934
rect 6380 21313 6408 27240
rect 7116 21585 7144 27240
rect 7760 22401 7788 27240
rect 7746 22392 7802 22401
rect 7746 22327 7802 22336
rect 7102 21576 7158 21585
rect 7102 21511 7158 21520
rect 6366 21304 6422 21313
rect 6366 21239 6422 21248
rect 5998 21168 6054 21177
rect 5998 21103 6054 21112
rect 4342 20896 4398 20905
rect 4342 20831 4398 20840
rect 8404 20497 8432 27240
rect 8944 23036 8996 23042
rect 8944 22978 8996 22984
rect 8956 22498 8984 22978
rect 8944 22492 8996 22498
rect 8944 22434 8996 22440
rect 9140 20633 9168 27240
rect 9312 22832 9364 22838
rect 9218 22800 9274 22809
rect 9312 22774 9364 22780
rect 9218 22735 9220 22744
rect 9272 22735 9274 22744
rect 9220 22706 9272 22712
rect 9324 22650 9352 22774
rect 9232 22622 9352 22650
rect 9232 22158 9260 22622
rect 9784 22537 9812 27240
rect 10520 25506 10548 27240
rect 10152 25478 10548 25506
rect 9956 22968 10008 22974
rect 10152 22945 10180 25478
rect 10289 25316 10585 25336
rect 10345 25314 10369 25316
rect 10425 25314 10449 25316
rect 10505 25314 10529 25316
rect 10367 25262 10369 25314
rect 10431 25262 10443 25314
rect 10505 25262 10507 25314
rect 10345 25260 10369 25262
rect 10425 25260 10449 25262
rect 10505 25260 10529 25262
rect 10289 25240 10585 25260
rect 10289 24228 10585 24248
rect 10345 24226 10369 24228
rect 10425 24226 10449 24228
rect 10505 24226 10529 24228
rect 10367 24174 10369 24226
rect 10431 24174 10443 24226
rect 10505 24174 10507 24226
rect 10345 24172 10369 24174
rect 10425 24172 10449 24174
rect 10505 24172 10529 24174
rect 10289 24152 10585 24172
rect 10968 23920 11020 23926
rect 10968 23862 11020 23868
rect 10876 23784 10928 23790
rect 10876 23726 10928 23732
rect 10888 23382 10916 23726
rect 10784 23376 10836 23382
rect 10784 23318 10836 23324
rect 10876 23376 10928 23382
rect 10876 23318 10928 23324
rect 10289 23140 10585 23160
rect 10345 23138 10369 23140
rect 10425 23138 10449 23140
rect 10505 23138 10529 23140
rect 10367 23086 10369 23138
rect 10431 23086 10443 23138
rect 10505 23086 10507 23138
rect 10345 23084 10369 23086
rect 10425 23084 10449 23086
rect 10505 23084 10529 23086
rect 10289 23064 10585 23084
rect 9956 22910 10008 22916
rect 10138 22936 10194 22945
rect 9770 22528 9826 22537
rect 9968 22498 9996 22910
rect 10138 22871 10194 22880
rect 9770 22463 9826 22472
rect 9956 22492 10008 22498
rect 9956 22434 10008 22440
rect 10796 22362 10824 23318
rect 10888 23217 10916 23318
rect 10874 23208 10930 23217
rect 10874 23143 10930 23152
rect 10980 22974 11008 23862
rect 11164 23625 11192 27240
rect 11150 23616 11206 23625
rect 11150 23551 11206 23560
rect 11428 23240 11480 23246
rect 11428 23182 11480 23188
rect 11060 23036 11112 23042
rect 11060 22978 11112 22984
rect 10968 22968 11020 22974
rect 10968 22910 11020 22916
rect 11072 22498 11100 22978
rect 11152 22900 11204 22906
rect 11152 22842 11204 22848
rect 11060 22492 11112 22498
rect 11060 22434 11112 22440
rect 10784 22356 10836 22362
rect 10784 22298 10836 22304
rect 9220 22152 9272 22158
rect 9220 22094 9272 22100
rect 9232 20769 9260 22094
rect 10289 22052 10585 22072
rect 10345 22050 10369 22052
rect 10425 22050 10449 22052
rect 10505 22050 10529 22052
rect 10367 21998 10369 22050
rect 10431 21998 10443 22050
rect 10505 21998 10507 22050
rect 10345 21996 10369 21998
rect 10425 21996 10449 21998
rect 10505 21996 10529 21998
rect 10289 21976 10585 21996
rect 10796 21954 10824 22298
rect 11164 22158 11192 22842
rect 11440 22838 11468 23182
rect 11900 23042 11928 27240
rect 12544 24305 12572 27240
rect 13188 24441 13216 27240
rect 13634 24568 13690 24577
rect 13634 24503 13690 24512
rect 13174 24432 13230 24441
rect 13174 24367 13230 24376
rect 12530 24296 12586 24305
rect 12530 24231 12586 24240
rect 13268 23920 13320 23926
rect 13268 23862 13320 23868
rect 13280 23194 13308 23862
rect 13358 23616 13414 23625
rect 13358 23551 13360 23560
rect 13412 23551 13414 23560
rect 13360 23522 13412 23528
rect 13360 23240 13412 23246
rect 13280 23188 13360 23194
rect 13280 23182 13412 23188
rect 13280 23166 13400 23182
rect 11888 23036 11940 23042
rect 11888 22978 11940 22984
rect 13372 22838 13400 23166
rect 13452 22968 13504 22974
rect 13452 22910 13504 22916
rect 11428 22832 11480 22838
rect 11428 22774 11480 22780
rect 13360 22832 13412 22838
rect 13360 22774 13412 22780
rect 11440 22294 11468 22774
rect 13372 22498 13400 22774
rect 13360 22492 13412 22498
rect 13360 22434 13412 22440
rect 11428 22288 11480 22294
rect 11428 22230 11480 22236
rect 11152 22152 11204 22158
rect 11152 22094 11204 22100
rect 10784 21948 10836 21954
rect 10784 21890 10836 21896
rect 10796 21410 10824 21890
rect 10784 21404 10836 21410
rect 10784 21346 10836 21352
rect 10692 21132 10744 21138
rect 10692 21074 10744 21080
rect 10289 20964 10585 20984
rect 10345 20962 10369 20964
rect 10425 20962 10449 20964
rect 10505 20962 10529 20964
rect 10367 20910 10369 20962
rect 10431 20910 10443 20962
rect 10505 20910 10507 20962
rect 10345 20908 10369 20910
rect 10425 20908 10449 20910
rect 10505 20908 10529 20910
rect 10289 20888 10585 20908
rect 10704 20905 10732 21074
rect 10690 20896 10746 20905
rect 10690 20831 10692 20840
rect 10744 20831 10746 20840
rect 10692 20802 10744 20808
rect 9218 20760 9274 20769
rect 9218 20695 9274 20704
rect 9126 20624 9182 20633
rect 9126 20559 9182 20568
rect 8390 20488 8446 20497
rect 5622 20420 5918 20440
rect 8390 20423 8446 20432
rect 5678 20418 5702 20420
rect 5758 20418 5782 20420
rect 5838 20418 5862 20420
rect 5700 20366 5702 20418
rect 5764 20366 5776 20418
rect 5838 20366 5840 20418
rect 5678 20364 5702 20366
rect 5758 20364 5782 20366
rect 5838 20364 5862 20366
rect 5622 20344 5918 20364
rect 10796 20186 10824 21346
rect 10968 20792 11020 20798
rect 10968 20734 11020 20740
rect 10980 20322 11008 20734
rect 11164 20730 11192 22094
rect 11440 21954 11468 22230
rect 13084 22152 13136 22158
rect 13084 22094 13136 22100
rect 13096 21954 13124 22094
rect 11428 21948 11480 21954
rect 11428 21890 11480 21896
rect 13084 21948 13136 21954
rect 13084 21890 13136 21896
rect 13464 21886 13492 22910
rect 13542 22256 13598 22265
rect 13542 22191 13598 22200
rect 13556 22158 13584 22191
rect 13544 22152 13596 22158
rect 13544 22094 13596 22100
rect 13452 21880 13504 21886
rect 13452 21822 13504 21828
rect 11242 21304 11298 21313
rect 11242 21239 11298 21248
rect 11256 20798 11284 21239
rect 11796 21064 11848 21070
rect 11796 21006 11848 21012
rect 13176 21064 13228 21070
rect 13176 21006 13228 21012
rect 11244 20792 11296 20798
rect 11244 20734 11296 20740
rect 11152 20724 11204 20730
rect 11152 20666 11204 20672
rect 10968 20316 11020 20322
rect 10968 20258 11020 20264
rect 10784 20180 10836 20186
rect 10784 20122 10836 20128
rect 10692 19976 10744 19982
rect 10690 19944 10692 19953
rect 11164 19953 11192 20666
rect 11808 20662 11836 21006
rect 12900 20860 12952 20866
rect 12900 20802 12952 20808
rect 12912 20662 12940 20802
rect 13188 20730 13216 21006
rect 13176 20724 13228 20730
rect 13176 20666 13228 20672
rect 11796 20656 11848 20662
rect 11796 20598 11848 20604
rect 12900 20656 12952 20662
rect 12900 20598 12952 20604
rect 12992 20656 13044 20662
rect 12992 20598 13044 20604
rect 11244 20180 11296 20186
rect 11244 20122 11296 20128
rect 10744 19944 10746 19953
rect 10289 19876 10585 19896
rect 10690 19879 10746 19888
rect 11150 19944 11206 19953
rect 11150 19879 11206 19888
rect 10345 19874 10369 19876
rect 10425 19874 10449 19876
rect 10505 19874 10529 19876
rect 10367 19822 10369 19874
rect 10431 19822 10443 19874
rect 10505 19822 10507 19874
rect 10345 19820 10369 19822
rect 10425 19820 10449 19822
rect 10505 19820 10529 19822
rect 10289 19800 10585 19820
rect 11256 19710 11284 20122
rect 11808 20118 11836 20598
rect 12912 20254 12940 20598
rect 13004 20322 13032 20598
rect 13188 20322 13216 20666
rect 13358 20488 13414 20497
rect 13358 20423 13414 20432
rect 12992 20316 13044 20322
rect 12992 20258 13044 20264
rect 13176 20316 13228 20322
rect 13176 20258 13228 20264
rect 12900 20248 12952 20254
rect 12900 20190 12952 20196
rect 11796 20112 11848 20118
rect 11796 20054 11848 20060
rect 11808 19778 11836 20054
rect 13004 19778 13032 20258
rect 13372 19778 13400 20423
rect 11796 19772 11848 19778
rect 11796 19714 11848 19720
rect 12348 19772 12400 19778
rect 12348 19714 12400 19720
rect 12992 19772 13044 19778
rect 12992 19714 13044 19720
rect 13360 19772 13412 19778
rect 13360 19714 13412 19720
rect 11244 19704 11296 19710
rect 11244 19646 11296 19652
rect 5622 19332 5918 19352
rect 5678 19330 5702 19332
rect 5758 19330 5782 19332
rect 5838 19330 5862 19332
rect 5700 19278 5702 19330
rect 5764 19278 5776 19330
rect 5838 19278 5840 19330
rect 5678 19276 5702 19278
rect 5758 19276 5782 19278
rect 5838 19276 5862 19278
rect 5622 19256 5918 19276
rect 11256 19234 11284 19646
rect 11244 19228 11296 19234
rect 11244 19170 11296 19176
rect 12072 19092 12124 19098
rect 12072 19034 12124 19040
rect 3698 18992 3754 19001
rect 3698 18927 3754 18936
rect 10289 18788 10585 18808
rect 10345 18786 10369 18788
rect 10425 18786 10449 18788
rect 10505 18786 10529 18788
rect 10367 18734 10369 18786
rect 10431 18734 10443 18786
rect 10505 18734 10507 18786
rect 10345 18732 10369 18734
rect 10425 18732 10449 18734
rect 10505 18732 10529 18734
rect 10289 18712 10585 18732
rect 2962 18584 3018 18593
rect 12084 18554 12112 19034
rect 12360 19030 12388 19714
rect 12348 19024 12400 19030
rect 12348 18966 12400 18972
rect 12360 18690 12388 18966
rect 13372 18690 13400 19714
rect 13544 19704 13596 19710
rect 13544 19646 13596 19652
rect 13556 18865 13584 19646
rect 13542 18856 13598 18865
rect 13542 18791 13598 18800
rect 12348 18684 12400 18690
rect 12348 18626 12400 18632
rect 13360 18684 13412 18690
rect 13360 18626 13412 18632
rect 13556 18554 13584 18791
rect 2962 18519 3018 18528
rect 12072 18548 12124 18554
rect 12072 18490 12124 18496
rect 13360 18548 13412 18554
rect 13360 18490 13412 18496
rect 13544 18548 13596 18554
rect 13544 18490 13596 18496
rect 13268 18480 13320 18486
rect 13268 18422 13320 18428
rect 5622 18244 5918 18264
rect 5678 18242 5702 18244
rect 5758 18242 5782 18244
rect 5838 18242 5862 18244
rect 5700 18190 5702 18242
rect 5764 18190 5776 18242
rect 5838 18190 5840 18242
rect 5678 18188 5702 18190
rect 5758 18188 5782 18190
rect 5838 18188 5862 18190
rect 5622 18168 5918 18188
rect 13280 17806 13308 18422
rect 13268 17800 13320 17806
rect 13268 17742 13320 17748
rect 10289 17700 10585 17720
rect 10345 17698 10369 17700
rect 10425 17698 10449 17700
rect 10505 17698 10529 17700
rect 10367 17646 10369 17698
rect 10431 17646 10443 17698
rect 10505 17646 10507 17698
rect 10345 17644 10369 17646
rect 10425 17644 10449 17646
rect 10505 17644 10529 17646
rect 10289 17624 10585 17644
rect 12164 17256 12216 17262
rect 12164 17198 12216 17204
rect 5622 17156 5918 17176
rect 5678 17154 5702 17156
rect 5758 17154 5782 17156
rect 5838 17154 5862 17156
rect 5700 17102 5702 17154
rect 5764 17102 5776 17154
rect 5838 17102 5840 17154
rect 5678 17100 5702 17102
rect 5758 17100 5782 17102
rect 5838 17100 5862 17102
rect 5622 17080 5918 17100
rect 12176 16922 12204 17198
rect 12164 16916 12216 16922
rect 12164 16858 12216 16864
rect 12624 16916 12676 16922
rect 12624 16858 12676 16864
rect 12256 16848 12308 16854
rect 11886 16816 11942 16825
rect 12256 16790 12308 16796
rect 11886 16751 11888 16760
rect 11940 16751 11942 16760
rect 11888 16722 11940 16728
rect 10289 16612 10585 16632
rect 10345 16610 10369 16612
rect 10425 16610 10449 16612
rect 10505 16610 10529 16612
rect 10367 16558 10369 16610
rect 10431 16558 10443 16610
rect 10505 16558 10507 16610
rect 10345 16556 10369 16558
rect 10425 16556 10449 16558
rect 10505 16556 10529 16558
rect 10289 16536 10585 16556
rect 12268 16514 12296 16790
rect 12256 16508 12308 16514
rect 12256 16450 12308 16456
rect 2318 16408 2374 16417
rect 2318 16343 2374 16352
rect 12440 16304 12492 16310
rect 1306 16272 1362 16281
rect 12440 16246 12492 16252
rect 1306 16207 1362 16216
rect 5622 16068 5918 16088
rect 5678 16066 5702 16068
rect 5758 16066 5782 16068
rect 5838 16066 5862 16068
rect 5700 16014 5702 16066
rect 5764 16014 5776 16066
rect 5838 16014 5840 16066
rect 5678 16012 5702 16014
rect 5758 16012 5782 16014
rect 5838 16012 5862 16014
rect 5622 15992 5918 16012
rect 12452 15766 12480 16246
rect 12440 15760 12492 15766
rect 12440 15702 12492 15708
rect 12452 15630 12480 15702
rect 12636 15698 12664 16858
rect 13372 16854 13400 18490
rect 13544 17052 13596 17058
rect 13544 16994 13596 17000
rect 13360 16848 13412 16854
rect 13360 16790 13412 16796
rect 13556 16514 13584 16994
rect 13544 16508 13596 16514
rect 13544 16450 13596 16456
rect 12624 15692 12676 15698
rect 12624 15634 12676 15640
rect 12440 15624 12492 15630
rect 12440 15566 12492 15572
rect 10289 15524 10585 15544
rect 10345 15522 10369 15524
rect 10425 15522 10449 15524
rect 10505 15522 10529 15524
rect 10367 15470 10369 15522
rect 10431 15470 10443 15522
rect 10505 15470 10507 15522
rect 10345 15468 10369 15470
rect 10425 15468 10449 15470
rect 10505 15468 10529 15470
rect 10289 15448 10585 15468
rect 12452 15222 12480 15566
rect 12716 15284 12768 15290
rect 12716 15226 12768 15232
rect 12440 15216 12492 15222
rect 12728 15193 12756 15226
rect 12440 15158 12492 15164
rect 12714 15184 12770 15193
rect 5622 14980 5918 15000
rect 5678 14978 5702 14980
rect 5758 14978 5782 14980
rect 5838 14978 5862 14980
rect 5700 14926 5702 14978
rect 5764 14926 5776 14978
rect 5838 14926 5840 14978
rect 5678 14924 5702 14926
rect 5758 14924 5782 14926
rect 5838 14924 5862 14926
rect 5622 14904 5918 14924
rect 12452 14542 12480 15158
rect 12714 15119 12770 15128
rect 12728 14882 12756 15119
rect 12716 14876 12768 14882
rect 12716 14818 12768 14824
rect 12440 14536 12492 14542
rect 12440 14478 12492 14484
rect 10289 14436 10585 14456
rect 10345 14434 10369 14436
rect 10425 14434 10449 14436
rect 10505 14434 10529 14436
rect 10367 14382 10369 14434
rect 10431 14382 10443 14434
rect 10505 14382 10507 14434
rect 10345 14380 10369 14382
rect 10425 14380 10449 14382
rect 10505 14380 10529 14382
rect 10289 14360 10585 14380
rect 5622 13892 5918 13912
rect 5678 13890 5702 13892
rect 5758 13890 5782 13892
rect 5838 13890 5862 13892
rect 5700 13838 5702 13890
rect 5764 13838 5776 13890
rect 5838 13838 5840 13890
rect 5678 13836 5702 13838
rect 5758 13836 5782 13838
rect 5838 13836 5862 13838
rect 5622 13816 5918 13836
rect 10289 13348 10585 13368
rect 10345 13346 10369 13348
rect 10425 13346 10449 13348
rect 10505 13346 10529 13348
rect 10367 13294 10369 13346
rect 10431 13294 10443 13346
rect 10505 13294 10507 13346
rect 10345 13292 10369 13294
rect 10425 13292 10449 13294
rect 10505 13292 10529 13294
rect 10289 13272 10585 13292
rect 5622 12804 5918 12824
rect 5678 12802 5702 12804
rect 5758 12802 5782 12804
rect 5838 12802 5862 12804
rect 5700 12750 5702 12802
rect 5764 12750 5776 12802
rect 5838 12750 5840 12802
rect 5678 12748 5702 12750
rect 5758 12748 5782 12750
rect 5838 12748 5862 12750
rect 5622 12728 5918 12748
rect 10289 12260 10585 12280
rect 10345 12258 10369 12260
rect 10425 12258 10449 12260
rect 10505 12258 10529 12260
rect 10367 12206 10369 12258
rect 10431 12206 10443 12258
rect 10505 12206 10507 12258
rect 10345 12204 10369 12206
rect 10425 12204 10449 12206
rect 10505 12204 10529 12206
rect 10289 12184 10585 12204
rect 5622 11716 5918 11736
rect 5678 11714 5702 11716
rect 5758 11714 5782 11716
rect 5838 11714 5862 11716
rect 5700 11662 5702 11714
rect 5764 11662 5776 11714
rect 5838 11662 5840 11714
rect 5678 11660 5702 11662
rect 5758 11660 5782 11662
rect 5838 11660 5862 11662
rect 5622 11640 5918 11660
rect 12452 11346 12480 14478
rect 13648 13250 13676 24503
rect 13820 23240 13872 23246
rect 13820 23182 13872 23188
rect 13832 22362 13860 23182
rect 13820 22356 13872 22362
rect 13820 22298 13872 22304
rect 13832 21954 13860 22298
rect 13820 21948 13872 21954
rect 13820 21890 13872 21896
rect 13728 20520 13780 20526
rect 13728 20462 13780 20468
rect 13740 20118 13768 20462
rect 13728 20112 13780 20118
rect 13728 20054 13780 20060
rect 13728 19568 13780 19574
rect 13728 19510 13780 19516
rect 13740 18894 13768 19510
rect 13924 19137 13952 27240
rect 14568 24577 14596 27240
rect 14956 24772 15252 24792
rect 15012 24770 15036 24772
rect 15092 24770 15116 24772
rect 15172 24770 15196 24772
rect 15034 24718 15036 24770
rect 15098 24718 15110 24770
rect 15172 24718 15174 24770
rect 15012 24716 15036 24718
rect 15092 24716 15116 24718
rect 15172 24716 15196 24718
rect 14956 24696 15252 24716
rect 14554 24568 14610 24577
rect 14554 24503 14610 24512
rect 14832 23988 14884 23994
rect 14832 23930 14884 23936
rect 14844 23897 14872 23930
rect 14830 23888 14886 23897
rect 14830 23823 14886 23832
rect 14188 23784 14240 23790
rect 14188 23726 14240 23732
rect 14200 23450 14228 23726
rect 14844 23586 14872 23823
rect 14956 23684 15252 23704
rect 15012 23682 15036 23684
rect 15092 23682 15116 23684
rect 15172 23682 15196 23684
rect 15034 23630 15036 23682
rect 15098 23630 15110 23682
rect 15172 23630 15174 23682
rect 15012 23628 15036 23630
rect 15092 23628 15116 23630
rect 15172 23628 15196 23630
rect 14956 23608 15252 23628
rect 14832 23580 14884 23586
rect 14832 23522 14884 23528
rect 14188 23444 14240 23450
rect 14188 23386 14240 23392
rect 14094 23208 14150 23217
rect 14094 23143 14150 23152
rect 14108 22362 14136 23143
rect 14200 22974 14228 23386
rect 14832 23240 14884 23246
rect 14738 23208 14794 23217
rect 14832 23182 14884 23188
rect 14738 23143 14794 23152
rect 14752 23042 14780 23143
rect 14740 23036 14792 23042
rect 14740 22978 14792 22984
rect 14188 22968 14240 22974
rect 14188 22910 14240 22916
rect 14738 22528 14794 22537
rect 14738 22463 14740 22472
rect 14792 22463 14794 22472
rect 14740 22434 14792 22440
rect 14096 22356 14148 22362
rect 14096 22298 14148 22304
rect 14108 21886 14136 22298
rect 14096 21880 14148 21886
rect 14096 21822 14148 21828
rect 14186 21304 14242 21313
rect 14186 21239 14188 21248
rect 14240 21239 14242 21248
rect 14188 21210 14240 21216
rect 14004 21200 14056 21206
rect 14004 21142 14056 21148
rect 14016 20866 14044 21142
rect 14004 20860 14056 20866
rect 14004 20802 14056 20808
rect 14372 20724 14424 20730
rect 14372 20666 14424 20672
rect 14384 20322 14412 20666
rect 14464 20656 14516 20662
rect 14464 20598 14516 20604
rect 14648 20656 14700 20662
rect 14648 20598 14700 20604
rect 14372 20316 14424 20322
rect 14372 20258 14424 20264
rect 14002 20080 14058 20089
rect 14002 20015 14004 20024
rect 14056 20015 14058 20024
rect 14004 19986 14056 19992
rect 14476 19778 14504 20598
rect 14660 20322 14688 20598
rect 14648 20316 14700 20322
rect 14648 20258 14700 20264
rect 14464 19772 14516 19778
rect 14464 19714 14516 19720
rect 14660 19710 14688 20258
rect 14740 19976 14792 19982
rect 14740 19918 14792 19924
rect 14648 19704 14700 19710
rect 14648 19646 14700 19652
rect 14752 19574 14780 19918
rect 14740 19568 14792 19574
rect 14740 19510 14792 19516
rect 13910 19128 13966 19137
rect 13910 19063 13966 19072
rect 14752 18894 14780 19510
rect 13728 18888 13780 18894
rect 13728 18830 13780 18836
rect 14740 18888 14792 18894
rect 14740 18830 14792 18836
rect 13740 18554 13768 18830
rect 13728 18548 13780 18554
rect 13728 18490 13780 18496
rect 13740 18146 13768 18490
rect 13728 18140 13780 18146
rect 13728 18082 13780 18088
rect 14752 17874 14780 18830
rect 14740 17868 14792 17874
rect 14740 17810 14792 17816
rect 13728 17800 13780 17806
rect 13728 17742 13780 17748
rect 14280 17800 14332 17806
rect 14280 17742 14332 17748
rect 13740 16718 13768 17742
rect 14292 17466 14320 17742
rect 14280 17460 14332 17466
rect 14280 17402 14332 17408
rect 14556 17392 14608 17398
rect 14094 17360 14150 17369
rect 14556 17334 14608 17340
rect 14740 17392 14792 17398
rect 14740 17334 14792 17340
rect 14094 17295 14096 17304
rect 14148 17295 14150 17304
rect 14096 17266 14148 17272
rect 14188 17256 14240 17262
rect 14188 17198 14240 17204
rect 14200 16922 14228 17198
rect 14568 17058 14596 17334
rect 14752 17058 14780 17334
rect 14556 17052 14608 17058
rect 14556 16994 14608 17000
rect 14740 17052 14792 17058
rect 14740 16994 14792 17000
rect 14188 16916 14240 16922
rect 14188 16858 14240 16864
rect 14004 16848 14056 16854
rect 14002 16816 14004 16825
rect 14056 16816 14058 16825
rect 14002 16751 14058 16760
rect 13728 16712 13780 16718
rect 13728 16654 13780 16660
rect 13740 16310 13768 16654
rect 14200 16446 14228 16858
rect 14188 16440 14240 16446
rect 14188 16382 14240 16388
rect 13728 16304 13780 16310
rect 13728 16246 13780 16252
rect 13740 15902 13768 16246
rect 14200 15970 14228 16382
rect 14188 15964 14240 15970
rect 14188 15906 14240 15912
rect 13728 15896 13780 15902
rect 13728 15838 13780 15844
rect 13820 15692 13872 15698
rect 13820 15634 13872 15640
rect 13832 15426 13860 15634
rect 14200 15426 14228 15906
rect 14844 15766 14872 23182
rect 14956 22596 15252 22616
rect 15012 22594 15036 22596
rect 15092 22594 15116 22596
rect 15172 22594 15196 22596
rect 15034 22542 15036 22594
rect 15098 22542 15110 22594
rect 15172 22542 15174 22594
rect 15012 22540 15036 22542
rect 15092 22540 15116 22542
rect 15172 22540 15196 22542
rect 14956 22520 15252 22540
rect 14956 21508 15252 21528
rect 15012 21506 15036 21508
rect 15092 21506 15116 21508
rect 15172 21506 15196 21508
rect 15034 21454 15036 21506
rect 15098 21454 15110 21506
rect 15172 21454 15174 21506
rect 15012 21452 15036 21454
rect 15092 21452 15116 21454
rect 15172 21452 15196 21454
rect 14956 21432 15252 21452
rect 14956 20420 15252 20440
rect 15012 20418 15036 20420
rect 15092 20418 15116 20420
rect 15172 20418 15196 20420
rect 15034 20366 15036 20418
rect 15098 20366 15110 20418
rect 15172 20366 15174 20418
rect 15012 20364 15036 20366
rect 15092 20364 15116 20366
rect 15172 20364 15196 20366
rect 14956 20344 15252 20364
rect 14956 19332 15252 19352
rect 15012 19330 15036 19332
rect 15092 19330 15116 19332
rect 15172 19330 15196 19332
rect 15034 19278 15036 19330
rect 15098 19278 15110 19330
rect 15172 19278 15174 19330
rect 15012 19276 15036 19278
rect 15092 19276 15116 19278
rect 15172 19276 15196 19278
rect 14956 19256 15252 19276
rect 14956 18244 15252 18264
rect 15012 18242 15036 18244
rect 15092 18242 15116 18244
rect 15172 18242 15196 18244
rect 15034 18190 15036 18242
rect 15098 18190 15110 18242
rect 15172 18190 15174 18242
rect 15012 18188 15036 18190
rect 15092 18188 15116 18190
rect 15172 18188 15196 18190
rect 14956 18168 15252 18188
rect 15304 17534 15332 27240
rect 15948 24538 15976 27240
rect 15384 24532 15436 24538
rect 15384 24474 15436 24480
rect 15936 24532 15988 24538
rect 15936 24474 15988 24480
rect 15292 17528 15344 17534
rect 15292 17470 15344 17476
rect 15108 17460 15160 17466
rect 15108 17402 15160 17408
rect 15120 17346 15148 17402
rect 15120 17318 15332 17346
rect 14956 17156 15252 17176
rect 15012 17154 15036 17156
rect 15092 17154 15116 17156
rect 15172 17154 15196 17156
rect 15034 17102 15036 17154
rect 15098 17102 15110 17154
rect 15172 17102 15174 17154
rect 15012 17100 15036 17102
rect 15092 17100 15116 17102
rect 15172 17100 15196 17102
rect 14956 17080 15252 17100
rect 15108 16916 15160 16922
rect 15108 16858 15160 16864
rect 15120 16514 15148 16858
rect 15108 16508 15160 16514
rect 15108 16450 15160 16456
rect 14956 16068 15252 16088
rect 15012 16066 15036 16068
rect 15092 16066 15116 16068
rect 15172 16066 15196 16068
rect 15034 16014 15036 16066
rect 15098 16014 15110 16066
rect 15172 16014 15174 16066
rect 15012 16012 15036 16014
rect 15092 16012 15116 16014
rect 15172 16012 15196 16014
rect 14956 15992 15252 16012
rect 15304 15970 15332 17318
rect 15292 15964 15344 15970
rect 15292 15906 15344 15912
rect 14832 15760 14884 15766
rect 14832 15702 14884 15708
rect 13820 15420 13872 15426
rect 13820 15362 13872 15368
rect 14188 15420 14240 15426
rect 14188 15362 14240 15368
rect 14956 14980 15252 15000
rect 15012 14978 15036 14980
rect 15092 14978 15116 14980
rect 15172 14978 15196 14980
rect 15034 14926 15036 14978
rect 15098 14926 15110 14978
rect 15172 14926 15174 14978
rect 15012 14924 15036 14926
rect 15092 14924 15116 14926
rect 15172 14924 15196 14926
rect 14956 14904 15252 14924
rect 14956 13892 15252 13912
rect 15012 13890 15036 13892
rect 15092 13890 15116 13892
rect 15172 13890 15196 13892
rect 15034 13838 15036 13890
rect 15098 13838 15110 13890
rect 15172 13838 15174 13890
rect 15012 13836 15036 13838
rect 15092 13836 15116 13838
rect 15172 13836 15196 13838
rect 14956 13816 15252 13836
rect 15396 13794 15424 24474
rect 16212 23920 16264 23926
rect 16212 23862 16264 23868
rect 16028 23784 16080 23790
rect 16028 23726 16080 23732
rect 16040 23314 16068 23726
rect 16028 23308 16080 23314
rect 16028 23250 16080 23256
rect 15476 22832 15528 22838
rect 15476 22774 15528 22780
rect 15488 22498 15516 22774
rect 15568 22696 15620 22702
rect 15568 22638 15620 22644
rect 15476 22492 15528 22498
rect 15476 22434 15528 22440
rect 15488 21954 15516 22434
rect 15580 22294 15608 22638
rect 16040 22362 16068 23250
rect 16224 23042 16252 23862
rect 16488 23376 16540 23382
rect 16488 23318 16540 23324
rect 16212 23036 16264 23042
rect 16212 22978 16264 22984
rect 16120 22696 16172 22702
rect 16118 22664 16120 22673
rect 16172 22664 16174 22673
rect 16118 22599 16174 22608
rect 16224 22498 16252 22978
rect 16212 22492 16264 22498
rect 16212 22434 16264 22440
rect 16028 22356 16080 22362
rect 16028 22298 16080 22304
rect 15568 22288 15620 22294
rect 15568 22230 15620 22236
rect 15844 22288 15896 22294
rect 15844 22230 15896 22236
rect 15476 21948 15528 21954
rect 15476 21890 15528 21896
rect 15568 21812 15620 21818
rect 15568 21754 15620 21760
rect 15752 21812 15804 21818
rect 15752 21754 15804 21760
rect 15580 21070 15608 21754
rect 15764 21274 15792 21754
rect 15752 21268 15804 21274
rect 15752 21210 15804 21216
rect 15568 21064 15620 21070
rect 15568 21006 15620 21012
rect 15580 19982 15608 21006
rect 15568 19976 15620 19982
rect 15568 19918 15620 19924
rect 15476 19704 15528 19710
rect 15476 19646 15528 19652
rect 15488 19234 15516 19646
rect 15476 19228 15528 19234
rect 15476 19170 15528 19176
rect 15488 18690 15516 19170
rect 15476 18684 15528 18690
rect 15476 18626 15528 18632
rect 15856 17618 15884 22230
rect 16040 21954 16068 22298
rect 16500 22294 16528 23318
rect 16488 22288 16540 22294
rect 16488 22230 16540 22236
rect 16028 21948 16080 21954
rect 16028 21890 16080 21896
rect 16396 20724 16448 20730
rect 16132 20662 16160 20693
rect 16396 20666 16448 20672
rect 16120 20656 16172 20662
rect 16118 20624 16120 20633
rect 16172 20624 16174 20633
rect 16118 20559 16174 20568
rect 16132 20322 16160 20559
rect 16120 20316 16172 20322
rect 16120 20258 16172 20264
rect 16408 19438 16436 20666
rect 16488 20588 16540 20594
rect 16488 20530 16540 20536
rect 16500 20050 16528 20530
rect 16488 20044 16540 20050
rect 16488 19986 16540 19992
rect 16500 19778 16528 19986
rect 16488 19772 16540 19778
rect 16488 19714 16540 19720
rect 16396 19432 16448 19438
rect 16396 19374 16448 19380
rect 15936 18344 15988 18350
rect 15936 18286 15988 18292
rect 15948 17942 15976 18286
rect 15936 17936 15988 17942
rect 15936 17878 15988 17884
rect 16396 17936 16448 17942
rect 16396 17878 16448 17884
rect 15856 17590 15976 17618
rect 15752 17528 15804 17534
rect 15752 17470 15804 17476
rect 15660 15624 15712 15630
rect 15660 15566 15712 15572
rect 15672 15426 15700 15566
rect 15660 15420 15712 15426
rect 15660 15362 15712 15368
rect 15384 13788 15436 13794
rect 15384 13730 15436 13736
rect 15476 13584 15528 13590
rect 15476 13526 15528 13532
rect 13636 13244 13688 13250
rect 13636 13186 13688 13192
rect 13452 13108 13504 13114
rect 13452 13050 13504 13056
rect 13464 12706 13492 13050
rect 14956 12804 15252 12824
rect 15012 12802 15036 12804
rect 15092 12802 15116 12804
rect 15172 12802 15196 12804
rect 15034 12750 15036 12802
rect 15098 12750 15110 12802
rect 15172 12750 15174 12802
rect 15012 12748 15036 12750
rect 15092 12748 15116 12750
rect 15172 12748 15196 12750
rect 14956 12728 15252 12748
rect 13452 12700 13504 12706
rect 13452 12642 13504 12648
rect 15488 12570 15516 13526
rect 15476 12564 15528 12570
rect 15476 12506 15528 12512
rect 12532 12496 12584 12502
rect 12532 12438 12584 12444
rect 15660 12496 15712 12502
rect 15660 12438 15712 12444
rect 12544 12162 12572 12438
rect 15672 12162 15700 12438
rect 12532 12156 12584 12162
rect 12532 12098 12584 12104
rect 15660 12156 15712 12162
rect 15660 12098 15712 12104
rect 13268 12020 13320 12026
rect 13268 11962 13320 11968
rect 12716 11816 12768 11822
rect 12716 11758 12768 11764
rect 12728 11414 12756 11758
rect 12716 11408 12768 11414
rect 12716 11350 12768 11356
rect 12440 11340 12492 11346
rect 12440 11282 12492 11288
rect 10289 11172 10585 11192
rect 10345 11170 10369 11172
rect 10425 11170 10449 11172
rect 10505 11170 10529 11172
rect 10367 11118 10369 11170
rect 10431 11118 10443 11170
rect 10505 11118 10507 11170
rect 10345 11116 10369 11118
rect 10425 11116 10449 11118
rect 10505 11116 10529 11118
rect 10289 11096 10585 11116
rect 5622 10628 5918 10648
rect 5678 10626 5702 10628
rect 5758 10626 5782 10628
rect 5838 10626 5862 10628
rect 5700 10574 5702 10626
rect 5764 10574 5776 10626
rect 5838 10574 5840 10626
rect 5678 10572 5702 10574
rect 5758 10572 5782 10574
rect 5838 10572 5862 10574
rect 5622 10552 5918 10572
rect 12452 10326 12480 11282
rect 12728 10530 12756 11350
rect 13280 11074 13308 11962
rect 13636 11952 13688 11958
rect 13636 11894 13688 11900
rect 14004 11952 14056 11958
rect 14004 11894 14056 11900
rect 13648 11074 13676 11894
rect 14016 11278 14044 11894
rect 14956 11716 15252 11736
rect 15012 11714 15036 11716
rect 15092 11714 15116 11716
rect 15172 11714 15196 11716
rect 15034 11662 15036 11714
rect 15098 11662 15110 11714
rect 15172 11662 15174 11714
rect 15012 11660 15036 11662
rect 15092 11660 15116 11662
rect 15172 11660 15196 11662
rect 14956 11640 15252 11660
rect 14556 11408 14608 11414
rect 14556 11350 14608 11356
rect 14004 11272 14056 11278
rect 14004 11214 14056 11220
rect 13268 11068 13320 11074
rect 13268 11010 13320 11016
rect 13636 11068 13688 11074
rect 13636 11010 13688 11016
rect 13648 10530 13676 11010
rect 14016 10938 14044 11214
rect 14004 10932 14056 10938
rect 14004 10874 14056 10880
rect 14464 10728 14516 10734
rect 14568 10682 14596 11350
rect 14740 11272 14792 11278
rect 14740 11214 14792 11220
rect 14752 11074 14780 11214
rect 14740 11068 14792 11074
rect 14740 11010 14792 11016
rect 14832 10932 14884 10938
rect 14832 10874 14884 10880
rect 14516 10676 14596 10682
rect 14464 10670 14596 10676
rect 14476 10654 14596 10670
rect 14568 10530 14596 10654
rect 14844 10530 14872 10874
rect 14956 10628 15252 10648
rect 15012 10626 15036 10628
rect 15092 10626 15116 10628
rect 15172 10626 15196 10628
rect 15034 10574 15036 10626
rect 15098 10574 15110 10626
rect 15172 10574 15174 10626
rect 15012 10572 15036 10574
rect 15092 10572 15116 10574
rect 15172 10572 15196 10574
rect 14956 10552 15252 10572
rect 12716 10524 12768 10530
rect 12716 10466 12768 10472
rect 13636 10524 13688 10530
rect 13636 10466 13688 10472
rect 14556 10524 14608 10530
rect 14556 10466 14608 10472
rect 14832 10524 14884 10530
rect 14832 10466 14884 10472
rect 10968 10320 11020 10326
rect 3422 10288 3478 10297
rect 3422 10223 3478 10232
rect 10782 10288 10838 10297
rect 10968 10262 11020 10268
rect 12440 10320 12492 10326
rect 12440 10262 12492 10268
rect 13818 10288 13874 10297
rect 10782 10223 10784 10232
rect 202 9744 258 9753
rect 202 9679 258 9688
rect 3436 6761 3464 10223
rect 10836 10223 10838 10232
rect 10784 10194 10836 10200
rect 10289 10084 10585 10104
rect 10345 10082 10369 10084
rect 10425 10082 10449 10084
rect 10505 10082 10529 10084
rect 10367 10030 10369 10082
rect 10431 10030 10443 10082
rect 10505 10030 10507 10082
rect 10345 10028 10369 10030
rect 10425 10028 10449 10030
rect 10505 10028 10529 10030
rect 10289 10008 10585 10028
rect 10980 9986 11008 10262
rect 13818 10223 13820 10232
rect 13872 10223 13874 10232
rect 13912 10252 13964 10258
rect 13820 10194 13872 10200
rect 13912 10194 13964 10200
rect 13924 9986 13952 10194
rect 10968 9980 11020 9986
rect 10968 9922 11020 9928
rect 13912 9980 13964 9986
rect 13912 9922 13964 9928
rect 13924 9753 13952 9922
rect 13910 9744 13966 9753
rect 13910 9679 13966 9688
rect 5622 9540 5918 9560
rect 5678 9538 5702 9540
rect 5758 9538 5782 9540
rect 5838 9538 5862 9540
rect 5700 9486 5702 9538
rect 5764 9486 5776 9538
rect 5838 9486 5840 9538
rect 5678 9484 5702 9486
rect 5758 9484 5782 9486
rect 5838 9484 5862 9486
rect 5622 9464 5918 9484
rect 14956 9540 15252 9560
rect 15012 9538 15036 9540
rect 15092 9538 15116 9540
rect 15172 9538 15196 9540
rect 15034 9486 15036 9538
rect 15098 9486 15110 9538
rect 15172 9486 15174 9538
rect 15012 9484 15036 9486
rect 15092 9484 15116 9486
rect 15172 9484 15196 9486
rect 14956 9464 15252 9484
rect 10289 8996 10585 9016
rect 10345 8994 10369 8996
rect 10425 8994 10449 8996
rect 10505 8994 10529 8996
rect 10367 8942 10369 8994
rect 10431 8942 10443 8994
rect 10505 8942 10507 8994
rect 10345 8940 10369 8942
rect 10425 8940 10449 8942
rect 10505 8940 10529 8942
rect 10289 8920 10585 8940
rect 5622 8452 5918 8472
rect 5678 8450 5702 8452
rect 5758 8450 5782 8452
rect 5838 8450 5862 8452
rect 5700 8398 5702 8450
rect 5764 8398 5776 8450
rect 5838 8398 5840 8450
rect 5678 8396 5702 8398
rect 5758 8396 5782 8398
rect 5838 8396 5862 8398
rect 5622 8376 5918 8396
rect 14956 8452 15252 8472
rect 15012 8450 15036 8452
rect 15092 8450 15116 8452
rect 15172 8450 15196 8452
rect 15034 8398 15036 8450
rect 15098 8398 15110 8450
rect 15172 8398 15174 8450
rect 15012 8396 15036 8398
rect 15092 8396 15116 8398
rect 15172 8396 15196 8398
rect 14956 8376 15252 8396
rect 10289 7908 10585 7928
rect 10345 7906 10369 7908
rect 10425 7906 10449 7908
rect 10505 7906 10529 7908
rect 10367 7854 10369 7906
rect 10431 7854 10443 7906
rect 10505 7854 10507 7906
rect 10345 7852 10369 7854
rect 10425 7852 10449 7854
rect 10505 7852 10529 7854
rect 10289 7832 10585 7852
rect 5622 7364 5918 7384
rect 5678 7362 5702 7364
rect 5758 7362 5782 7364
rect 5838 7362 5862 7364
rect 5700 7310 5702 7362
rect 5764 7310 5776 7362
rect 5838 7310 5840 7362
rect 5678 7308 5702 7310
rect 5758 7308 5782 7310
rect 5838 7308 5862 7310
rect 5622 7288 5918 7308
rect 14956 7364 15252 7384
rect 15012 7362 15036 7364
rect 15092 7362 15116 7364
rect 15172 7362 15196 7364
rect 15034 7310 15036 7362
rect 15098 7310 15110 7362
rect 15172 7310 15174 7362
rect 15012 7308 15036 7310
rect 15092 7308 15116 7310
rect 15172 7308 15196 7310
rect 14956 7288 15252 7308
rect 10289 6820 10585 6840
rect 10345 6818 10369 6820
rect 10425 6818 10449 6820
rect 10505 6818 10529 6820
rect 10367 6766 10369 6818
rect 10431 6766 10443 6818
rect 10505 6766 10507 6818
rect 10345 6764 10369 6766
rect 10425 6764 10449 6766
rect 10505 6764 10529 6766
rect 3422 6752 3478 6761
rect 10289 6744 10585 6764
rect 3422 6687 3478 6696
rect 5622 6276 5918 6296
rect 5678 6274 5702 6276
rect 5758 6274 5782 6276
rect 5838 6274 5862 6276
rect 5700 6222 5702 6274
rect 5764 6222 5776 6274
rect 5838 6222 5840 6274
rect 5678 6220 5702 6222
rect 5758 6220 5782 6222
rect 5838 6220 5862 6222
rect 5622 6200 5918 6220
rect 14956 6276 15252 6296
rect 15012 6274 15036 6276
rect 15092 6274 15116 6276
rect 15172 6274 15196 6276
rect 15034 6222 15036 6274
rect 15098 6222 15110 6274
rect 15172 6222 15174 6274
rect 15012 6220 15036 6222
rect 15092 6220 15116 6222
rect 15172 6220 15196 6222
rect 14956 6200 15252 6220
rect 10289 5732 10585 5752
rect 10345 5730 10369 5732
rect 10425 5730 10449 5732
rect 10505 5730 10529 5732
rect 10367 5678 10369 5730
rect 10431 5678 10443 5730
rect 10505 5678 10507 5730
rect 10345 5676 10369 5678
rect 10425 5676 10449 5678
rect 10505 5676 10529 5678
rect 10289 5656 10585 5676
rect 5622 5188 5918 5208
rect 5678 5186 5702 5188
rect 5758 5186 5782 5188
rect 5838 5186 5862 5188
rect 5700 5134 5702 5186
rect 5764 5134 5776 5186
rect 5838 5134 5840 5186
rect 5678 5132 5702 5134
rect 5758 5132 5782 5134
rect 5838 5132 5862 5134
rect 5622 5112 5918 5132
rect 14956 5188 15252 5208
rect 15012 5186 15036 5188
rect 15092 5186 15116 5188
rect 15172 5186 15196 5188
rect 15034 5134 15036 5186
rect 15098 5134 15110 5186
rect 15172 5134 15174 5186
rect 15012 5132 15036 5134
rect 15092 5132 15116 5134
rect 15172 5132 15196 5134
rect 14956 5112 15252 5132
rect 15764 5090 15792 17470
rect 15844 17460 15896 17466
rect 15844 17402 15896 17408
rect 15856 16446 15884 17402
rect 15948 16825 15976 17590
rect 16212 17460 16264 17466
rect 16212 17402 16264 17408
rect 15934 16816 15990 16825
rect 15934 16751 15990 16760
rect 16224 16514 16252 17402
rect 16408 17398 16436 17878
rect 16396 17392 16448 17398
rect 16396 17334 16448 17340
rect 16408 17058 16436 17334
rect 16396 17052 16448 17058
rect 16396 16994 16448 17000
rect 16408 16514 16436 16994
rect 16212 16508 16264 16514
rect 16212 16450 16264 16456
rect 16396 16508 16448 16514
rect 16396 16450 16448 16456
rect 15844 16440 15896 16446
rect 15842 16408 15844 16417
rect 15896 16408 15898 16417
rect 15842 16343 15898 16352
rect 16394 16272 16450 16281
rect 16394 16207 16450 16216
rect 15844 15828 15896 15834
rect 15844 15770 15896 15776
rect 15856 15358 15884 15770
rect 16304 15760 16356 15766
rect 16302 15728 16304 15737
rect 16356 15728 16358 15737
rect 16302 15663 16358 15672
rect 16408 15426 16436 16207
rect 16396 15420 16448 15426
rect 16396 15362 16448 15368
rect 15844 15352 15896 15358
rect 15844 15294 15896 15300
rect 16396 15284 16448 15290
rect 16396 15226 16448 15232
rect 16028 14604 16080 14610
rect 16028 14546 16080 14552
rect 16040 14066 16068 14546
rect 16408 14338 16436 15226
rect 16396 14332 16448 14338
rect 16396 14274 16448 14280
rect 16120 14196 16172 14202
rect 16120 14138 16172 14144
rect 16028 14060 16080 14066
rect 16028 14002 16080 14008
rect 16132 13794 16160 14138
rect 16120 13788 16172 13794
rect 16120 13730 16172 13736
rect 16028 12020 16080 12026
rect 16028 11962 16080 11968
rect 15936 11952 15988 11958
rect 15936 11894 15988 11900
rect 15948 9986 15976 11894
rect 16040 11074 16068 11962
rect 16396 11952 16448 11958
rect 16396 11894 16448 11900
rect 16304 11408 16356 11414
rect 16304 11350 16356 11356
rect 16028 11068 16080 11074
rect 16028 11010 16080 11016
rect 16316 10326 16344 11350
rect 16408 11278 16436 11894
rect 16488 11340 16540 11346
rect 16488 11282 16540 11288
rect 16396 11272 16448 11278
rect 16396 11214 16448 11220
rect 16408 11006 16436 11214
rect 16396 11000 16448 11006
rect 16396 10942 16448 10948
rect 16408 10530 16436 10942
rect 16396 10524 16448 10530
rect 16396 10466 16448 10472
rect 16304 10320 16356 10326
rect 16304 10262 16356 10268
rect 16396 10252 16448 10258
rect 16396 10194 16448 10200
rect 15936 9980 15988 9986
rect 15936 9922 15988 9928
rect 16028 9844 16080 9850
rect 16028 9786 16080 9792
rect 16040 9102 16068 9786
rect 16408 9782 16436 10194
rect 16500 9782 16528 11282
rect 16396 9776 16448 9782
rect 16396 9718 16448 9724
rect 16488 9776 16540 9782
rect 16488 9718 16540 9724
rect 16408 9481 16436 9718
rect 16394 9472 16450 9481
rect 16500 9442 16528 9718
rect 16394 9407 16396 9416
rect 16448 9407 16450 9416
rect 16488 9436 16540 9442
rect 16396 9378 16448 9384
rect 16488 9378 16540 9384
rect 16028 9096 16080 9102
rect 16028 9038 16080 9044
rect 16040 5401 16068 9038
rect 16592 6602 16620 27240
rect 17224 23240 17276 23246
rect 17224 23182 17276 23188
rect 17236 22770 17264 23182
rect 17224 22764 17276 22770
rect 17224 22706 17276 22712
rect 17236 22226 17264 22706
rect 17224 22220 17276 22226
rect 17224 22162 17276 22168
rect 16856 21064 16908 21070
rect 16856 21006 16908 21012
rect 17132 21064 17184 21070
rect 17132 21006 17184 21012
rect 16868 19030 16896 21006
rect 17144 20866 17172 21006
rect 17132 20860 17184 20866
rect 17132 20802 17184 20808
rect 17040 19432 17092 19438
rect 17040 19374 17092 19380
rect 16856 19024 16908 19030
rect 16856 18966 16908 18972
rect 17052 18729 17080 19374
rect 17038 18720 17094 18729
rect 17038 18655 17094 18664
rect 17052 17466 17080 18655
rect 17328 18434 17356 27240
rect 17684 21268 17736 21274
rect 17684 21210 17736 21216
rect 17696 20322 17724 21210
rect 17684 20316 17736 20322
rect 17684 20258 17736 20264
rect 17590 19944 17646 19953
rect 17590 19879 17646 19888
rect 17236 18406 17356 18434
rect 17040 17460 17092 17466
rect 17040 17402 17092 17408
rect 17040 16848 17092 16854
rect 17040 16790 17092 16796
rect 16856 15284 16908 15290
rect 16856 15226 16908 15232
rect 16868 14270 16896 15226
rect 16948 15216 17000 15222
rect 16946 15184 16948 15193
rect 17000 15184 17002 15193
rect 16946 15119 17002 15128
rect 16960 14882 16988 15119
rect 16948 14876 17000 14882
rect 16948 14818 17000 14824
rect 17052 14354 17080 16790
rect 17130 15864 17186 15873
rect 17130 15799 17132 15808
rect 17184 15799 17186 15808
rect 17132 15770 17184 15776
rect 16960 14326 17080 14354
rect 16856 14264 16908 14270
rect 16856 14206 16908 14212
rect 16868 13794 16896 14206
rect 16960 14134 16988 14326
rect 16948 14128 17000 14134
rect 16948 14070 17000 14076
rect 16960 13833 16988 14070
rect 16946 13824 17002 13833
rect 16856 13788 16908 13794
rect 16946 13759 17002 13768
rect 16856 13730 16908 13736
rect 16960 13726 16988 13759
rect 16948 13720 17000 13726
rect 16948 13662 17000 13668
rect 17236 13250 17264 18406
rect 17316 18344 17368 18350
rect 17316 18286 17368 18292
rect 17328 17806 17356 18286
rect 17316 17800 17368 17806
rect 17316 17742 17368 17748
rect 17328 17058 17356 17742
rect 17316 17052 17368 17058
rect 17316 16994 17368 17000
rect 17604 16990 17632 19879
rect 17776 17256 17828 17262
rect 17776 17198 17828 17204
rect 17788 17058 17816 17198
rect 17776 17052 17828 17058
rect 17776 16994 17828 17000
rect 17592 16984 17644 16990
rect 17592 16926 17644 16932
rect 17868 16780 17920 16786
rect 17868 16722 17920 16728
rect 17776 16712 17828 16718
rect 17776 16654 17828 16660
rect 17788 16446 17816 16654
rect 17880 16514 17908 16722
rect 17868 16508 17920 16514
rect 17868 16450 17920 16456
rect 17684 16440 17736 16446
rect 17684 16382 17736 16388
rect 17776 16440 17828 16446
rect 17776 16382 17828 16388
rect 17696 15698 17724 16382
rect 17684 15692 17736 15698
rect 17684 15634 17736 15640
rect 17316 15624 17368 15630
rect 17316 15566 17368 15572
rect 17328 14338 17356 15566
rect 17316 14332 17368 14338
rect 17316 14274 17368 14280
rect 17328 13658 17356 14274
rect 17776 14128 17828 14134
rect 17776 14070 17828 14076
rect 17788 13697 17816 14070
rect 17774 13688 17830 13697
rect 17316 13652 17368 13658
rect 17774 13623 17776 13632
rect 17316 13594 17368 13600
rect 17828 13623 17830 13632
rect 17776 13594 17828 13600
rect 17500 13584 17552 13590
rect 17498 13552 17500 13561
rect 17552 13552 17554 13561
rect 17498 13487 17554 13496
rect 17788 13250 17816 13594
rect 17224 13244 17276 13250
rect 17224 13186 17276 13192
rect 17776 13244 17828 13250
rect 17776 13186 17828 13192
rect 16764 13108 16816 13114
rect 16764 13050 16816 13056
rect 16776 12570 16804 13050
rect 16764 12564 16816 12570
rect 16764 12506 16816 12512
rect 16856 10524 16908 10530
rect 16856 10466 16908 10472
rect 16868 10326 16896 10466
rect 16856 10320 16908 10326
rect 16856 10262 16908 10268
rect 17972 7282 18000 27240
rect 18708 27138 18736 27240
rect 18340 27110 18736 27138
rect 18052 23308 18104 23314
rect 18052 23250 18104 23256
rect 18064 22294 18092 23250
rect 18340 22378 18368 27110
rect 19352 24470 19380 27240
rect 19622 25316 19918 25336
rect 19678 25314 19702 25316
rect 19758 25314 19782 25316
rect 19838 25314 19862 25316
rect 19700 25262 19702 25314
rect 19764 25262 19776 25314
rect 19838 25262 19840 25314
rect 19678 25260 19702 25262
rect 19758 25260 19782 25262
rect 19838 25260 19862 25262
rect 19622 25240 19918 25260
rect 19340 24464 19392 24470
rect 19340 24406 19392 24412
rect 19156 24328 19208 24334
rect 19156 24270 19208 24276
rect 19168 23994 19196 24270
rect 19622 24228 19918 24248
rect 19678 24226 19702 24228
rect 19758 24226 19782 24228
rect 19838 24226 19862 24228
rect 19700 24174 19702 24226
rect 19764 24174 19776 24226
rect 19838 24174 19840 24226
rect 19678 24172 19702 24174
rect 19758 24172 19782 24174
rect 19838 24172 19862 24174
rect 19622 24152 19918 24172
rect 19156 23988 19208 23994
rect 19156 23930 19208 23936
rect 18420 23784 18472 23790
rect 18420 23726 18472 23732
rect 18604 23784 18656 23790
rect 18604 23726 18656 23732
rect 18432 23382 18460 23726
rect 18420 23376 18472 23382
rect 18420 23318 18472 23324
rect 18432 22770 18460 23318
rect 18616 23042 18644 23726
rect 19064 23308 19116 23314
rect 19064 23250 19116 23256
rect 18604 23036 18656 23042
rect 18604 22978 18656 22984
rect 18788 22968 18840 22974
rect 18510 22936 18566 22945
rect 18788 22910 18840 22916
rect 18510 22871 18512 22880
rect 18564 22871 18566 22880
rect 18512 22842 18564 22848
rect 18420 22764 18472 22770
rect 18420 22706 18472 22712
rect 18432 22498 18460 22706
rect 18420 22492 18472 22498
rect 18420 22434 18472 22440
rect 18524 22430 18552 22842
rect 18512 22424 18564 22430
rect 18340 22350 18460 22378
rect 18512 22366 18564 22372
rect 18052 22288 18104 22294
rect 18052 22230 18104 22236
rect 18326 21848 18382 21857
rect 18052 21812 18104 21818
rect 18326 21783 18328 21792
rect 18052 21754 18104 21760
rect 18380 21783 18382 21792
rect 18328 21754 18380 21760
rect 18064 21342 18092 21754
rect 18052 21336 18104 21342
rect 18052 21278 18104 21284
rect 18064 20866 18092 21278
rect 18328 21064 18380 21070
rect 18328 21006 18380 21012
rect 18052 20860 18104 20866
rect 18052 20802 18104 20808
rect 18052 19976 18104 19982
rect 18052 19918 18104 19924
rect 18064 18486 18092 19918
rect 18052 18480 18104 18486
rect 18052 18422 18104 18428
rect 18064 17874 18092 18422
rect 18052 17868 18104 17874
rect 18052 17810 18104 17816
rect 18052 16508 18104 16514
rect 18052 16450 18104 16456
rect 18064 16417 18092 16450
rect 18050 16408 18106 16417
rect 18050 16343 18106 16352
rect 18236 15760 18288 15766
rect 18340 15737 18368 21006
rect 18236 15702 18288 15708
rect 18326 15728 18382 15737
rect 18248 15426 18276 15702
rect 18326 15663 18382 15672
rect 18236 15420 18288 15426
rect 18236 15362 18288 15368
rect 18248 14762 18276 15362
rect 18248 14734 18368 14762
rect 18340 14678 18368 14734
rect 18328 14672 18380 14678
rect 18328 14614 18380 14620
rect 18328 12360 18380 12366
rect 18328 12302 18380 12308
rect 18236 11952 18288 11958
rect 18236 11894 18288 11900
rect 18248 11550 18276 11894
rect 18340 11618 18368 12302
rect 18328 11612 18380 11618
rect 18328 11554 18380 11560
rect 18236 11544 18288 11550
rect 18236 11486 18288 11492
rect 18432 7577 18460 22350
rect 18800 21954 18828 22910
rect 19076 22906 19104 23250
rect 19168 23042 19196 23930
rect 19432 23920 19484 23926
rect 19430 23888 19432 23897
rect 19484 23888 19486 23897
rect 19430 23823 19486 23832
rect 19340 23784 19392 23790
rect 19340 23726 19392 23732
rect 19248 23580 19300 23586
rect 19248 23522 19300 23528
rect 19156 23036 19208 23042
rect 19156 22978 19208 22984
rect 19260 22974 19288 23522
rect 19248 22968 19300 22974
rect 19248 22910 19300 22916
rect 19064 22900 19116 22906
rect 19064 22842 19116 22848
rect 19352 22294 19380 23726
rect 19444 23518 19472 23823
rect 19432 23512 19484 23518
rect 19432 23454 19484 23460
rect 19444 23042 19472 23454
rect 19622 23140 19918 23160
rect 19678 23138 19702 23140
rect 19758 23138 19782 23140
rect 19838 23138 19862 23140
rect 19700 23086 19702 23138
rect 19764 23086 19776 23138
rect 19838 23086 19840 23138
rect 19678 23084 19702 23086
rect 19758 23084 19782 23086
rect 19838 23084 19862 23086
rect 19622 23064 19918 23084
rect 19432 23036 19484 23042
rect 19432 22978 19484 22984
rect 19798 22936 19854 22945
rect 19798 22871 19854 22880
rect 19812 22362 19840 22871
rect 19800 22356 19852 22362
rect 19800 22298 19852 22304
rect 19340 22288 19392 22294
rect 19340 22230 19392 22236
rect 19352 21954 19380 22230
rect 19622 22052 19918 22072
rect 19678 22050 19702 22052
rect 19758 22050 19782 22052
rect 19838 22050 19862 22052
rect 19700 21998 19702 22050
rect 19764 21998 19776 22050
rect 19838 21998 19840 22050
rect 19678 21996 19702 21998
rect 19758 21996 19782 21998
rect 19838 21996 19862 21998
rect 19622 21976 19918 21996
rect 18788 21948 18840 21954
rect 18788 21890 18840 21896
rect 19340 21948 19392 21954
rect 19340 21890 19392 21896
rect 18694 21168 18750 21177
rect 18694 21103 18696 21112
rect 18748 21103 18750 21112
rect 18696 21074 18748 21080
rect 18696 20656 18748 20662
rect 18696 20598 18748 20604
rect 18512 20044 18564 20050
rect 18512 19986 18564 19992
rect 18524 19778 18552 19986
rect 18708 19982 18736 20598
rect 18696 19976 18748 19982
rect 18696 19918 18748 19924
rect 18512 19772 18564 19778
rect 18512 19714 18564 19720
rect 18800 17466 18828 21890
rect 19246 21712 19302 21721
rect 19246 21647 19248 21656
rect 19300 21647 19302 21656
rect 19248 21618 19300 21624
rect 19260 21274 19288 21618
rect 19248 21268 19300 21274
rect 19248 21210 19300 21216
rect 19156 21200 19208 21206
rect 19156 21142 19208 21148
rect 19168 21070 19196 21142
rect 18880 21064 18932 21070
rect 18880 21006 18932 21012
rect 19156 21064 19208 21070
rect 19156 21006 19208 21012
rect 18892 20866 18920 21006
rect 18880 20860 18932 20866
rect 18880 20802 18932 20808
rect 19260 20798 19288 21210
rect 19622 20964 19918 20984
rect 19678 20962 19702 20964
rect 19758 20962 19782 20964
rect 19838 20962 19862 20964
rect 19700 20910 19702 20962
rect 19764 20910 19776 20962
rect 19838 20910 19840 20962
rect 19678 20908 19702 20910
rect 19758 20908 19782 20910
rect 19838 20908 19862 20910
rect 19430 20896 19486 20905
rect 19340 20860 19392 20866
rect 19622 20888 19918 20908
rect 19430 20831 19432 20840
rect 19340 20802 19392 20808
rect 19484 20831 19486 20840
rect 19432 20802 19484 20808
rect 19248 20792 19300 20798
rect 19248 20734 19300 20740
rect 19352 20186 19380 20802
rect 19340 20180 19392 20186
rect 19444 20168 19472 20802
rect 19524 20180 19576 20186
rect 19444 20140 19524 20168
rect 19340 20122 19392 20128
rect 19524 20122 19576 20128
rect 18972 19976 19024 19982
rect 18972 19918 19024 19924
rect 18984 19642 19012 19918
rect 19622 19876 19918 19896
rect 19678 19874 19702 19876
rect 19758 19874 19782 19876
rect 19838 19874 19862 19876
rect 19700 19822 19702 19874
rect 19764 19822 19776 19874
rect 19838 19822 19840 19874
rect 19678 19820 19702 19822
rect 19758 19820 19782 19822
rect 19838 19820 19862 19822
rect 19622 19800 19918 19820
rect 19798 19672 19854 19681
rect 18972 19636 19024 19642
rect 18972 19578 19024 19584
rect 19524 19636 19576 19642
rect 19798 19607 19800 19616
rect 19524 19578 19576 19584
rect 19852 19607 19854 19616
rect 19800 19578 19852 19584
rect 19340 19432 19392 19438
rect 19340 19374 19392 19380
rect 19352 18894 19380 19374
rect 19536 19234 19564 19578
rect 19524 19228 19576 19234
rect 19524 19170 19576 19176
rect 19524 19024 19576 19030
rect 19524 18966 19576 18972
rect 19064 18888 19116 18894
rect 19064 18830 19116 18836
rect 19248 18888 19300 18894
rect 19340 18888 19392 18894
rect 19248 18830 19300 18836
rect 19338 18856 19340 18865
rect 19392 18856 19394 18865
rect 19076 18593 19104 18830
rect 19062 18584 19118 18593
rect 19062 18519 19118 18528
rect 19260 18457 19288 18830
rect 19338 18791 19394 18800
rect 19246 18448 19302 18457
rect 19246 18383 19302 18392
rect 19248 18344 19300 18350
rect 19248 18286 19300 18292
rect 19260 17874 19288 18286
rect 19536 18146 19564 18966
rect 19622 18788 19918 18808
rect 19678 18786 19702 18788
rect 19758 18786 19782 18788
rect 19838 18786 19862 18788
rect 19700 18734 19702 18786
rect 19764 18734 19776 18786
rect 19838 18734 19840 18786
rect 19678 18732 19702 18734
rect 19758 18732 19782 18734
rect 19838 18732 19862 18734
rect 19622 18712 19918 18732
rect 19524 18140 19576 18146
rect 19524 18082 19576 18088
rect 19248 17868 19300 17874
rect 19248 17810 19300 17816
rect 19156 17596 19208 17602
rect 19156 17538 19208 17544
rect 18788 17460 18840 17466
rect 18788 17402 18840 17408
rect 18512 17256 18564 17262
rect 18512 17198 18564 17204
rect 18524 16514 18552 17198
rect 18800 16718 18828 17402
rect 19168 17058 19196 17538
rect 19260 17466 19288 17810
rect 19536 17534 19564 18082
rect 19622 17700 19918 17720
rect 19678 17698 19702 17700
rect 19758 17698 19782 17700
rect 19838 17698 19862 17700
rect 19700 17646 19702 17698
rect 19764 17646 19776 17698
rect 19838 17646 19840 17698
rect 19678 17644 19702 17646
rect 19758 17644 19782 17646
rect 19838 17644 19862 17646
rect 19622 17624 19918 17644
rect 19524 17528 19576 17534
rect 19524 17470 19576 17476
rect 19248 17460 19300 17466
rect 19248 17402 19300 17408
rect 19156 17052 19208 17058
rect 19156 16994 19208 17000
rect 18788 16712 18840 16718
rect 18788 16654 18840 16660
rect 18512 16508 18564 16514
rect 18512 16450 18564 16456
rect 18524 15970 18552 16450
rect 18604 16304 18656 16310
rect 18604 16246 18656 16252
rect 18512 15964 18564 15970
rect 18512 15906 18564 15912
rect 18616 15902 18644 16246
rect 18604 15896 18656 15902
rect 18604 15838 18656 15844
rect 18800 13561 18828 16654
rect 19064 16440 19116 16446
rect 19064 16382 19116 16388
rect 19076 15970 19104 16382
rect 19260 16310 19288 17402
rect 19622 16612 19918 16632
rect 19678 16610 19702 16612
rect 19758 16610 19782 16612
rect 19838 16610 19862 16612
rect 19700 16558 19702 16610
rect 19764 16558 19776 16610
rect 19838 16558 19840 16610
rect 19678 16556 19702 16558
rect 19758 16556 19782 16558
rect 19838 16556 19862 16558
rect 19622 16536 19918 16556
rect 19248 16304 19300 16310
rect 19248 16246 19300 16252
rect 19064 15964 19116 15970
rect 19064 15906 19116 15912
rect 19622 15524 19918 15544
rect 19678 15522 19702 15524
rect 19758 15522 19782 15524
rect 19838 15522 19862 15524
rect 19700 15470 19702 15522
rect 19764 15470 19776 15522
rect 19838 15470 19840 15522
rect 19678 15468 19702 15470
rect 19758 15468 19782 15470
rect 19838 15468 19862 15470
rect 19622 15448 19918 15468
rect 19156 15216 19208 15222
rect 19154 15184 19156 15193
rect 19208 15184 19210 15193
rect 19154 15119 19210 15128
rect 19168 14610 19196 15119
rect 19156 14604 19208 14610
rect 19156 14546 19208 14552
rect 19168 14338 19196 14546
rect 19340 14536 19392 14542
rect 19340 14478 19392 14484
rect 19156 14332 19208 14338
rect 19156 14274 19208 14280
rect 19352 13697 19380 14478
rect 19622 14436 19918 14456
rect 19678 14434 19702 14436
rect 19758 14434 19782 14436
rect 19838 14434 19862 14436
rect 19700 14382 19702 14434
rect 19764 14382 19776 14434
rect 19838 14382 19840 14434
rect 19678 14380 19702 14382
rect 19758 14380 19782 14382
rect 19838 14380 19862 14382
rect 19622 14360 19918 14380
rect 19338 13688 19394 13697
rect 19338 13623 19394 13632
rect 18786 13552 18842 13561
rect 18786 13487 18842 13496
rect 19622 13348 19918 13368
rect 19678 13346 19702 13348
rect 19758 13346 19782 13348
rect 19838 13346 19862 13348
rect 19700 13294 19702 13346
rect 19764 13294 19776 13346
rect 19838 13294 19840 13346
rect 19678 13292 19702 13294
rect 19758 13292 19782 13294
rect 19838 13292 19862 13294
rect 19622 13272 19918 13292
rect 19984 12360 20036 12366
rect 19984 12302 20036 12308
rect 19622 12260 19918 12280
rect 19678 12258 19702 12260
rect 19758 12258 19782 12260
rect 19838 12258 19862 12260
rect 19700 12206 19702 12258
rect 19764 12206 19776 12258
rect 19838 12206 19840 12258
rect 19678 12204 19702 12206
rect 19758 12204 19782 12206
rect 19838 12204 19862 12206
rect 19622 12184 19918 12204
rect 19996 12026 20024 12302
rect 19984 12020 20036 12026
rect 19984 11962 20036 11968
rect 18788 11816 18840 11822
rect 18788 11758 18840 11764
rect 18800 11482 18828 11758
rect 19996 11618 20024 11962
rect 19984 11612 20036 11618
rect 19984 11554 20036 11560
rect 18788 11476 18840 11482
rect 18788 11418 18840 11424
rect 18512 10932 18564 10938
rect 18512 10874 18564 10880
rect 18696 10932 18748 10938
rect 18696 10874 18748 10880
rect 18524 10841 18552 10874
rect 18510 10832 18566 10841
rect 18510 10767 18566 10776
rect 18708 10258 18736 10874
rect 18696 10252 18748 10258
rect 18696 10194 18748 10200
rect 18800 9986 18828 11418
rect 18880 11340 18932 11346
rect 18880 11282 18932 11288
rect 18892 11074 18920 11282
rect 19524 11272 19576 11278
rect 19524 11214 19576 11220
rect 18880 11068 18932 11074
rect 18880 11010 18932 11016
rect 18878 10832 18934 10841
rect 18878 10767 18934 10776
rect 18892 10530 18920 10767
rect 18880 10524 18932 10530
rect 18880 10466 18932 10472
rect 19248 10184 19300 10190
rect 19248 10126 19300 10132
rect 19260 10002 19288 10126
rect 18788 9980 18840 9986
rect 18788 9922 18840 9928
rect 19156 9980 19208 9986
rect 19260 9974 19472 10002
rect 19536 9986 19564 11214
rect 19622 11172 19918 11192
rect 19678 11170 19702 11172
rect 19758 11170 19782 11172
rect 19838 11170 19862 11172
rect 19700 11118 19702 11170
rect 19764 11118 19776 11170
rect 19838 11118 19840 11170
rect 19678 11116 19702 11118
rect 19758 11116 19782 11118
rect 19838 11116 19862 11118
rect 19622 11096 19918 11116
rect 19622 10084 19918 10104
rect 19678 10082 19702 10084
rect 19758 10082 19782 10084
rect 19838 10082 19862 10084
rect 19700 10030 19702 10082
rect 19764 10030 19776 10082
rect 19838 10030 19840 10082
rect 19678 10028 19702 10030
rect 19758 10028 19782 10030
rect 19838 10028 19862 10030
rect 19622 10008 19918 10028
rect 19156 9922 19208 9928
rect 18880 9844 18932 9850
rect 18880 9786 18932 9792
rect 18892 9102 18920 9786
rect 19168 9481 19196 9922
rect 19444 9782 19472 9974
rect 19524 9980 19576 9986
rect 19524 9922 19576 9928
rect 19432 9776 19484 9782
rect 19432 9718 19484 9724
rect 19154 9472 19210 9481
rect 19154 9407 19156 9416
rect 19208 9407 19210 9416
rect 19156 9378 19208 9384
rect 19168 9347 19196 9378
rect 19444 9374 19472 9718
rect 19432 9368 19484 9374
rect 20088 9345 20116 27240
rect 20732 24538 20760 27240
rect 20720 24532 20772 24538
rect 20720 24474 20772 24480
rect 20444 24464 20496 24470
rect 20444 24406 20496 24412
rect 20352 23988 20404 23994
rect 20352 23930 20404 23936
rect 20364 23586 20392 23930
rect 20352 23580 20404 23586
rect 20352 23522 20404 23528
rect 20168 17460 20220 17466
rect 20168 17402 20220 17408
rect 20180 17058 20208 17402
rect 20168 17052 20220 17058
rect 20168 16994 20220 17000
rect 20168 15284 20220 15290
rect 20168 15226 20220 15232
rect 20180 14785 20208 15226
rect 20166 14776 20222 14785
rect 20166 14711 20222 14720
rect 20180 14338 20208 14711
rect 20168 14332 20220 14338
rect 20168 14274 20220 14280
rect 20260 12700 20312 12706
rect 20260 12642 20312 12648
rect 20272 10938 20300 12642
rect 20260 10932 20312 10938
rect 20260 10874 20312 10880
rect 20272 10841 20300 10874
rect 20258 10832 20314 10841
rect 20258 10767 20314 10776
rect 19432 9310 19484 9316
rect 20074 9336 20130 9345
rect 20074 9271 20130 9280
rect 18880 9096 18932 9102
rect 20456 9073 20484 24406
rect 21178 24024 21234 24033
rect 21178 23959 21234 23968
rect 21192 23926 21220 23959
rect 21180 23920 21232 23926
rect 21180 23862 21232 23868
rect 21192 23586 21220 23862
rect 21180 23580 21232 23586
rect 21180 23522 21232 23528
rect 20720 23444 20772 23450
rect 20720 23386 20772 23392
rect 20732 22922 20760 23386
rect 20994 23344 21050 23353
rect 20994 23279 21050 23288
rect 20640 22906 20852 22922
rect 20628 22900 20852 22906
rect 20680 22894 20852 22900
rect 20628 22842 20680 22848
rect 20640 22498 20668 22842
rect 20720 22696 20772 22702
rect 20720 22638 20772 22644
rect 20628 22492 20680 22498
rect 20628 22434 20680 22440
rect 20732 21721 20760 22638
rect 20718 21712 20774 21721
rect 20640 21670 20718 21698
rect 20640 20322 20668 21670
rect 20718 21647 20774 21656
rect 20824 21206 20852 22894
rect 21008 21970 21036 23279
rect 21088 22900 21140 22906
rect 21088 22842 21140 22848
rect 21100 22498 21128 22842
rect 21088 22492 21140 22498
rect 21088 22434 21140 22440
rect 21100 22158 21128 22434
rect 21088 22152 21140 22158
rect 21088 22094 21140 22100
rect 21008 21942 21128 21970
rect 20812 21200 20864 21206
rect 20732 21148 20812 21154
rect 20732 21142 20864 21148
rect 20732 21126 20852 21142
rect 20732 21070 20760 21126
rect 20824 21077 20852 21126
rect 20720 21064 20772 21070
rect 20720 21006 20772 21012
rect 20732 20730 20760 21006
rect 20720 20724 20772 20730
rect 20720 20666 20772 20672
rect 20628 20316 20680 20322
rect 20628 20258 20680 20264
rect 20628 18888 20680 18894
rect 20628 18830 20680 18836
rect 20640 18706 20668 18830
rect 20640 18678 20852 18706
rect 20720 18072 20772 18078
rect 20720 18014 20772 18020
rect 20732 17754 20760 18014
rect 20640 17726 20760 17754
rect 20640 17534 20668 17726
rect 20536 17528 20588 17534
rect 20536 17470 20588 17476
rect 20628 17528 20680 17534
rect 20628 17470 20680 17476
rect 20548 17058 20576 17470
rect 20536 17052 20588 17058
rect 20536 16994 20588 17000
rect 20640 15986 20668 17470
rect 20640 15970 20760 15986
rect 20640 15964 20772 15970
rect 20640 15958 20720 15964
rect 20720 15906 20772 15912
rect 20732 15193 20760 15906
rect 20824 15290 20852 18678
rect 20996 17868 21048 17874
rect 20996 17810 21048 17816
rect 20904 17800 20956 17806
rect 20902 17768 20904 17777
rect 20956 17768 20958 17777
rect 20902 17703 20958 17712
rect 21008 16922 21036 17810
rect 20996 16916 21048 16922
rect 20996 16858 21048 16864
rect 20812 15284 20864 15290
rect 20812 15226 20864 15232
rect 20718 15184 20774 15193
rect 20718 15119 20774 15128
rect 20732 14882 20760 15119
rect 20720 14876 20772 14882
rect 20720 14818 20772 14824
rect 20732 13674 20760 14818
rect 21100 14338 21128 21942
rect 21180 21132 21232 21138
rect 21180 21074 21232 21080
rect 21192 20798 21220 21074
rect 21180 20792 21232 20798
rect 21180 20734 21232 20740
rect 21376 20610 21404 27240
rect 21548 26436 21600 26442
rect 21548 26378 21600 26384
rect 21560 23450 21588 26378
rect 21640 24532 21692 24538
rect 21640 24474 21692 24480
rect 21548 23444 21600 23450
rect 21548 23386 21600 23392
rect 21376 20582 21496 20610
rect 21270 19128 21326 19137
rect 21270 19063 21326 19072
rect 21180 18548 21232 18554
rect 21180 18490 21232 18496
rect 21192 18078 21220 18490
rect 21180 18072 21232 18078
rect 21180 18014 21232 18020
rect 21284 15358 21312 19063
rect 21362 18448 21418 18457
rect 21362 18383 21418 18392
rect 21376 17942 21404 18383
rect 21364 17936 21416 17942
rect 21364 17878 21416 17884
rect 21272 15352 21324 15358
rect 21272 15294 21324 15300
rect 21180 15080 21232 15086
rect 21180 15022 21232 15028
rect 21192 14610 21220 15022
rect 21180 14604 21232 14610
rect 21180 14546 21232 14552
rect 21088 14332 21140 14338
rect 21088 14274 21140 14280
rect 21192 13998 21220 14546
rect 21284 14270 21312 15294
rect 21272 14264 21324 14270
rect 21272 14206 21324 14212
rect 21364 14196 21416 14202
rect 21364 14138 21416 14144
rect 21180 13992 21232 13998
rect 21180 13934 21232 13940
rect 20640 13646 20760 13674
rect 21376 13658 21404 14138
rect 21364 13652 21416 13658
rect 20640 13114 20668 13646
rect 21364 13594 21416 13600
rect 20720 13584 20772 13590
rect 20720 13526 20772 13532
rect 20628 13108 20680 13114
rect 20628 13050 20680 13056
rect 20640 12706 20668 13050
rect 20628 12700 20680 12706
rect 20628 12642 20680 12648
rect 20732 12162 20760 13526
rect 20812 13176 20864 13182
rect 20812 13118 20864 13124
rect 20720 12156 20772 12162
rect 20720 12098 20772 12104
rect 20824 11890 20852 13118
rect 20996 12904 21048 12910
rect 20996 12846 21048 12852
rect 21008 12502 21036 12846
rect 20996 12496 21048 12502
rect 20996 12438 21048 12444
rect 20904 11952 20956 11958
rect 20904 11894 20956 11900
rect 20812 11884 20864 11890
rect 20812 11826 20864 11832
rect 20916 11618 20944 11894
rect 20904 11612 20956 11618
rect 20904 11554 20956 11560
rect 20916 11074 20944 11554
rect 21008 11482 21036 12438
rect 20996 11476 21048 11482
rect 20996 11418 21048 11424
rect 21270 11376 21326 11385
rect 21270 11311 21272 11320
rect 21324 11311 21326 11320
rect 21272 11282 21324 11288
rect 20904 11068 20956 11074
rect 20904 11010 20956 11016
rect 21364 11000 21416 11006
rect 21364 10942 21416 10948
rect 20996 10932 21048 10938
rect 20996 10874 21048 10880
rect 21008 10530 21036 10874
rect 21376 10530 21404 10942
rect 21468 10569 21496 20582
rect 21652 20066 21680 24474
rect 22112 23994 22140 27240
rect 22560 24464 22612 24470
rect 22558 24432 22560 24441
rect 22612 24432 22614 24441
rect 22558 24367 22614 24376
rect 22100 23988 22152 23994
rect 22100 23930 22152 23936
rect 22284 23920 22336 23926
rect 22284 23862 22336 23868
rect 22008 23784 22060 23790
rect 22008 23726 22060 23732
rect 22020 22344 22048 23726
rect 22296 23314 22324 23862
rect 22756 23353 22784 27240
rect 23492 27138 23520 27240
rect 23492 27110 23704 27138
rect 23570 26880 23626 26889
rect 23570 26815 23626 26824
rect 23386 26200 23442 26209
rect 23386 26135 23442 26144
rect 22836 25076 22888 25082
rect 22836 25018 22888 25024
rect 22848 24606 22876 25018
rect 22836 24600 22888 24606
rect 22834 24568 22836 24577
rect 22888 24568 22890 24577
rect 22834 24503 22890 24512
rect 22848 24477 22876 24503
rect 23400 24334 23428 26135
rect 23584 25218 23612 26815
rect 23572 25212 23624 25218
rect 23572 25154 23624 25160
rect 23388 24328 23440 24334
rect 23388 24270 23440 24276
rect 23388 23988 23440 23994
rect 23388 23930 23440 23936
rect 23572 23988 23624 23994
rect 23572 23930 23624 23936
rect 22742 23344 22798 23353
rect 22284 23308 22336 23314
rect 22742 23279 22798 23288
rect 23296 23308 23348 23314
rect 22284 23250 22336 23256
rect 23296 23250 23348 23256
rect 22020 22316 22232 22344
rect 22204 22226 22232 22316
rect 22008 22220 22060 22226
rect 22008 22162 22060 22168
rect 22192 22220 22244 22226
rect 22192 22162 22244 22168
rect 22020 21954 22048 22162
rect 22008 21948 22060 21954
rect 22008 21890 22060 21896
rect 22296 21410 22324 23250
rect 22928 23240 22980 23246
rect 22928 23182 22980 23188
rect 22940 22362 22968 23182
rect 22928 22356 22980 22362
rect 22928 22298 22980 22304
rect 23308 22242 23336 23250
rect 23400 22702 23428 23930
rect 23584 23246 23612 23930
rect 23676 23314 23704 27110
rect 23952 26442 23980 27359
rect 24122 27240 24178 27720
rect 24766 27240 24822 27720
rect 25502 27240 25558 27720
rect 26146 27240 26202 27720
rect 26882 27240 26938 27720
rect 27526 27240 27582 27720
rect 23940 26436 23992 26442
rect 23940 26378 23992 26384
rect 24136 24554 24164 27240
rect 24780 25778 24808 27240
rect 24688 25750 24808 25778
rect 24289 24772 24585 24792
rect 24345 24770 24369 24772
rect 24425 24770 24449 24772
rect 24505 24770 24529 24772
rect 24367 24718 24369 24770
rect 24431 24718 24443 24770
rect 24505 24718 24507 24770
rect 24345 24716 24369 24718
rect 24425 24716 24449 24718
rect 24505 24716 24529 24718
rect 24289 24696 24585 24716
rect 23952 24526 24164 24554
rect 23664 23308 23716 23314
rect 23664 23250 23716 23256
rect 23572 23240 23624 23246
rect 23848 23240 23900 23246
rect 23572 23182 23624 23188
rect 23662 23208 23718 23217
rect 23584 22809 23612 23182
rect 23848 23182 23900 23188
rect 23662 23143 23718 23152
rect 23570 22800 23626 22809
rect 23570 22735 23626 22744
rect 23388 22696 23440 22702
rect 23388 22638 23440 22644
rect 23572 22696 23624 22702
rect 23572 22638 23624 22644
rect 23584 22242 23612 22638
rect 23676 22498 23704 23143
rect 23756 22900 23808 22906
rect 23756 22842 23808 22848
rect 23664 22492 23716 22498
rect 23664 22434 23716 22440
rect 23768 22430 23796 22842
rect 23756 22424 23808 22430
rect 23756 22366 23808 22372
rect 23860 22265 23888 23182
rect 23846 22256 23902 22265
rect 23308 22214 23428 22242
rect 23584 22214 23796 22242
rect 22376 22152 22428 22158
rect 22376 22094 22428 22100
rect 23296 22152 23348 22158
rect 23296 22094 23348 22100
rect 23400 22106 23428 22214
rect 22388 21886 22416 22094
rect 22376 21880 22428 21886
rect 23308 21857 23336 22094
rect 23400 22078 23612 22106
rect 22376 21822 22428 21828
rect 23294 21848 23350 21857
rect 23294 21783 23350 21792
rect 22284 21404 22336 21410
rect 22284 21346 22336 21352
rect 22100 21200 22152 21206
rect 22100 21142 22152 21148
rect 22006 21032 22062 21041
rect 22006 20967 22062 20976
rect 22020 20866 22048 20967
rect 22008 20860 22060 20866
rect 22008 20802 22060 20808
rect 22112 20186 22140 21142
rect 23204 21064 23256 21070
rect 23204 21006 23256 21012
rect 23480 21064 23532 21070
rect 23480 21006 23532 21012
rect 22192 20860 22244 20866
rect 22192 20802 22244 20808
rect 22100 20180 22152 20186
rect 22100 20122 22152 20128
rect 21652 20038 21772 20066
rect 21640 19976 21692 19982
rect 21640 19918 21692 19924
rect 21548 18616 21600 18622
rect 21548 18558 21600 18564
rect 21560 18010 21588 18558
rect 21548 18004 21600 18010
rect 21548 17946 21600 17952
rect 21560 17602 21588 17946
rect 21548 17596 21600 17602
rect 21548 17538 21600 17544
rect 21652 16825 21680 19918
rect 21638 16816 21694 16825
rect 21638 16751 21694 16760
rect 21652 16378 21680 16751
rect 21640 16372 21692 16378
rect 21640 16314 21692 16320
rect 21652 15630 21680 16314
rect 21640 15624 21692 15630
rect 21640 15566 21692 15572
rect 21454 10560 21510 10569
rect 20996 10524 21048 10530
rect 20996 10466 21048 10472
rect 21364 10524 21416 10530
rect 21454 10495 21510 10504
rect 21364 10466 21416 10472
rect 18880 9038 18932 9044
rect 20442 9064 20498 9073
rect 18892 7713 18920 9038
rect 19622 8996 19918 9016
rect 20442 8999 20498 9008
rect 19678 8994 19702 8996
rect 19758 8994 19782 8996
rect 19838 8994 19862 8996
rect 19700 8942 19702 8994
rect 19764 8942 19776 8994
rect 19838 8942 19840 8994
rect 19678 8940 19702 8942
rect 19758 8940 19782 8942
rect 19838 8940 19862 8942
rect 19622 8920 19918 8940
rect 19622 7908 19918 7928
rect 19678 7906 19702 7908
rect 19758 7906 19782 7908
rect 19838 7906 19862 7908
rect 19700 7854 19702 7906
rect 19764 7854 19776 7906
rect 19838 7854 19840 7906
rect 19678 7852 19702 7854
rect 19758 7852 19782 7854
rect 19838 7852 19862 7854
rect 19622 7832 19918 7852
rect 18878 7704 18934 7713
rect 18878 7639 18934 7648
rect 18418 7568 18474 7577
rect 18418 7503 18474 7512
rect 17880 7266 18000 7282
rect 17868 7260 18000 7266
rect 17920 7254 18000 7260
rect 17868 7202 17920 7208
rect 18234 7160 18290 7169
rect 18234 7095 18236 7104
rect 18288 7095 18290 7104
rect 18236 7066 18288 7072
rect 19622 6820 19918 6840
rect 19678 6818 19702 6820
rect 19758 6818 19782 6820
rect 19838 6818 19862 6820
rect 19700 6766 19702 6818
rect 19764 6766 19776 6818
rect 19838 6766 19840 6818
rect 19678 6764 19702 6766
rect 19758 6764 19782 6766
rect 19838 6764 19862 6766
rect 19622 6744 19918 6764
rect 16500 6574 16620 6602
rect 16500 6178 16528 6574
rect 16488 6172 16540 6178
rect 16488 6114 16540 6120
rect 16946 5936 17002 5945
rect 16946 5871 16948 5880
rect 17000 5871 17002 5880
rect 16948 5842 17000 5848
rect 19622 5732 19918 5752
rect 19678 5730 19702 5732
rect 19758 5730 19782 5732
rect 19838 5730 19862 5732
rect 19700 5678 19702 5730
rect 19764 5678 19776 5730
rect 19838 5678 19840 5730
rect 19678 5676 19702 5678
rect 19758 5676 19782 5678
rect 19838 5676 19862 5678
rect 19622 5656 19918 5676
rect 16026 5392 16082 5401
rect 16026 5327 16082 5336
rect 15752 5084 15804 5090
rect 15752 5026 15804 5032
rect 15934 4984 15990 4993
rect 15934 4919 15936 4928
rect 15988 4919 15990 4928
rect 15936 4890 15988 4896
rect 10289 4644 10585 4664
rect 10345 4642 10369 4644
rect 10425 4642 10449 4644
rect 10505 4642 10529 4644
rect 10367 4590 10369 4642
rect 10431 4590 10443 4642
rect 10505 4590 10507 4642
rect 10345 4588 10369 4590
rect 10425 4588 10449 4590
rect 10505 4588 10529 4590
rect 10289 4568 10585 4588
rect 19622 4644 19918 4664
rect 19678 4642 19702 4644
rect 19758 4642 19782 4644
rect 19838 4642 19862 4644
rect 19700 4590 19702 4642
rect 19764 4590 19776 4642
rect 19838 4590 19840 4642
rect 19678 4588 19702 4590
rect 19758 4588 19782 4590
rect 19838 4588 19862 4590
rect 19622 4568 19918 4588
rect 5622 4100 5918 4120
rect 5678 4098 5702 4100
rect 5758 4098 5782 4100
rect 5838 4098 5862 4100
rect 5700 4046 5702 4098
rect 5764 4046 5776 4098
rect 5838 4046 5840 4098
rect 5678 4044 5702 4046
rect 5758 4044 5782 4046
rect 5838 4044 5862 4046
rect 5622 4024 5918 4044
rect 14956 4100 15252 4120
rect 15012 4098 15036 4100
rect 15092 4098 15116 4100
rect 15172 4098 15196 4100
rect 15034 4046 15036 4098
rect 15098 4046 15110 4098
rect 15172 4046 15174 4098
rect 15012 4044 15036 4046
rect 15092 4044 15116 4046
rect 15172 4044 15196 4046
rect 14956 4024 15252 4044
rect 21652 3769 21680 15566
rect 21744 10025 21772 20038
rect 22204 19982 22232 20802
rect 22466 20760 22522 20769
rect 22466 20695 22468 20704
rect 22520 20695 22522 20704
rect 22468 20666 22520 20672
rect 22480 20338 22508 20666
rect 22652 20520 22704 20526
rect 22652 20462 22704 20468
rect 22388 20322 22508 20338
rect 22376 20316 22508 20322
rect 22428 20310 22508 20316
rect 22376 20258 22428 20264
rect 22376 20180 22428 20186
rect 22376 20122 22428 20128
rect 22388 20050 22416 20122
rect 22664 20118 22692 20462
rect 22652 20112 22704 20118
rect 22652 20054 22704 20060
rect 22376 20044 22428 20050
rect 22376 19986 22428 19992
rect 22192 19976 22244 19982
rect 22192 19918 22244 19924
rect 22388 19778 22416 19986
rect 22376 19772 22428 19778
rect 22376 19714 22428 19720
rect 22664 19710 22692 20054
rect 23216 19778 23244 21006
rect 23204 19772 23256 19778
rect 23204 19714 23256 19720
rect 22652 19704 22704 19710
rect 22652 19646 22704 19652
rect 23492 19642 23520 21006
rect 23480 19636 23532 19642
rect 23480 19578 23532 19584
rect 22008 19024 22060 19030
rect 22008 18966 22060 18972
rect 22282 18992 22338 19001
rect 21916 18888 21968 18894
rect 21916 18830 21968 18836
rect 21928 18593 21956 18830
rect 21914 18584 21970 18593
rect 21914 18519 21970 18528
rect 22020 18350 22048 18966
rect 22282 18927 22284 18936
rect 22336 18927 22338 18936
rect 22284 18898 22336 18904
rect 22376 18888 22428 18894
rect 22376 18830 22428 18836
rect 23388 18888 23440 18894
rect 23388 18830 23440 18836
rect 22388 18486 22416 18830
rect 22376 18480 22428 18486
rect 22376 18422 22428 18428
rect 22008 18344 22060 18350
rect 22008 18286 22060 18292
rect 22468 18344 22520 18350
rect 22468 18286 22520 18292
rect 22480 17942 22508 18286
rect 22468 17936 22520 17942
rect 22468 17878 22520 17884
rect 23112 17936 23164 17942
rect 23112 17878 23164 17884
rect 23124 17602 23152 17878
rect 23112 17596 23164 17602
rect 23112 17538 23164 17544
rect 23400 17482 23428 18830
rect 23480 18480 23532 18486
rect 23480 18422 23532 18428
rect 23492 17602 23520 18422
rect 23480 17596 23532 17602
rect 23480 17538 23532 17544
rect 23400 17454 23520 17482
rect 21824 16508 21876 16514
rect 21824 16450 21876 16456
rect 21836 14649 21864 16450
rect 21916 16304 21968 16310
rect 21916 16246 21968 16252
rect 21928 15766 21956 16246
rect 22376 16168 22428 16174
rect 22376 16110 22428 16116
rect 21916 15760 21968 15766
rect 21916 15702 21968 15708
rect 21928 15426 21956 15702
rect 22388 15698 22416 16110
rect 22376 15692 22428 15698
rect 22376 15634 22428 15640
rect 21916 15420 21968 15426
rect 21916 15362 21968 15368
rect 22008 15284 22060 15290
rect 22008 15226 22060 15232
rect 22020 15034 22048 15226
rect 22020 15006 22140 15034
rect 21822 14640 21878 14649
rect 21822 14575 21878 14584
rect 22008 13992 22060 13998
rect 22112 13980 22140 15006
rect 22388 14542 22416 15634
rect 23492 15630 23520 17454
rect 23584 15834 23612 22078
rect 23768 21410 23796 22214
rect 23846 22191 23902 22200
rect 23848 21608 23900 21614
rect 23848 21550 23900 21556
rect 23756 21404 23808 21410
rect 23756 21346 23808 21352
rect 23756 21268 23808 21274
rect 23756 21210 23808 21216
rect 23768 20798 23796 21210
rect 23860 21070 23888 21550
rect 23848 21064 23900 21070
rect 23846 21032 23848 21041
rect 23900 21032 23902 21041
rect 23846 20967 23902 20976
rect 23756 20792 23808 20798
rect 23756 20734 23808 20740
rect 23664 20656 23716 20662
rect 23664 20598 23716 20604
rect 23676 20050 23704 20598
rect 23768 20322 23796 20734
rect 23756 20316 23808 20322
rect 23756 20258 23808 20264
rect 23756 20180 23808 20186
rect 23756 20122 23808 20128
rect 23664 20044 23716 20050
rect 23664 19986 23716 19992
rect 23664 18344 23716 18350
rect 23664 18286 23716 18292
rect 23676 17466 23704 18286
rect 23664 17460 23716 17466
rect 23664 17402 23716 17408
rect 23768 17346 23796 20122
rect 23848 19636 23900 19642
rect 23848 19578 23900 19584
rect 23860 19234 23888 19578
rect 23848 19228 23900 19234
rect 23848 19170 23900 19176
rect 23846 17768 23902 17777
rect 23846 17703 23902 17712
rect 23676 17318 23796 17346
rect 23572 15828 23624 15834
rect 23572 15770 23624 15776
rect 22928 15624 22980 15630
rect 22928 15566 22980 15572
rect 23480 15624 23532 15630
rect 23480 15566 23532 15572
rect 22940 14814 22968 15566
rect 23480 15284 23532 15290
rect 23480 15226 23532 15232
rect 23492 14898 23520 15226
rect 23676 15170 23704 17318
rect 23754 17224 23810 17233
rect 23754 17159 23810 17168
rect 23768 15902 23796 17159
rect 23860 17058 23888 17703
rect 23848 17052 23900 17058
rect 23848 16994 23900 17000
rect 23860 16854 23888 16994
rect 23848 16848 23900 16854
rect 23848 16790 23900 16796
rect 23846 16408 23902 16417
rect 23846 16343 23848 16352
rect 23900 16343 23902 16352
rect 23848 16314 23900 16320
rect 23860 15970 23888 16314
rect 23848 15964 23900 15970
rect 23848 15906 23900 15912
rect 23756 15896 23808 15902
rect 23756 15838 23808 15844
rect 23848 15828 23900 15834
rect 23848 15770 23900 15776
rect 23756 15624 23808 15630
rect 23756 15566 23808 15572
rect 23400 14882 23520 14898
rect 23388 14876 23520 14882
rect 23440 14870 23520 14876
rect 23584 15142 23704 15170
rect 23388 14818 23440 14824
rect 22928 14808 22980 14814
rect 22926 14776 22928 14785
rect 22980 14776 22982 14785
rect 22926 14711 22982 14720
rect 22376 14536 22428 14542
rect 22376 14478 22428 14484
rect 23400 14338 23428 14818
rect 23478 14640 23534 14649
rect 23478 14575 23480 14584
rect 23532 14575 23534 14584
rect 23480 14546 23532 14552
rect 23388 14332 23440 14338
rect 23388 14274 23440 14280
rect 23584 14218 23612 15142
rect 23664 15080 23716 15086
rect 23664 15022 23716 15028
rect 23676 14678 23704 15022
rect 23664 14672 23716 14678
rect 23664 14614 23716 14620
rect 23676 14338 23704 14614
rect 23664 14332 23716 14338
rect 23664 14274 23716 14280
rect 23584 14190 23704 14218
rect 22284 13992 22336 13998
rect 22112 13952 22284 13980
rect 22008 13934 22060 13940
rect 22284 13934 22336 13940
rect 22020 13250 22048 13934
rect 22008 13244 22060 13250
rect 22008 13186 22060 13192
rect 21916 12360 21968 12366
rect 21916 12302 21968 12308
rect 21928 11958 21956 12302
rect 21916 11952 21968 11958
rect 21916 11894 21968 11900
rect 21928 11618 21956 11894
rect 21916 11612 21968 11618
rect 21916 11554 21968 11560
rect 22192 11476 22244 11482
rect 22192 11418 22244 11424
rect 22204 11074 22232 11418
rect 22192 11068 22244 11074
rect 22192 11010 22244 11016
rect 21730 10016 21786 10025
rect 21730 9951 21786 9960
rect 21638 3760 21694 3769
rect 21638 3695 21694 3704
rect 10289 3556 10585 3576
rect 10345 3554 10369 3556
rect 10425 3554 10449 3556
rect 10505 3554 10529 3556
rect 10367 3502 10369 3554
rect 10431 3502 10443 3554
rect 10505 3502 10507 3554
rect 10345 3500 10369 3502
rect 10425 3500 10449 3502
rect 10505 3500 10529 3502
rect 10289 3480 10585 3500
rect 19622 3556 19918 3576
rect 19678 3554 19702 3556
rect 19758 3554 19782 3556
rect 19838 3554 19862 3556
rect 19700 3502 19702 3554
rect 19764 3502 19776 3554
rect 19838 3502 19840 3554
rect 19678 3500 19702 3502
rect 19758 3500 19782 3502
rect 19838 3500 19862 3502
rect 19622 3480 19918 3500
rect 5622 3012 5918 3032
rect 5678 3010 5702 3012
rect 5758 3010 5782 3012
rect 5838 3010 5862 3012
rect 5700 2958 5702 3010
rect 5764 2958 5776 3010
rect 5838 2958 5840 3010
rect 5678 2956 5702 2958
rect 5758 2956 5782 2958
rect 5838 2956 5862 2958
rect 5622 2936 5918 2956
rect 14956 3012 15252 3032
rect 15012 3010 15036 3012
rect 15092 3010 15116 3012
rect 15172 3010 15196 3012
rect 15034 2958 15036 3010
rect 15098 2958 15110 3010
rect 15172 2958 15174 3010
rect 15012 2956 15036 2958
rect 15092 2956 15116 2958
rect 15172 2956 15196 2958
rect 14956 2936 15252 2956
rect 10289 2468 10585 2488
rect 10345 2466 10369 2468
rect 10425 2466 10449 2468
rect 10505 2466 10529 2468
rect 10367 2414 10369 2466
rect 10431 2414 10443 2466
rect 10505 2414 10507 2466
rect 10345 2412 10369 2414
rect 10425 2412 10449 2414
rect 10505 2412 10529 2414
rect 10289 2392 10585 2412
rect 19622 2468 19918 2488
rect 19678 2466 19702 2468
rect 19758 2466 19782 2468
rect 19838 2466 19862 2468
rect 19700 2414 19702 2466
rect 19764 2414 19776 2466
rect 19838 2414 19840 2466
rect 19678 2412 19702 2414
rect 19758 2412 19782 2414
rect 19838 2412 19862 2414
rect 19622 2392 19918 2412
rect 22296 2409 22324 13934
rect 23570 13824 23626 13833
rect 23676 13794 23704 14190
rect 23570 13759 23626 13768
rect 23664 13788 23716 13794
rect 23478 10560 23534 10569
rect 23478 10495 23480 10504
rect 23532 10495 23534 10504
rect 23480 10466 23532 10472
rect 23478 3760 23534 3769
rect 23478 3695 23534 3704
rect 22282 2400 22338 2409
rect 22282 2335 22338 2344
rect 5622 1924 5918 1944
rect 5678 1922 5702 1924
rect 5758 1922 5782 1924
rect 5838 1922 5862 1924
rect 5700 1870 5702 1922
rect 5764 1870 5776 1922
rect 5838 1870 5840 1922
rect 5678 1868 5702 1870
rect 5758 1868 5782 1870
rect 5838 1868 5862 1870
rect 5622 1848 5918 1868
rect 14956 1924 15252 1944
rect 15012 1922 15036 1924
rect 15092 1922 15116 1924
rect 15172 1922 15196 1924
rect 15034 1870 15036 1922
rect 15098 1870 15110 1922
rect 15172 1870 15174 1922
rect 15012 1868 15036 1870
rect 15092 1868 15116 1870
rect 15172 1868 15196 1870
rect 14956 1848 15252 1868
rect 23492 1185 23520 3695
rect 23584 3225 23612 13759
rect 23664 13730 23716 13736
rect 23768 13674 23796 15566
rect 23676 13646 23796 13674
rect 23570 3216 23626 3225
rect 23570 3151 23626 3160
rect 23570 2400 23626 2409
rect 23570 2335 23626 2344
rect 23478 1176 23534 1185
rect 23478 1111 23534 1120
rect 23584 97 23612 2335
rect 23676 641 23704 13646
rect 23754 13552 23810 13561
rect 23754 13487 23810 13496
rect 23768 7266 23796 13487
rect 23860 12586 23888 15770
rect 23952 12706 23980 24526
rect 24124 24464 24176 24470
rect 24124 24406 24176 24412
rect 24032 22832 24084 22838
rect 24032 22774 24084 22780
rect 24044 20225 24072 22774
rect 24136 22673 24164 24406
rect 24289 23684 24585 23704
rect 24345 23682 24369 23684
rect 24425 23682 24449 23684
rect 24505 23682 24529 23684
rect 24367 23630 24369 23682
rect 24431 23630 24443 23682
rect 24505 23630 24507 23682
rect 24345 23628 24369 23630
rect 24425 23628 24449 23630
rect 24505 23628 24529 23630
rect 24289 23608 24585 23628
rect 24122 22664 24178 22673
rect 24122 22599 24178 22608
rect 24289 22596 24585 22616
rect 24345 22594 24369 22596
rect 24425 22594 24449 22596
rect 24505 22594 24529 22596
rect 24367 22542 24369 22594
rect 24431 22542 24443 22594
rect 24505 22542 24507 22594
rect 24345 22540 24369 22542
rect 24425 22540 24449 22542
rect 24505 22540 24529 22542
rect 24289 22520 24585 22540
rect 24582 22392 24638 22401
rect 24582 22327 24638 22336
rect 24596 22294 24624 22327
rect 24584 22288 24636 22294
rect 24584 22230 24636 22236
rect 24688 21818 24716 25750
rect 24766 25656 24822 25665
rect 24766 25591 24822 25600
rect 24780 25218 24808 25591
rect 24768 25212 24820 25218
rect 24768 25154 24820 25160
rect 25134 25112 25190 25121
rect 24768 25076 24820 25082
rect 25134 25047 25190 25056
rect 24768 25018 24820 25024
rect 24780 24334 24808 25018
rect 25148 24674 25176 25047
rect 25136 24668 25188 24674
rect 25136 24610 25188 24616
rect 24952 24464 25004 24470
rect 24952 24406 25004 24412
rect 25134 24432 25190 24441
rect 24768 24328 24820 24334
rect 24768 24270 24820 24276
rect 24780 24062 24808 24270
rect 24768 24056 24820 24062
rect 24768 23998 24820 24004
rect 24860 23988 24912 23994
rect 24860 23930 24912 23936
rect 24766 23752 24822 23761
rect 24766 23687 24822 23696
rect 24780 22242 24808 23687
rect 24872 23246 24900 23930
rect 24964 23450 24992 24406
rect 25134 24367 25190 24376
rect 25320 24396 25372 24402
rect 25148 24130 25176 24367
rect 25320 24338 25372 24344
rect 25136 24124 25188 24130
rect 25136 24066 25188 24072
rect 24952 23444 25004 23450
rect 24952 23386 25004 23392
rect 25332 23382 25360 24338
rect 25516 24010 25544 27240
rect 25686 24568 25742 24577
rect 25686 24503 25742 24512
rect 25424 23982 25544 24010
rect 25424 23761 25452 23982
rect 25502 23888 25558 23897
rect 25502 23823 25558 23832
rect 25410 23752 25466 23761
rect 25410 23687 25466 23696
rect 25516 23586 25544 23823
rect 25504 23580 25556 23586
rect 25504 23522 25556 23528
rect 25320 23376 25372 23382
rect 25320 23318 25372 23324
rect 24860 23240 24912 23246
rect 24860 23182 24912 23188
rect 24872 22945 24900 23182
rect 24858 22936 24914 22945
rect 24858 22871 24914 22880
rect 24952 22900 25004 22906
rect 24952 22842 25004 22848
rect 24964 22498 24992 22842
rect 25136 22696 25188 22702
rect 25134 22664 25136 22673
rect 25188 22664 25190 22673
rect 25134 22599 25190 22608
rect 24952 22492 25004 22498
rect 24952 22434 25004 22440
rect 25504 22492 25556 22498
rect 25504 22434 25556 22440
rect 24780 22214 24900 22242
rect 24768 22152 24820 22158
rect 24766 22120 24768 22129
rect 24820 22120 24822 22129
rect 24766 22055 24822 22064
rect 24676 21812 24728 21818
rect 24676 21754 24728 21760
rect 24124 21744 24176 21750
rect 24124 21686 24176 21692
rect 24216 21744 24268 21750
rect 24872 21698 24900 22214
rect 24216 21686 24268 21692
rect 24136 21585 24164 21686
rect 24122 21576 24178 21585
rect 24122 21511 24178 21520
rect 24136 21410 24164 21511
rect 24124 21404 24176 21410
rect 24124 21346 24176 21352
rect 24124 20792 24176 20798
rect 24124 20734 24176 20740
rect 24136 20322 24164 20734
rect 24124 20316 24176 20322
rect 24124 20258 24176 20264
rect 24030 20216 24086 20225
rect 24030 20151 24086 20160
rect 24136 19658 24164 20258
rect 24044 19630 24164 19658
rect 24044 18690 24072 19630
rect 24124 19568 24176 19574
rect 24124 19510 24176 19516
rect 24136 19030 24164 19510
rect 24124 19024 24176 19030
rect 24124 18966 24176 18972
rect 24032 18684 24084 18690
rect 24032 18626 24084 18632
rect 24124 18616 24176 18622
rect 24124 18558 24176 18564
rect 24032 18548 24084 18554
rect 24032 18490 24084 18496
rect 24044 17602 24072 18490
rect 24136 18146 24164 18558
rect 24124 18140 24176 18146
rect 24124 18082 24176 18088
rect 24032 17596 24084 17602
rect 24032 17538 24084 17544
rect 24044 16990 24072 17538
rect 24124 17460 24176 17466
rect 24124 17402 24176 17408
rect 24136 17058 24164 17402
rect 24124 17052 24176 17058
rect 24124 16994 24176 17000
rect 24032 16984 24084 16990
rect 24032 16926 24084 16932
rect 24122 15728 24178 15737
rect 24122 15663 24178 15672
rect 24136 15426 24164 15663
rect 24124 15420 24176 15426
rect 24124 15362 24176 15368
rect 24032 15148 24084 15154
rect 24032 15090 24084 15096
rect 24044 14542 24072 15090
rect 24136 14882 24164 15362
rect 24124 14876 24176 14882
rect 24124 14818 24176 14824
rect 24032 14536 24084 14542
rect 24032 14478 24084 14484
rect 24044 14338 24072 14478
rect 24122 14368 24178 14377
rect 24032 14332 24084 14338
rect 24122 14303 24178 14312
rect 24032 14274 24084 14280
rect 24032 14060 24084 14066
rect 24032 14002 24084 14008
rect 24044 12722 24072 14002
rect 24136 13794 24164 14303
rect 24124 13788 24176 13794
rect 24124 13730 24176 13736
rect 24136 13590 24164 13730
rect 24124 13584 24176 13590
rect 24124 13526 24176 13532
rect 24228 13250 24256 21686
rect 24688 21670 24900 21698
rect 24289 21508 24585 21528
rect 24345 21506 24369 21508
rect 24425 21506 24449 21508
rect 24505 21506 24529 21508
rect 24367 21454 24369 21506
rect 24431 21454 24443 21506
rect 24505 21454 24507 21506
rect 24345 21452 24369 21454
rect 24425 21452 24449 21454
rect 24505 21452 24529 21454
rect 24289 21432 24585 21452
rect 24289 20420 24585 20440
rect 24345 20418 24369 20420
rect 24425 20418 24449 20420
rect 24505 20418 24529 20420
rect 24367 20366 24369 20418
rect 24431 20366 24443 20418
rect 24505 20366 24507 20418
rect 24345 20364 24369 20366
rect 24425 20364 24449 20366
rect 24505 20364 24529 20366
rect 24289 20344 24585 20364
rect 24289 19332 24585 19352
rect 24345 19330 24369 19332
rect 24425 19330 24449 19332
rect 24505 19330 24529 19332
rect 24367 19278 24369 19330
rect 24431 19278 24443 19330
rect 24505 19278 24507 19330
rect 24345 19276 24369 19278
rect 24425 19276 24449 19278
rect 24505 19276 24529 19278
rect 24289 19256 24585 19276
rect 24289 18244 24585 18264
rect 24345 18242 24369 18244
rect 24425 18242 24449 18244
rect 24505 18242 24529 18244
rect 24367 18190 24369 18242
rect 24431 18190 24443 18242
rect 24505 18190 24507 18242
rect 24345 18188 24369 18190
rect 24425 18188 24449 18190
rect 24505 18188 24529 18190
rect 24289 18168 24585 18188
rect 24289 17156 24585 17176
rect 24345 17154 24369 17156
rect 24425 17154 24449 17156
rect 24505 17154 24529 17156
rect 24367 17102 24369 17154
rect 24431 17102 24443 17154
rect 24505 17102 24507 17154
rect 24345 17100 24369 17102
rect 24425 17100 24449 17102
rect 24505 17100 24529 17102
rect 24289 17080 24585 17100
rect 24289 16068 24585 16088
rect 24345 16066 24369 16068
rect 24425 16066 24449 16068
rect 24505 16066 24529 16068
rect 24367 16014 24369 16066
rect 24431 16014 24443 16066
rect 24505 16014 24507 16066
rect 24345 16012 24369 16014
rect 24425 16012 24449 16014
rect 24505 16012 24529 16014
rect 24289 15992 24585 16012
rect 24289 14980 24585 15000
rect 24345 14978 24369 14980
rect 24425 14978 24449 14980
rect 24505 14978 24529 14980
rect 24367 14926 24369 14978
rect 24431 14926 24443 14978
rect 24505 14926 24507 14978
rect 24345 14924 24369 14926
rect 24425 14924 24449 14926
rect 24505 14924 24529 14926
rect 24289 14904 24585 14924
rect 24308 14536 24360 14542
rect 24308 14478 24360 14484
rect 24320 14066 24348 14478
rect 24308 14060 24360 14066
rect 24308 14002 24360 14008
rect 24289 13892 24585 13912
rect 24345 13890 24369 13892
rect 24425 13890 24449 13892
rect 24505 13890 24529 13892
rect 24367 13838 24369 13890
rect 24431 13838 24443 13890
rect 24505 13838 24507 13890
rect 24345 13836 24369 13838
rect 24425 13836 24449 13838
rect 24505 13836 24529 13838
rect 24289 13816 24585 13836
rect 24688 13794 24716 21670
rect 24768 21608 24820 21614
rect 24768 21550 24820 21556
rect 24780 21449 24808 21550
rect 24766 21440 24822 21449
rect 24766 21375 24822 21384
rect 24768 21336 24820 21342
rect 25516 21313 25544 22434
rect 24768 21278 24820 21284
rect 25502 21304 25558 21313
rect 24780 19794 24808 21278
rect 25502 21239 25558 21248
rect 24952 21200 25004 21206
rect 24952 21142 25004 21148
rect 24858 20216 24914 20225
rect 24858 20151 24914 20160
rect 24872 20118 24900 20151
rect 24860 20112 24912 20118
rect 24964 20089 24992 21142
rect 25136 21064 25188 21070
rect 25136 21006 25188 21012
rect 25148 20905 25176 21006
rect 25134 20896 25190 20905
rect 25134 20831 25190 20840
rect 25318 20352 25374 20361
rect 25318 20287 25374 20296
rect 24860 20054 24912 20060
rect 24950 20080 25006 20089
rect 24950 20015 25006 20024
rect 25044 19976 25096 19982
rect 25044 19918 25096 19924
rect 24780 19766 24992 19794
rect 24858 19672 24914 19681
rect 24858 19607 24860 19616
rect 24912 19607 24914 19616
rect 24860 19578 24912 19584
rect 24872 19234 24900 19578
rect 24860 19228 24912 19234
rect 24860 19170 24912 19176
rect 24766 19128 24822 19137
rect 24766 19063 24822 19072
rect 24780 18894 24808 19063
rect 24768 18888 24820 18894
rect 24768 18830 24820 18836
rect 24860 17868 24912 17874
rect 24860 17810 24912 17816
rect 24872 17754 24900 17810
rect 24780 17726 24900 17754
rect 24780 17534 24808 17726
rect 24964 17618 24992 19766
rect 25056 19681 25084 19918
rect 25332 19778 25360 20287
rect 25320 19772 25372 19778
rect 25320 19714 25372 19720
rect 25042 19672 25098 19681
rect 25042 19607 25098 19616
rect 25228 18548 25280 18554
rect 25228 18490 25280 18496
rect 25240 17874 25268 18490
rect 25410 18448 25466 18457
rect 25410 18383 25412 18392
rect 25464 18383 25466 18392
rect 25412 18354 25464 18360
rect 25594 17904 25650 17913
rect 25228 17868 25280 17874
rect 25594 17839 25650 17848
rect 25228 17810 25280 17816
rect 24872 17590 24992 17618
rect 25608 17602 25636 17839
rect 25596 17596 25648 17602
rect 24768 17528 24820 17534
rect 24768 17470 24820 17476
rect 24872 17346 24900 17590
rect 25596 17538 25648 17544
rect 25412 17460 25464 17466
rect 25412 17402 25464 17408
rect 24780 17318 24900 17346
rect 24780 16360 24808 17318
rect 25424 16922 25452 17402
rect 25502 17360 25558 17369
rect 25502 17295 25558 17304
rect 25516 17058 25544 17295
rect 25504 17052 25556 17058
rect 25504 16994 25556 17000
rect 25412 16916 25464 16922
rect 25412 16858 25464 16864
rect 25320 16848 25372 16854
rect 25320 16790 25372 16796
rect 25332 16446 25360 16790
rect 25410 16680 25466 16689
rect 25410 16615 25466 16624
rect 25424 16514 25452 16615
rect 25412 16508 25464 16514
rect 25412 16450 25464 16456
rect 25320 16440 25372 16446
rect 25320 16382 25372 16388
rect 25228 16372 25280 16378
rect 24780 16332 24900 16360
rect 24766 16272 24822 16281
rect 24766 16207 24822 16216
rect 24780 14202 24808 16207
rect 24768 14196 24820 14202
rect 24768 14138 24820 14144
rect 24676 13788 24728 13794
rect 24676 13730 24728 13736
rect 24780 13658 24808 14138
rect 24768 13652 24820 13658
rect 24768 13594 24820 13600
rect 24872 13538 24900 16332
rect 25228 16314 25280 16320
rect 25240 15970 25268 16314
rect 25318 16136 25374 16145
rect 25318 16071 25374 16080
rect 25228 15964 25280 15970
rect 25228 15906 25280 15912
rect 25136 15284 25188 15290
rect 25136 15226 25188 15232
rect 25148 14814 25176 15226
rect 25332 14882 25360 16071
rect 25502 15456 25558 15465
rect 25502 15391 25558 15400
rect 25412 15216 25464 15222
rect 25412 15158 25464 15164
rect 25320 14876 25372 14882
rect 25320 14818 25372 14824
rect 25136 14808 25188 14814
rect 25136 14750 25188 14756
rect 25044 14672 25096 14678
rect 25044 14614 25096 14620
rect 25056 14338 25084 14614
rect 25044 14332 25096 14338
rect 25044 14274 25096 14280
rect 25424 14202 25452 15158
rect 25516 14338 25544 15391
rect 25594 14912 25650 14921
rect 25594 14847 25650 14856
rect 25504 14332 25556 14338
rect 25504 14274 25556 14280
rect 25412 14196 25464 14202
rect 25412 14138 25464 14144
rect 25424 13794 25452 14138
rect 25412 13788 25464 13794
rect 25412 13730 25464 13736
rect 25226 13688 25282 13697
rect 25226 13623 25228 13632
rect 25280 13623 25282 13632
rect 25228 13594 25280 13600
rect 24780 13510 24900 13538
rect 24216 13244 24268 13250
rect 24216 13186 24268 13192
rect 24582 13144 24638 13153
rect 24582 13079 24584 13088
rect 24636 13079 24638 13088
rect 24584 13050 24636 13056
rect 24596 12994 24624 13050
rect 24596 12966 24716 12994
rect 24289 12804 24585 12824
rect 24345 12802 24369 12804
rect 24425 12802 24449 12804
rect 24505 12802 24529 12804
rect 24367 12750 24369 12802
rect 24431 12750 24443 12802
rect 24505 12750 24507 12802
rect 24345 12748 24369 12750
rect 24425 12748 24449 12750
rect 24505 12748 24529 12750
rect 24289 12728 24585 12748
rect 23940 12700 23992 12706
rect 24044 12694 24164 12722
rect 24688 12706 24716 12966
rect 23940 12642 23992 12648
rect 23860 12558 24072 12586
rect 23848 12428 23900 12434
rect 23848 12370 23900 12376
rect 23756 7260 23808 7266
rect 23756 7202 23808 7208
rect 23860 2409 23888 12370
rect 24044 12162 24072 12558
rect 24136 12434 24164 12694
rect 24676 12700 24728 12706
rect 24676 12642 24728 12648
rect 24398 12600 24454 12609
rect 24398 12535 24400 12544
rect 24452 12535 24454 12544
rect 24400 12506 24452 12512
rect 24124 12428 24176 12434
rect 24124 12370 24176 12376
rect 24032 12156 24084 12162
rect 24032 12098 24084 12104
rect 24400 12020 24452 12026
rect 24400 11962 24452 11968
rect 24412 11929 24440 11962
rect 24398 11920 24454 11929
rect 24398 11855 24454 11864
rect 24674 11920 24730 11929
rect 24674 11855 24730 11864
rect 24289 11716 24585 11736
rect 24345 11714 24369 11716
rect 24425 11714 24449 11716
rect 24505 11714 24529 11716
rect 24367 11662 24369 11714
rect 24431 11662 24443 11714
rect 24505 11662 24507 11714
rect 24345 11660 24369 11662
rect 24425 11660 24449 11662
rect 24505 11660 24529 11662
rect 24289 11640 24585 11660
rect 24688 11618 24716 11855
rect 24676 11612 24728 11618
rect 24676 11554 24728 11560
rect 24780 11074 24808 13510
rect 25608 12706 25636 14847
rect 25596 12700 25648 12706
rect 25596 12642 25648 12648
rect 25700 12366 25728 24503
rect 26160 20186 26188 27240
rect 26896 24577 26924 27240
rect 26882 24568 26938 24577
rect 26882 24503 26938 24512
rect 26148 20180 26200 20186
rect 26148 20122 26200 20128
rect 26332 17460 26384 17466
rect 26332 17402 26384 17408
rect 26344 17058 26372 17402
rect 26332 17052 26384 17058
rect 26332 16994 26384 17000
rect 27540 16990 27568 27240
rect 26240 16984 26292 16990
rect 26240 16926 26292 16932
rect 27528 16984 27580 16990
rect 27528 16926 27580 16932
rect 25688 12360 25740 12366
rect 25688 12302 25740 12308
rect 24768 11068 24820 11074
rect 24768 11010 24820 11016
rect 24676 10932 24728 10938
rect 24676 10874 24728 10880
rect 24688 10705 24716 10874
rect 24674 10696 24730 10705
rect 24289 10628 24585 10648
rect 24674 10631 24730 10640
rect 24345 10626 24369 10628
rect 24425 10626 24449 10628
rect 24505 10626 24529 10628
rect 24367 10574 24369 10626
rect 24431 10574 24443 10626
rect 24505 10574 24507 10626
rect 24345 10572 24369 10574
rect 24425 10572 24449 10574
rect 24505 10572 24529 10574
rect 24289 10552 24585 10572
rect 24688 10462 24716 10631
rect 24676 10456 24728 10462
rect 24676 10398 24728 10404
rect 24122 10288 24178 10297
rect 24122 10223 24178 10232
rect 23940 7260 23992 7266
rect 23940 7202 23992 7208
rect 23846 2400 23902 2409
rect 23846 2335 23902 2344
rect 23952 2137 23980 7202
rect 24136 4313 24164 10223
rect 25228 10184 25280 10190
rect 25226 10152 25228 10161
rect 25280 10152 25282 10161
rect 25226 10087 25282 10096
rect 24766 10016 24822 10025
rect 24766 9951 24768 9960
rect 24820 9951 24822 9960
rect 24768 9922 24820 9928
rect 24676 9844 24728 9850
rect 24676 9786 24728 9792
rect 24688 9617 24716 9786
rect 24674 9608 24730 9617
rect 24289 9540 24585 9560
rect 24674 9543 24730 9552
rect 25226 9608 25282 9617
rect 25226 9543 25282 9552
rect 24345 9538 24369 9540
rect 24425 9538 24449 9540
rect 24505 9538 24529 9540
rect 24367 9486 24369 9538
rect 24431 9486 24443 9538
rect 24505 9486 24507 9538
rect 24345 9484 24369 9486
rect 24425 9484 24449 9486
rect 24505 9484 24529 9486
rect 24289 9464 24585 9484
rect 25240 9374 25268 9543
rect 24768 9368 24820 9374
rect 24766 9336 24768 9345
rect 25228 9368 25280 9374
rect 24820 9336 24822 9345
rect 25228 9310 25280 9316
rect 24766 9271 24822 9280
rect 24492 9096 24544 9102
rect 24492 9038 24544 9044
rect 24766 9064 24822 9073
rect 24504 8937 24532 9038
rect 24766 8999 24822 9008
rect 24490 8928 24546 8937
rect 24780 8898 24808 8999
rect 24490 8863 24546 8872
rect 24768 8892 24820 8898
rect 24768 8834 24820 8840
rect 24676 8756 24728 8762
rect 24676 8698 24728 8704
rect 24289 8452 24585 8472
rect 24345 8450 24369 8452
rect 24425 8450 24449 8452
rect 24505 8450 24529 8452
rect 24367 8398 24369 8450
rect 24431 8398 24443 8450
rect 24505 8398 24507 8450
rect 24345 8396 24369 8398
rect 24425 8396 24449 8398
rect 24505 8396 24529 8398
rect 24289 8376 24585 8396
rect 24688 8393 24716 8698
rect 24674 8384 24730 8393
rect 24674 8319 24676 8328
rect 24728 8319 24730 8328
rect 24676 8290 24728 8296
rect 24214 7704 24270 7713
rect 24214 7639 24270 7648
rect 24582 7704 24638 7713
rect 24582 7639 24584 7648
rect 24228 6625 24256 7639
rect 24636 7639 24638 7648
rect 24584 7610 24636 7616
rect 24596 7554 24624 7610
rect 24766 7568 24822 7577
rect 24596 7526 24716 7554
rect 24289 7364 24585 7384
rect 24345 7362 24369 7364
rect 24425 7362 24449 7364
rect 24505 7362 24529 7364
rect 24367 7310 24369 7362
rect 24431 7310 24443 7362
rect 24505 7310 24507 7362
rect 24345 7308 24369 7310
rect 24425 7308 24449 7310
rect 24505 7308 24529 7310
rect 24289 7288 24585 7308
rect 24688 7266 24716 7526
rect 24766 7503 24768 7512
rect 24820 7503 24822 7512
rect 24768 7474 24820 7480
rect 24676 7260 24728 7266
rect 24676 7202 24728 7208
rect 24214 6616 24270 6625
rect 24214 6551 24270 6560
rect 24289 6276 24585 6296
rect 24345 6274 24369 6276
rect 24425 6274 24449 6276
rect 24505 6274 24529 6276
rect 24367 6222 24369 6274
rect 24431 6222 24443 6274
rect 24505 6222 24507 6274
rect 24345 6220 24369 6222
rect 24425 6220 24449 6222
rect 24505 6220 24529 6222
rect 24289 6200 24585 6220
rect 24289 5188 24585 5208
rect 24345 5186 24369 5188
rect 24425 5186 24449 5188
rect 24505 5186 24529 5188
rect 24367 5134 24369 5186
rect 24431 5134 24443 5186
rect 24505 5134 24507 5186
rect 24345 5132 24369 5134
rect 24425 5132 24449 5134
rect 24505 5132 24529 5134
rect 24289 5112 24585 5132
rect 24122 4304 24178 4313
rect 24122 4239 24178 4248
rect 24289 4100 24585 4120
rect 24345 4098 24369 4100
rect 24425 4098 24449 4100
rect 24505 4098 24529 4100
rect 24367 4046 24369 4098
rect 24431 4046 24443 4098
rect 24505 4046 24507 4098
rect 24345 4044 24369 4046
rect 24425 4044 24449 4046
rect 24505 4044 24529 4046
rect 24289 4024 24585 4044
rect 26252 3769 26280 16926
rect 24766 3760 24822 3769
rect 24766 3695 24822 3704
rect 26238 3760 26294 3769
rect 26238 3695 26294 3704
rect 24780 3662 24808 3695
rect 24768 3656 24820 3662
rect 25228 3656 25280 3662
rect 24768 3598 24820 3604
rect 25226 3624 25228 3633
rect 25280 3624 25282 3633
rect 25226 3559 25282 3568
rect 24289 3012 24585 3032
rect 24345 3010 24369 3012
rect 24425 3010 24449 3012
rect 24505 3010 24529 3012
rect 24367 2958 24369 3010
rect 24431 2958 24443 3010
rect 24505 2958 24507 3010
rect 24345 2956 24369 2958
rect 24425 2956 24449 2958
rect 24505 2956 24529 2958
rect 24289 2936 24585 2956
rect 23938 2128 23994 2137
rect 23938 2063 23994 2072
rect 24289 1924 24585 1944
rect 24345 1922 24369 1924
rect 24425 1922 24449 1924
rect 24505 1922 24529 1924
rect 24367 1870 24369 1922
rect 24431 1870 24443 1922
rect 24505 1870 24507 1922
rect 24345 1868 24369 1870
rect 24425 1868 24449 1870
rect 24505 1868 24529 1870
rect 24289 1848 24585 1868
rect 23662 632 23718 641
rect 23662 567 23718 576
rect 23570 88 23626 97
rect 23570 23 23626 32
<< via2 >>
rect 23938 27368 23994 27424
rect 1582 16760 1638 16816
rect 5622 24770 5678 24772
rect 5702 24770 5758 24772
rect 5782 24770 5838 24772
rect 5862 24770 5918 24772
rect 5622 24718 5648 24770
rect 5648 24718 5678 24770
rect 5702 24718 5712 24770
rect 5712 24718 5758 24770
rect 5782 24718 5828 24770
rect 5828 24718 5838 24770
rect 5862 24718 5892 24770
rect 5892 24718 5918 24770
rect 5622 24716 5678 24718
rect 5702 24716 5758 24718
rect 5782 24716 5838 24718
rect 5862 24716 5918 24718
rect 4986 23968 5042 24024
rect 5622 23682 5678 23684
rect 5702 23682 5758 23684
rect 5782 23682 5838 23684
rect 5862 23682 5918 23684
rect 5622 23630 5648 23682
rect 5648 23630 5678 23682
rect 5702 23630 5712 23682
rect 5712 23630 5758 23682
rect 5782 23630 5828 23682
rect 5828 23630 5838 23682
rect 5862 23630 5892 23682
rect 5892 23630 5918 23682
rect 5622 23628 5678 23630
rect 5702 23628 5758 23630
rect 5782 23628 5838 23630
rect 5862 23628 5918 23630
rect 5622 22594 5678 22596
rect 5702 22594 5758 22596
rect 5782 22594 5838 22596
rect 5862 22594 5918 22596
rect 5622 22542 5648 22594
rect 5648 22542 5678 22594
rect 5702 22542 5712 22594
rect 5712 22542 5758 22594
rect 5782 22542 5828 22594
rect 5828 22542 5838 22594
rect 5862 22542 5892 22594
rect 5892 22542 5918 22594
rect 5622 22540 5678 22542
rect 5702 22540 5758 22542
rect 5782 22540 5838 22542
rect 5862 22540 5918 22542
rect 5622 21506 5678 21508
rect 5702 21506 5758 21508
rect 5782 21506 5838 21508
rect 5862 21506 5918 21508
rect 5622 21454 5648 21506
rect 5648 21454 5678 21506
rect 5702 21454 5712 21506
rect 5712 21454 5758 21506
rect 5782 21454 5828 21506
rect 5828 21454 5838 21506
rect 5862 21454 5892 21506
rect 5892 21454 5918 21506
rect 5622 21452 5678 21454
rect 5702 21452 5758 21454
rect 5782 21452 5838 21454
rect 5862 21452 5918 21454
rect 7746 22336 7802 22392
rect 7102 21520 7158 21576
rect 6366 21248 6422 21304
rect 5998 21112 6054 21168
rect 4342 20840 4398 20896
rect 9218 22764 9274 22800
rect 9218 22744 9220 22764
rect 9220 22744 9272 22764
rect 9272 22744 9274 22764
rect 10289 25314 10345 25316
rect 10369 25314 10425 25316
rect 10449 25314 10505 25316
rect 10529 25314 10585 25316
rect 10289 25262 10315 25314
rect 10315 25262 10345 25314
rect 10369 25262 10379 25314
rect 10379 25262 10425 25314
rect 10449 25262 10495 25314
rect 10495 25262 10505 25314
rect 10529 25262 10559 25314
rect 10559 25262 10585 25314
rect 10289 25260 10345 25262
rect 10369 25260 10425 25262
rect 10449 25260 10505 25262
rect 10529 25260 10585 25262
rect 10289 24226 10345 24228
rect 10369 24226 10425 24228
rect 10449 24226 10505 24228
rect 10529 24226 10585 24228
rect 10289 24174 10315 24226
rect 10315 24174 10345 24226
rect 10369 24174 10379 24226
rect 10379 24174 10425 24226
rect 10449 24174 10495 24226
rect 10495 24174 10505 24226
rect 10529 24174 10559 24226
rect 10559 24174 10585 24226
rect 10289 24172 10345 24174
rect 10369 24172 10425 24174
rect 10449 24172 10505 24174
rect 10529 24172 10585 24174
rect 10289 23138 10345 23140
rect 10369 23138 10425 23140
rect 10449 23138 10505 23140
rect 10529 23138 10585 23140
rect 10289 23086 10315 23138
rect 10315 23086 10345 23138
rect 10369 23086 10379 23138
rect 10379 23086 10425 23138
rect 10449 23086 10495 23138
rect 10495 23086 10505 23138
rect 10529 23086 10559 23138
rect 10559 23086 10585 23138
rect 10289 23084 10345 23086
rect 10369 23084 10425 23086
rect 10449 23084 10505 23086
rect 10529 23084 10585 23086
rect 9770 22472 9826 22528
rect 10138 22880 10194 22936
rect 10874 23152 10930 23208
rect 11150 23560 11206 23616
rect 10289 22050 10345 22052
rect 10369 22050 10425 22052
rect 10449 22050 10505 22052
rect 10529 22050 10585 22052
rect 10289 21998 10315 22050
rect 10315 21998 10345 22050
rect 10369 21998 10379 22050
rect 10379 21998 10425 22050
rect 10449 21998 10495 22050
rect 10495 21998 10505 22050
rect 10529 21998 10559 22050
rect 10559 21998 10585 22050
rect 10289 21996 10345 21998
rect 10369 21996 10425 21998
rect 10449 21996 10505 21998
rect 10529 21996 10585 21998
rect 13634 24512 13690 24568
rect 13174 24376 13230 24432
rect 12530 24240 12586 24296
rect 13358 23580 13414 23616
rect 13358 23560 13360 23580
rect 13360 23560 13412 23580
rect 13412 23560 13414 23580
rect 10289 20962 10345 20964
rect 10369 20962 10425 20964
rect 10449 20962 10505 20964
rect 10529 20962 10585 20964
rect 10289 20910 10315 20962
rect 10315 20910 10345 20962
rect 10369 20910 10379 20962
rect 10379 20910 10425 20962
rect 10449 20910 10495 20962
rect 10495 20910 10505 20962
rect 10529 20910 10559 20962
rect 10559 20910 10585 20962
rect 10289 20908 10345 20910
rect 10369 20908 10425 20910
rect 10449 20908 10505 20910
rect 10529 20908 10585 20910
rect 10690 20860 10746 20896
rect 10690 20840 10692 20860
rect 10692 20840 10744 20860
rect 10744 20840 10746 20860
rect 9218 20704 9274 20760
rect 9126 20568 9182 20624
rect 8390 20432 8446 20488
rect 5622 20418 5678 20420
rect 5702 20418 5758 20420
rect 5782 20418 5838 20420
rect 5862 20418 5918 20420
rect 5622 20366 5648 20418
rect 5648 20366 5678 20418
rect 5702 20366 5712 20418
rect 5712 20366 5758 20418
rect 5782 20366 5828 20418
rect 5828 20366 5838 20418
rect 5862 20366 5892 20418
rect 5892 20366 5918 20418
rect 5622 20364 5678 20366
rect 5702 20364 5758 20366
rect 5782 20364 5838 20366
rect 5862 20364 5918 20366
rect 13542 22200 13598 22256
rect 11242 21248 11298 21304
rect 10690 19924 10692 19944
rect 10692 19924 10744 19944
rect 10744 19924 10746 19944
rect 10690 19888 10746 19924
rect 11150 19888 11206 19944
rect 10289 19874 10345 19876
rect 10369 19874 10425 19876
rect 10449 19874 10505 19876
rect 10529 19874 10585 19876
rect 10289 19822 10315 19874
rect 10315 19822 10345 19874
rect 10369 19822 10379 19874
rect 10379 19822 10425 19874
rect 10449 19822 10495 19874
rect 10495 19822 10505 19874
rect 10529 19822 10559 19874
rect 10559 19822 10585 19874
rect 10289 19820 10345 19822
rect 10369 19820 10425 19822
rect 10449 19820 10505 19822
rect 10529 19820 10585 19822
rect 13358 20432 13414 20488
rect 5622 19330 5678 19332
rect 5702 19330 5758 19332
rect 5782 19330 5838 19332
rect 5862 19330 5918 19332
rect 5622 19278 5648 19330
rect 5648 19278 5678 19330
rect 5702 19278 5712 19330
rect 5712 19278 5758 19330
rect 5782 19278 5828 19330
rect 5828 19278 5838 19330
rect 5862 19278 5892 19330
rect 5892 19278 5918 19330
rect 5622 19276 5678 19278
rect 5702 19276 5758 19278
rect 5782 19276 5838 19278
rect 5862 19276 5918 19278
rect 3698 18936 3754 18992
rect 10289 18786 10345 18788
rect 10369 18786 10425 18788
rect 10449 18786 10505 18788
rect 10529 18786 10585 18788
rect 10289 18734 10315 18786
rect 10315 18734 10345 18786
rect 10369 18734 10379 18786
rect 10379 18734 10425 18786
rect 10449 18734 10495 18786
rect 10495 18734 10505 18786
rect 10529 18734 10559 18786
rect 10559 18734 10585 18786
rect 10289 18732 10345 18734
rect 10369 18732 10425 18734
rect 10449 18732 10505 18734
rect 10529 18732 10585 18734
rect 2962 18528 3018 18584
rect 13542 18800 13598 18856
rect 5622 18242 5678 18244
rect 5702 18242 5758 18244
rect 5782 18242 5838 18244
rect 5862 18242 5918 18244
rect 5622 18190 5648 18242
rect 5648 18190 5678 18242
rect 5702 18190 5712 18242
rect 5712 18190 5758 18242
rect 5782 18190 5828 18242
rect 5828 18190 5838 18242
rect 5862 18190 5892 18242
rect 5892 18190 5918 18242
rect 5622 18188 5678 18190
rect 5702 18188 5758 18190
rect 5782 18188 5838 18190
rect 5862 18188 5918 18190
rect 10289 17698 10345 17700
rect 10369 17698 10425 17700
rect 10449 17698 10505 17700
rect 10529 17698 10585 17700
rect 10289 17646 10315 17698
rect 10315 17646 10345 17698
rect 10369 17646 10379 17698
rect 10379 17646 10425 17698
rect 10449 17646 10495 17698
rect 10495 17646 10505 17698
rect 10529 17646 10559 17698
rect 10559 17646 10585 17698
rect 10289 17644 10345 17646
rect 10369 17644 10425 17646
rect 10449 17644 10505 17646
rect 10529 17644 10585 17646
rect 5622 17154 5678 17156
rect 5702 17154 5758 17156
rect 5782 17154 5838 17156
rect 5862 17154 5918 17156
rect 5622 17102 5648 17154
rect 5648 17102 5678 17154
rect 5702 17102 5712 17154
rect 5712 17102 5758 17154
rect 5782 17102 5828 17154
rect 5828 17102 5838 17154
rect 5862 17102 5892 17154
rect 5892 17102 5918 17154
rect 5622 17100 5678 17102
rect 5702 17100 5758 17102
rect 5782 17100 5838 17102
rect 5862 17100 5918 17102
rect 11886 16780 11942 16816
rect 11886 16760 11888 16780
rect 11888 16760 11940 16780
rect 11940 16760 11942 16780
rect 10289 16610 10345 16612
rect 10369 16610 10425 16612
rect 10449 16610 10505 16612
rect 10529 16610 10585 16612
rect 10289 16558 10315 16610
rect 10315 16558 10345 16610
rect 10369 16558 10379 16610
rect 10379 16558 10425 16610
rect 10449 16558 10495 16610
rect 10495 16558 10505 16610
rect 10529 16558 10559 16610
rect 10559 16558 10585 16610
rect 10289 16556 10345 16558
rect 10369 16556 10425 16558
rect 10449 16556 10505 16558
rect 10529 16556 10585 16558
rect 2318 16352 2374 16408
rect 1306 16216 1362 16272
rect 5622 16066 5678 16068
rect 5702 16066 5758 16068
rect 5782 16066 5838 16068
rect 5862 16066 5918 16068
rect 5622 16014 5648 16066
rect 5648 16014 5678 16066
rect 5702 16014 5712 16066
rect 5712 16014 5758 16066
rect 5782 16014 5828 16066
rect 5828 16014 5838 16066
rect 5862 16014 5892 16066
rect 5892 16014 5918 16066
rect 5622 16012 5678 16014
rect 5702 16012 5758 16014
rect 5782 16012 5838 16014
rect 5862 16012 5918 16014
rect 10289 15522 10345 15524
rect 10369 15522 10425 15524
rect 10449 15522 10505 15524
rect 10529 15522 10585 15524
rect 10289 15470 10315 15522
rect 10315 15470 10345 15522
rect 10369 15470 10379 15522
rect 10379 15470 10425 15522
rect 10449 15470 10495 15522
rect 10495 15470 10505 15522
rect 10529 15470 10559 15522
rect 10559 15470 10585 15522
rect 10289 15468 10345 15470
rect 10369 15468 10425 15470
rect 10449 15468 10505 15470
rect 10529 15468 10585 15470
rect 5622 14978 5678 14980
rect 5702 14978 5758 14980
rect 5782 14978 5838 14980
rect 5862 14978 5918 14980
rect 5622 14926 5648 14978
rect 5648 14926 5678 14978
rect 5702 14926 5712 14978
rect 5712 14926 5758 14978
rect 5782 14926 5828 14978
rect 5828 14926 5838 14978
rect 5862 14926 5892 14978
rect 5892 14926 5918 14978
rect 5622 14924 5678 14926
rect 5702 14924 5758 14926
rect 5782 14924 5838 14926
rect 5862 14924 5918 14926
rect 12714 15128 12770 15184
rect 10289 14434 10345 14436
rect 10369 14434 10425 14436
rect 10449 14434 10505 14436
rect 10529 14434 10585 14436
rect 10289 14382 10315 14434
rect 10315 14382 10345 14434
rect 10369 14382 10379 14434
rect 10379 14382 10425 14434
rect 10449 14382 10495 14434
rect 10495 14382 10505 14434
rect 10529 14382 10559 14434
rect 10559 14382 10585 14434
rect 10289 14380 10345 14382
rect 10369 14380 10425 14382
rect 10449 14380 10505 14382
rect 10529 14380 10585 14382
rect 5622 13890 5678 13892
rect 5702 13890 5758 13892
rect 5782 13890 5838 13892
rect 5862 13890 5918 13892
rect 5622 13838 5648 13890
rect 5648 13838 5678 13890
rect 5702 13838 5712 13890
rect 5712 13838 5758 13890
rect 5782 13838 5828 13890
rect 5828 13838 5838 13890
rect 5862 13838 5892 13890
rect 5892 13838 5918 13890
rect 5622 13836 5678 13838
rect 5702 13836 5758 13838
rect 5782 13836 5838 13838
rect 5862 13836 5918 13838
rect 10289 13346 10345 13348
rect 10369 13346 10425 13348
rect 10449 13346 10505 13348
rect 10529 13346 10585 13348
rect 10289 13294 10315 13346
rect 10315 13294 10345 13346
rect 10369 13294 10379 13346
rect 10379 13294 10425 13346
rect 10449 13294 10495 13346
rect 10495 13294 10505 13346
rect 10529 13294 10559 13346
rect 10559 13294 10585 13346
rect 10289 13292 10345 13294
rect 10369 13292 10425 13294
rect 10449 13292 10505 13294
rect 10529 13292 10585 13294
rect 5622 12802 5678 12804
rect 5702 12802 5758 12804
rect 5782 12802 5838 12804
rect 5862 12802 5918 12804
rect 5622 12750 5648 12802
rect 5648 12750 5678 12802
rect 5702 12750 5712 12802
rect 5712 12750 5758 12802
rect 5782 12750 5828 12802
rect 5828 12750 5838 12802
rect 5862 12750 5892 12802
rect 5892 12750 5918 12802
rect 5622 12748 5678 12750
rect 5702 12748 5758 12750
rect 5782 12748 5838 12750
rect 5862 12748 5918 12750
rect 10289 12258 10345 12260
rect 10369 12258 10425 12260
rect 10449 12258 10505 12260
rect 10529 12258 10585 12260
rect 10289 12206 10315 12258
rect 10315 12206 10345 12258
rect 10369 12206 10379 12258
rect 10379 12206 10425 12258
rect 10449 12206 10495 12258
rect 10495 12206 10505 12258
rect 10529 12206 10559 12258
rect 10559 12206 10585 12258
rect 10289 12204 10345 12206
rect 10369 12204 10425 12206
rect 10449 12204 10505 12206
rect 10529 12204 10585 12206
rect 5622 11714 5678 11716
rect 5702 11714 5758 11716
rect 5782 11714 5838 11716
rect 5862 11714 5918 11716
rect 5622 11662 5648 11714
rect 5648 11662 5678 11714
rect 5702 11662 5712 11714
rect 5712 11662 5758 11714
rect 5782 11662 5828 11714
rect 5828 11662 5838 11714
rect 5862 11662 5892 11714
rect 5892 11662 5918 11714
rect 5622 11660 5678 11662
rect 5702 11660 5758 11662
rect 5782 11660 5838 11662
rect 5862 11660 5918 11662
rect 14956 24770 15012 24772
rect 15036 24770 15092 24772
rect 15116 24770 15172 24772
rect 15196 24770 15252 24772
rect 14956 24718 14982 24770
rect 14982 24718 15012 24770
rect 15036 24718 15046 24770
rect 15046 24718 15092 24770
rect 15116 24718 15162 24770
rect 15162 24718 15172 24770
rect 15196 24718 15226 24770
rect 15226 24718 15252 24770
rect 14956 24716 15012 24718
rect 15036 24716 15092 24718
rect 15116 24716 15172 24718
rect 15196 24716 15252 24718
rect 14554 24512 14610 24568
rect 14830 23832 14886 23888
rect 14956 23682 15012 23684
rect 15036 23682 15092 23684
rect 15116 23682 15172 23684
rect 15196 23682 15252 23684
rect 14956 23630 14982 23682
rect 14982 23630 15012 23682
rect 15036 23630 15046 23682
rect 15046 23630 15092 23682
rect 15116 23630 15162 23682
rect 15162 23630 15172 23682
rect 15196 23630 15226 23682
rect 15226 23630 15252 23682
rect 14956 23628 15012 23630
rect 15036 23628 15092 23630
rect 15116 23628 15172 23630
rect 15196 23628 15252 23630
rect 14094 23152 14150 23208
rect 14738 23152 14794 23208
rect 14738 22492 14794 22528
rect 14738 22472 14740 22492
rect 14740 22472 14792 22492
rect 14792 22472 14794 22492
rect 14186 21268 14242 21304
rect 14186 21248 14188 21268
rect 14188 21248 14240 21268
rect 14240 21248 14242 21268
rect 14002 20044 14058 20080
rect 14002 20024 14004 20044
rect 14004 20024 14056 20044
rect 14056 20024 14058 20044
rect 13910 19072 13966 19128
rect 14094 17324 14150 17360
rect 14094 17304 14096 17324
rect 14096 17304 14148 17324
rect 14148 17304 14150 17324
rect 14002 16796 14004 16816
rect 14004 16796 14056 16816
rect 14056 16796 14058 16816
rect 14002 16760 14058 16796
rect 14956 22594 15012 22596
rect 15036 22594 15092 22596
rect 15116 22594 15172 22596
rect 15196 22594 15252 22596
rect 14956 22542 14982 22594
rect 14982 22542 15012 22594
rect 15036 22542 15046 22594
rect 15046 22542 15092 22594
rect 15116 22542 15162 22594
rect 15162 22542 15172 22594
rect 15196 22542 15226 22594
rect 15226 22542 15252 22594
rect 14956 22540 15012 22542
rect 15036 22540 15092 22542
rect 15116 22540 15172 22542
rect 15196 22540 15252 22542
rect 14956 21506 15012 21508
rect 15036 21506 15092 21508
rect 15116 21506 15172 21508
rect 15196 21506 15252 21508
rect 14956 21454 14982 21506
rect 14982 21454 15012 21506
rect 15036 21454 15046 21506
rect 15046 21454 15092 21506
rect 15116 21454 15162 21506
rect 15162 21454 15172 21506
rect 15196 21454 15226 21506
rect 15226 21454 15252 21506
rect 14956 21452 15012 21454
rect 15036 21452 15092 21454
rect 15116 21452 15172 21454
rect 15196 21452 15252 21454
rect 14956 20418 15012 20420
rect 15036 20418 15092 20420
rect 15116 20418 15172 20420
rect 15196 20418 15252 20420
rect 14956 20366 14982 20418
rect 14982 20366 15012 20418
rect 15036 20366 15046 20418
rect 15046 20366 15092 20418
rect 15116 20366 15162 20418
rect 15162 20366 15172 20418
rect 15196 20366 15226 20418
rect 15226 20366 15252 20418
rect 14956 20364 15012 20366
rect 15036 20364 15092 20366
rect 15116 20364 15172 20366
rect 15196 20364 15252 20366
rect 14956 19330 15012 19332
rect 15036 19330 15092 19332
rect 15116 19330 15172 19332
rect 15196 19330 15252 19332
rect 14956 19278 14982 19330
rect 14982 19278 15012 19330
rect 15036 19278 15046 19330
rect 15046 19278 15092 19330
rect 15116 19278 15162 19330
rect 15162 19278 15172 19330
rect 15196 19278 15226 19330
rect 15226 19278 15252 19330
rect 14956 19276 15012 19278
rect 15036 19276 15092 19278
rect 15116 19276 15172 19278
rect 15196 19276 15252 19278
rect 14956 18242 15012 18244
rect 15036 18242 15092 18244
rect 15116 18242 15172 18244
rect 15196 18242 15252 18244
rect 14956 18190 14982 18242
rect 14982 18190 15012 18242
rect 15036 18190 15046 18242
rect 15046 18190 15092 18242
rect 15116 18190 15162 18242
rect 15162 18190 15172 18242
rect 15196 18190 15226 18242
rect 15226 18190 15252 18242
rect 14956 18188 15012 18190
rect 15036 18188 15092 18190
rect 15116 18188 15172 18190
rect 15196 18188 15252 18190
rect 14956 17154 15012 17156
rect 15036 17154 15092 17156
rect 15116 17154 15172 17156
rect 15196 17154 15252 17156
rect 14956 17102 14982 17154
rect 14982 17102 15012 17154
rect 15036 17102 15046 17154
rect 15046 17102 15092 17154
rect 15116 17102 15162 17154
rect 15162 17102 15172 17154
rect 15196 17102 15226 17154
rect 15226 17102 15252 17154
rect 14956 17100 15012 17102
rect 15036 17100 15092 17102
rect 15116 17100 15172 17102
rect 15196 17100 15252 17102
rect 14956 16066 15012 16068
rect 15036 16066 15092 16068
rect 15116 16066 15172 16068
rect 15196 16066 15252 16068
rect 14956 16014 14982 16066
rect 14982 16014 15012 16066
rect 15036 16014 15046 16066
rect 15046 16014 15092 16066
rect 15116 16014 15162 16066
rect 15162 16014 15172 16066
rect 15196 16014 15226 16066
rect 15226 16014 15252 16066
rect 14956 16012 15012 16014
rect 15036 16012 15092 16014
rect 15116 16012 15172 16014
rect 15196 16012 15252 16014
rect 14956 14978 15012 14980
rect 15036 14978 15092 14980
rect 15116 14978 15172 14980
rect 15196 14978 15252 14980
rect 14956 14926 14982 14978
rect 14982 14926 15012 14978
rect 15036 14926 15046 14978
rect 15046 14926 15092 14978
rect 15116 14926 15162 14978
rect 15162 14926 15172 14978
rect 15196 14926 15226 14978
rect 15226 14926 15252 14978
rect 14956 14924 15012 14926
rect 15036 14924 15092 14926
rect 15116 14924 15172 14926
rect 15196 14924 15252 14926
rect 14956 13890 15012 13892
rect 15036 13890 15092 13892
rect 15116 13890 15172 13892
rect 15196 13890 15252 13892
rect 14956 13838 14982 13890
rect 14982 13838 15012 13890
rect 15036 13838 15046 13890
rect 15046 13838 15092 13890
rect 15116 13838 15162 13890
rect 15162 13838 15172 13890
rect 15196 13838 15226 13890
rect 15226 13838 15252 13890
rect 14956 13836 15012 13838
rect 15036 13836 15092 13838
rect 15116 13836 15172 13838
rect 15196 13836 15252 13838
rect 16118 22644 16120 22664
rect 16120 22644 16172 22664
rect 16172 22644 16174 22664
rect 16118 22608 16174 22644
rect 16118 20604 16120 20624
rect 16120 20604 16172 20624
rect 16172 20604 16174 20624
rect 16118 20568 16174 20604
rect 14956 12802 15012 12804
rect 15036 12802 15092 12804
rect 15116 12802 15172 12804
rect 15196 12802 15252 12804
rect 14956 12750 14982 12802
rect 14982 12750 15012 12802
rect 15036 12750 15046 12802
rect 15046 12750 15092 12802
rect 15116 12750 15162 12802
rect 15162 12750 15172 12802
rect 15196 12750 15226 12802
rect 15226 12750 15252 12802
rect 14956 12748 15012 12750
rect 15036 12748 15092 12750
rect 15116 12748 15172 12750
rect 15196 12748 15252 12750
rect 10289 11170 10345 11172
rect 10369 11170 10425 11172
rect 10449 11170 10505 11172
rect 10529 11170 10585 11172
rect 10289 11118 10315 11170
rect 10315 11118 10345 11170
rect 10369 11118 10379 11170
rect 10379 11118 10425 11170
rect 10449 11118 10495 11170
rect 10495 11118 10505 11170
rect 10529 11118 10559 11170
rect 10559 11118 10585 11170
rect 10289 11116 10345 11118
rect 10369 11116 10425 11118
rect 10449 11116 10505 11118
rect 10529 11116 10585 11118
rect 5622 10626 5678 10628
rect 5702 10626 5758 10628
rect 5782 10626 5838 10628
rect 5862 10626 5918 10628
rect 5622 10574 5648 10626
rect 5648 10574 5678 10626
rect 5702 10574 5712 10626
rect 5712 10574 5758 10626
rect 5782 10574 5828 10626
rect 5828 10574 5838 10626
rect 5862 10574 5892 10626
rect 5892 10574 5918 10626
rect 5622 10572 5678 10574
rect 5702 10572 5758 10574
rect 5782 10572 5838 10574
rect 5862 10572 5918 10574
rect 14956 11714 15012 11716
rect 15036 11714 15092 11716
rect 15116 11714 15172 11716
rect 15196 11714 15252 11716
rect 14956 11662 14982 11714
rect 14982 11662 15012 11714
rect 15036 11662 15046 11714
rect 15046 11662 15092 11714
rect 15116 11662 15162 11714
rect 15162 11662 15172 11714
rect 15196 11662 15226 11714
rect 15226 11662 15252 11714
rect 14956 11660 15012 11662
rect 15036 11660 15092 11662
rect 15116 11660 15172 11662
rect 15196 11660 15252 11662
rect 14956 10626 15012 10628
rect 15036 10626 15092 10628
rect 15116 10626 15172 10628
rect 15196 10626 15252 10628
rect 14956 10574 14982 10626
rect 14982 10574 15012 10626
rect 15036 10574 15046 10626
rect 15046 10574 15092 10626
rect 15116 10574 15162 10626
rect 15162 10574 15172 10626
rect 15196 10574 15226 10626
rect 15226 10574 15252 10626
rect 14956 10572 15012 10574
rect 15036 10572 15092 10574
rect 15116 10572 15172 10574
rect 15196 10572 15252 10574
rect 3422 10232 3478 10288
rect 10782 10252 10838 10288
rect 10782 10232 10784 10252
rect 10784 10232 10836 10252
rect 10836 10232 10838 10252
rect 202 9688 258 9744
rect 10289 10082 10345 10084
rect 10369 10082 10425 10084
rect 10449 10082 10505 10084
rect 10529 10082 10585 10084
rect 10289 10030 10315 10082
rect 10315 10030 10345 10082
rect 10369 10030 10379 10082
rect 10379 10030 10425 10082
rect 10449 10030 10495 10082
rect 10495 10030 10505 10082
rect 10529 10030 10559 10082
rect 10559 10030 10585 10082
rect 10289 10028 10345 10030
rect 10369 10028 10425 10030
rect 10449 10028 10505 10030
rect 10529 10028 10585 10030
rect 13818 10252 13874 10288
rect 13818 10232 13820 10252
rect 13820 10232 13872 10252
rect 13872 10232 13874 10252
rect 13910 9688 13966 9744
rect 5622 9538 5678 9540
rect 5702 9538 5758 9540
rect 5782 9538 5838 9540
rect 5862 9538 5918 9540
rect 5622 9486 5648 9538
rect 5648 9486 5678 9538
rect 5702 9486 5712 9538
rect 5712 9486 5758 9538
rect 5782 9486 5828 9538
rect 5828 9486 5838 9538
rect 5862 9486 5892 9538
rect 5892 9486 5918 9538
rect 5622 9484 5678 9486
rect 5702 9484 5758 9486
rect 5782 9484 5838 9486
rect 5862 9484 5918 9486
rect 14956 9538 15012 9540
rect 15036 9538 15092 9540
rect 15116 9538 15172 9540
rect 15196 9538 15252 9540
rect 14956 9486 14982 9538
rect 14982 9486 15012 9538
rect 15036 9486 15046 9538
rect 15046 9486 15092 9538
rect 15116 9486 15162 9538
rect 15162 9486 15172 9538
rect 15196 9486 15226 9538
rect 15226 9486 15252 9538
rect 14956 9484 15012 9486
rect 15036 9484 15092 9486
rect 15116 9484 15172 9486
rect 15196 9484 15252 9486
rect 10289 8994 10345 8996
rect 10369 8994 10425 8996
rect 10449 8994 10505 8996
rect 10529 8994 10585 8996
rect 10289 8942 10315 8994
rect 10315 8942 10345 8994
rect 10369 8942 10379 8994
rect 10379 8942 10425 8994
rect 10449 8942 10495 8994
rect 10495 8942 10505 8994
rect 10529 8942 10559 8994
rect 10559 8942 10585 8994
rect 10289 8940 10345 8942
rect 10369 8940 10425 8942
rect 10449 8940 10505 8942
rect 10529 8940 10585 8942
rect 5622 8450 5678 8452
rect 5702 8450 5758 8452
rect 5782 8450 5838 8452
rect 5862 8450 5918 8452
rect 5622 8398 5648 8450
rect 5648 8398 5678 8450
rect 5702 8398 5712 8450
rect 5712 8398 5758 8450
rect 5782 8398 5828 8450
rect 5828 8398 5838 8450
rect 5862 8398 5892 8450
rect 5892 8398 5918 8450
rect 5622 8396 5678 8398
rect 5702 8396 5758 8398
rect 5782 8396 5838 8398
rect 5862 8396 5918 8398
rect 14956 8450 15012 8452
rect 15036 8450 15092 8452
rect 15116 8450 15172 8452
rect 15196 8450 15252 8452
rect 14956 8398 14982 8450
rect 14982 8398 15012 8450
rect 15036 8398 15046 8450
rect 15046 8398 15092 8450
rect 15116 8398 15162 8450
rect 15162 8398 15172 8450
rect 15196 8398 15226 8450
rect 15226 8398 15252 8450
rect 14956 8396 15012 8398
rect 15036 8396 15092 8398
rect 15116 8396 15172 8398
rect 15196 8396 15252 8398
rect 10289 7906 10345 7908
rect 10369 7906 10425 7908
rect 10449 7906 10505 7908
rect 10529 7906 10585 7908
rect 10289 7854 10315 7906
rect 10315 7854 10345 7906
rect 10369 7854 10379 7906
rect 10379 7854 10425 7906
rect 10449 7854 10495 7906
rect 10495 7854 10505 7906
rect 10529 7854 10559 7906
rect 10559 7854 10585 7906
rect 10289 7852 10345 7854
rect 10369 7852 10425 7854
rect 10449 7852 10505 7854
rect 10529 7852 10585 7854
rect 5622 7362 5678 7364
rect 5702 7362 5758 7364
rect 5782 7362 5838 7364
rect 5862 7362 5918 7364
rect 5622 7310 5648 7362
rect 5648 7310 5678 7362
rect 5702 7310 5712 7362
rect 5712 7310 5758 7362
rect 5782 7310 5828 7362
rect 5828 7310 5838 7362
rect 5862 7310 5892 7362
rect 5892 7310 5918 7362
rect 5622 7308 5678 7310
rect 5702 7308 5758 7310
rect 5782 7308 5838 7310
rect 5862 7308 5918 7310
rect 14956 7362 15012 7364
rect 15036 7362 15092 7364
rect 15116 7362 15172 7364
rect 15196 7362 15252 7364
rect 14956 7310 14982 7362
rect 14982 7310 15012 7362
rect 15036 7310 15046 7362
rect 15046 7310 15092 7362
rect 15116 7310 15162 7362
rect 15162 7310 15172 7362
rect 15196 7310 15226 7362
rect 15226 7310 15252 7362
rect 14956 7308 15012 7310
rect 15036 7308 15092 7310
rect 15116 7308 15172 7310
rect 15196 7308 15252 7310
rect 10289 6818 10345 6820
rect 10369 6818 10425 6820
rect 10449 6818 10505 6820
rect 10529 6818 10585 6820
rect 10289 6766 10315 6818
rect 10315 6766 10345 6818
rect 10369 6766 10379 6818
rect 10379 6766 10425 6818
rect 10449 6766 10495 6818
rect 10495 6766 10505 6818
rect 10529 6766 10559 6818
rect 10559 6766 10585 6818
rect 10289 6764 10345 6766
rect 10369 6764 10425 6766
rect 10449 6764 10505 6766
rect 10529 6764 10585 6766
rect 3422 6696 3478 6752
rect 5622 6274 5678 6276
rect 5702 6274 5758 6276
rect 5782 6274 5838 6276
rect 5862 6274 5918 6276
rect 5622 6222 5648 6274
rect 5648 6222 5678 6274
rect 5702 6222 5712 6274
rect 5712 6222 5758 6274
rect 5782 6222 5828 6274
rect 5828 6222 5838 6274
rect 5862 6222 5892 6274
rect 5892 6222 5918 6274
rect 5622 6220 5678 6222
rect 5702 6220 5758 6222
rect 5782 6220 5838 6222
rect 5862 6220 5918 6222
rect 14956 6274 15012 6276
rect 15036 6274 15092 6276
rect 15116 6274 15172 6276
rect 15196 6274 15252 6276
rect 14956 6222 14982 6274
rect 14982 6222 15012 6274
rect 15036 6222 15046 6274
rect 15046 6222 15092 6274
rect 15116 6222 15162 6274
rect 15162 6222 15172 6274
rect 15196 6222 15226 6274
rect 15226 6222 15252 6274
rect 14956 6220 15012 6222
rect 15036 6220 15092 6222
rect 15116 6220 15172 6222
rect 15196 6220 15252 6222
rect 10289 5730 10345 5732
rect 10369 5730 10425 5732
rect 10449 5730 10505 5732
rect 10529 5730 10585 5732
rect 10289 5678 10315 5730
rect 10315 5678 10345 5730
rect 10369 5678 10379 5730
rect 10379 5678 10425 5730
rect 10449 5678 10495 5730
rect 10495 5678 10505 5730
rect 10529 5678 10559 5730
rect 10559 5678 10585 5730
rect 10289 5676 10345 5678
rect 10369 5676 10425 5678
rect 10449 5676 10505 5678
rect 10529 5676 10585 5678
rect 5622 5186 5678 5188
rect 5702 5186 5758 5188
rect 5782 5186 5838 5188
rect 5862 5186 5918 5188
rect 5622 5134 5648 5186
rect 5648 5134 5678 5186
rect 5702 5134 5712 5186
rect 5712 5134 5758 5186
rect 5782 5134 5828 5186
rect 5828 5134 5838 5186
rect 5862 5134 5892 5186
rect 5892 5134 5918 5186
rect 5622 5132 5678 5134
rect 5702 5132 5758 5134
rect 5782 5132 5838 5134
rect 5862 5132 5918 5134
rect 14956 5186 15012 5188
rect 15036 5186 15092 5188
rect 15116 5186 15172 5188
rect 15196 5186 15252 5188
rect 14956 5134 14982 5186
rect 14982 5134 15012 5186
rect 15036 5134 15046 5186
rect 15046 5134 15092 5186
rect 15116 5134 15162 5186
rect 15162 5134 15172 5186
rect 15196 5134 15226 5186
rect 15226 5134 15252 5186
rect 14956 5132 15012 5134
rect 15036 5132 15092 5134
rect 15116 5132 15172 5134
rect 15196 5132 15252 5134
rect 15934 16760 15990 16816
rect 15842 16388 15844 16408
rect 15844 16388 15896 16408
rect 15896 16388 15898 16408
rect 15842 16352 15898 16388
rect 16394 16216 16450 16272
rect 16302 15708 16304 15728
rect 16304 15708 16356 15728
rect 16356 15708 16358 15728
rect 16302 15672 16358 15708
rect 16394 9436 16450 9472
rect 16394 9416 16396 9436
rect 16396 9416 16448 9436
rect 16448 9416 16450 9436
rect 17038 18664 17094 18720
rect 17590 19888 17646 19944
rect 16946 15164 16948 15184
rect 16948 15164 17000 15184
rect 17000 15164 17002 15184
rect 16946 15128 17002 15164
rect 17130 15828 17186 15864
rect 17130 15808 17132 15828
rect 17132 15808 17184 15828
rect 17184 15808 17186 15828
rect 16946 13768 17002 13824
rect 17774 13652 17830 13688
rect 17774 13632 17776 13652
rect 17776 13632 17828 13652
rect 17828 13632 17830 13652
rect 17498 13532 17500 13552
rect 17500 13532 17552 13552
rect 17552 13532 17554 13552
rect 17498 13496 17554 13532
rect 19622 25314 19678 25316
rect 19702 25314 19758 25316
rect 19782 25314 19838 25316
rect 19862 25314 19918 25316
rect 19622 25262 19648 25314
rect 19648 25262 19678 25314
rect 19702 25262 19712 25314
rect 19712 25262 19758 25314
rect 19782 25262 19828 25314
rect 19828 25262 19838 25314
rect 19862 25262 19892 25314
rect 19892 25262 19918 25314
rect 19622 25260 19678 25262
rect 19702 25260 19758 25262
rect 19782 25260 19838 25262
rect 19862 25260 19918 25262
rect 19622 24226 19678 24228
rect 19702 24226 19758 24228
rect 19782 24226 19838 24228
rect 19862 24226 19918 24228
rect 19622 24174 19648 24226
rect 19648 24174 19678 24226
rect 19702 24174 19712 24226
rect 19712 24174 19758 24226
rect 19782 24174 19828 24226
rect 19828 24174 19838 24226
rect 19862 24174 19892 24226
rect 19892 24174 19918 24226
rect 19622 24172 19678 24174
rect 19702 24172 19758 24174
rect 19782 24172 19838 24174
rect 19862 24172 19918 24174
rect 18510 22900 18566 22936
rect 18510 22880 18512 22900
rect 18512 22880 18564 22900
rect 18564 22880 18566 22900
rect 18326 21812 18382 21848
rect 18326 21792 18328 21812
rect 18328 21792 18380 21812
rect 18380 21792 18382 21812
rect 18050 16352 18106 16408
rect 18326 15672 18382 15728
rect 19430 23868 19432 23888
rect 19432 23868 19484 23888
rect 19484 23868 19486 23888
rect 19430 23832 19486 23868
rect 19622 23138 19678 23140
rect 19702 23138 19758 23140
rect 19782 23138 19838 23140
rect 19862 23138 19918 23140
rect 19622 23086 19648 23138
rect 19648 23086 19678 23138
rect 19702 23086 19712 23138
rect 19712 23086 19758 23138
rect 19782 23086 19828 23138
rect 19828 23086 19838 23138
rect 19862 23086 19892 23138
rect 19892 23086 19918 23138
rect 19622 23084 19678 23086
rect 19702 23084 19758 23086
rect 19782 23084 19838 23086
rect 19862 23084 19918 23086
rect 19798 22880 19854 22936
rect 19622 22050 19678 22052
rect 19702 22050 19758 22052
rect 19782 22050 19838 22052
rect 19862 22050 19918 22052
rect 19622 21998 19648 22050
rect 19648 21998 19678 22050
rect 19702 21998 19712 22050
rect 19712 21998 19758 22050
rect 19782 21998 19828 22050
rect 19828 21998 19838 22050
rect 19862 21998 19892 22050
rect 19892 21998 19918 22050
rect 19622 21996 19678 21998
rect 19702 21996 19758 21998
rect 19782 21996 19838 21998
rect 19862 21996 19918 21998
rect 18694 21132 18750 21168
rect 18694 21112 18696 21132
rect 18696 21112 18748 21132
rect 18748 21112 18750 21132
rect 19246 21676 19302 21712
rect 19246 21656 19248 21676
rect 19248 21656 19300 21676
rect 19300 21656 19302 21676
rect 19622 20962 19678 20964
rect 19702 20962 19758 20964
rect 19782 20962 19838 20964
rect 19862 20962 19918 20964
rect 19622 20910 19648 20962
rect 19648 20910 19678 20962
rect 19702 20910 19712 20962
rect 19712 20910 19758 20962
rect 19782 20910 19828 20962
rect 19828 20910 19838 20962
rect 19862 20910 19892 20962
rect 19892 20910 19918 20962
rect 19622 20908 19678 20910
rect 19702 20908 19758 20910
rect 19782 20908 19838 20910
rect 19862 20908 19918 20910
rect 19430 20860 19486 20896
rect 19430 20840 19432 20860
rect 19432 20840 19484 20860
rect 19484 20840 19486 20860
rect 19622 19874 19678 19876
rect 19702 19874 19758 19876
rect 19782 19874 19838 19876
rect 19862 19874 19918 19876
rect 19622 19822 19648 19874
rect 19648 19822 19678 19874
rect 19702 19822 19712 19874
rect 19712 19822 19758 19874
rect 19782 19822 19828 19874
rect 19828 19822 19838 19874
rect 19862 19822 19892 19874
rect 19892 19822 19918 19874
rect 19622 19820 19678 19822
rect 19702 19820 19758 19822
rect 19782 19820 19838 19822
rect 19862 19820 19918 19822
rect 19798 19636 19854 19672
rect 19798 19616 19800 19636
rect 19800 19616 19852 19636
rect 19852 19616 19854 19636
rect 19338 18836 19340 18856
rect 19340 18836 19392 18856
rect 19392 18836 19394 18856
rect 19062 18528 19118 18584
rect 19338 18800 19394 18836
rect 19246 18392 19302 18448
rect 19622 18786 19678 18788
rect 19702 18786 19758 18788
rect 19782 18786 19838 18788
rect 19862 18786 19918 18788
rect 19622 18734 19648 18786
rect 19648 18734 19678 18786
rect 19702 18734 19712 18786
rect 19712 18734 19758 18786
rect 19782 18734 19828 18786
rect 19828 18734 19838 18786
rect 19862 18734 19892 18786
rect 19892 18734 19918 18786
rect 19622 18732 19678 18734
rect 19702 18732 19758 18734
rect 19782 18732 19838 18734
rect 19862 18732 19918 18734
rect 19622 17698 19678 17700
rect 19702 17698 19758 17700
rect 19782 17698 19838 17700
rect 19862 17698 19918 17700
rect 19622 17646 19648 17698
rect 19648 17646 19678 17698
rect 19702 17646 19712 17698
rect 19712 17646 19758 17698
rect 19782 17646 19828 17698
rect 19828 17646 19838 17698
rect 19862 17646 19892 17698
rect 19892 17646 19918 17698
rect 19622 17644 19678 17646
rect 19702 17644 19758 17646
rect 19782 17644 19838 17646
rect 19862 17644 19918 17646
rect 19622 16610 19678 16612
rect 19702 16610 19758 16612
rect 19782 16610 19838 16612
rect 19862 16610 19918 16612
rect 19622 16558 19648 16610
rect 19648 16558 19678 16610
rect 19702 16558 19712 16610
rect 19712 16558 19758 16610
rect 19782 16558 19828 16610
rect 19828 16558 19838 16610
rect 19862 16558 19892 16610
rect 19892 16558 19918 16610
rect 19622 16556 19678 16558
rect 19702 16556 19758 16558
rect 19782 16556 19838 16558
rect 19862 16556 19918 16558
rect 19622 15522 19678 15524
rect 19702 15522 19758 15524
rect 19782 15522 19838 15524
rect 19862 15522 19918 15524
rect 19622 15470 19648 15522
rect 19648 15470 19678 15522
rect 19702 15470 19712 15522
rect 19712 15470 19758 15522
rect 19782 15470 19828 15522
rect 19828 15470 19838 15522
rect 19862 15470 19892 15522
rect 19892 15470 19918 15522
rect 19622 15468 19678 15470
rect 19702 15468 19758 15470
rect 19782 15468 19838 15470
rect 19862 15468 19918 15470
rect 19154 15164 19156 15184
rect 19156 15164 19208 15184
rect 19208 15164 19210 15184
rect 19154 15128 19210 15164
rect 19622 14434 19678 14436
rect 19702 14434 19758 14436
rect 19782 14434 19838 14436
rect 19862 14434 19918 14436
rect 19622 14382 19648 14434
rect 19648 14382 19678 14434
rect 19702 14382 19712 14434
rect 19712 14382 19758 14434
rect 19782 14382 19828 14434
rect 19828 14382 19838 14434
rect 19862 14382 19892 14434
rect 19892 14382 19918 14434
rect 19622 14380 19678 14382
rect 19702 14380 19758 14382
rect 19782 14380 19838 14382
rect 19862 14380 19918 14382
rect 19338 13632 19394 13688
rect 18786 13496 18842 13552
rect 19622 13346 19678 13348
rect 19702 13346 19758 13348
rect 19782 13346 19838 13348
rect 19862 13346 19918 13348
rect 19622 13294 19648 13346
rect 19648 13294 19678 13346
rect 19702 13294 19712 13346
rect 19712 13294 19758 13346
rect 19782 13294 19828 13346
rect 19828 13294 19838 13346
rect 19862 13294 19892 13346
rect 19892 13294 19918 13346
rect 19622 13292 19678 13294
rect 19702 13292 19758 13294
rect 19782 13292 19838 13294
rect 19862 13292 19918 13294
rect 19622 12258 19678 12260
rect 19702 12258 19758 12260
rect 19782 12258 19838 12260
rect 19862 12258 19918 12260
rect 19622 12206 19648 12258
rect 19648 12206 19678 12258
rect 19702 12206 19712 12258
rect 19712 12206 19758 12258
rect 19782 12206 19828 12258
rect 19828 12206 19838 12258
rect 19862 12206 19892 12258
rect 19892 12206 19918 12258
rect 19622 12204 19678 12206
rect 19702 12204 19758 12206
rect 19782 12204 19838 12206
rect 19862 12204 19918 12206
rect 18510 10776 18566 10832
rect 18878 10776 18934 10832
rect 19622 11170 19678 11172
rect 19702 11170 19758 11172
rect 19782 11170 19838 11172
rect 19862 11170 19918 11172
rect 19622 11118 19648 11170
rect 19648 11118 19678 11170
rect 19702 11118 19712 11170
rect 19712 11118 19758 11170
rect 19782 11118 19828 11170
rect 19828 11118 19838 11170
rect 19862 11118 19892 11170
rect 19892 11118 19918 11170
rect 19622 11116 19678 11118
rect 19702 11116 19758 11118
rect 19782 11116 19838 11118
rect 19862 11116 19918 11118
rect 19622 10082 19678 10084
rect 19702 10082 19758 10084
rect 19782 10082 19838 10084
rect 19862 10082 19918 10084
rect 19622 10030 19648 10082
rect 19648 10030 19678 10082
rect 19702 10030 19712 10082
rect 19712 10030 19758 10082
rect 19782 10030 19828 10082
rect 19828 10030 19838 10082
rect 19862 10030 19892 10082
rect 19892 10030 19918 10082
rect 19622 10028 19678 10030
rect 19702 10028 19758 10030
rect 19782 10028 19838 10030
rect 19862 10028 19918 10030
rect 19154 9436 19210 9472
rect 19154 9416 19156 9436
rect 19156 9416 19208 9436
rect 19208 9416 19210 9436
rect 20166 14720 20222 14776
rect 20258 10776 20314 10832
rect 20074 9280 20130 9336
rect 21178 23968 21234 24024
rect 20994 23288 21050 23344
rect 20718 21656 20774 21712
rect 20902 17748 20904 17768
rect 20904 17748 20956 17768
rect 20956 17748 20958 17768
rect 20902 17712 20958 17748
rect 20718 15128 20774 15184
rect 21270 19072 21326 19128
rect 21362 18392 21418 18448
rect 21270 11340 21326 11376
rect 21270 11320 21272 11340
rect 21272 11320 21324 11340
rect 21324 11320 21326 11340
rect 22558 24412 22560 24432
rect 22560 24412 22612 24432
rect 22612 24412 22614 24432
rect 22558 24376 22614 24412
rect 23570 26824 23626 26880
rect 23386 26144 23442 26200
rect 22834 24548 22836 24568
rect 22836 24548 22888 24568
rect 22888 24548 22890 24568
rect 22834 24512 22890 24548
rect 22742 23288 22798 23344
rect 24289 24770 24345 24772
rect 24369 24770 24425 24772
rect 24449 24770 24505 24772
rect 24529 24770 24585 24772
rect 24289 24718 24315 24770
rect 24315 24718 24345 24770
rect 24369 24718 24379 24770
rect 24379 24718 24425 24770
rect 24449 24718 24495 24770
rect 24495 24718 24505 24770
rect 24529 24718 24559 24770
rect 24559 24718 24585 24770
rect 24289 24716 24345 24718
rect 24369 24716 24425 24718
rect 24449 24716 24505 24718
rect 24529 24716 24585 24718
rect 23662 23152 23718 23208
rect 23570 22744 23626 22800
rect 23294 21792 23350 21848
rect 22006 20976 22062 21032
rect 21638 16760 21694 16816
rect 21454 10504 21510 10560
rect 20442 9008 20498 9064
rect 19622 8994 19678 8996
rect 19702 8994 19758 8996
rect 19782 8994 19838 8996
rect 19862 8994 19918 8996
rect 19622 8942 19648 8994
rect 19648 8942 19678 8994
rect 19702 8942 19712 8994
rect 19712 8942 19758 8994
rect 19782 8942 19828 8994
rect 19828 8942 19838 8994
rect 19862 8942 19892 8994
rect 19892 8942 19918 8994
rect 19622 8940 19678 8942
rect 19702 8940 19758 8942
rect 19782 8940 19838 8942
rect 19862 8940 19918 8942
rect 19622 7906 19678 7908
rect 19702 7906 19758 7908
rect 19782 7906 19838 7908
rect 19862 7906 19918 7908
rect 19622 7854 19648 7906
rect 19648 7854 19678 7906
rect 19702 7854 19712 7906
rect 19712 7854 19758 7906
rect 19782 7854 19828 7906
rect 19828 7854 19838 7906
rect 19862 7854 19892 7906
rect 19892 7854 19918 7906
rect 19622 7852 19678 7854
rect 19702 7852 19758 7854
rect 19782 7852 19838 7854
rect 19862 7852 19918 7854
rect 18878 7648 18934 7704
rect 18418 7512 18474 7568
rect 18234 7124 18290 7160
rect 18234 7104 18236 7124
rect 18236 7104 18288 7124
rect 18288 7104 18290 7124
rect 19622 6818 19678 6820
rect 19702 6818 19758 6820
rect 19782 6818 19838 6820
rect 19862 6818 19918 6820
rect 19622 6766 19648 6818
rect 19648 6766 19678 6818
rect 19702 6766 19712 6818
rect 19712 6766 19758 6818
rect 19782 6766 19828 6818
rect 19828 6766 19838 6818
rect 19862 6766 19892 6818
rect 19892 6766 19918 6818
rect 19622 6764 19678 6766
rect 19702 6764 19758 6766
rect 19782 6764 19838 6766
rect 19862 6764 19918 6766
rect 16946 5900 17002 5936
rect 16946 5880 16948 5900
rect 16948 5880 17000 5900
rect 17000 5880 17002 5900
rect 19622 5730 19678 5732
rect 19702 5730 19758 5732
rect 19782 5730 19838 5732
rect 19862 5730 19918 5732
rect 19622 5678 19648 5730
rect 19648 5678 19678 5730
rect 19702 5678 19712 5730
rect 19712 5678 19758 5730
rect 19782 5678 19828 5730
rect 19828 5678 19838 5730
rect 19862 5678 19892 5730
rect 19892 5678 19918 5730
rect 19622 5676 19678 5678
rect 19702 5676 19758 5678
rect 19782 5676 19838 5678
rect 19862 5676 19918 5678
rect 16026 5336 16082 5392
rect 15934 4948 15990 4984
rect 15934 4928 15936 4948
rect 15936 4928 15988 4948
rect 15988 4928 15990 4948
rect 10289 4642 10345 4644
rect 10369 4642 10425 4644
rect 10449 4642 10505 4644
rect 10529 4642 10585 4644
rect 10289 4590 10315 4642
rect 10315 4590 10345 4642
rect 10369 4590 10379 4642
rect 10379 4590 10425 4642
rect 10449 4590 10495 4642
rect 10495 4590 10505 4642
rect 10529 4590 10559 4642
rect 10559 4590 10585 4642
rect 10289 4588 10345 4590
rect 10369 4588 10425 4590
rect 10449 4588 10505 4590
rect 10529 4588 10585 4590
rect 19622 4642 19678 4644
rect 19702 4642 19758 4644
rect 19782 4642 19838 4644
rect 19862 4642 19918 4644
rect 19622 4590 19648 4642
rect 19648 4590 19678 4642
rect 19702 4590 19712 4642
rect 19712 4590 19758 4642
rect 19782 4590 19828 4642
rect 19828 4590 19838 4642
rect 19862 4590 19892 4642
rect 19892 4590 19918 4642
rect 19622 4588 19678 4590
rect 19702 4588 19758 4590
rect 19782 4588 19838 4590
rect 19862 4588 19918 4590
rect 5622 4098 5678 4100
rect 5702 4098 5758 4100
rect 5782 4098 5838 4100
rect 5862 4098 5918 4100
rect 5622 4046 5648 4098
rect 5648 4046 5678 4098
rect 5702 4046 5712 4098
rect 5712 4046 5758 4098
rect 5782 4046 5828 4098
rect 5828 4046 5838 4098
rect 5862 4046 5892 4098
rect 5892 4046 5918 4098
rect 5622 4044 5678 4046
rect 5702 4044 5758 4046
rect 5782 4044 5838 4046
rect 5862 4044 5918 4046
rect 14956 4098 15012 4100
rect 15036 4098 15092 4100
rect 15116 4098 15172 4100
rect 15196 4098 15252 4100
rect 14956 4046 14982 4098
rect 14982 4046 15012 4098
rect 15036 4046 15046 4098
rect 15046 4046 15092 4098
rect 15116 4046 15162 4098
rect 15162 4046 15172 4098
rect 15196 4046 15226 4098
rect 15226 4046 15252 4098
rect 14956 4044 15012 4046
rect 15036 4044 15092 4046
rect 15116 4044 15172 4046
rect 15196 4044 15252 4046
rect 22466 20724 22522 20760
rect 22466 20704 22468 20724
rect 22468 20704 22520 20724
rect 22520 20704 22522 20724
rect 21914 18528 21970 18584
rect 22282 18956 22338 18992
rect 22282 18936 22284 18956
rect 22284 18936 22336 18956
rect 22336 18936 22338 18956
rect 21822 14584 21878 14640
rect 23846 22200 23902 22256
rect 23846 21012 23848 21032
rect 23848 21012 23900 21032
rect 23900 21012 23902 21032
rect 23846 20976 23902 21012
rect 23846 17712 23902 17768
rect 23754 17168 23810 17224
rect 23846 16372 23902 16408
rect 23846 16352 23848 16372
rect 23848 16352 23900 16372
rect 23900 16352 23902 16372
rect 22926 14756 22928 14776
rect 22928 14756 22980 14776
rect 22980 14756 22982 14776
rect 22926 14720 22982 14756
rect 23478 14604 23534 14640
rect 23478 14584 23480 14604
rect 23480 14584 23532 14604
rect 23532 14584 23534 14604
rect 21730 9960 21786 10016
rect 21638 3704 21694 3760
rect 10289 3554 10345 3556
rect 10369 3554 10425 3556
rect 10449 3554 10505 3556
rect 10529 3554 10585 3556
rect 10289 3502 10315 3554
rect 10315 3502 10345 3554
rect 10369 3502 10379 3554
rect 10379 3502 10425 3554
rect 10449 3502 10495 3554
rect 10495 3502 10505 3554
rect 10529 3502 10559 3554
rect 10559 3502 10585 3554
rect 10289 3500 10345 3502
rect 10369 3500 10425 3502
rect 10449 3500 10505 3502
rect 10529 3500 10585 3502
rect 19622 3554 19678 3556
rect 19702 3554 19758 3556
rect 19782 3554 19838 3556
rect 19862 3554 19918 3556
rect 19622 3502 19648 3554
rect 19648 3502 19678 3554
rect 19702 3502 19712 3554
rect 19712 3502 19758 3554
rect 19782 3502 19828 3554
rect 19828 3502 19838 3554
rect 19862 3502 19892 3554
rect 19892 3502 19918 3554
rect 19622 3500 19678 3502
rect 19702 3500 19758 3502
rect 19782 3500 19838 3502
rect 19862 3500 19918 3502
rect 5622 3010 5678 3012
rect 5702 3010 5758 3012
rect 5782 3010 5838 3012
rect 5862 3010 5918 3012
rect 5622 2958 5648 3010
rect 5648 2958 5678 3010
rect 5702 2958 5712 3010
rect 5712 2958 5758 3010
rect 5782 2958 5828 3010
rect 5828 2958 5838 3010
rect 5862 2958 5892 3010
rect 5892 2958 5918 3010
rect 5622 2956 5678 2958
rect 5702 2956 5758 2958
rect 5782 2956 5838 2958
rect 5862 2956 5918 2958
rect 14956 3010 15012 3012
rect 15036 3010 15092 3012
rect 15116 3010 15172 3012
rect 15196 3010 15252 3012
rect 14956 2958 14982 3010
rect 14982 2958 15012 3010
rect 15036 2958 15046 3010
rect 15046 2958 15092 3010
rect 15116 2958 15162 3010
rect 15162 2958 15172 3010
rect 15196 2958 15226 3010
rect 15226 2958 15252 3010
rect 14956 2956 15012 2958
rect 15036 2956 15092 2958
rect 15116 2956 15172 2958
rect 15196 2956 15252 2958
rect 10289 2466 10345 2468
rect 10369 2466 10425 2468
rect 10449 2466 10505 2468
rect 10529 2466 10585 2468
rect 10289 2414 10315 2466
rect 10315 2414 10345 2466
rect 10369 2414 10379 2466
rect 10379 2414 10425 2466
rect 10449 2414 10495 2466
rect 10495 2414 10505 2466
rect 10529 2414 10559 2466
rect 10559 2414 10585 2466
rect 10289 2412 10345 2414
rect 10369 2412 10425 2414
rect 10449 2412 10505 2414
rect 10529 2412 10585 2414
rect 19622 2466 19678 2468
rect 19702 2466 19758 2468
rect 19782 2466 19838 2468
rect 19862 2466 19918 2468
rect 19622 2414 19648 2466
rect 19648 2414 19678 2466
rect 19702 2414 19712 2466
rect 19712 2414 19758 2466
rect 19782 2414 19828 2466
rect 19828 2414 19838 2466
rect 19862 2414 19892 2466
rect 19892 2414 19918 2466
rect 19622 2412 19678 2414
rect 19702 2412 19758 2414
rect 19782 2412 19838 2414
rect 19862 2412 19918 2414
rect 23570 13768 23626 13824
rect 23478 10524 23534 10560
rect 23478 10504 23480 10524
rect 23480 10504 23532 10524
rect 23532 10504 23534 10524
rect 23478 3704 23534 3760
rect 22282 2344 22338 2400
rect 5622 1922 5678 1924
rect 5702 1922 5758 1924
rect 5782 1922 5838 1924
rect 5862 1922 5918 1924
rect 5622 1870 5648 1922
rect 5648 1870 5678 1922
rect 5702 1870 5712 1922
rect 5712 1870 5758 1922
rect 5782 1870 5828 1922
rect 5828 1870 5838 1922
rect 5862 1870 5892 1922
rect 5892 1870 5918 1922
rect 5622 1868 5678 1870
rect 5702 1868 5758 1870
rect 5782 1868 5838 1870
rect 5862 1868 5918 1870
rect 14956 1922 15012 1924
rect 15036 1922 15092 1924
rect 15116 1922 15172 1924
rect 15196 1922 15252 1924
rect 14956 1870 14982 1922
rect 14982 1870 15012 1922
rect 15036 1870 15046 1922
rect 15046 1870 15092 1922
rect 15116 1870 15162 1922
rect 15162 1870 15172 1922
rect 15196 1870 15226 1922
rect 15226 1870 15252 1922
rect 14956 1868 15012 1870
rect 15036 1868 15092 1870
rect 15116 1868 15172 1870
rect 15196 1868 15252 1870
rect 23570 3160 23626 3216
rect 23570 2344 23626 2400
rect 23478 1120 23534 1176
rect 23754 13496 23810 13552
rect 24289 23682 24345 23684
rect 24369 23682 24425 23684
rect 24449 23682 24505 23684
rect 24529 23682 24585 23684
rect 24289 23630 24315 23682
rect 24315 23630 24345 23682
rect 24369 23630 24379 23682
rect 24379 23630 24425 23682
rect 24449 23630 24495 23682
rect 24495 23630 24505 23682
rect 24529 23630 24559 23682
rect 24559 23630 24585 23682
rect 24289 23628 24345 23630
rect 24369 23628 24425 23630
rect 24449 23628 24505 23630
rect 24529 23628 24585 23630
rect 24122 22608 24178 22664
rect 24289 22594 24345 22596
rect 24369 22594 24425 22596
rect 24449 22594 24505 22596
rect 24529 22594 24585 22596
rect 24289 22542 24315 22594
rect 24315 22542 24345 22594
rect 24369 22542 24379 22594
rect 24379 22542 24425 22594
rect 24449 22542 24495 22594
rect 24495 22542 24505 22594
rect 24529 22542 24559 22594
rect 24559 22542 24585 22594
rect 24289 22540 24345 22542
rect 24369 22540 24425 22542
rect 24449 22540 24505 22542
rect 24529 22540 24585 22542
rect 24582 22336 24638 22392
rect 24766 25600 24822 25656
rect 25134 25056 25190 25112
rect 24766 23696 24822 23752
rect 25134 24376 25190 24432
rect 25686 24512 25742 24568
rect 25502 23832 25558 23888
rect 25410 23696 25466 23752
rect 24858 22880 24914 22936
rect 25134 22644 25136 22664
rect 25136 22644 25188 22664
rect 25188 22644 25190 22664
rect 25134 22608 25190 22644
rect 24766 22100 24768 22120
rect 24768 22100 24820 22120
rect 24820 22100 24822 22120
rect 24766 22064 24822 22100
rect 24122 21520 24178 21576
rect 24030 20160 24086 20216
rect 24122 15672 24178 15728
rect 24122 14312 24178 14368
rect 24289 21506 24345 21508
rect 24369 21506 24425 21508
rect 24449 21506 24505 21508
rect 24529 21506 24585 21508
rect 24289 21454 24315 21506
rect 24315 21454 24345 21506
rect 24369 21454 24379 21506
rect 24379 21454 24425 21506
rect 24449 21454 24495 21506
rect 24495 21454 24505 21506
rect 24529 21454 24559 21506
rect 24559 21454 24585 21506
rect 24289 21452 24345 21454
rect 24369 21452 24425 21454
rect 24449 21452 24505 21454
rect 24529 21452 24585 21454
rect 24289 20418 24345 20420
rect 24369 20418 24425 20420
rect 24449 20418 24505 20420
rect 24529 20418 24585 20420
rect 24289 20366 24315 20418
rect 24315 20366 24345 20418
rect 24369 20366 24379 20418
rect 24379 20366 24425 20418
rect 24449 20366 24495 20418
rect 24495 20366 24505 20418
rect 24529 20366 24559 20418
rect 24559 20366 24585 20418
rect 24289 20364 24345 20366
rect 24369 20364 24425 20366
rect 24449 20364 24505 20366
rect 24529 20364 24585 20366
rect 24289 19330 24345 19332
rect 24369 19330 24425 19332
rect 24449 19330 24505 19332
rect 24529 19330 24585 19332
rect 24289 19278 24315 19330
rect 24315 19278 24345 19330
rect 24369 19278 24379 19330
rect 24379 19278 24425 19330
rect 24449 19278 24495 19330
rect 24495 19278 24505 19330
rect 24529 19278 24559 19330
rect 24559 19278 24585 19330
rect 24289 19276 24345 19278
rect 24369 19276 24425 19278
rect 24449 19276 24505 19278
rect 24529 19276 24585 19278
rect 24289 18242 24345 18244
rect 24369 18242 24425 18244
rect 24449 18242 24505 18244
rect 24529 18242 24585 18244
rect 24289 18190 24315 18242
rect 24315 18190 24345 18242
rect 24369 18190 24379 18242
rect 24379 18190 24425 18242
rect 24449 18190 24495 18242
rect 24495 18190 24505 18242
rect 24529 18190 24559 18242
rect 24559 18190 24585 18242
rect 24289 18188 24345 18190
rect 24369 18188 24425 18190
rect 24449 18188 24505 18190
rect 24529 18188 24585 18190
rect 24289 17154 24345 17156
rect 24369 17154 24425 17156
rect 24449 17154 24505 17156
rect 24529 17154 24585 17156
rect 24289 17102 24315 17154
rect 24315 17102 24345 17154
rect 24369 17102 24379 17154
rect 24379 17102 24425 17154
rect 24449 17102 24495 17154
rect 24495 17102 24505 17154
rect 24529 17102 24559 17154
rect 24559 17102 24585 17154
rect 24289 17100 24345 17102
rect 24369 17100 24425 17102
rect 24449 17100 24505 17102
rect 24529 17100 24585 17102
rect 24289 16066 24345 16068
rect 24369 16066 24425 16068
rect 24449 16066 24505 16068
rect 24529 16066 24585 16068
rect 24289 16014 24315 16066
rect 24315 16014 24345 16066
rect 24369 16014 24379 16066
rect 24379 16014 24425 16066
rect 24449 16014 24495 16066
rect 24495 16014 24505 16066
rect 24529 16014 24559 16066
rect 24559 16014 24585 16066
rect 24289 16012 24345 16014
rect 24369 16012 24425 16014
rect 24449 16012 24505 16014
rect 24529 16012 24585 16014
rect 24289 14978 24345 14980
rect 24369 14978 24425 14980
rect 24449 14978 24505 14980
rect 24529 14978 24585 14980
rect 24289 14926 24315 14978
rect 24315 14926 24345 14978
rect 24369 14926 24379 14978
rect 24379 14926 24425 14978
rect 24449 14926 24495 14978
rect 24495 14926 24505 14978
rect 24529 14926 24559 14978
rect 24559 14926 24585 14978
rect 24289 14924 24345 14926
rect 24369 14924 24425 14926
rect 24449 14924 24505 14926
rect 24529 14924 24585 14926
rect 24289 13890 24345 13892
rect 24369 13890 24425 13892
rect 24449 13890 24505 13892
rect 24529 13890 24585 13892
rect 24289 13838 24315 13890
rect 24315 13838 24345 13890
rect 24369 13838 24379 13890
rect 24379 13838 24425 13890
rect 24449 13838 24495 13890
rect 24495 13838 24505 13890
rect 24529 13838 24559 13890
rect 24559 13838 24585 13890
rect 24289 13836 24345 13838
rect 24369 13836 24425 13838
rect 24449 13836 24505 13838
rect 24529 13836 24585 13838
rect 24766 21384 24822 21440
rect 25502 21248 25558 21304
rect 24858 20160 24914 20216
rect 25134 20840 25190 20896
rect 25318 20296 25374 20352
rect 24950 20024 25006 20080
rect 24858 19636 24914 19672
rect 24858 19616 24860 19636
rect 24860 19616 24912 19636
rect 24912 19616 24914 19636
rect 24766 19072 24822 19128
rect 25042 19616 25098 19672
rect 25410 18412 25466 18448
rect 25410 18392 25412 18412
rect 25412 18392 25464 18412
rect 25464 18392 25466 18412
rect 25594 17848 25650 17904
rect 25502 17304 25558 17360
rect 25410 16624 25466 16680
rect 24766 16216 24822 16272
rect 25318 16080 25374 16136
rect 25502 15400 25558 15456
rect 25594 14856 25650 14912
rect 25226 13652 25282 13688
rect 25226 13632 25228 13652
rect 25228 13632 25280 13652
rect 25280 13632 25282 13652
rect 24582 13108 24638 13144
rect 24582 13088 24584 13108
rect 24584 13088 24636 13108
rect 24636 13088 24638 13108
rect 24289 12802 24345 12804
rect 24369 12802 24425 12804
rect 24449 12802 24505 12804
rect 24529 12802 24585 12804
rect 24289 12750 24315 12802
rect 24315 12750 24345 12802
rect 24369 12750 24379 12802
rect 24379 12750 24425 12802
rect 24449 12750 24495 12802
rect 24495 12750 24505 12802
rect 24529 12750 24559 12802
rect 24559 12750 24585 12802
rect 24289 12748 24345 12750
rect 24369 12748 24425 12750
rect 24449 12748 24505 12750
rect 24529 12748 24585 12750
rect 24398 12564 24454 12600
rect 24398 12544 24400 12564
rect 24400 12544 24452 12564
rect 24452 12544 24454 12564
rect 24398 11864 24454 11920
rect 24674 11864 24730 11920
rect 24289 11714 24345 11716
rect 24369 11714 24425 11716
rect 24449 11714 24505 11716
rect 24529 11714 24585 11716
rect 24289 11662 24315 11714
rect 24315 11662 24345 11714
rect 24369 11662 24379 11714
rect 24379 11662 24425 11714
rect 24449 11662 24495 11714
rect 24495 11662 24505 11714
rect 24529 11662 24559 11714
rect 24559 11662 24585 11714
rect 24289 11660 24345 11662
rect 24369 11660 24425 11662
rect 24449 11660 24505 11662
rect 24529 11660 24585 11662
rect 26882 24512 26938 24568
rect 24674 10640 24730 10696
rect 24289 10626 24345 10628
rect 24369 10626 24425 10628
rect 24449 10626 24505 10628
rect 24529 10626 24585 10628
rect 24289 10574 24315 10626
rect 24315 10574 24345 10626
rect 24369 10574 24379 10626
rect 24379 10574 24425 10626
rect 24449 10574 24495 10626
rect 24495 10574 24505 10626
rect 24529 10574 24559 10626
rect 24559 10574 24585 10626
rect 24289 10572 24345 10574
rect 24369 10572 24425 10574
rect 24449 10572 24505 10574
rect 24529 10572 24585 10574
rect 24122 10232 24178 10288
rect 23846 2344 23902 2400
rect 25226 10132 25228 10152
rect 25228 10132 25280 10152
rect 25280 10132 25282 10152
rect 25226 10096 25282 10132
rect 24766 9980 24822 10016
rect 24766 9960 24768 9980
rect 24768 9960 24820 9980
rect 24820 9960 24822 9980
rect 24674 9552 24730 9608
rect 25226 9552 25282 9608
rect 24289 9538 24345 9540
rect 24369 9538 24425 9540
rect 24449 9538 24505 9540
rect 24529 9538 24585 9540
rect 24289 9486 24315 9538
rect 24315 9486 24345 9538
rect 24369 9486 24379 9538
rect 24379 9486 24425 9538
rect 24449 9486 24495 9538
rect 24495 9486 24505 9538
rect 24529 9486 24559 9538
rect 24559 9486 24585 9538
rect 24289 9484 24345 9486
rect 24369 9484 24425 9486
rect 24449 9484 24505 9486
rect 24529 9484 24585 9486
rect 24766 9316 24768 9336
rect 24768 9316 24820 9336
rect 24820 9316 24822 9336
rect 24766 9280 24822 9316
rect 24766 9008 24822 9064
rect 24490 8872 24546 8928
rect 24289 8450 24345 8452
rect 24369 8450 24425 8452
rect 24449 8450 24505 8452
rect 24529 8450 24585 8452
rect 24289 8398 24315 8450
rect 24315 8398 24345 8450
rect 24369 8398 24379 8450
rect 24379 8398 24425 8450
rect 24449 8398 24495 8450
rect 24495 8398 24505 8450
rect 24529 8398 24559 8450
rect 24559 8398 24585 8450
rect 24289 8396 24345 8398
rect 24369 8396 24425 8398
rect 24449 8396 24505 8398
rect 24529 8396 24585 8398
rect 24674 8348 24730 8384
rect 24674 8328 24676 8348
rect 24676 8328 24728 8348
rect 24728 8328 24730 8348
rect 24214 7648 24270 7704
rect 24582 7668 24638 7704
rect 24582 7648 24584 7668
rect 24584 7648 24636 7668
rect 24636 7648 24638 7668
rect 24289 7362 24345 7364
rect 24369 7362 24425 7364
rect 24449 7362 24505 7364
rect 24529 7362 24585 7364
rect 24289 7310 24315 7362
rect 24315 7310 24345 7362
rect 24369 7310 24379 7362
rect 24379 7310 24425 7362
rect 24449 7310 24495 7362
rect 24495 7310 24505 7362
rect 24529 7310 24559 7362
rect 24559 7310 24585 7362
rect 24289 7308 24345 7310
rect 24369 7308 24425 7310
rect 24449 7308 24505 7310
rect 24529 7308 24585 7310
rect 24766 7532 24822 7568
rect 24766 7512 24768 7532
rect 24768 7512 24820 7532
rect 24820 7512 24822 7532
rect 24214 6560 24270 6616
rect 24289 6274 24345 6276
rect 24369 6274 24425 6276
rect 24449 6274 24505 6276
rect 24529 6274 24585 6276
rect 24289 6222 24315 6274
rect 24315 6222 24345 6274
rect 24369 6222 24379 6274
rect 24379 6222 24425 6274
rect 24449 6222 24495 6274
rect 24495 6222 24505 6274
rect 24529 6222 24559 6274
rect 24559 6222 24585 6274
rect 24289 6220 24345 6222
rect 24369 6220 24425 6222
rect 24449 6220 24505 6222
rect 24529 6220 24585 6222
rect 24289 5186 24345 5188
rect 24369 5186 24425 5188
rect 24449 5186 24505 5188
rect 24529 5186 24585 5188
rect 24289 5134 24315 5186
rect 24315 5134 24345 5186
rect 24369 5134 24379 5186
rect 24379 5134 24425 5186
rect 24449 5134 24495 5186
rect 24495 5134 24505 5186
rect 24529 5134 24559 5186
rect 24559 5134 24585 5186
rect 24289 5132 24345 5134
rect 24369 5132 24425 5134
rect 24449 5132 24505 5134
rect 24529 5132 24585 5134
rect 24122 4248 24178 4304
rect 24289 4098 24345 4100
rect 24369 4098 24425 4100
rect 24449 4098 24505 4100
rect 24529 4098 24585 4100
rect 24289 4046 24315 4098
rect 24315 4046 24345 4098
rect 24369 4046 24379 4098
rect 24379 4046 24425 4098
rect 24449 4046 24495 4098
rect 24495 4046 24505 4098
rect 24529 4046 24559 4098
rect 24559 4046 24585 4098
rect 24289 4044 24345 4046
rect 24369 4044 24425 4046
rect 24449 4044 24505 4046
rect 24529 4044 24585 4046
rect 24766 3704 24822 3760
rect 26238 3704 26294 3760
rect 25226 3604 25228 3624
rect 25228 3604 25280 3624
rect 25280 3604 25282 3624
rect 25226 3568 25282 3604
rect 24289 3010 24345 3012
rect 24369 3010 24425 3012
rect 24449 3010 24505 3012
rect 24529 3010 24585 3012
rect 24289 2958 24315 3010
rect 24315 2958 24345 3010
rect 24369 2958 24379 3010
rect 24379 2958 24425 3010
rect 24449 2958 24495 3010
rect 24495 2958 24505 3010
rect 24529 2958 24559 3010
rect 24559 2958 24585 3010
rect 24289 2956 24345 2958
rect 24369 2956 24425 2958
rect 24449 2956 24505 2958
rect 24529 2956 24585 2958
rect 23938 2072 23994 2128
rect 24289 1922 24345 1924
rect 24369 1922 24425 1924
rect 24449 1922 24505 1924
rect 24529 1922 24585 1924
rect 24289 1870 24315 1922
rect 24315 1870 24345 1922
rect 24369 1870 24379 1922
rect 24379 1870 24425 1922
rect 24449 1870 24495 1922
rect 24495 1870 24505 1922
rect 24529 1870 24559 1922
rect 24559 1870 24585 1922
rect 24289 1868 24345 1870
rect 24369 1868 24425 1870
rect 24449 1868 24505 1870
rect 24529 1868 24585 1870
rect 23662 576 23718 632
rect 23570 32 23626 88
<< metal3 >>
rect 23933 27426 23999 27429
rect 27520 27426 28000 27456
rect 23933 27424 28000 27426
rect 23933 27368 23938 27424
rect 23994 27368 28000 27424
rect 23933 27366 28000 27368
rect 23933 27363 23999 27366
rect 27520 27336 28000 27366
rect 23565 26882 23631 26885
rect 27520 26882 28000 26912
rect 23565 26880 28000 26882
rect 23565 26824 23570 26880
rect 23626 26824 28000 26880
rect 23565 26822 28000 26824
rect 23565 26819 23631 26822
rect 27520 26792 28000 26822
rect 23381 26202 23447 26205
rect 27520 26202 28000 26232
rect 23381 26200 28000 26202
rect 23381 26144 23386 26200
rect 23442 26144 28000 26200
rect 23381 26142 28000 26144
rect 23381 26139 23447 26142
rect 27520 26112 28000 26142
rect 24761 25658 24827 25661
rect 27520 25658 28000 25688
rect 24761 25656 28000 25658
rect 24761 25600 24766 25656
rect 24822 25600 28000 25656
rect 24761 25598 28000 25600
rect 24761 25595 24827 25598
rect 27520 25568 28000 25598
rect 10277 25320 10597 25321
rect 10277 25256 10285 25320
rect 10349 25256 10365 25320
rect 10429 25256 10445 25320
rect 10509 25256 10525 25320
rect 10589 25256 10597 25320
rect 10277 25255 10597 25256
rect 19610 25320 19930 25321
rect 19610 25256 19618 25320
rect 19682 25256 19698 25320
rect 19762 25256 19778 25320
rect 19842 25256 19858 25320
rect 19922 25256 19930 25320
rect 19610 25255 19930 25256
rect 25129 25114 25195 25117
rect 27520 25114 28000 25144
rect 25129 25112 28000 25114
rect 25129 25056 25134 25112
rect 25190 25056 28000 25112
rect 25129 25054 28000 25056
rect 25129 25051 25195 25054
rect 27520 25024 28000 25054
rect 5610 24776 5930 24777
rect 5610 24712 5618 24776
rect 5682 24712 5698 24776
rect 5762 24712 5778 24776
rect 5842 24712 5858 24776
rect 5922 24712 5930 24776
rect 5610 24711 5930 24712
rect 14944 24776 15264 24777
rect 14944 24712 14952 24776
rect 15016 24712 15032 24776
rect 15096 24712 15112 24776
rect 15176 24712 15192 24776
rect 15256 24712 15264 24776
rect 14944 24711 15264 24712
rect 24277 24776 24597 24777
rect 24277 24712 24285 24776
rect 24349 24712 24365 24776
rect 24429 24712 24445 24776
rect 24509 24712 24525 24776
rect 24589 24712 24597 24776
rect 24277 24711 24597 24712
rect 13629 24570 13695 24573
rect 14549 24570 14615 24573
rect 22829 24570 22895 24573
rect 13629 24568 14615 24570
rect 13629 24512 13634 24568
rect 13690 24512 14554 24568
rect 14610 24512 14615 24568
rect 13629 24510 14615 24512
rect 13629 24507 13695 24510
rect 14549 24507 14615 24510
rect 17542 24568 22895 24570
rect 17542 24512 22834 24568
rect 22890 24512 22895 24568
rect 17542 24510 22895 24512
rect 13169 24434 13235 24437
rect 17542 24434 17602 24510
rect 22829 24507 22895 24510
rect 25681 24570 25747 24573
rect 26877 24570 26943 24573
rect 25681 24568 26943 24570
rect 25681 24512 25686 24568
rect 25742 24512 26882 24568
rect 26938 24512 26943 24568
rect 25681 24510 26943 24512
rect 25681 24507 25747 24510
rect 26877 24507 26943 24510
rect 22553 24434 22619 24437
rect 13169 24432 17602 24434
rect 13169 24376 13174 24432
rect 13230 24376 17602 24432
rect 13169 24374 17602 24376
rect 17726 24432 22619 24434
rect 17726 24376 22558 24432
rect 22614 24376 22619 24432
rect 17726 24374 22619 24376
rect 13169 24371 13235 24374
rect 12525 24298 12591 24301
rect 17726 24298 17786 24374
rect 22553 24371 22619 24374
rect 25129 24434 25195 24437
rect 27520 24434 28000 24464
rect 25129 24432 28000 24434
rect 25129 24376 25134 24432
rect 25190 24376 28000 24432
rect 25129 24374 28000 24376
rect 25129 24371 25195 24374
rect 27520 24344 28000 24374
rect 12525 24296 17786 24298
rect 12525 24240 12530 24296
rect 12586 24240 17786 24296
rect 12525 24238 17786 24240
rect 12525 24235 12591 24238
rect 10277 24232 10597 24233
rect 10277 24168 10285 24232
rect 10349 24168 10365 24232
rect 10429 24168 10445 24232
rect 10509 24168 10525 24232
rect 10589 24168 10597 24232
rect 10277 24167 10597 24168
rect 19610 24232 19930 24233
rect 19610 24168 19618 24232
rect 19682 24168 19698 24232
rect 19762 24168 19778 24232
rect 19842 24168 19858 24232
rect 19922 24168 19930 24232
rect 19610 24167 19930 24168
rect 4981 24026 5047 24029
rect 21173 24026 21239 24029
rect 4981 24024 21239 24026
rect 4981 23968 4986 24024
rect 5042 23968 21178 24024
rect 21234 23968 21239 24024
rect 4981 23966 21239 23968
rect 4981 23963 5047 23966
rect 21173 23963 21239 23966
rect 14825 23890 14891 23893
rect 19425 23890 19491 23893
rect 14825 23888 19491 23890
rect 14825 23832 14830 23888
rect 14886 23832 19430 23888
rect 19486 23832 19491 23888
rect 14825 23830 19491 23832
rect 14825 23827 14891 23830
rect 19425 23827 19491 23830
rect 25497 23890 25563 23893
rect 27520 23890 28000 23920
rect 25497 23888 28000 23890
rect 25497 23832 25502 23888
rect 25558 23832 28000 23888
rect 25497 23830 28000 23832
rect 25497 23827 25563 23830
rect 27520 23800 28000 23830
rect 24761 23754 24827 23757
rect 25405 23754 25471 23757
rect 24761 23752 25471 23754
rect 24761 23696 24766 23752
rect 24822 23696 25410 23752
rect 25466 23696 25471 23752
rect 24761 23694 25471 23696
rect 24761 23691 24827 23694
rect 25405 23691 25471 23694
rect 5610 23688 5930 23689
rect 5610 23624 5618 23688
rect 5682 23624 5698 23688
rect 5762 23624 5778 23688
rect 5842 23624 5858 23688
rect 5922 23624 5930 23688
rect 5610 23623 5930 23624
rect 14944 23688 15264 23689
rect 14944 23624 14952 23688
rect 15016 23624 15032 23688
rect 15096 23624 15112 23688
rect 15176 23624 15192 23688
rect 15256 23624 15264 23688
rect 14944 23623 15264 23624
rect 24277 23688 24597 23689
rect 24277 23624 24285 23688
rect 24349 23624 24365 23688
rect 24429 23624 24445 23688
rect 24509 23624 24525 23688
rect 24589 23624 24597 23688
rect 24277 23623 24597 23624
rect 11145 23618 11211 23621
rect 13353 23618 13419 23621
rect 11145 23616 13419 23618
rect 11145 23560 11150 23616
rect 11206 23560 13358 23616
rect 13414 23560 13419 23616
rect 11145 23558 13419 23560
rect 11145 23555 11211 23558
rect 13353 23555 13419 23558
rect 20989 23346 21055 23349
rect 22737 23346 22803 23349
rect 20989 23344 22803 23346
rect 20989 23288 20994 23344
rect 21050 23288 22742 23344
rect 22798 23288 22803 23344
rect 20989 23286 22803 23288
rect 20989 23283 21055 23286
rect 22737 23283 22803 23286
rect 10869 23210 10935 23213
rect 14089 23210 14155 23213
rect 14733 23210 14799 23213
rect 10869 23208 14799 23210
rect 10869 23152 10874 23208
rect 10930 23152 14094 23208
rect 14150 23152 14738 23208
rect 14794 23152 14799 23208
rect 10869 23150 14799 23152
rect 10869 23147 10935 23150
rect 14089 23147 14155 23150
rect 14733 23147 14799 23150
rect 23657 23210 23723 23213
rect 27520 23210 28000 23240
rect 23657 23208 28000 23210
rect 23657 23152 23662 23208
rect 23718 23152 28000 23208
rect 23657 23150 28000 23152
rect 23657 23147 23723 23150
rect 10277 23144 10597 23145
rect 10277 23080 10285 23144
rect 10349 23080 10365 23144
rect 10429 23080 10445 23144
rect 10509 23080 10525 23144
rect 10589 23080 10597 23144
rect 10277 23079 10597 23080
rect 19610 23144 19930 23145
rect 19610 23080 19618 23144
rect 19682 23080 19698 23144
rect 19762 23080 19778 23144
rect 19842 23080 19858 23144
rect 19922 23080 19930 23144
rect 27520 23120 28000 23150
rect 19610 23079 19930 23080
rect 10133 22938 10199 22941
rect 18505 22938 18571 22941
rect 10133 22936 18571 22938
rect 10133 22880 10138 22936
rect 10194 22880 18510 22936
rect 18566 22880 18571 22936
rect 10133 22878 18571 22880
rect 10133 22875 10199 22878
rect 18505 22875 18571 22878
rect 19793 22938 19859 22941
rect 24853 22938 24919 22941
rect 19793 22936 24919 22938
rect 19793 22880 19798 22936
rect 19854 22880 24858 22936
rect 24914 22880 24919 22936
rect 19793 22878 24919 22880
rect 19793 22875 19859 22878
rect 24853 22875 24919 22878
rect 9213 22802 9279 22805
rect 23565 22802 23631 22805
rect 9213 22800 23631 22802
rect 9213 22744 9218 22800
rect 9274 22744 23570 22800
rect 23626 22744 23631 22800
rect 9213 22742 23631 22744
rect 9213 22739 9279 22742
rect 23565 22739 23631 22742
rect 16113 22666 16179 22669
rect 24117 22666 24183 22669
rect 16113 22664 24183 22666
rect 16113 22608 16118 22664
rect 16174 22608 24122 22664
rect 24178 22608 24183 22664
rect 16113 22606 24183 22608
rect 16113 22603 16179 22606
rect 24117 22603 24183 22606
rect 25129 22666 25195 22669
rect 27520 22666 28000 22696
rect 25129 22664 28000 22666
rect 25129 22608 25134 22664
rect 25190 22608 28000 22664
rect 25129 22606 28000 22608
rect 25129 22603 25195 22606
rect 5610 22600 5930 22601
rect 5610 22536 5618 22600
rect 5682 22536 5698 22600
rect 5762 22536 5778 22600
rect 5842 22536 5858 22600
rect 5922 22536 5930 22600
rect 5610 22535 5930 22536
rect 14944 22600 15264 22601
rect 14944 22536 14952 22600
rect 15016 22536 15032 22600
rect 15096 22536 15112 22600
rect 15176 22536 15192 22600
rect 15256 22536 15264 22600
rect 14944 22535 15264 22536
rect 24277 22600 24597 22601
rect 24277 22536 24285 22600
rect 24349 22536 24365 22600
rect 24429 22536 24445 22600
rect 24509 22536 24525 22600
rect 24589 22536 24597 22600
rect 27520 22576 28000 22606
rect 24277 22535 24597 22536
rect 9765 22530 9831 22533
rect 14733 22530 14799 22533
rect 9765 22528 14799 22530
rect 9765 22472 9770 22528
rect 9826 22472 14738 22528
rect 14794 22472 14799 22528
rect 9765 22470 14799 22472
rect 9765 22467 9831 22470
rect 14733 22467 14799 22470
rect 7741 22394 7807 22397
rect 24577 22394 24643 22397
rect 7741 22392 24643 22394
rect 7741 22336 7746 22392
rect 7802 22336 24582 22392
rect 24638 22336 24643 22392
rect 7741 22334 24643 22336
rect 7741 22331 7807 22334
rect 24577 22331 24643 22334
rect 13537 22258 13603 22261
rect 23841 22258 23907 22261
rect 13537 22256 23907 22258
rect 13537 22200 13542 22256
rect 13598 22200 23846 22256
rect 23902 22200 23907 22256
rect 13537 22198 23907 22200
rect 13537 22195 13603 22198
rect 23841 22195 23907 22198
rect 24761 22122 24827 22125
rect 27520 22122 28000 22152
rect 24761 22120 28000 22122
rect 24761 22064 24766 22120
rect 24822 22064 28000 22120
rect 24761 22062 28000 22064
rect 24761 22059 24827 22062
rect 10277 22056 10597 22057
rect 10277 21992 10285 22056
rect 10349 21992 10365 22056
rect 10429 21992 10445 22056
rect 10509 21992 10525 22056
rect 10589 21992 10597 22056
rect 10277 21991 10597 21992
rect 19610 22056 19930 22057
rect 19610 21992 19618 22056
rect 19682 21992 19698 22056
rect 19762 21992 19778 22056
rect 19842 21992 19858 22056
rect 19922 21992 19930 22056
rect 27520 22032 28000 22062
rect 19610 21991 19930 21992
rect 18321 21850 18387 21853
rect 23289 21850 23355 21853
rect 14782 21790 15394 21850
rect 7097 21578 7163 21581
rect 14782 21578 14842 21790
rect 7097 21576 14842 21578
rect 7097 21520 7102 21576
rect 7158 21520 14842 21576
rect 7097 21518 14842 21520
rect 15334 21578 15394 21790
rect 18321 21848 23355 21850
rect 18321 21792 18326 21848
rect 18382 21792 23294 21848
rect 23350 21792 23355 21848
rect 18321 21790 23355 21792
rect 18321 21787 18387 21790
rect 23289 21787 23355 21790
rect 19241 21714 19307 21717
rect 20713 21714 20779 21717
rect 19241 21712 20779 21714
rect 19241 21656 19246 21712
rect 19302 21656 20718 21712
rect 20774 21656 20779 21712
rect 19241 21654 20779 21656
rect 19241 21651 19307 21654
rect 20713 21651 20779 21654
rect 24117 21578 24183 21581
rect 15334 21576 24183 21578
rect 15334 21520 24122 21576
rect 24178 21520 24183 21576
rect 15334 21518 24183 21520
rect 7097 21515 7163 21518
rect 24117 21515 24183 21518
rect 5610 21512 5930 21513
rect 5610 21448 5618 21512
rect 5682 21448 5698 21512
rect 5762 21448 5778 21512
rect 5842 21448 5858 21512
rect 5922 21448 5930 21512
rect 5610 21447 5930 21448
rect 14944 21512 15264 21513
rect 14944 21448 14952 21512
rect 15016 21448 15032 21512
rect 15096 21448 15112 21512
rect 15176 21448 15192 21512
rect 15256 21448 15264 21512
rect 14944 21447 15264 21448
rect 24277 21512 24597 21513
rect 24277 21448 24285 21512
rect 24349 21448 24365 21512
rect 24429 21448 24445 21512
rect 24509 21448 24525 21512
rect 24589 21448 24597 21512
rect 24277 21447 24597 21448
rect 24761 21442 24827 21445
rect 27520 21442 28000 21472
rect 24761 21440 28000 21442
rect 24761 21384 24766 21440
rect 24822 21384 28000 21440
rect 24761 21382 28000 21384
rect 24761 21379 24827 21382
rect 27520 21352 28000 21382
rect 6361 21306 6427 21309
rect 11237 21306 11303 21309
rect 6361 21304 11303 21306
rect 6361 21248 6366 21304
rect 6422 21248 11242 21304
rect 11298 21248 11303 21304
rect 6361 21246 11303 21248
rect 6361 21243 6427 21246
rect 11237 21243 11303 21246
rect 14181 21306 14247 21309
rect 25497 21306 25563 21309
rect 14181 21304 25563 21306
rect 14181 21248 14186 21304
rect 14242 21248 25502 21304
rect 25558 21248 25563 21304
rect 14181 21246 25563 21248
rect 14181 21243 14247 21246
rect 25497 21243 25563 21246
rect 5993 21170 6059 21173
rect 18689 21170 18755 21173
rect 5993 21168 18755 21170
rect 5993 21112 5998 21168
rect 6054 21112 18694 21168
rect 18750 21112 18755 21168
rect 5993 21110 18755 21112
rect 5993 21107 6059 21110
rect 18689 21107 18755 21110
rect 22001 21034 22067 21037
rect 23841 21034 23907 21037
rect 22001 21032 23907 21034
rect 22001 20976 22006 21032
rect 22062 20976 23846 21032
rect 23902 20976 23907 21032
rect 22001 20974 23907 20976
rect 22001 20971 22067 20974
rect 23841 20971 23907 20974
rect 10277 20968 10597 20969
rect 10277 20904 10285 20968
rect 10349 20904 10365 20968
rect 10429 20904 10445 20968
rect 10509 20904 10525 20968
rect 10589 20904 10597 20968
rect 10277 20903 10597 20904
rect 19610 20968 19930 20969
rect 19610 20904 19618 20968
rect 19682 20904 19698 20968
rect 19762 20904 19778 20968
rect 19842 20904 19858 20968
rect 19922 20904 19930 20968
rect 19610 20903 19930 20904
rect 4337 20898 4403 20901
rect 10685 20898 10751 20901
rect 19425 20898 19491 20901
rect 4337 20896 10058 20898
rect 4337 20840 4342 20896
rect 4398 20840 10058 20896
rect 4337 20838 10058 20840
rect 4337 20835 4403 20838
rect 0 20762 480 20792
rect 9213 20762 9279 20765
rect 0 20760 9279 20762
rect 0 20704 9218 20760
rect 9274 20704 9279 20760
rect 0 20702 9279 20704
rect 9998 20762 10058 20838
rect 10685 20896 19491 20898
rect 10685 20840 10690 20896
rect 10746 20840 19430 20896
rect 19486 20840 19491 20896
rect 10685 20838 19491 20840
rect 10685 20835 10751 20838
rect 19425 20835 19491 20838
rect 25129 20898 25195 20901
rect 27520 20898 28000 20928
rect 25129 20896 28000 20898
rect 25129 20840 25134 20896
rect 25190 20840 28000 20896
rect 25129 20838 28000 20840
rect 25129 20835 25195 20838
rect 27520 20808 28000 20838
rect 22461 20762 22527 20765
rect 9998 20760 22527 20762
rect 9998 20704 22466 20760
rect 22522 20704 22527 20760
rect 9998 20702 22527 20704
rect 0 20672 480 20702
rect 9213 20699 9279 20702
rect 22461 20699 22527 20702
rect 9121 20626 9187 20629
rect 16113 20626 16179 20629
rect 9121 20624 16179 20626
rect 9121 20568 9126 20624
rect 9182 20568 16118 20624
rect 16174 20568 16179 20624
rect 9121 20566 16179 20568
rect 9121 20563 9187 20566
rect 16113 20563 16179 20566
rect 8385 20490 8451 20493
rect 13353 20490 13419 20493
rect 8385 20488 13419 20490
rect 8385 20432 8390 20488
rect 8446 20432 13358 20488
rect 13414 20432 13419 20488
rect 8385 20430 13419 20432
rect 8385 20427 8451 20430
rect 13353 20427 13419 20430
rect 5610 20424 5930 20425
rect 5610 20360 5618 20424
rect 5682 20360 5698 20424
rect 5762 20360 5778 20424
rect 5842 20360 5858 20424
rect 5922 20360 5930 20424
rect 5610 20359 5930 20360
rect 14944 20424 15264 20425
rect 14944 20360 14952 20424
rect 15016 20360 15032 20424
rect 15096 20360 15112 20424
rect 15176 20360 15192 20424
rect 15256 20360 15264 20424
rect 14944 20359 15264 20360
rect 24277 20424 24597 20425
rect 24277 20360 24285 20424
rect 24349 20360 24365 20424
rect 24429 20360 24445 20424
rect 24509 20360 24525 20424
rect 24589 20360 24597 20424
rect 24277 20359 24597 20360
rect 25313 20354 25379 20357
rect 27520 20354 28000 20384
rect 25313 20352 28000 20354
rect 25313 20296 25318 20352
rect 25374 20296 28000 20352
rect 25313 20294 28000 20296
rect 25313 20291 25379 20294
rect 27520 20264 28000 20294
rect 24025 20218 24091 20221
rect 24853 20218 24919 20221
rect 24025 20216 24919 20218
rect 24025 20160 24030 20216
rect 24086 20160 24858 20216
rect 24914 20160 24919 20216
rect 24025 20158 24919 20160
rect 24025 20155 24091 20158
rect 24853 20155 24919 20158
rect 13997 20082 14063 20085
rect 24945 20082 25011 20085
rect 13997 20080 25011 20082
rect 13997 20024 14002 20080
rect 14058 20024 24950 20080
rect 25006 20024 25011 20080
rect 13997 20022 25011 20024
rect 13997 20019 14063 20022
rect 24945 20019 25011 20022
rect 10685 19946 10751 19949
rect 11145 19946 11211 19949
rect 17585 19946 17651 19949
rect 10685 19944 17651 19946
rect 10685 19888 10690 19944
rect 10746 19888 11150 19944
rect 11206 19888 17590 19944
rect 17646 19888 17651 19944
rect 10685 19886 17651 19888
rect 10685 19883 10751 19886
rect 11145 19883 11211 19886
rect 17585 19883 17651 19886
rect 10277 19880 10597 19881
rect 10277 19816 10285 19880
rect 10349 19816 10365 19880
rect 10429 19816 10445 19880
rect 10509 19816 10525 19880
rect 10589 19816 10597 19880
rect 10277 19815 10597 19816
rect 19610 19880 19930 19881
rect 19610 19816 19618 19880
rect 19682 19816 19698 19880
rect 19762 19816 19778 19880
rect 19842 19816 19858 19880
rect 19922 19816 19930 19880
rect 19610 19815 19930 19816
rect 19793 19674 19859 19677
rect 24853 19674 24919 19677
rect 19793 19672 24919 19674
rect 19793 19616 19798 19672
rect 19854 19616 24858 19672
rect 24914 19616 24919 19672
rect 19793 19614 24919 19616
rect 19793 19611 19859 19614
rect 24853 19611 24919 19614
rect 25037 19674 25103 19677
rect 27520 19674 28000 19704
rect 25037 19672 28000 19674
rect 25037 19616 25042 19672
rect 25098 19616 28000 19672
rect 25037 19614 28000 19616
rect 25037 19611 25103 19614
rect 27520 19584 28000 19614
rect 5610 19336 5930 19337
rect 5610 19272 5618 19336
rect 5682 19272 5698 19336
rect 5762 19272 5778 19336
rect 5842 19272 5858 19336
rect 5922 19272 5930 19336
rect 5610 19271 5930 19272
rect 14944 19336 15264 19337
rect 14944 19272 14952 19336
rect 15016 19272 15032 19336
rect 15096 19272 15112 19336
rect 15176 19272 15192 19336
rect 15256 19272 15264 19336
rect 14944 19271 15264 19272
rect 24277 19336 24597 19337
rect 24277 19272 24285 19336
rect 24349 19272 24365 19336
rect 24429 19272 24445 19336
rect 24509 19272 24525 19336
rect 24589 19272 24597 19336
rect 24277 19271 24597 19272
rect 13905 19130 13971 19133
rect 21265 19130 21331 19133
rect 13905 19128 21331 19130
rect 13905 19072 13910 19128
rect 13966 19072 21270 19128
rect 21326 19072 21331 19128
rect 13905 19070 21331 19072
rect 13905 19067 13971 19070
rect 21265 19067 21331 19070
rect 24761 19130 24827 19133
rect 27520 19130 28000 19160
rect 24761 19128 28000 19130
rect 24761 19072 24766 19128
rect 24822 19072 28000 19128
rect 24761 19070 28000 19072
rect 24761 19067 24827 19070
rect 27520 19040 28000 19070
rect 3693 18994 3759 18997
rect 22277 18994 22343 18997
rect 3693 18992 22343 18994
rect 3693 18936 3698 18992
rect 3754 18936 22282 18992
rect 22338 18936 22343 18992
rect 3693 18934 22343 18936
rect 3693 18931 3759 18934
rect 22277 18931 22343 18934
rect 13537 18858 13603 18861
rect 19333 18858 19399 18861
rect 13537 18856 19399 18858
rect 13537 18800 13542 18856
rect 13598 18800 19338 18856
rect 19394 18800 19399 18856
rect 13537 18798 19399 18800
rect 13537 18795 13603 18798
rect 19333 18795 19399 18798
rect 10277 18792 10597 18793
rect 10277 18728 10285 18792
rect 10349 18728 10365 18792
rect 10429 18728 10445 18792
rect 10509 18728 10525 18792
rect 10589 18728 10597 18792
rect 10277 18727 10597 18728
rect 19610 18792 19930 18793
rect 19610 18728 19618 18792
rect 19682 18728 19698 18792
rect 19762 18728 19778 18792
rect 19842 18728 19858 18792
rect 19922 18728 19930 18792
rect 19610 18727 19930 18728
rect 17033 18722 17099 18725
rect 17033 18720 19258 18722
rect 17033 18664 17038 18720
rect 17094 18664 19258 18720
rect 17033 18662 19258 18664
rect 17033 18659 17099 18662
rect 2957 18586 3023 18589
rect 19057 18586 19123 18589
rect 2957 18584 19123 18586
rect 2957 18528 2962 18584
rect 3018 18528 19062 18584
rect 19118 18528 19123 18584
rect 2957 18526 19123 18528
rect 19198 18586 19258 18662
rect 21909 18586 21975 18589
rect 19198 18584 21975 18586
rect 19198 18528 21914 18584
rect 21970 18528 21975 18584
rect 19198 18526 21975 18528
rect 2957 18523 3023 18526
rect 19057 18523 19123 18526
rect 21909 18523 21975 18526
rect 19241 18450 19307 18453
rect 21357 18450 21423 18453
rect 19241 18448 21423 18450
rect 19241 18392 19246 18448
rect 19302 18392 21362 18448
rect 21418 18392 21423 18448
rect 19241 18390 21423 18392
rect 19241 18387 19307 18390
rect 21357 18387 21423 18390
rect 25405 18450 25471 18453
rect 27520 18450 28000 18480
rect 25405 18448 28000 18450
rect 25405 18392 25410 18448
rect 25466 18392 28000 18448
rect 25405 18390 28000 18392
rect 25405 18387 25471 18390
rect 27520 18360 28000 18390
rect 5610 18248 5930 18249
rect 5610 18184 5618 18248
rect 5682 18184 5698 18248
rect 5762 18184 5778 18248
rect 5842 18184 5858 18248
rect 5922 18184 5930 18248
rect 5610 18183 5930 18184
rect 14944 18248 15264 18249
rect 14944 18184 14952 18248
rect 15016 18184 15032 18248
rect 15096 18184 15112 18248
rect 15176 18184 15192 18248
rect 15256 18184 15264 18248
rect 14944 18183 15264 18184
rect 24277 18248 24597 18249
rect 24277 18184 24285 18248
rect 24349 18184 24365 18248
rect 24429 18184 24445 18248
rect 24509 18184 24525 18248
rect 24589 18184 24597 18248
rect 24277 18183 24597 18184
rect 25589 17906 25655 17909
rect 27520 17906 28000 17936
rect 25589 17904 28000 17906
rect 25589 17848 25594 17904
rect 25650 17848 28000 17904
rect 25589 17846 28000 17848
rect 25589 17843 25655 17846
rect 27520 17816 28000 17846
rect 20897 17770 20963 17773
rect 23841 17770 23907 17773
rect 20897 17768 23907 17770
rect 20897 17712 20902 17768
rect 20958 17712 23846 17768
rect 23902 17712 23907 17768
rect 20897 17710 23907 17712
rect 20897 17707 20963 17710
rect 23841 17707 23907 17710
rect 10277 17704 10597 17705
rect 10277 17640 10285 17704
rect 10349 17640 10365 17704
rect 10429 17640 10445 17704
rect 10509 17640 10525 17704
rect 10589 17640 10597 17704
rect 10277 17639 10597 17640
rect 19610 17704 19930 17705
rect 19610 17640 19618 17704
rect 19682 17640 19698 17704
rect 19762 17640 19778 17704
rect 19842 17640 19858 17704
rect 19922 17640 19930 17704
rect 19610 17639 19930 17640
rect 14089 17362 14155 17365
rect 25497 17362 25563 17365
rect 27520 17362 28000 17392
rect 14089 17360 18154 17362
rect 14089 17304 14094 17360
rect 14150 17304 18154 17360
rect 14089 17302 18154 17304
rect 14089 17299 14155 17302
rect 18094 17226 18154 17302
rect 25497 17360 28000 17362
rect 25497 17304 25502 17360
rect 25558 17304 28000 17360
rect 25497 17302 28000 17304
rect 25497 17299 25563 17302
rect 27520 17272 28000 17302
rect 23749 17226 23815 17229
rect 18094 17224 23815 17226
rect 18094 17168 23754 17224
rect 23810 17168 23815 17224
rect 18094 17166 23815 17168
rect 23749 17163 23815 17166
rect 5610 17160 5930 17161
rect 5610 17096 5618 17160
rect 5682 17096 5698 17160
rect 5762 17096 5778 17160
rect 5842 17096 5858 17160
rect 5922 17096 5930 17160
rect 5610 17095 5930 17096
rect 14944 17160 15264 17161
rect 14944 17096 14952 17160
rect 15016 17096 15032 17160
rect 15096 17096 15112 17160
rect 15176 17096 15192 17160
rect 15256 17096 15264 17160
rect 14944 17095 15264 17096
rect 24277 17160 24597 17161
rect 24277 17096 24285 17160
rect 24349 17096 24365 17160
rect 24429 17096 24445 17160
rect 24509 17096 24525 17160
rect 24589 17096 24597 17160
rect 24277 17095 24597 17096
rect 1577 16818 1643 16821
rect 11881 16818 11947 16821
rect 1577 16816 11947 16818
rect 1577 16760 1582 16816
rect 1638 16760 11886 16816
rect 11942 16760 11947 16816
rect 1577 16758 11947 16760
rect 1577 16755 1643 16758
rect 11881 16755 11947 16758
rect 13997 16818 14063 16821
rect 15929 16818 15995 16821
rect 21633 16818 21699 16821
rect 13997 16816 21699 16818
rect 13997 16760 14002 16816
rect 14058 16760 15934 16816
rect 15990 16760 21638 16816
rect 21694 16760 21699 16816
rect 13997 16758 21699 16760
rect 13997 16755 14063 16758
rect 15929 16755 15995 16758
rect 21633 16755 21699 16758
rect 25405 16682 25471 16685
rect 27520 16682 28000 16712
rect 25405 16680 28000 16682
rect 25405 16624 25410 16680
rect 25466 16624 28000 16680
rect 25405 16622 28000 16624
rect 25405 16619 25471 16622
rect 10277 16616 10597 16617
rect 10277 16552 10285 16616
rect 10349 16552 10365 16616
rect 10429 16552 10445 16616
rect 10509 16552 10525 16616
rect 10589 16552 10597 16616
rect 10277 16551 10597 16552
rect 19610 16616 19930 16617
rect 19610 16552 19618 16616
rect 19682 16552 19698 16616
rect 19762 16552 19778 16616
rect 19842 16552 19858 16616
rect 19922 16552 19930 16616
rect 27520 16592 28000 16622
rect 19610 16551 19930 16552
rect 2313 16410 2379 16413
rect 15837 16410 15903 16413
rect 2313 16408 15903 16410
rect 2313 16352 2318 16408
rect 2374 16352 15842 16408
rect 15898 16352 15903 16408
rect 2313 16350 15903 16352
rect 2313 16347 2379 16350
rect 15837 16347 15903 16350
rect 18045 16410 18111 16413
rect 23841 16410 23907 16413
rect 18045 16408 23907 16410
rect 18045 16352 18050 16408
rect 18106 16352 23846 16408
rect 23902 16352 23907 16408
rect 18045 16350 23907 16352
rect 18045 16347 18111 16350
rect 23841 16347 23907 16350
rect 1301 16274 1367 16277
rect 16389 16274 16455 16277
rect 24761 16274 24827 16277
rect 1301 16272 11714 16274
rect 1301 16216 1306 16272
rect 1362 16216 11714 16272
rect 1301 16214 11714 16216
rect 1301 16211 1367 16214
rect 5610 16072 5930 16073
rect 5610 16008 5618 16072
rect 5682 16008 5698 16072
rect 5762 16008 5778 16072
rect 5842 16008 5858 16072
rect 5922 16008 5930 16072
rect 5610 16007 5930 16008
rect 11654 15866 11714 16214
rect 16389 16272 24827 16274
rect 16389 16216 16394 16272
rect 16450 16216 24766 16272
rect 24822 16216 24827 16272
rect 16389 16214 24827 16216
rect 16389 16211 16455 16214
rect 24761 16211 24827 16214
rect 25313 16138 25379 16141
rect 27520 16138 28000 16168
rect 25313 16136 28000 16138
rect 25313 16080 25318 16136
rect 25374 16080 28000 16136
rect 25313 16078 28000 16080
rect 25313 16075 25379 16078
rect 14944 16072 15264 16073
rect 14944 16008 14952 16072
rect 15016 16008 15032 16072
rect 15096 16008 15112 16072
rect 15176 16008 15192 16072
rect 15256 16008 15264 16072
rect 14944 16007 15264 16008
rect 24277 16072 24597 16073
rect 24277 16008 24285 16072
rect 24349 16008 24365 16072
rect 24429 16008 24445 16072
rect 24509 16008 24525 16072
rect 24589 16008 24597 16072
rect 27520 16048 28000 16078
rect 24277 16007 24597 16008
rect 17125 15866 17191 15869
rect 11654 15864 17191 15866
rect 11654 15808 17130 15864
rect 17186 15808 17191 15864
rect 11654 15806 17191 15808
rect 17125 15803 17191 15806
rect 16297 15730 16363 15733
rect 18321 15730 18387 15733
rect 24117 15730 24183 15733
rect 16297 15728 24183 15730
rect 16297 15672 16302 15728
rect 16358 15672 18326 15728
rect 18382 15672 24122 15728
rect 24178 15672 24183 15728
rect 16297 15670 24183 15672
rect 16297 15667 16363 15670
rect 18321 15667 18387 15670
rect 24117 15667 24183 15670
rect 10277 15528 10597 15529
rect 10277 15464 10285 15528
rect 10349 15464 10365 15528
rect 10429 15464 10445 15528
rect 10509 15464 10525 15528
rect 10589 15464 10597 15528
rect 10277 15463 10597 15464
rect 19610 15528 19930 15529
rect 19610 15464 19618 15528
rect 19682 15464 19698 15528
rect 19762 15464 19778 15528
rect 19842 15464 19858 15528
rect 19922 15464 19930 15528
rect 19610 15463 19930 15464
rect 25497 15458 25563 15461
rect 27520 15458 28000 15488
rect 25497 15456 28000 15458
rect 25497 15400 25502 15456
rect 25558 15400 28000 15456
rect 25497 15398 28000 15400
rect 25497 15395 25563 15398
rect 27520 15368 28000 15398
rect 12709 15186 12775 15189
rect 16941 15186 17007 15189
rect 12709 15184 17007 15186
rect 12709 15128 12714 15184
rect 12770 15128 16946 15184
rect 17002 15128 17007 15184
rect 12709 15126 17007 15128
rect 12709 15123 12775 15126
rect 16941 15123 17007 15126
rect 19149 15186 19215 15189
rect 20713 15186 20779 15189
rect 19149 15184 20779 15186
rect 19149 15128 19154 15184
rect 19210 15128 20718 15184
rect 20774 15128 20779 15184
rect 19149 15126 20779 15128
rect 19149 15123 19215 15126
rect 20713 15123 20779 15126
rect 5610 14984 5930 14985
rect 5610 14920 5618 14984
rect 5682 14920 5698 14984
rect 5762 14920 5778 14984
rect 5842 14920 5858 14984
rect 5922 14920 5930 14984
rect 5610 14919 5930 14920
rect 14944 14984 15264 14985
rect 14944 14920 14952 14984
rect 15016 14920 15032 14984
rect 15096 14920 15112 14984
rect 15176 14920 15192 14984
rect 15256 14920 15264 14984
rect 14944 14919 15264 14920
rect 24277 14984 24597 14985
rect 24277 14920 24285 14984
rect 24349 14920 24365 14984
rect 24429 14920 24445 14984
rect 24509 14920 24525 14984
rect 24589 14920 24597 14984
rect 24277 14919 24597 14920
rect 25589 14914 25655 14917
rect 27520 14914 28000 14944
rect 25589 14912 28000 14914
rect 25589 14856 25594 14912
rect 25650 14856 28000 14912
rect 25589 14854 28000 14856
rect 25589 14851 25655 14854
rect 27520 14824 28000 14854
rect 20161 14778 20227 14781
rect 22921 14778 22987 14781
rect 20161 14776 22987 14778
rect 20161 14720 20166 14776
rect 20222 14720 22926 14776
rect 22982 14720 22987 14776
rect 20161 14718 22987 14720
rect 20161 14715 20227 14718
rect 22921 14715 22987 14718
rect 21817 14642 21883 14645
rect 23473 14642 23539 14645
rect 21817 14640 23539 14642
rect 21817 14584 21822 14640
rect 21878 14584 23478 14640
rect 23534 14584 23539 14640
rect 21817 14582 23539 14584
rect 21817 14579 21883 14582
rect 23473 14579 23539 14582
rect 10277 14440 10597 14441
rect 10277 14376 10285 14440
rect 10349 14376 10365 14440
rect 10429 14376 10445 14440
rect 10509 14376 10525 14440
rect 10589 14376 10597 14440
rect 10277 14375 10597 14376
rect 19610 14440 19930 14441
rect 19610 14376 19618 14440
rect 19682 14376 19698 14440
rect 19762 14376 19778 14440
rect 19842 14376 19858 14440
rect 19922 14376 19930 14440
rect 19610 14375 19930 14376
rect 24117 14370 24183 14373
rect 27520 14370 28000 14400
rect 24117 14368 28000 14370
rect 24117 14312 24122 14368
rect 24178 14312 28000 14368
rect 24117 14310 28000 14312
rect 24117 14307 24183 14310
rect 27520 14280 28000 14310
rect 5610 13896 5930 13897
rect 5610 13832 5618 13896
rect 5682 13832 5698 13896
rect 5762 13832 5778 13896
rect 5842 13832 5858 13896
rect 5922 13832 5930 13896
rect 5610 13831 5930 13832
rect 14944 13896 15264 13897
rect 14944 13832 14952 13896
rect 15016 13832 15032 13896
rect 15096 13832 15112 13896
rect 15176 13832 15192 13896
rect 15256 13832 15264 13896
rect 14944 13831 15264 13832
rect 24277 13896 24597 13897
rect 24277 13832 24285 13896
rect 24349 13832 24365 13896
rect 24429 13832 24445 13896
rect 24509 13832 24525 13896
rect 24589 13832 24597 13896
rect 24277 13831 24597 13832
rect 16941 13826 17007 13829
rect 23565 13826 23631 13829
rect 16941 13824 23631 13826
rect 16941 13768 16946 13824
rect 17002 13768 23570 13824
rect 23626 13768 23631 13824
rect 16941 13766 23631 13768
rect 16941 13763 17007 13766
rect 23565 13763 23631 13766
rect 17769 13690 17835 13693
rect 19333 13690 19399 13693
rect 17769 13688 19399 13690
rect 17769 13632 17774 13688
rect 17830 13632 19338 13688
rect 19394 13632 19399 13688
rect 17769 13630 19399 13632
rect 17769 13627 17835 13630
rect 19333 13627 19399 13630
rect 25221 13690 25287 13693
rect 27520 13690 28000 13720
rect 25221 13688 28000 13690
rect 25221 13632 25226 13688
rect 25282 13632 28000 13688
rect 25221 13630 28000 13632
rect 25221 13627 25287 13630
rect 27520 13600 28000 13630
rect 17493 13554 17559 13557
rect 18781 13554 18847 13557
rect 23749 13554 23815 13557
rect 17493 13552 23815 13554
rect 17493 13496 17498 13552
rect 17554 13496 18786 13552
rect 18842 13496 23754 13552
rect 23810 13496 23815 13552
rect 17493 13494 23815 13496
rect 17493 13491 17559 13494
rect 18781 13491 18847 13494
rect 23749 13491 23815 13494
rect 10277 13352 10597 13353
rect 10277 13288 10285 13352
rect 10349 13288 10365 13352
rect 10429 13288 10445 13352
rect 10509 13288 10525 13352
rect 10589 13288 10597 13352
rect 10277 13287 10597 13288
rect 19610 13352 19930 13353
rect 19610 13288 19618 13352
rect 19682 13288 19698 13352
rect 19762 13288 19778 13352
rect 19842 13288 19858 13352
rect 19922 13288 19930 13352
rect 19610 13287 19930 13288
rect 24577 13146 24643 13149
rect 27520 13146 28000 13176
rect 24577 13144 28000 13146
rect 24577 13088 24582 13144
rect 24638 13088 28000 13144
rect 24577 13086 28000 13088
rect 24577 13083 24643 13086
rect 27520 13056 28000 13086
rect 5610 12808 5930 12809
rect 5610 12744 5618 12808
rect 5682 12744 5698 12808
rect 5762 12744 5778 12808
rect 5842 12744 5858 12808
rect 5922 12744 5930 12808
rect 5610 12743 5930 12744
rect 14944 12808 15264 12809
rect 14944 12744 14952 12808
rect 15016 12744 15032 12808
rect 15096 12744 15112 12808
rect 15176 12744 15192 12808
rect 15256 12744 15264 12808
rect 14944 12743 15264 12744
rect 24277 12808 24597 12809
rect 24277 12744 24285 12808
rect 24349 12744 24365 12808
rect 24429 12744 24445 12808
rect 24509 12744 24525 12808
rect 24589 12744 24597 12808
rect 24277 12743 24597 12744
rect 24393 12602 24459 12605
rect 27520 12602 28000 12632
rect 24393 12600 28000 12602
rect 24393 12544 24398 12600
rect 24454 12544 28000 12600
rect 24393 12542 28000 12544
rect 24393 12539 24459 12542
rect 27520 12512 28000 12542
rect 10277 12264 10597 12265
rect 10277 12200 10285 12264
rect 10349 12200 10365 12264
rect 10429 12200 10445 12264
rect 10509 12200 10525 12264
rect 10589 12200 10597 12264
rect 10277 12199 10597 12200
rect 19610 12264 19930 12265
rect 19610 12200 19618 12264
rect 19682 12200 19698 12264
rect 19762 12200 19778 12264
rect 19842 12200 19858 12264
rect 19922 12200 19930 12264
rect 19610 12199 19930 12200
rect 24393 11922 24459 11925
rect 24669 11922 24735 11925
rect 27520 11922 28000 11952
rect 24393 11920 28000 11922
rect 24393 11864 24398 11920
rect 24454 11864 24674 11920
rect 24730 11864 28000 11920
rect 24393 11862 28000 11864
rect 24393 11859 24459 11862
rect 24669 11859 24735 11862
rect 27520 11832 28000 11862
rect 5610 11720 5930 11721
rect 5610 11656 5618 11720
rect 5682 11656 5698 11720
rect 5762 11656 5778 11720
rect 5842 11656 5858 11720
rect 5922 11656 5930 11720
rect 5610 11655 5930 11656
rect 14944 11720 15264 11721
rect 14944 11656 14952 11720
rect 15016 11656 15032 11720
rect 15096 11656 15112 11720
rect 15176 11656 15192 11720
rect 15256 11656 15264 11720
rect 14944 11655 15264 11656
rect 24277 11720 24597 11721
rect 24277 11656 24285 11720
rect 24349 11656 24365 11720
rect 24429 11656 24445 11720
rect 24509 11656 24525 11720
rect 24589 11656 24597 11720
rect 24277 11655 24597 11656
rect 21265 11378 21331 11381
rect 27520 11378 28000 11408
rect 21265 11376 28000 11378
rect 21265 11320 21270 11376
rect 21326 11320 28000 11376
rect 21265 11318 28000 11320
rect 21265 11315 21331 11318
rect 27520 11288 28000 11318
rect 10277 11176 10597 11177
rect 10277 11112 10285 11176
rect 10349 11112 10365 11176
rect 10429 11112 10445 11176
rect 10509 11112 10525 11176
rect 10589 11112 10597 11176
rect 10277 11111 10597 11112
rect 19610 11176 19930 11177
rect 19610 11112 19618 11176
rect 19682 11112 19698 11176
rect 19762 11112 19778 11176
rect 19842 11112 19858 11176
rect 19922 11112 19930 11176
rect 19610 11111 19930 11112
rect 18505 10834 18571 10837
rect 18873 10834 18939 10837
rect 20253 10834 20319 10837
rect 18505 10832 20319 10834
rect 18505 10776 18510 10832
rect 18566 10776 18878 10832
rect 18934 10776 20258 10832
rect 20314 10776 20319 10832
rect 18505 10774 20319 10776
rect 18505 10771 18571 10774
rect 18873 10771 18939 10774
rect 20253 10771 20319 10774
rect 24669 10698 24735 10701
rect 27520 10698 28000 10728
rect 24669 10696 28000 10698
rect 24669 10640 24674 10696
rect 24730 10640 28000 10696
rect 24669 10638 28000 10640
rect 24669 10635 24735 10638
rect 5610 10632 5930 10633
rect 5610 10568 5618 10632
rect 5682 10568 5698 10632
rect 5762 10568 5778 10632
rect 5842 10568 5858 10632
rect 5922 10568 5930 10632
rect 5610 10567 5930 10568
rect 14944 10632 15264 10633
rect 14944 10568 14952 10632
rect 15016 10568 15032 10632
rect 15096 10568 15112 10632
rect 15176 10568 15192 10632
rect 15256 10568 15264 10632
rect 14944 10567 15264 10568
rect 24277 10632 24597 10633
rect 24277 10568 24285 10632
rect 24349 10568 24365 10632
rect 24429 10568 24445 10632
rect 24509 10568 24525 10632
rect 24589 10568 24597 10632
rect 27520 10608 28000 10638
rect 24277 10567 24597 10568
rect 21449 10562 21515 10565
rect 23473 10562 23539 10565
rect 21449 10560 23539 10562
rect 21449 10504 21454 10560
rect 21510 10504 23478 10560
rect 23534 10504 23539 10560
rect 21449 10502 23539 10504
rect 21449 10499 21515 10502
rect 23473 10499 23539 10502
rect 3417 10290 3483 10293
rect 10777 10290 10843 10293
rect 3417 10288 10843 10290
rect 3417 10232 3422 10288
rect 3478 10232 10782 10288
rect 10838 10232 10843 10288
rect 3417 10230 10843 10232
rect 3417 10227 3483 10230
rect 10777 10227 10843 10230
rect 13813 10290 13879 10293
rect 24117 10290 24183 10293
rect 13813 10288 24183 10290
rect 13813 10232 13818 10288
rect 13874 10232 24122 10288
rect 24178 10232 24183 10288
rect 13813 10230 24183 10232
rect 13813 10227 13879 10230
rect 24117 10227 24183 10230
rect 25221 10154 25287 10157
rect 27520 10154 28000 10184
rect 25221 10152 28000 10154
rect 25221 10096 25226 10152
rect 25282 10096 28000 10152
rect 25221 10094 28000 10096
rect 25221 10091 25287 10094
rect 10277 10088 10597 10089
rect 10277 10024 10285 10088
rect 10349 10024 10365 10088
rect 10429 10024 10445 10088
rect 10509 10024 10525 10088
rect 10589 10024 10597 10088
rect 10277 10023 10597 10024
rect 19610 10088 19930 10089
rect 19610 10024 19618 10088
rect 19682 10024 19698 10088
rect 19762 10024 19778 10088
rect 19842 10024 19858 10088
rect 19922 10024 19930 10088
rect 27520 10064 28000 10094
rect 19610 10023 19930 10024
rect 21725 10018 21791 10021
rect 24761 10018 24827 10021
rect 21725 10016 24827 10018
rect 21725 9960 21730 10016
rect 21786 9960 24766 10016
rect 24822 9960 24827 10016
rect 21725 9958 24827 9960
rect 21725 9955 21791 9958
rect 24761 9955 24827 9958
rect 197 9746 263 9749
rect 13905 9746 13971 9749
rect 197 9744 13971 9746
rect 197 9688 202 9744
rect 258 9688 13910 9744
rect 13966 9688 13971 9744
rect 197 9686 13971 9688
rect 197 9683 263 9686
rect 13905 9683 13971 9686
rect 24669 9610 24735 9613
rect 25221 9610 25287 9613
rect 27520 9610 28000 9640
rect 24669 9608 28000 9610
rect 24669 9552 24674 9608
rect 24730 9552 25226 9608
rect 25282 9552 28000 9608
rect 24669 9550 28000 9552
rect 24669 9547 24735 9550
rect 25221 9547 25287 9550
rect 5610 9544 5930 9545
rect 5610 9480 5618 9544
rect 5682 9480 5698 9544
rect 5762 9480 5778 9544
rect 5842 9480 5858 9544
rect 5922 9480 5930 9544
rect 5610 9479 5930 9480
rect 14944 9544 15264 9545
rect 14944 9480 14952 9544
rect 15016 9480 15032 9544
rect 15096 9480 15112 9544
rect 15176 9480 15192 9544
rect 15256 9480 15264 9544
rect 14944 9479 15264 9480
rect 24277 9544 24597 9545
rect 24277 9480 24285 9544
rect 24349 9480 24365 9544
rect 24429 9480 24445 9544
rect 24509 9480 24525 9544
rect 24589 9480 24597 9544
rect 27520 9520 28000 9550
rect 24277 9479 24597 9480
rect 16389 9474 16455 9477
rect 19149 9474 19215 9477
rect 16389 9472 19215 9474
rect 16389 9416 16394 9472
rect 16450 9416 19154 9472
rect 19210 9416 19215 9472
rect 16389 9414 19215 9416
rect 16389 9411 16455 9414
rect 19149 9411 19215 9414
rect 20069 9338 20135 9341
rect 24761 9338 24827 9341
rect 20069 9336 24827 9338
rect 20069 9280 20074 9336
rect 20130 9280 24766 9336
rect 24822 9280 24827 9336
rect 20069 9278 24827 9280
rect 20069 9275 20135 9278
rect 24761 9275 24827 9278
rect 20437 9066 20503 9069
rect 24761 9066 24827 9069
rect 20437 9064 24827 9066
rect 20437 9008 20442 9064
rect 20498 9008 24766 9064
rect 24822 9008 24827 9064
rect 20437 9006 24827 9008
rect 20437 9003 20503 9006
rect 24761 9003 24827 9006
rect 10277 9000 10597 9001
rect 10277 8936 10285 9000
rect 10349 8936 10365 9000
rect 10429 8936 10445 9000
rect 10509 8936 10525 9000
rect 10589 8936 10597 9000
rect 10277 8935 10597 8936
rect 19610 9000 19930 9001
rect 19610 8936 19618 9000
rect 19682 8936 19698 9000
rect 19762 8936 19778 9000
rect 19842 8936 19858 9000
rect 19922 8936 19930 9000
rect 19610 8935 19930 8936
rect 24485 8930 24551 8933
rect 27520 8930 28000 8960
rect 24485 8928 28000 8930
rect 24485 8872 24490 8928
rect 24546 8872 28000 8928
rect 24485 8870 28000 8872
rect 24485 8867 24551 8870
rect 27520 8840 28000 8870
rect 5610 8456 5930 8457
rect 5610 8392 5618 8456
rect 5682 8392 5698 8456
rect 5762 8392 5778 8456
rect 5842 8392 5858 8456
rect 5922 8392 5930 8456
rect 5610 8391 5930 8392
rect 14944 8456 15264 8457
rect 14944 8392 14952 8456
rect 15016 8392 15032 8456
rect 15096 8392 15112 8456
rect 15176 8392 15192 8456
rect 15256 8392 15264 8456
rect 14944 8391 15264 8392
rect 24277 8456 24597 8457
rect 24277 8392 24285 8456
rect 24349 8392 24365 8456
rect 24429 8392 24445 8456
rect 24509 8392 24525 8456
rect 24589 8392 24597 8456
rect 24277 8391 24597 8392
rect 24669 8386 24735 8389
rect 27520 8386 28000 8416
rect 24669 8384 28000 8386
rect 24669 8328 24674 8384
rect 24730 8328 28000 8384
rect 24669 8326 28000 8328
rect 24669 8323 24735 8326
rect 27520 8296 28000 8326
rect 10277 7912 10597 7913
rect 10277 7848 10285 7912
rect 10349 7848 10365 7912
rect 10429 7848 10445 7912
rect 10509 7848 10525 7912
rect 10589 7848 10597 7912
rect 10277 7847 10597 7848
rect 19610 7912 19930 7913
rect 19610 7848 19618 7912
rect 19682 7848 19698 7912
rect 19762 7848 19778 7912
rect 19842 7848 19858 7912
rect 19922 7848 19930 7912
rect 19610 7847 19930 7848
rect 18873 7706 18939 7709
rect 24209 7706 24275 7709
rect 18873 7704 24275 7706
rect 18873 7648 18878 7704
rect 18934 7648 24214 7704
rect 24270 7648 24275 7704
rect 18873 7646 24275 7648
rect 18873 7643 18939 7646
rect 24209 7643 24275 7646
rect 24577 7706 24643 7709
rect 27520 7706 28000 7736
rect 24577 7704 28000 7706
rect 24577 7648 24582 7704
rect 24638 7648 28000 7704
rect 24577 7646 28000 7648
rect 24577 7643 24643 7646
rect 27520 7616 28000 7646
rect 18413 7570 18479 7573
rect 24761 7570 24827 7573
rect 18413 7568 24827 7570
rect 18413 7512 18418 7568
rect 18474 7512 24766 7568
rect 24822 7512 24827 7568
rect 18413 7510 24827 7512
rect 18413 7507 18479 7510
rect 24761 7507 24827 7510
rect 5610 7368 5930 7369
rect 5610 7304 5618 7368
rect 5682 7304 5698 7368
rect 5762 7304 5778 7368
rect 5842 7304 5858 7368
rect 5922 7304 5930 7368
rect 5610 7303 5930 7304
rect 14944 7368 15264 7369
rect 14944 7304 14952 7368
rect 15016 7304 15032 7368
rect 15096 7304 15112 7368
rect 15176 7304 15192 7368
rect 15256 7304 15264 7368
rect 14944 7303 15264 7304
rect 24277 7368 24597 7369
rect 24277 7304 24285 7368
rect 24349 7304 24365 7368
rect 24429 7304 24445 7368
rect 24509 7304 24525 7368
rect 24589 7304 24597 7368
rect 24277 7303 24597 7304
rect 18229 7162 18295 7165
rect 27520 7162 28000 7192
rect 18229 7160 28000 7162
rect 18229 7104 18234 7160
rect 18290 7104 28000 7160
rect 18229 7102 28000 7104
rect 18229 7099 18295 7102
rect 27520 7072 28000 7102
rect 10277 6824 10597 6825
rect 0 6754 480 6784
rect 10277 6760 10285 6824
rect 10349 6760 10365 6824
rect 10429 6760 10445 6824
rect 10509 6760 10525 6824
rect 10589 6760 10597 6824
rect 10277 6759 10597 6760
rect 19610 6824 19930 6825
rect 19610 6760 19618 6824
rect 19682 6760 19698 6824
rect 19762 6760 19778 6824
rect 19842 6760 19858 6824
rect 19922 6760 19930 6824
rect 19610 6759 19930 6760
rect 3417 6754 3483 6757
rect 0 6752 3483 6754
rect 0 6696 3422 6752
rect 3478 6696 3483 6752
rect 0 6694 3483 6696
rect 0 6664 480 6694
rect 3417 6691 3483 6694
rect 24209 6618 24275 6621
rect 27520 6618 28000 6648
rect 24209 6616 28000 6618
rect 24209 6560 24214 6616
rect 24270 6560 28000 6616
rect 24209 6558 28000 6560
rect 24209 6555 24275 6558
rect 27520 6528 28000 6558
rect 5610 6280 5930 6281
rect 5610 6216 5618 6280
rect 5682 6216 5698 6280
rect 5762 6216 5778 6280
rect 5842 6216 5858 6280
rect 5922 6216 5930 6280
rect 5610 6215 5930 6216
rect 14944 6280 15264 6281
rect 14944 6216 14952 6280
rect 15016 6216 15032 6280
rect 15096 6216 15112 6280
rect 15176 6216 15192 6280
rect 15256 6216 15264 6280
rect 14944 6215 15264 6216
rect 24277 6280 24597 6281
rect 24277 6216 24285 6280
rect 24349 6216 24365 6280
rect 24429 6216 24445 6280
rect 24509 6216 24525 6280
rect 24589 6216 24597 6280
rect 24277 6215 24597 6216
rect 16941 5938 17007 5941
rect 27520 5938 28000 5968
rect 16941 5936 28000 5938
rect 16941 5880 16946 5936
rect 17002 5880 28000 5936
rect 16941 5878 28000 5880
rect 16941 5875 17007 5878
rect 27520 5848 28000 5878
rect 10277 5736 10597 5737
rect 10277 5672 10285 5736
rect 10349 5672 10365 5736
rect 10429 5672 10445 5736
rect 10509 5672 10525 5736
rect 10589 5672 10597 5736
rect 10277 5671 10597 5672
rect 19610 5736 19930 5737
rect 19610 5672 19618 5736
rect 19682 5672 19698 5736
rect 19762 5672 19778 5736
rect 19842 5672 19858 5736
rect 19922 5672 19930 5736
rect 19610 5671 19930 5672
rect 16021 5394 16087 5397
rect 27520 5394 28000 5424
rect 16021 5392 28000 5394
rect 16021 5336 16026 5392
rect 16082 5336 28000 5392
rect 16021 5334 28000 5336
rect 16021 5331 16087 5334
rect 27520 5304 28000 5334
rect 5610 5192 5930 5193
rect 5610 5128 5618 5192
rect 5682 5128 5698 5192
rect 5762 5128 5778 5192
rect 5842 5128 5858 5192
rect 5922 5128 5930 5192
rect 5610 5127 5930 5128
rect 14944 5192 15264 5193
rect 14944 5128 14952 5192
rect 15016 5128 15032 5192
rect 15096 5128 15112 5192
rect 15176 5128 15192 5192
rect 15256 5128 15264 5192
rect 14944 5127 15264 5128
rect 24277 5192 24597 5193
rect 24277 5128 24285 5192
rect 24349 5128 24365 5192
rect 24429 5128 24445 5192
rect 24509 5128 24525 5192
rect 24589 5128 24597 5192
rect 24277 5127 24597 5128
rect 15929 4986 15995 4989
rect 15929 4984 27538 4986
rect 15929 4928 15934 4984
rect 15990 4928 27538 4984
rect 15929 4926 27538 4928
rect 15929 4923 15995 4926
rect 27478 4880 27538 4926
rect 27478 4790 28000 4880
rect 27520 4760 28000 4790
rect 10277 4648 10597 4649
rect 10277 4584 10285 4648
rect 10349 4584 10365 4648
rect 10429 4584 10445 4648
rect 10509 4584 10525 4648
rect 10589 4584 10597 4648
rect 10277 4583 10597 4584
rect 19610 4648 19930 4649
rect 19610 4584 19618 4648
rect 19682 4584 19698 4648
rect 19762 4584 19778 4648
rect 19842 4584 19858 4648
rect 19922 4584 19930 4648
rect 19610 4583 19930 4584
rect 24117 4306 24183 4309
rect 24117 4304 24778 4306
rect 24117 4248 24122 4304
rect 24178 4248 24778 4304
rect 24117 4246 24778 4248
rect 24117 4243 24183 4246
rect 24718 4170 24778 4246
rect 27520 4170 28000 4200
rect 24718 4110 28000 4170
rect 5610 4104 5930 4105
rect 5610 4040 5618 4104
rect 5682 4040 5698 4104
rect 5762 4040 5778 4104
rect 5842 4040 5858 4104
rect 5922 4040 5930 4104
rect 5610 4039 5930 4040
rect 14944 4104 15264 4105
rect 14944 4040 14952 4104
rect 15016 4040 15032 4104
rect 15096 4040 15112 4104
rect 15176 4040 15192 4104
rect 15256 4040 15264 4104
rect 14944 4039 15264 4040
rect 24277 4104 24597 4105
rect 24277 4040 24285 4104
rect 24349 4040 24365 4104
rect 24429 4040 24445 4104
rect 24509 4040 24525 4104
rect 24589 4040 24597 4104
rect 27520 4080 28000 4110
rect 24277 4039 24597 4040
rect 21633 3762 21699 3765
rect 23473 3762 23539 3765
rect 21633 3760 23539 3762
rect 21633 3704 21638 3760
rect 21694 3704 23478 3760
rect 23534 3704 23539 3760
rect 21633 3702 23539 3704
rect 21633 3699 21699 3702
rect 23473 3699 23539 3702
rect 24761 3762 24827 3765
rect 26233 3762 26299 3765
rect 24761 3760 26299 3762
rect 24761 3704 24766 3760
rect 24822 3704 26238 3760
rect 26294 3704 26299 3760
rect 24761 3702 26299 3704
rect 24761 3699 24827 3702
rect 26233 3699 26299 3702
rect 25221 3626 25287 3629
rect 27520 3626 28000 3656
rect 25221 3624 28000 3626
rect 25221 3568 25226 3624
rect 25282 3568 28000 3624
rect 25221 3566 28000 3568
rect 25221 3563 25287 3566
rect 10277 3560 10597 3561
rect 10277 3496 10285 3560
rect 10349 3496 10365 3560
rect 10429 3496 10445 3560
rect 10509 3496 10525 3560
rect 10589 3496 10597 3560
rect 10277 3495 10597 3496
rect 19610 3560 19930 3561
rect 19610 3496 19618 3560
rect 19682 3496 19698 3560
rect 19762 3496 19778 3560
rect 19842 3496 19858 3560
rect 19922 3496 19930 3560
rect 27520 3536 28000 3566
rect 19610 3495 19930 3496
rect 23565 3218 23631 3221
rect 23565 3216 25698 3218
rect 23565 3160 23570 3216
rect 23626 3160 25698 3216
rect 23565 3158 25698 3160
rect 23565 3155 23631 3158
rect 5610 3016 5930 3017
rect 5610 2952 5618 3016
rect 5682 2952 5698 3016
rect 5762 2952 5778 3016
rect 5842 2952 5858 3016
rect 5922 2952 5930 3016
rect 5610 2951 5930 2952
rect 14944 3016 15264 3017
rect 14944 2952 14952 3016
rect 15016 2952 15032 3016
rect 15096 2952 15112 3016
rect 15176 2952 15192 3016
rect 15256 2952 15264 3016
rect 14944 2951 15264 2952
rect 24277 3016 24597 3017
rect 24277 2952 24285 3016
rect 24349 2952 24365 3016
rect 24429 2952 24445 3016
rect 24509 2952 24525 3016
rect 24589 2952 24597 3016
rect 24277 2951 24597 2952
rect 25638 2946 25698 3158
rect 27520 2946 28000 2976
rect 25638 2886 28000 2946
rect 27520 2856 28000 2886
rect 10277 2472 10597 2473
rect 10277 2408 10285 2472
rect 10349 2408 10365 2472
rect 10429 2408 10445 2472
rect 10509 2408 10525 2472
rect 10589 2408 10597 2472
rect 10277 2407 10597 2408
rect 19610 2472 19930 2473
rect 19610 2408 19618 2472
rect 19682 2408 19698 2472
rect 19762 2408 19778 2472
rect 19842 2408 19858 2472
rect 19922 2408 19930 2472
rect 19610 2407 19930 2408
rect 22277 2402 22343 2405
rect 23565 2402 23631 2405
rect 22277 2400 23631 2402
rect 22277 2344 22282 2400
rect 22338 2344 23570 2400
rect 23626 2344 23631 2400
rect 22277 2342 23631 2344
rect 22277 2339 22343 2342
rect 23565 2339 23631 2342
rect 23841 2402 23907 2405
rect 27520 2402 28000 2432
rect 23841 2400 28000 2402
rect 23841 2344 23846 2400
rect 23902 2344 28000 2400
rect 23841 2342 28000 2344
rect 23841 2339 23907 2342
rect 27520 2312 28000 2342
rect 23933 2130 23999 2133
rect 23933 2128 27538 2130
rect 23933 2072 23938 2128
rect 23994 2072 27538 2128
rect 23933 2070 27538 2072
rect 23933 2067 23999 2070
rect 5610 1928 5930 1929
rect 5610 1864 5618 1928
rect 5682 1864 5698 1928
rect 5762 1864 5778 1928
rect 5842 1864 5858 1928
rect 5922 1864 5930 1928
rect 5610 1863 5930 1864
rect 14944 1928 15264 1929
rect 14944 1864 14952 1928
rect 15016 1864 15032 1928
rect 15096 1864 15112 1928
rect 15176 1864 15192 1928
rect 15256 1864 15264 1928
rect 14944 1863 15264 1864
rect 24277 1928 24597 1929
rect 24277 1864 24285 1928
rect 24349 1864 24365 1928
rect 24429 1864 24445 1928
rect 24509 1864 24525 1928
rect 24589 1864 24597 1928
rect 24277 1863 24597 1864
rect 27478 1888 27538 2070
rect 27478 1798 28000 1888
rect 27520 1768 28000 1798
rect 23473 1178 23539 1181
rect 27520 1178 28000 1208
rect 23473 1176 28000 1178
rect 23473 1120 23478 1176
rect 23534 1120 28000 1176
rect 23473 1118 28000 1120
rect 23473 1115 23539 1118
rect 27520 1088 28000 1118
rect 23657 634 23723 637
rect 27520 634 28000 664
rect 23657 632 28000 634
rect 23657 576 23662 632
rect 23718 576 28000 632
rect 23657 574 28000 576
rect 23657 571 23723 574
rect 27520 544 28000 574
rect 23565 90 23631 93
rect 27520 90 28000 120
rect 23565 88 28000 90
rect 23565 32 23570 88
rect 23626 32 28000 88
rect 23565 30 28000 32
rect 23565 27 23631 30
rect 27520 0 28000 30
<< via3 >>
rect 10285 25316 10349 25320
rect 10285 25260 10289 25316
rect 10289 25260 10345 25316
rect 10345 25260 10349 25316
rect 10285 25256 10349 25260
rect 10365 25316 10429 25320
rect 10365 25260 10369 25316
rect 10369 25260 10425 25316
rect 10425 25260 10429 25316
rect 10365 25256 10429 25260
rect 10445 25316 10509 25320
rect 10445 25260 10449 25316
rect 10449 25260 10505 25316
rect 10505 25260 10509 25316
rect 10445 25256 10509 25260
rect 10525 25316 10589 25320
rect 10525 25260 10529 25316
rect 10529 25260 10585 25316
rect 10585 25260 10589 25316
rect 10525 25256 10589 25260
rect 19618 25316 19682 25320
rect 19618 25260 19622 25316
rect 19622 25260 19678 25316
rect 19678 25260 19682 25316
rect 19618 25256 19682 25260
rect 19698 25316 19762 25320
rect 19698 25260 19702 25316
rect 19702 25260 19758 25316
rect 19758 25260 19762 25316
rect 19698 25256 19762 25260
rect 19778 25316 19842 25320
rect 19778 25260 19782 25316
rect 19782 25260 19838 25316
rect 19838 25260 19842 25316
rect 19778 25256 19842 25260
rect 19858 25316 19922 25320
rect 19858 25260 19862 25316
rect 19862 25260 19918 25316
rect 19918 25260 19922 25316
rect 19858 25256 19922 25260
rect 5618 24772 5682 24776
rect 5618 24716 5622 24772
rect 5622 24716 5678 24772
rect 5678 24716 5682 24772
rect 5618 24712 5682 24716
rect 5698 24772 5762 24776
rect 5698 24716 5702 24772
rect 5702 24716 5758 24772
rect 5758 24716 5762 24772
rect 5698 24712 5762 24716
rect 5778 24772 5842 24776
rect 5778 24716 5782 24772
rect 5782 24716 5838 24772
rect 5838 24716 5842 24772
rect 5778 24712 5842 24716
rect 5858 24772 5922 24776
rect 5858 24716 5862 24772
rect 5862 24716 5918 24772
rect 5918 24716 5922 24772
rect 5858 24712 5922 24716
rect 14952 24772 15016 24776
rect 14952 24716 14956 24772
rect 14956 24716 15012 24772
rect 15012 24716 15016 24772
rect 14952 24712 15016 24716
rect 15032 24772 15096 24776
rect 15032 24716 15036 24772
rect 15036 24716 15092 24772
rect 15092 24716 15096 24772
rect 15032 24712 15096 24716
rect 15112 24772 15176 24776
rect 15112 24716 15116 24772
rect 15116 24716 15172 24772
rect 15172 24716 15176 24772
rect 15112 24712 15176 24716
rect 15192 24772 15256 24776
rect 15192 24716 15196 24772
rect 15196 24716 15252 24772
rect 15252 24716 15256 24772
rect 15192 24712 15256 24716
rect 24285 24772 24349 24776
rect 24285 24716 24289 24772
rect 24289 24716 24345 24772
rect 24345 24716 24349 24772
rect 24285 24712 24349 24716
rect 24365 24772 24429 24776
rect 24365 24716 24369 24772
rect 24369 24716 24425 24772
rect 24425 24716 24429 24772
rect 24365 24712 24429 24716
rect 24445 24772 24509 24776
rect 24445 24716 24449 24772
rect 24449 24716 24505 24772
rect 24505 24716 24509 24772
rect 24445 24712 24509 24716
rect 24525 24772 24589 24776
rect 24525 24716 24529 24772
rect 24529 24716 24585 24772
rect 24585 24716 24589 24772
rect 24525 24712 24589 24716
rect 10285 24228 10349 24232
rect 10285 24172 10289 24228
rect 10289 24172 10345 24228
rect 10345 24172 10349 24228
rect 10285 24168 10349 24172
rect 10365 24228 10429 24232
rect 10365 24172 10369 24228
rect 10369 24172 10425 24228
rect 10425 24172 10429 24228
rect 10365 24168 10429 24172
rect 10445 24228 10509 24232
rect 10445 24172 10449 24228
rect 10449 24172 10505 24228
rect 10505 24172 10509 24228
rect 10445 24168 10509 24172
rect 10525 24228 10589 24232
rect 10525 24172 10529 24228
rect 10529 24172 10585 24228
rect 10585 24172 10589 24228
rect 10525 24168 10589 24172
rect 19618 24228 19682 24232
rect 19618 24172 19622 24228
rect 19622 24172 19678 24228
rect 19678 24172 19682 24228
rect 19618 24168 19682 24172
rect 19698 24228 19762 24232
rect 19698 24172 19702 24228
rect 19702 24172 19758 24228
rect 19758 24172 19762 24228
rect 19698 24168 19762 24172
rect 19778 24228 19842 24232
rect 19778 24172 19782 24228
rect 19782 24172 19838 24228
rect 19838 24172 19842 24228
rect 19778 24168 19842 24172
rect 19858 24228 19922 24232
rect 19858 24172 19862 24228
rect 19862 24172 19918 24228
rect 19918 24172 19922 24228
rect 19858 24168 19922 24172
rect 5618 23684 5682 23688
rect 5618 23628 5622 23684
rect 5622 23628 5678 23684
rect 5678 23628 5682 23684
rect 5618 23624 5682 23628
rect 5698 23684 5762 23688
rect 5698 23628 5702 23684
rect 5702 23628 5758 23684
rect 5758 23628 5762 23684
rect 5698 23624 5762 23628
rect 5778 23684 5842 23688
rect 5778 23628 5782 23684
rect 5782 23628 5838 23684
rect 5838 23628 5842 23684
rect 5778 23624 5842 23628
rect 5858 23684 5922 23688
rect 5858 23628 5862 23684
rect 5862 23628 5918 23684
rect 5918 23628 5922 23684
rect 5858 23624 5922 23628
rect 14952 23684 15016 23688
rect 14952 23628 14956 23684
rect 14956 23628 15012 23684
rect 15012 23628 15016 23684
rect 14952 23624 15016 23628
rect 15032 23684 15096 23688
rect 15032 23628 15036 23684
rect 15036 23628 15092 23684
rect 15092 23628 15096 23684
rect 15032 23624 15096 23628
rect 15112 23684 15176 23688
rect 15112 23628 15116 23684
rect 15116 23628 15172 23684
rect 15172 23628 15176 23684
rect 15112 23624 15176 23628
rect 15192 23684 15256 23688
rect 15192 23628 15196 23684
rect 15196 23628 15252 23684
rect 15252 23628 15256 23684
rect 15192 23624 15256 23628
rect 24285 23684 24349 23688
rect 24285 23628 24289 23684
rect 24289 23628 24345 23684
rect 24345 23628 24349 23684
rect 24285 23624 24349 23628
rect 24365 23684 24429 23688
rect 24365 23628 24369 23684
rect 24369 23628 24425 23684
rect 24425 23628 24429 23684
rect 24365 23624 24429 23628
rect 24445 23684 24509 23688
rect 24445 23628 24449 23684
rect 24449 23628 24505 23684
rect 24505 23628 24509 23684
rect 24445 23624 24509 23628
rect 24525 23684 24589 23688
rect 24525 23628 24529 23684
rect 24529 23628 24585 23684
rect 24585 23628 24589 23684
rect 24525 23624 24589 23628
rect 10285 23140 10349 23144
rect 10285 23084 10289 23140
rect 10289 23084 10345 23140
rect 10345 23084 10349 23140
rect 10285 23080 10349 23084
rect 10365 23140 10429 23144
rect 10365 23084 10369 23140
rect 10369 23084 10425 23140
rect 10425 23084 10429 23140
rect 10365 23080 10429 23084
rect 10445 23140 10509 23144
rect 10445 23084 10449 23140
rect 10449 23084 10505 23140
rect 10505 23084 10509 23140
rect 10445 23080 10509 23084
rect 10525 23140 10589 23144
rect 10525 23084 10529 23140
rect 10529 23084 10585 23140
rect 10585 23084 10589 23140
rect 10525 23080 10589 23084
rect 19618 23140 19682 23144
rect 19618 23084 19622 23140
rect 19622 23084 19678 23140
rect 19678 23084 19682 23140
rect 19618 23080 19682 23084
rect 19698 23140 19762 23144
rect 19698 23084 19702 23140
rect 19702 23084 19758 23140
rect 19758 23084 19762 23140
rect 19698 23080 19762 23084
rect 19778 23140 19842 23144
rect 19778 23084 19782 23140
rect 19782 23084 19838 23140
rect 19838 23084 19842 23140
rect 19778 23080 19842 23084
rect 19858 23140 19922 23144
rect 19858 23084 19862 23140
rect 19862 23084 19918 23140
rect 19918 23084 19922 23140
rect 19858 23080 19922 23084
rect 5618 22596 5682 22600
rect 5618 22540 5622 22596
rect 5622 22540 5678 22596
rect 5678 22540 5682 22596
rect 5618 22536 5682 22540
rect 5698 22596 5762 22600
rect 5698 22540 5702 22596
rect 5702 22540 5758 22596
rect 5758 22540 5762 22596
rect 5698 22536 5762 22540
rect 5778 22596 5842 22600
rect 5778 22540 5782 22596
rect 5782 22540 5838 22596
rect 5838 22540 5842 22596
rect 5778 22536 5842 22540
rect 5858 22596 5922 22600
rect 5858 22540 5862 22596
rect 5862 22540 5918 22596
rect 5918 22540 5922 22596
rect 5858 22536 5922 22540
rect 14952 22596 15016 22600
rect 14952 22540 14956 22596
rect 14956 22540 15012 22596
rect 15012 22540 15016 22596
rect 14952 22536 15016 22540
rect 15032 22596 15096 22600
rect 15032 22540 15036 22596
rect 15036 22540 15092 22596
rect 15092 22540 15096 22596
rect 15032 22536 15096 22540
rect 15112 22596 15176 22600
rect 15112 22540 15116 22596
rect 15116 22540 15172 22596
rect 15172 22540 15176 22596
rect 15112 22536 15176 22540
rect 15192 22596 15256 22600
rect 15192 22540 15196 22596
rect 15196 22540 15252 22596
rect 15252 22540 15256 22596
rect 15192 22536 15256 22540
rect 24285 22596 24349 22600
rect 24285 22540 24289 22596
rect 24289 22540 24345 22596
rect 24345 22540 24349 22596
rect 24285 22536 24349 22540
rect 24365 22596 24429 22600
rect 24365 22540 24369 22596
rect 24369 22540 24425 22596
rect 24425 22540 24429 22596
rect 24365 22536 24429 22540
rect 24445 22596 24509 22600
rect 24445 22540 24449 22596
rect 24449 22540 24505 22596
rect 24505 22540 24509 22596
rect 24445 22536 24509 22540
rect 24525 22596 24589 22600
rect 24525 22540 24529 22596
rect 24529 22540 24585 22596
rect 24585 22540 24589 22596
rect 24525 22536 24589 22540
rect 10285 22052 10349 22056
rect 10285 21996 10289 22052
rect 10289 21996 10345 22052
rect 10345 21996 10349 22052
rect 10285 21992 10349 21996
rect 10365 22052 10429 22056
rect 10365 21996 10369 22052
rect 10369 21996 10425 22052
rect 10425 21996 10429 22052
rect 10365 21992 10429 21996
rect 10445 22052 10509 22056
rect 10445 21996 10449 22052
rect 10449 21996 10505 22052
rect 10505 21996 10509 22052
rect 10445 21992 10509 21996
rect 10525 22052 10589 22056
rect 10525 21996 10529 22052
rect 10529 21996 10585 22052
rect 10585 21996 10589 22052
rect 10525 21992 10589 21996
rect 19618 22052 19682 22056
rect 19618 21996 19622 22052
rect 19622 21996 19678 22052
rect 19678 21996 19682 22052
rect 19618 21992 19682 21996
rect 19698 22052 19762 22056
rect 19698 21996 19702 22052
rect 19702 21996 19758 22052
rect 19758 21996 19762 22052
rect 19698 21992 19762 21996
rect 19778 22052 19842 22056
rect 19778 21996 19782 22052
rect 19782 21996 19838 22052
rect 19838 21996 19842 22052
rect 19778 21992 19842 21996
rect 19858 22052 19922 22056
rect 19858 21996 19862 22052
rect 19862 21996 19918 22052
rect 19918 21996 19922 22052
rect 19858 21992 19922 21996
rect 5618 21508 5682 21512
rect 5618 21452 5622 21508
rect 5622 21452 5678 21508
rect 5678 21452 5682 21508
rect 5618 21448 5682 21452
rect 5698 21508 5762 21512
rect 5698 21452 5702 21508
rect 5702 21452 5758 21508
rect 5758 21452 5762 21508
rect 5698 21448 5762 21452
rect 5778 21508 5842 21512
rect 5778 21452 5782 21508
rect 5782 21452 5838 21508
rect 5838 21452 5842 21508
rect 5778 21448 5842 21452
rect 5858 21508 5922 21512
rect 5858 21452 5862 21508
rect 5862 21452 5918 21508
rect 5918 21452 5922 21508
rect 5858 21448 5922 21452
rect 14952 21508 15016 21512
rect 14952 21452 14956 21508
rect 14956 21452 15012 21508
rect 15012 21452 15016 21508
rect 14952 21448 15016 21452
rect 15032 21508 15096 21512
rect 15032 21452 15036 21508
rect 15036 21452 15092 21508
rect 15092 21452 15096 21508
rect 15032 21448 15096 21452
rect 15112 21508 15176 21512
rect 15112 21452 15116 21508
rect 15116 21452 15172 21508
rect 15172 21452 15176 21508
rect 15112 21448 15176 21452
rect 15192 21508 15256 21512
rect 15192 21452 15196 21508
rect 15196 21452 15252 21508
rect 15252 21452 15256 21508
rect 15192 21448 15256 21452
rect 24285 21508 24349 21512
rect 24285 21452 24289 21508
rect 24289 21452 24345 21508
rect 24345 21452 24349 21508
rect 24285 21448 24349 21452
rect 24365 21508 24429 21512
rect 24365 21452 24369 21508
rect 24369 21452 24425 21508
rect 24425 21452 24429 21508
rect 24365 21448 24429 21452
rect 24445 21508 24509 21512
rect 24445 21452 24449 21508
rect 24449 21452 24505 21508
rect 24505 21452 24509 21508
rect 24445 21448 24509 21452
rect 24525 21508 24589 21512
rect 24525 21452 24529 21508
rect 24529 21452 24585 21508
rect 24585 21452 24589 21508
rect 24525 21448 24589 21452
rect 10285 20964 10349 20968
rect 10285 20908 10289 20964
rect 10289 20908 10345 20964
rect 10345 20908 10349 20964
rect 10285 20904 10349 20908
rect 10365 20964 10429 20968
rect 10365 20908 10369 20964
rect 10369 20908 10425 20964
rect 10425 20908 10429 20964
rect 10365 20904 10429 20908
rect 10445 20964 10509 20968
rect 10445 20908 10449 20964
rect 10449 20908 10505 20964
rect 10505 20908 10509 20964
rect 10445 20904 10509 20908
rect 10525 20964 10589 20968
rect 10525 20908 10529 20964
rect 10529 20908 10585 20964
rect 10585 20908 10589 20964
rect 10525 20904 10589 20908
rect 19618 20964 19682 20968
rect 19618 20908 19622 20964
rect 19622 20908 19678 20964
rect 19678 20908 19682 20964
rect 19618 20904 19682 20908
rect 19698 20964 19762 20968
rect 19698 20908 19702 20964
rect 19702 20908 19758 20964
rect 19758 20908 19762 20964
rect 19698 20904 19762 20908
rect 19778 20964 19842 20968
rect 19778 20908 19782 20964
rect 19782 20908 19838 20964
rect 19838 20908 19842 20964
rect 19778 20904 19842 20908
rect 19858 20964 19922 20968
rect 19858 20908 19862 20964
rect 19862 20908 19918 20964
rect 19918 20908 19922 20964
rect 19858 20904 19922 20908
rect 5618 20420 5682 20424
rect 5618 20364 5622 20420
rect 5622 20364 5678 20420
rect 5678 20364 5682 20420
rect 5618 20360 5682 20364
rect 5698 20420 5762 20424
rect 5698 20364 5702 20420
rect 5702 20364 5758 20420
rect 5758 20364 5762 20420
rect 5698 20360 5762 20364
rect 5778 20420 5842 20424
rect 5778 20364 5782 20420
rect 5782 20364 5838 20420
rect 5838 20364 5842 20420
rect 5778 20360 5842 20364
rect 5858 20420 5922 20424
rect 5858 20364 5862 20420
rect 5862 20364 5918 20420
rect 5918 20364 5922 20420
rect 5858 20360 5922 20364
rect 14952 20420 15016 20424
rect 14952 20364 14956 20420
rect 14956 20364 15012 20420
rect 15012 20364 15016 20420
rect 14952 20360 15016 20364
rect 15032 20420 15096 20424
rect 15032 20364 15036 20420
rect 15036 20364 15092 20420
rect 15092 20364 15096 20420
rect 15032 20360 15096 20364
rect 15112 20420 15176 20424
rect 15112 20364 15116 20420
rect 15116 20364 15172 20420
rect 15172 20364 15176 20420
rect 15112 20360 15176 20364
rect 15192 20420 15256 20424
rect 15192 20364 15196 20420
rect 15196 20364 15252 20420
rect 15252 20364 15256 20420
rect 15192 20360 15256 20364
rect 24285 20420 24349 20424
rect 24285 20364 24289 20420
rect 24289 20364 24345 20420
rect 24345 20364 24349 20420
rect 24285 20360 24349 20364
rect 24365 20420 24429 20424
rect 24365 20364 24369 20420
rect 24369 20364 24425 20420
rect 24425 20364 24429 20420
rect 24365 20360 24429 20364
rect 24445 20420 24509 20424
rect 24445 20364 24449 20420
rect 24449 20364 24505 20420
rect 24505 20364 24509 20420
rect 24445 20360 24509 20364
rect 24525 20420 24589 20424
rect 24525 20364 24529 20420
rect 24529 20364 24585 20420
rect 24585 20364 24589 20420
rect 24525 20360 24589 20364
rect 10285 19876 10349 19880
rect 10285 19820 10289 19876
rect 10289 19820 10345 19876
rect 10345 19820 10349 19876
rect 10285 19816 10349 19820
rect 10365 19876 10429 19880
rect 10365 19820 10369 19876
rect 10369 19820 10425 19876
rect 10425 19820 10429 19876
rect 10365 19816 10429 19820
rect 10445 19876 10509 19880
rect 10445 19820 10449 19876
rect 10449 19820 10505 19876
rect 10505 19820 10509 19876
rect 10445 19816 10509 19820
rect 10525 19876 10589 19880
rect 10525 19820 10529 19876
rect 10529 19820 10585 19876
rect 10585 19820 10589 19876
rect 10525 19816 10589 19820
rect 19618 19876 19682 19880
rect 19618 19820 19622 19876
rect 19622 19820 19678 19876
rect 19678 19820 19682 19876
rect 19618 19816 19682 19820
rect 19698 19876 19762 19880
rect 19698 19820 19702 19876
rect 19702 19820 19758 19876
rect 19758 19820 19762 19876
rect 19698 19816 19762 19820
rect 19778 19876 19842 19880
rect 19778 19820 19782 19876
rect 19782 19820 19838 19876
rect 19838 19820 19842 19876
rect 19778 19816 19842 19820
rect 19858 19876 19922 19880
rect 19858 19820 19862 19876
rect 19862 19820 19918 19876
rect 19918 19820 19922 19876
rect 19858 19816 19922 19820
rect 5618 19332 5682 19336
rect 5618 19276 5622 19332
rect 5622 19276 5678 19332
rect 5678 19276 5682 19332
rect 5618 19272 5682 19276
rect 5698 19332 5762 19336
rect 5698 19276 5702 19332
rect 5702 19276 5758 19332
rect 5758 19276 5762 19332
rect 5698 19272 5762 19276
rect 5778 19332 5842 19336
rect 5778 19276 5782 19332
rect 5782 19276 5838 19332
rect 5838 19276 5842 19332
rect 5778 19272 5842 19276
rect 5858 19332 5922 19336
rect 5858 19276 5862 19332
rect 5862 19276 5918 19332
rect 5918 19276 5922 19332
rect 5858 19272 5922 19276
rect 14952 19332 15016 19336
rect 14952 19276 14956 19332
rect 14956 19276 15012 19332
rect 15012 19276 15016 19332
rect 14952 19272 15016 19276
rect 15032 19332 15096 19336
rect 15032 19276 15036 19332
rect 15036 19276 15092 19332
rect 15092 19276 15096 19332
rect 15032 19272 15096 19276
rect 15112 19332 15176 19336
rect 15112 19276 15116 19332
rect 15116 19276 15172 19332
rect 15172 19276 15176 19332
rect 15112 19272 15176 19276
rect 15192 19332 15256 19336
rect 15192 19276 15196 19332
rect 15196 19276 15252 19332
rect 15252 19276 15256 19332
rect 15192 19272 15256 19276
rect 24285 19332 24349 19336
rect 24285 19276 24289 19332
rect 24289 19276 24345 19332
rect 24345 19276 24349 19332
rect 24285 19272 24349 19276
rect 24365 19332 24429 19336
rect 24365 19276 24369 19332
rect 24369 19276 24425 19332
rect 24425 19276 24429 19332
rect 24365 19272 24429 19276
rect 24445 19332 24509 19336
rect 24445 19276 24449 19332
rect 24449 19276 24505 19332
rect 24505 19276 24509 19332
rect 24445 19272 24509 19276
rect 24525 19332 24589 19336
rect 24525 19276 24529 19332
rect 24529 19276 24585 19332
rect 24585 19276 24589 19332
rect 24525 19272 24589 19276
rect 10285 18788 10349 18792
rect 10285 18732 10289 18788
rect 10289 18732 10345 18788
rect 10345 18732 10349 18788
rect 10285 18728 10349 18732
rect 10365 18788 10429 18792
rect 10365 18732 10369 18788
rect 10369 18732 10425 18788
rect 10425 18732 10429 18788
rect 10365 18728 10429 18732
rect 10445 18788 10509 18792
rect 10445 18732 10449 18788
rect 10449 18732 10505 18788
rect 10505 18732 10509 18788
rect 10445 18728 10509 18732
rect 10525 18788 10589 18792
rect 10525 18732 10529 18788
rect 10529 18732 10585 18788
rect 10585 18732 10589 18788
rect 10525 18728 10589 18732
rect 19618 18788 19682 18792
rect 19618 18732 19622 18788
rect 19622 18732 19678 18788
rect 19678 18732 19682 18788
rect 19618 18728 19682 18732
rect 19698 18788 19762 18792
rect 19698 18732 19702 18788
rect 19702 18732 19758 18788
rect 19758 18732 19762 18788
rect 19698 18728 19762 18732
rect 19778 18788 19842 18792
rect 19778 18732 19782 18788
rect 19782 18732 19838 18788
rect 19838 18732 19842 18788
rect 19778 18728 19842 18732
rect 19858 18788 19922 18792
rect 19858 18732 19862 18788
rect 19862 18732 19918 18788
rect 19918 18732 19922 18788
rect 19858 18728 19922 18732
rect 5618 18244 5682 18248
rect 5618 18188 5622 18244
rect 5622 18188 5678 18244
rect 5678 18188 5682 18244
rect 5618 18184 5682 18188
rect 5698 18244 5762 18248
rect 5698 18188 5702 18244
rect 5702 18188 5758 18244
rect 5758 18188 5762 18244
rect 5698 18184 5762 18188
rect 5778 18244 5842 18248
rect 5778 18188 5782 18244
rect 5782 18188 5838 18244
rect 5838 18188 5842 18244
rect 5778 18184 5842 18188
rect 5858 18244 5922 18248
rect 5858 18188 5862 18244
rect 5862 18188 5918 18244
rect 5918 18188 5922 18244
rect 5858 18184 5922 18188
rect 14952 18244 15016 18248
rect 14952 18188 14956 18244
rect 14956 18188 15012 18244
rect 15012 18188 15016 18244
rect 14952 18184 15016 18188
rect 15032 18244 15096 18248
rect 15032 18188 15036 18244
rect 15036 18188 15092 18244
rect 15092 18188 15096 18244
rect 15032 18184 15096 18188
rect 15112 18244 15176 18248
rect 15112 18188 15116 18244
rect 15116 18188 15172 18244
rect 15172 18188 15176 18244
rect 15112 18184 15176 18188
rect 15192 18244 15256 18248
rect 15192 18188 15196 18244
rect 15196 18188 15252 18244
rect 15252 18188 15256 18244
rect 15192 18184 15256 18188
rect 24285 18244 24349 18248
rect 24285 18188 24289 18244
rect 24289 18188 24345 18244
rect 24345 18188 24349 18244
rect 24285 18184 24349 18188
rect 24365 18244 24429 18248
rect 24365 18188 24369 18244
rect 24369 18188 24425 18244
rect 24425 18188 24429 18244
rect 24365 18184 24429 18188
rect 24445 18244 24509 18248
rect 24445 18188 24449 18244
rect 24449 18188 24505 18244
rect 24505 18188 24509 18244
rect 24445 18184 24509 18188
rect 24525 18244 24589 18248
rect 24525 18188 24529 18244
rect 24529 18188 24585 18244
rect 24585 18188 24589 18244
rect 24525 18184 24589 18188
rect 10285 17700 10349 17704
rect 10285 17644 10289 17700
rect 10289 17644 10345 17700
rect 10345 17644 10349 17700
rect 10285 17640 10349 17644
rect 10365 17700 10429 17704
rect 10365 17644 10369 17700
rect 10369 17644 10425 17700
rect 10425 17644 10429 17700
rect 10365 17640 10429 17644
rect 10445 17700 10509 17704
rect 10445 17644 10449 17700
rect 10449 17644 10505 17700
rect 10505 17644 10509 17700
rect 10445 17640 10509 17644
rect 10525 17700 10589 17704
rect 10525 17644 10529 17700
rect 10529 17644 10585 17700
rect 10585 17644 10589 17700
rect 10525 17640 10589 17644
rect 19618 17700 19682 17704
rect 19618 17644 19622 17700
rect 19622 17644 19678 17700
rect 19678 17644 19682 17700
rect 19618 17640 19682 17644
rect 19698 17700 19762 17704
rect 19698 17644 19702 17700
rect 19702 17644 19758 17700
rect 19758 17644 19762 17700
rect 19698 17640 19762 17644
rect 19778 17700 19842 17704
rect 19778 17644 19782 17700
rect 19782 17644 19838 17700
rect 19838 17644 19842 17700
rect 19778 17640 19842 17644
rect 19858 17700 19922 17704
rect 19858 17644 19862 17700
rect 19862 17644 19918 17700
rect 19918 17644 19922 17700
rect 19858 17640 19922 17644
rect 5618 17156 5682 17160
rect 5618 17100 5622 17156
rect 5622 17100 5678 17156
rect 5678 17100 5682 17156
rect 5618 17096 5682 17100
rect 5698 17156 5762 17160
rect 5698 17100 5702 17156
rect 5702 17100 5758 17156
rect 5758 17100 5762 17156
rect 5698 17096 5762 17100
rect 5778 17156 5842 17160
rect 5778 17100 5782 17156
rect 5782 17100 5838 17156
rect 5838 17100 5842 17156
rect 5778 17096 5842 17100
rect 5858 17156 5922 17160
rect 5858 17100 5862 17156
rect 5862 17100 5918 17156
rect 5918 17100 5922 17156
rect 5858 17096 5922 17100
rect 14952 17156 15016 17160
rect 14952 17100 14956 17156
rect 14956 17100 15012 17156
rect 15012 17100 15016 17156
rect 14952 17096 15016 17100
rect 15032 17156 15096 17160
rect 15032 17100 15036 17156
rect 15036 17100 15092 17156
rect 15092 17100 15096 17156
rect 15032 17096 15096 17100
rect 15112 17156 15176 17160
rect 15112 17100 15116 17156
rect 15116 17100 15172 17156
rect 15172 17100 15176 17156
rect 15112 17096 15176 17100
rect 15192 17156 15256 17160
rect 15192 17100 15196 17156
rect 15196 17100 15252 17156
rect 15252 17100 15256 17156
rect 15192 17096 15256 17100
rect 24285 17156 24349 17160
rect 24285 17100 24289 17156
rect 24289 17100 24345 17156
rect 24345 17100 24349 17156
rect 24285 17096 24349 17100
rect 24365 17156 24429 17160
rect 24365 17100 24369 17156
rect 24369 17100 24425 17156
rect 24425 17100 24429 17156
rect 24365 17096 24429 17100
rect 24445 17156 24509 17160
rect 24445 17100 24449 17156
rect 24449 17100 24505 17156
rect 24505 17100 24509 17156
rect 24445 17096 24509 17100
rect 24525 17156 24589 17160
rect 24525 17100 24529 17156
rect 24529 17100 24585 17156
rect 24585 17100 24589 17156
rect 24525 17096 24589 17100
rect 10285 16612 10349 16616
rect 10285 16556 10289 16612
rect 10289 16556 10345 16612
rect 10345 16556 10349 16612
rect 10285 16552 10349 16556
rect 10365 16612 10429 16616
rect 10365 16556 10369 16612
rect 10369 16556 10425 16612
rect 10425 16556 10429 16612
rect 10365 16552 10429 16556
rect 10445 16612 10509 16616
rect 10445 16556 10449 16612
rect 10449 16556 10505 16612
rect 10505 16556 10509 16612
rect 10445 16552 10509 16556
rect 10525 16612 10589 16616
rect 10525 16556 10529 16612
rect 10529 16556 10585 16612
rect 10585 16556 10589 16612
rect 10525 16552 10589 16556
rect 19618 16612 19682 16616
rect 19618 16556 19622 16612
rect 19622 16556 19678 16612
rect 19678 16556 19682 16612
rect 19618 16552 19682 16556
rect 19698 16612 19762 16616
rect 19698 16556 19702 16612
rect 19702 16556 19758 16612
rect 19758 16556 19762 16612
rect 19698 16552 19762 16556
rect 19778 16612 19842 16616
rect 19778 16556 19782 16612
rect 19782 16556 19838 16612
rect 19838 16556 19842 16612
rect 19778 16552 19842 16556
rect 19858 16612 19922 16616
rect 19858 16556 19862 16612
rect 19862 16556 19918 16612
rect 19918 16556 19922 16612
rect 19858 16552 19922 16556
rect 5618 16068 5682 16072
rect 5618 16012 5622 16068
rect 5622 16012 5678 16068
rect 5678 16012 5682 16068
rect 5618 16008 5682 16012
rect 5698 16068 5762 16072
rect 5698 16012 5702 16068
rect 5702 16012 5758 16068
rect 5758 16012 5762 16068
rect 5698 16008 5762 16012
rect 5778 16068 5842 16072
rect 5778 16012 5782 16068
rect 5782 16012 5838 16068
rect 5838 16012 5842 16068
rect 5778 16008 5842 16012
rect 5858 16068 5922 16072
rect 5858 16012 5862 16068
rect 5862 16012 5918 16068
rect 5918 16012 5922 16068
rect 5858 16008 5922 16012
rect 14952 16068 15016 16072
rect 14952 16012 14956 16068
rect 14956 16012 15012 16068
rect 15012 16012 15016 16068
rect 14952 16008 15016 16012
rect 15032 16068 15096 16072
rect 15032 16012 15036 16068
rect 15036 16012 15092 16068
rect 15092 16012 15096 16068
rect 15032 16008 15096 16012
rect 15112 16068 15176 16072
rect 15112 16012 15116 16068
rect 15116 16012 15172 16068
rect 15172 16012 15176 16068
rect 15112 16008 15176 16012
rect 15192 16068 15256 16072
rect 15192 16012 15196 16068
rect 15196 16012 15252 16068
rect 15252 16012 15256 16068
rect 15192 16008 15256 16012
rect 24285 16068 24349 16072
rect 24285 16012 24289 16068
rect 24289 16012 24345 16068
rect 24345 16012 24349 16068
rect 24285 16008 24349 16012
rect 24365 16068 24429 16072
rect 24365 16012 24369 16068
rect 24369 16012 24425 16068
rect 24425 16012 24429 16068
rect 24365 16008 24429 16012
rect 24445 16068 24509 16072
rect 24445 16012 24449 16068
rect 24449 16012 24505 16068
rect 24505 16012 24509 16068
rect 24445 16008 24509 16012
rect 24525 16068 24589 16072
rect 24525 16012 24529 16068
rect 24529 16012 24585 16068
rect 24585 16012 24589 16068
rect 24525 16008 24589 16012
rect 10285 15524 10349 15528
rect 10285 15468 10289 15524
rect 10289 15468 10345 15524
rect 10345 15468 10349 15524
rect 10285 15464 10349 15468
rect 10365 15524 10429 15528
rect 10365 15468 10369 15524
rect 10369 15468 10425 15524
rect 10425 15468 10429 15524
rect 10365 15464 10429 15468
rect 10445 15524 10509 15528
rect 10445 15468 10449 15524
rect 10449 15468 10505 15524
rect 10505 15468 10509 15524
rect 10445 15464 10509 15468
rect 10525 15524 10589 15528
rect 10525 15468 10529 15524
rect 10529 15468 10585 15524
rect 10585 15468 10589 15524
rect 10525 15464 10589 15468
rect 19618 15524 19682 15528
rect 19618 15468 19622 15524
rect 19622 15468 19678 15524
rect 19678 15468 19682 15524
rect 19618 15464 19682 15468
rect 19698 15524 19762 15528
rect 19698 15468 19702 15524
rect 19702 15468 19758 15524
rect 19758 15468 19762 15524
rect 19698 15464 19762 15468
rect 19778 15524 19842 15528
rect 19778 15468 19782 15524
rect 19782 15468 19838 15524
rect 19838 15468 19842 15524
rect 19778 15464 19842 15468
rect 19858 15524 19922 15528
rect 19858 15468 19862 15524
rect 19862 15468 19918 15524
rect 19918 15468 19922 15524
rect 19858 15464 19922 15468
rect 5618 14980 5682 14984
rect 5618 14924 5622 14980
rect 5622 14924 5678 14980
rect 5678 14924 5682 14980
rect 5618 14920 5682 14924
rect 5698 14980 5762 14984
rect 5698 14924 5702 14980
rect 5702 14924 5758 14980
rect 5758 14924 5762 14980
rect 5698 14920 5762 14924
rect 5778 14980 5842 14984
rect 5778 14924 5782 14980
rect 5782 14924 5838 14980
rect 5838 14924 5842 14980
rect 5778 14920 5842 14924
rect 5858 14980 5922 14984
rect 5858 14924 5862 14980
rect 5862 14924 5918 14980
rect 5918 14924 5922 14980
rect 5858 14920 5922 14924
rect 14952 14980 15016 14984
rect 14952 14924 14956 14980
rect 14956 14924 15012 14980
rect 15012 14924 15016 14980
rect 14952 14920 15016 14924
rect 15032 14980 15096 14984
rect 15032 14924 15036 14980
rect 15036 14924 15092 14980
rect 15092 14924 15096 14980
rect 15032 14920 15096 14924
rect 15112 14980 15176 14984
rect 15112 14924 15116 14980
rect 15116 14924 15172 14980
rect 15172 14924 15176 14980
rect 15112 14920 15176 14924
rect 15192 14980 15256 14984
rect 15192 14924 15196 14980
rect 15196 14924 15252 14980
rect 15252 14924 15256 14980
rect 15192 14920 15256 14924
rect 24285 14980 24349 14984
rect 24285 14924 24289 14980
rect 24289 14924 24345 14980
rect 24345 14924 24349 14980
rect 24285 14920 24349 14924
rect 24365 14980 24429 14984
rect 24365 14924 24369 14980
rect 24369 14924 24425 14980
rect 24425 14924 24429 14980
rect 24365 14920 24429 14924
rect 24445 14980 24509 14984
rect 24445 14924 24449 14980
rect 24449 14924 24505 14980
rect 24505 14924 24509 14980
rect 24445 14920 24509 14924
rect 24525 14980 24589 14984
rect 24525 14924 24529 14980
rect 24529 14924 24585 14980
rect 24585 14924 24589 14980
rect 24525 14920 24589 14924
rect 10285 14436 10349 14440
rect 10285 14380 10289 14436
rect 10289 14380 10345 14436
rect 10345 14380 10349 14436
rect 10285 14376 10349 14380
rect 10365 14436 10429 14440
rect 10365 14380 10369 14436
rect 10369 14380 10425 14436
rect 10425 14380 10429 14436
rect 10365 14376 10429 14380
rect 10445 14436 10509 14440
rect 10445 14380 10449 14436
rect 10449 14380 10505 14436
rect 10505 14380 10509 14436
rect 10445 14376 10509 14380
rect 10525 14436 10589 14440
rect 10525 14380 10529 14436
rect 10529 14380 10585 14436
rect 10585 14380 10589 14436
rect 10525 14376 10589 14380
rect 19618 14436 19682 14440
rect 19618 14380 19622 14436
rect 19622 14380 19678 14436
rect 19678 14380 19682 14436
rect 19618 14376 19682 14380
rect 19698 14436 19762 14440
rect 19698 14380 19702 14436
rect 19702 14380 19758 14436
rect 19758 14380 19762 14436
rect 19698 14376 19762 14380
rect 19778 14436 19842 14440
rect 19778 14380 19782 14436
rect 19782 14380 19838 14436
rect 19838 14380 19842 14436
rect 19778 14376 19842 14380
rect 19858 14436 19922 14440
rect 19858 14380 19862 14436
rect 19862 14380 19918 14436
rect 19918 14380 19922 14436
rect 19858 14376 19922 14380
rect 5618 13892 5682 13896
rect 5618 13836 5622 13892
rect 5622 13836 5678 13892
rect 5678 13836 5682 13892
rect 5618 13832 5682 13836
rect 5698 13892 5762 13896
rect 5698 13836 5702 13892
rect 5702 13836 5758 13892
rect 5758 13836 5762 13892
rect 5698 13832 5762 13836
rect 5778 13892 5842 13896
rect 5778 13836 5782 13892
rect 5782 13836 5838 13892
rect 5838 13836 5842 13892
rect 5778 13832 5842 13836
rect 5858 13892 5922 13896
rect 5858 13836 5862 13892
rect 5862 13836 5918 13892
rect 5918 13836 5922 13892
rect 5858 13832 5922 13836
rect 14952 13892 15016 13896
rect 14952 13836 14956 13892
rect 14956 13836 15012 13892
rect 15012 13836 15016 13892
rect 14952 13832 15016 13836
rect 15032 13892 15096 13896
rect 15032 13836 15036 13892
rect 15036 13836 15092 13892
rect 15092 13836 15096 13892
rect 15032 13832 15096 13836
rect 15112 13892 15176 13896
rect 15112 13836 15116 13892
rect 15116 13836 15172 13892
rect 15172 13836 15176 13892
rect 15112 13832 15176 13836
rect 15192 13892 15256 13896
rect 15192 13836 15196 13892
rect 15196 13836 15252 13892
rect 15252 13836 15256 13892
rect 15192 13832 15256 13836
rect 24285 13892 24349 13896
rect 24285 13836 24289 13892
rect 24289 13836 24345 13892
rect 24345 13836 24349 13892
rect 24285 13832 24349 13836
rect 24365 13892 24429 13896
rect 24365 13836 24369 13892
rect 24369 13836 24425 13892
rect 24425 13836 24429 13892
rect 24365 13832 24429 13836
rect 24445 13892 24509 13896
rect 24445 13836 24449 13892
rect 24449 13836 24505 13892
rect 24505 13836 24509 13892
rect 24445 13832 24509 13836
rect 24525 13892 24589 13896
rect 24525 13836 24529 13892
rect 24529 13836 24585 13892
rect 24585 13836 24589 13892
rect 24525 13832 24589 13836
rect 10285 13348 10349 13352
rect 10285 13292 10289 13348
rect 10289 13292 10345 13348
rect 10345 13292 10349 13348
rect 10285 13288 10349 13292
rect 10365 13348 10429 13352
rect 10365 13292 10369 13348
rect 10369 13292 10425 13348
rect 10425 13292 10429 13348
rect 10365 13288 10429 13292
rect 10445 13348 10509 13352
rect 10445 13292 10449 13348
rect 10449 13292 10505 13348
rect 10505 13292 10509 13348
rect 10445 13288 10509 13292
rect 10525 13348 10589 13352
rect 10525 13292 10529 13348
rect 10529 13292 10585 13348
rect 10585 13292 10589 13348
rect 10525 13288 10589 13292
rect 19618 13348 19682 13352
rect 19618 13292 19622 13348
rect 19622 13292 19678 13348
rect 19678 13292 19682 13348
rect 19618 13288 19682 13292
rect 19698 13348 19762 13352
rect 19698 13292 19702 13348
rect 19702 13292 19758 13348
rect 19758 13292 19762 13348
rect 19698 13288 19762 13292
rect 19778 13348 19842 13352
rect 19778 13292 19782 13348
rect 19782 13292 19838 13348
rect 19838 13292 19842 13348
rect 19778 13288 19842 13292
rect 19858 13348 19922 13352
rect 19858 13292 19862 13348
rect 19862 13292 19918 13348
rect 19918 13292 19922 13348
rect 19858 13288 19922 13292
rect 5618 12804 5682 12808
rect 5618 12748 5622 12804
rect 5622 12748 5678 12804
rect 5678 12748 5682 12804
rect 5618 12744 5682 12748
rect 5698 12804 5762 12808
rect 5698 12748 5702 12804
rect 5702 12748 5758 12804
rect 5758 12748 5762 12804
rect 5698 12744 5762 12748
rect 5778 12804 5842 12808
rect 5778 12748 5782 12804
rect 5782 12748 5838 12804
rect 5838 12748 5842 12804
rect 5778 12744 5842 12748
rect 5858 12804 5922 12808
rect 5858 12748 5862 12804
rect 5862 12748 5918 12804
rect 5918 12748 5922 12804
rect 5858 12744 5922 12748
rect 14952 12804 15016 12808
rect 14952 12748 14956 12804
rect 14956 12748 15012 12804
rect 15012 12748 15016 12804
rect 14952 12744 15016 12748
rect 15032 12804 15096 12808
rect 15032 12748 15036 12804
rect 15036 12748 15092 12804
rect 15092 12748 15096 12804
rect 15032 12744 15096 12748
rect 15112 12804 15176 12808
rect 15112 12748 15116 12804
rect 15116 12748 15172 12804
rect 15172 12748 15176 12804
rect 15112 12744 15176 12748
rect 15192 12804 15256 12808
rect 15192 12748 15196 12804
rect 15196 12748 15252 12804
rect 15252 12748 15256 12804
rect 15192 12744 15256 12748
rect 24285 12804 24349 12808
rect 24285 12748 24289 12804
rect 24289 12748 24345 12804
rect 24345 12748 24349 12804
rect 24285 12744 24349 12748
rect 24365 12804 24429 12808
rect 24365 12748 24369 12804
rect 24369 12748 24425 12804
rect 24425 12748 24429 12804
rect 24365 12744 24429 12748
rect 24445 12804 24509 12808
rect 24445 12748 24449 12804
rect 24449 12748 24505 12804
rect 24505 12748 24509 12804
rect 24445 12744 24509 12748
rect 24525 12804 24589 12808
rect 24525 12748 24529 12804
rect 24529 12748 24585 12804
rect 24585 12748 24589 12804
rect 24525 12744 24589 12748
rect 10285 12260 10349 12264
rect 10285 12204 10289 12260
rect 10289 12204 10345 12260
rect 10345 12204 10349 12260
rect 10285 12200 10349 12204
rect 10365 12260 10429 12264
rect 10365 12204 10369 12260
rect 10369 12204 10425 12260
rect 10425 12204 10429 12260
rect 10365 12200 10429 12204
rect 10445 12260 10509 12264
rect 10445 12204 10449 12260
rect 10449 12204 10505 12260
rect 10505 12204 10509 12260
rect 10445 12200 10509 12204
rect 10525 12260 10589 12264
rect 10525 12204 10529 12260
rect 10529 12204 10585 12260
rect 10585 12204 10589 12260
rect 10525 12200 10589 12204
rect 19618 12260 19682 12264
rect 19618 12204 19622 12260
rect 19622 12204 19678 12260
rect 19678 12204 19682 12260
rect 19618 12200 19682 12204
rect 19698 12260 19762 12264
rect 19698 12204 19702 12260
rect 19702 12204 19758 12260
rect 19758 12204 19762 12260
rect 19698 12200 19762 12204
rect 19778 12260 19842 12264
rect 19778 12204 19782 12260
rect 19782 12204 19838 12260
rect 19838 12204 19842 12260
rect 19778 12200 19842 12204
rect 19858 12260 19922 12264
rect 19858 12204 19862 12260
rect 19862 12204 19918 12260
rect 19918 12204 19922 12260
rect 19858 12200 19922 12204
rect 5618 11716 5682 11720
rect 5618 11660 5622 11716
rect 5622 11660 5678 11716
rect 5678 11660 5682 11716
rect 5618 11656 5682 11660
rect 5698 11716 5762 11720
rect 5698 11660 5702 11716
rect 5702 11660 5758 11716
rect 5758 11660 5762 11716
rect 5698 11656 5762 11660
rect 5778 11716 5842 11720
rect 5778 11660 5782 11716
rect 5782 11660 5838 11716
rect 5838 11660 5842 11716
rect 5778 11656 5842 11660
rect 5858 11716 5922 11720
rect 5858 11660 5862 11716
rect 5862 11660 5918 11716
rect 5918 11660 5922 11716
rect 5858 11656 5922 11660
rect 14952 11716 15016 11720
rect 14952 11660 14956 11716
rect 14956 11660 15012 11716
rect 15012 11660 15016 11716
rect 14952 11656 15016 11660
rect 15032 11716 15096 11720
rect 15032 11660 15036 11716
rect 15036 11660 15092 11716
rect 15092 11660 15096 11716
rect 15032 11656 15096 11660
rect 15112 11716 15176 11720
rect 15112 11660 15116 11716
rect 15116 11660 15172 11716
rect 15172 11660 15176 11716
rect 15112 11656 15176 11660
rect 15192 11716 15256 11720
rect 15192 11660 15196 11716
rect 15196 11660 15252 11716
rect 15252 11660 15256 11716
rect 15192 11656 15256 11660
rect 24285 11716 24349 11720
rect 24285 11660 24289 11716
rect 24289 11660 24345 11716
rect 24345 11660 24349 11716
rect 24285 11656 24349 11660
rect 24365 11716 24429 11720
rect 24365 11660 24369 11716
rect 24369 11660 24425 11716
rect 24425 11660 24429 11716
rect 24365 11656 24429 11660
rect 24445 11716 24509 11720
rect 24445 11660 24449 11716
rect 24449 11660 24505 11716
rect 24505 11660 24509 11716
rect 24445 11656 24509 11660
rect 24525 11716 24589 11720
rect 24525 11660 24529 11716
rect 24529 11660 24585 11716
rect 24585 11660 24589 11716
rect 24525 11656 24589 11660
rect 10285 11172 10349 11176
rect 10285 11116 10289 11172
rect 10289 11116 10345 11172
rect 10345 11116 10349 11172
rect 10285 11112 10349 11116
rect 10365 11172 10429 11176
rect 10365 11116 10369 11172
rect 10369 11116 10425 11172
rect 10425 11116 10429 11172
rect 10365 11112 10429 11116
rect 10445 11172 10509 11176
rect 10445 11116 10449 11172
rect 10449 11116 10505 11172
rect 10505 11116 10509 11172
rect 10445 11112 10509 11116
rect 10525 11172 10589 11176
rect 10525 11116 10529 11172
rect 10529 11116 10585 11172
rect 10585 11116 10589 11172
rect 10525 11112 10589 11116
rect 19618 11172 19682 11176
rect 19618 11116 19622 11172
rect 19622 11116 19678 11172
rect 19678 11116 19682 11172
rect 19618 11112 19682 11116
rect 19698 11172 19762 11176
rect 19698 11116 19702 11172
rect 19702 11116 19758 11172
rect 19758 11116 19762 11172
rect 19698 11112 19762 11116
rect 19778 11172 19842 11176
rect 19778 11116 19782 11172
rect 19782 11116 19838 11172
rect 19838 11116 19842 11172
rect 19778 11112 19842 11116
rect 19858 11172 19922 11176
rect 19858 11116 19862 11172
rect 19862 11116 19918 11172
rect 19918 11116 19922 11172
rect 19858 11112 19922 11116
rect 5618 10628 5682 10632
rect 5618 10572 5622 10628
rect 5622 10572 5678 10628
rect 5678 10572 5682 10628
rect 5618 10568 5682 10572
rect 5698 10628 5762 10632
rect 5698 10572 5702 10628
rect 5702 10572 5758 10628
rect 5758 10572 5762 10628
rect 5698 10568 5762 10572
rect 5778 10628 5842 10632
rect 5778 10572 5782 10628
rect 5782 10572 5838 10628
rect 5838 10572 5842 10628
rect 5778 10568 5842 10572
rect 5858 10628 5922 10632
rect 5858 10572 5862 10628
rect 5862 10572 5918 10628
rect 5918 10572 5922 10628
rect 5858 10568 5922 10572
rect 14952 10628 15016 10632
rect 14952 10572 14956 10628
rect 14956 10572 15012 10628
rect 15012 10572 15016 10628
rect 14952 10568 15016 10572
rect 15032 10628 15096 10632
rect 15032 10572 15036 10628
rect 15036 10572 15092 10628
rect 15092 10572 15096 10628
rect 15032 10568 15096 10572
rect 15112 10628 15176 10632
rect 15112 10572 15116 10628
rect 15116 10572 15172 10628
rect 15172 10572 15176 10628
rect 15112 10568 15176 10572
rect 15192 10628 15256 10632
rect 15192 10572 15196 10628
rect 15196 10572 15252 10628
rect 15252 10572 15256 10628
rect 15192 10568 15256 10572
rect 24285 10628 24349 10632
rect 24285 10572 24289 10628
rect 24289 10572 24345 10628
rect 24345 10572 24349 10628
rect 24285 10568 24349 10572
rect 24365 10628 24429 10632
rect 24365 10572 24369 10628
rect 24369 10572 24425 10628
rect 24425 10572 24429 10628
rect 24365 10568 24429 10572
rect 24445 10628 24509 10632
rect 24445 10572 24449 10628
rect 24449 10572 24505 10628
rect 24505 10572 24509 10628
rect 24445 10568 24509 10572
rect 24525 10628 24589 10632
rect 24525 10572 24529 10628
rect 24529 10572 24585 10628
rect 24585 10572 24589 10628
rect 24525 10568 24589 10572
rect 10285 10084 10349 10088
rect 10285 10028 10289 10084
rect 10289 10028 10345 10084
rect 10345 10028 10349 10084
rect 10285 10024 10349 10028
rect 10365 10084 10429 10088
rect 10365 10028 10369 10084
rect 10369 10028 10425 10084
rect 10425 10028 10429 10084
rect 10365 10024 10429 10028
rect 10445 10084 10509 10088
rect 10445 10028 10449 10084
rect 10449 10028 10505 10084
rect 10505 10028 10509 10084
rect 10445 10024 10509 10028
rect 10525 10084 10589 10088
rect 10525 10028 10529 10084
rect 10529 10028 10585 10084
rect 10585 10028 10589 10084
rect 10525 10024 10589 10028
rect 19618 10084 19682 10088
rect 19618 10028 19622 10084
rect 19622 10028 19678 10084
rect 19678 10028 19682 10084
rect 19618 10024 19682 10028
rect 19698 10084 19762 10088
rect 19698 10028 19702 10084
rect 19702 10028 19758 10084
rect 19758 10028 19762 10084
rect 19698 10024 19762 10028
rect 19778 10084 19842 10088
rect 19778 10028 19782 10084
rect 19782 10028 19838 10084
rect 19838 10028 19842 10084
rect 19778 10024 19842 10028
rect 19858 10084 19922 10088
rect 19858 10028 19862 10084
rect 19862 10028 19918 10084
rect 19918 10028 19922 10084
rect 19858 10024 19922 10028
rect 5618 9540 5682 9544
rect 5618 9484 5622 9540
rect 5622 9484 5678 9540
rect 5678 9484 5682 9540
rect 5618 9480 5682 9484
rect 5698 9540 5762 9544
rect 5698 9484 5702 9540
rect 5702 9484 5758 9540
rect 5758 9484 5762 9540
rect 5698 9480 5762 9484
rect 5778 9540 5842 9544
rect 5778 9484 5782 9540
rect 5782 9484 5838 9540
rect 5838 9484 5842 9540
rect 5778 9480 5842 9484
rect 5858 9540 5922 9544
rect 5858 9484 5862 9540
rect 5862 9484 5918 9540
rect 5918 9484 5922 9540
rect 5858 9480 5922 9484
rect 14952 9540 15016 9544
rect 14952 9484 14956 9540
rect 14956 9484 15012 9540
rect 15012 9484 15016 9540
rect 14952 9480 15016 9484
rect 15032 9540 15096 9544
rect 15032 9484 15036 9540
rect 15036 9484 15092 9540
rect 15092 9484 15096 9540
rect 15032 9480 15096 9484
rect 15112 9540 15176 9544
rect 15112 9484 15116 9540
rect 15116 9484 15172 9540
rect 15172 9484 15176 9540
rect 15112 9480 15176 9484
rect 15192 9540 15256 9544
rect 15192 9484 15196 9540
rect 15196 9484 15252 9540
rect 15252 9484 15256 9540
rect 15192 9480 15256 9484
rect 24285 9540 24349 9544
rect 24285 9484 24289 9540
rect 24289 9484 24345 9540
rect 24345 9484 24349 9540
rect 24285 9480 24349 9484
rect 24365 9540 24429 9544
rect 24365 9484 24369 9540
rect 24369 9484 24425 9540
rect 24425 9484 24429 9540
rect 24365 9480 24429 9484
rect 24445 9540 24509 9544
rect 24445 9484 24449 9540
rect 24449 9484 24505 9540
rect 24505 9484 24509 9540
rect 24445 9480 24509 9484
rect 24525 9540 24589 9544
rect 24525 9484 24529 9540
rect 24529 9484 24585 9540
rect 24585 9484 24589 9540
rect 24525 9480 24589 9484
rect 10285 8996 10349 9000
rect 10285 8940 10289 8996
rect 10289 8940 10345 8996
rect 10345 8940 10349 8996
rect 10285 8936 10349 8940
rect 10365 8996 10429 9000
rect 10365 8940 10369 8996
rect 10369 8940 10425 8996
rect 10425 8940 10429 8996
rect 10365 8936 10429 8940
rect 10445 8996 10509 9000
rect 10445 8940 10449 8996
rect 10449 8940 10505 8996
rect 10505 8940 10509 8996
rect 10445 8936 10509 8940
rect 10525 8996 10589 9000
rect 10525 8940 10529 8996
rect 10529 8940 10585 8996
rect 10585 8940 10589 8996
rect 10525 8936 10589 8940
rect 19618 8996 19682 9000
rect 19618 8940 19622 8996
rect 19622 8940 19678 8996
rect 19678 8940 19682 8996
rect 19618 8936 19682 8940
rect 19698 8996 19762 9000
rect 19698 8940 19702 8996
rect 19702 8940 19758 8996
rect 19758 8940 19762 8996
rect 19698 8936 19762 8940
rect 19778 8996 19842 9000
rect 19778 8940 19782 8996
rect 19782 8940 19838 8996
rect 19838 8940 19842 8996
rect 19778 8936 19842 8940
rect 19858 8996 19922 9000
rect 19858 8940 19862 8996
rect 19862 8940 19918 8996
rect 19918 8940 19922 8996
rect 19858 8936 19922 8940
rect 5618 8452 5682 8456
rect 5618 8396 5622 8452
rect 5622 8396 5678 8452
rect 5678 8396 5682 8452
rect 5618 8392 5682 8396
rect 5698 8452 5762 8456
rect 5698 8396 5702 8452
rect 5702 8396 5758 8452
rect 5758 8396 5762 8452
rect 5698 8392 5762 8396
rect 5778 8452 5842 8456
rect 5778 8396 5782 8452
rect 5782 8396 5838 8452
rect 5838 8396 5842 8452
rect 5778 8392 5842 8396
rect 5858 8452 5922 8456
rect 5858 8396 5862 8452
rect 5862 8396 5918 8452
rect 5918 8396 5922 8452
rect 5858 8392 5922 8396
rect 14952 8452 15016 8456
rect 14952 8396 14956 8452
rect 14956 8396 15012 8452
rect 15012 8396 15016 8452
rect 14952 8392 15016 8396
rect 15032 8452 15096 8456
rect 15032 8396 15036 8452
rect 15036 8396 15092 8452
rect 15092 8396 15096 8452
rect 15032 8392 15096 8396
rect 15112 8452 15176 8456
rect 15112 8396 15116 8452
rect 15116 8396 15172 8452
rect 15172 8396 15176 8452
rect 15112 8392 15176 8396
rect 15192 8452 15256 8456
rect 15192 8396 15196 8452
rect 15196 8396 15252 8452
rect 15252 8396 15256 8452
rect 15192 8392 15256 8396
rect 24285 8452 24349 8456
rect 24285 8396 24289 8452
rect 24289 8396 24345 8452
rect 24345 8396 24349 8452
rect 24285 8392 24349 8396
rect 24365 8452 24429 8456
rect 24365 8396 24369 8452
rect 24369 8396 24425 8452
rect 24425 8396 24429 8452
rect 24365 8392 24429 8396
rect 24445 8452 24509 8456
rect 24445 8396 24449 8452
rect 24449 8396 24505 8452
rect 24505 8396 24509 8452
rect 24445 8392 24509 8396
rect 24525 8452 24589 8456
rect 24525 8396 24529 8452
rect 24529 8396 24585 8452
rect 24585 8396 24589 8452
rect 24525 8392 24589 8396
rect 10285 7908 10349 7912
rect 10285 7852 10289 7908
rect 10289 7852 10345 7908
rect 10345 7852 10349 7908
rect 10285 7848 10349 7852
rect 10365 7908 10429 7912
rect 10365 7852 10369 7908
rect 10369 7852 10425 7908
rect 10425 7852 10429 7908
rect 10365 7848 10429 7852
rect 10445 7908 10509 7912
rect 10445 7852 10449 7908
rect 10449 7852 10505 7908
rect 10505 7852 10509 7908
rect 10445 7848 10509 7852
rect 10525 7908 10589 7912
rect 10525 7852 10529 7908
rect 10529 7852 10585 7908
rect 10585 7852 10589 7908
rect 10525 7848 10589 7852
rect 19618 7908 19682 7912
rect 19618 7852 19622 7908
rect 19622 7852 19678 7908
rect 19678 7852 19682 7908
rect 19618 7848 19682 7852
rect 19698 7908 19762 7912
rect 19698 7852 19702 7908
rect 19702 7852 19758 7908
rect 19758 7852 19762 7908
rect 19698 7848 19762 7852
rect 19778 7908 19842 7912
rect 19778 7852 19782 7908
rect 19782 7852 19838 7908
rect 19838 7852 19842 7908
rect 19778 7848 19842 7852
rect 19858 7908 19922 7912
rect 19858 7852 19862 7908
rect 19862 7852 19918 7908
rect 19918 7852 19922 7908
rect 19858 7848 19922 7852
rect 5618 7364 5682 7368
rect 5618 7308 5622 7364
rect 5622 7308 5678 7364
rect 5678 7308 5682 7364
rect 5618 7304 5682 7308
rect 5698 7364 5762 7368
rect 5698 7308 5702 7364
rect 5702 7308 5758 7364
rect 5758 7308 5762 7364
rect 5698 7304 5762 7308
rect 5778 7364 5842 7368
rect 5778 7308 5782 7364
rect 5782 7308 5838 7364
rect 5838 7308 5842 7364
rect 5778 7304 5842 7308
rect 5858 7364 5922 7368
rect 5858 7308 5862 7364
rect 5862 7308 5918 7364
rect 5918 7308 5922 7364
rect 5858 7304 5922 7308
rect 14952 7364 15016 7368
rect 14952 7308 14956 7364
rect 14956 7308 15012 7364
rect 15012 7308 15016 7364
rect 14952 7304 15016 7308
rect 15032 7364 15096 7368
rect 15032 7308 15036 7364
rect 15036 7308 15092 7364
rect 15092 7308 15096 7364
rect 15032 7304 15096 7308
rect 15112 7364 15176 7368
rect 15112 7308 15116 7364
rect 15116 7308 15172 7364
rect 15172 7308 15176 7364
rect 15112 7304 15176 7308
rect 15192 7364 15256 7368
rect 15192 7308 15196 7364
rect 15196 7308 15252 7364
rect 15252 7308 15256 7364
rect 15192 7304 15256 7308
rect 24285 7364 24349 7368
rect 24285 7308 24289 7364
rect 24289 7308 24345 7364
rect 24345 7308 24349 7364
rect 24285 7304 24349 7308
rect 24365 7364 24429 7368
rect 24365 7308 24369 7364
rect 24369 7308 24425 7364
rect 24425 7308 24429 7364
rect 24365 7304 24429 7308
rect 24445 7364 24509 7368
rect 24445 7308 24449 7364
rect 24449 7308 24505 7364
rect 24505 7308 24509 7364
rect 24445 7304 24509 7308
rect 24525 7364 24589 7368
rect 24525 7308 24529 7364
rect 24529 7308 24585 7364
rect 24585 7308 24589 7364
rect 24525 7304 24589 7308
rect 10285 6820 10349 6824
rect 10285 6764 10289 6820
rect 10289 6764 10345 6820
rect 10345 6764 10349 6820
rect 10285 6760 10349 6764
rect 10365 6820 10429 6824
rect 10365 6764 10369 6820
rect 10369 6764 10425 6820
rect 10425 6764 10429 6820
rect 10365 6760 10429 6764
rect 10445 6820 10509 6824
rect 10445 6764 10449 6820
rect 10449 6764 10505 6820
rect 10505 6764 10509 6820
rect 10445 6760 10509 6764
rect 10525 6820 10589 6824
rect 10525 6764 10529 6820
rect 10529 6764 10585 6820
rect 10585 6764 10589 6820
rect 10525 6760 10589 6764
rect 19618 6820 19682 6824
rect 19618 6764 19622 6820
rect 19622 6764 19678 6820
rect 19678 6764 19682 6820
rect 19618 6760 19682 6764
rect 19698 6820 19762 6824
rect 19698 6764 19702 6820
rect 19702 6764 19758 6820
rect 19758 6764 19762 6820
rect 19698 6760 19762 6764
rect 19778 6820 19842 6824
rect 19778 6764 19782 6820
rect 19782 6764 19838 6820
rect 19838 6764 19842 6820
rect 19778 6760 19842 6764
rect 19858 6820 19922 6824
rect 19858 6764 19862 6820
rect 19862 6764 19918 6820
rect 19918 6764 19922 6820
rect 19858 6760 19922 6764
rect 5618 6276 5682 6280
rect 5618 6220 5622 6276
rect 5622 6220 5678 6276
rect 5678 6220 5682 6276
rect 5618 6216 5682 6220
rect 5698 6276 5762 6280
rect 5698 6220 5702 6276
rect 5702 6220 5758 6276
rect 5758 6220 5762 6276
rect 5698 6216 5762 6220
rect 5778 6276 5842 6280
rect 5778 6220 5782 6276
rect 5782 6220 5838 6276
rect 5838 6220 5842 6276
rect 5778 6216 5842 6220
rect 5858 6276 5922 6280
rect 5858 6220 5862 6276
rect 5862 6220 5918 6276
rect 5918 6220 5922 6276
rect 5858 6216 5922 6220
rect 14952 6276 15016 6280
rect 14952 6220 14956 6276
rect 14956 6220 15012 6276
rect 15012 6220 15016 6276
rect 14952 6216 15016 6220
rect 15032 6276 15096 6280
rect 15032 6220 15036 6276
rect 15036 6220 15092 6276
rect 15092 6220 15096 6276
rect 15032 6216 15096 6220
rect 15112 6276 15176 6280
rect 15112 6220 15116 6276
rect 15116 6220 15172 6276
rect 15172 6220 15176 6276
rect 15112 6216 15176 6220
rect 15192 6276 15256 6280
rect 15192 6220 15196 6276
rect 15196 6220 15252 6276
rect 15252 6220 15256 6276
rect 15192 6216 15256 6220
rect 24285 6276 24349 6280
rect 24285 6220 24289 6276
rect 24289 6220 24345 6276
rect 24345 6220 24349 6276
rect 24285 6216 24349 6220
rect 24365 6276 24429 6280
rect 24365 6220 24369 6276
rect 24369 6220 24425 6276
rect 24425 6220 24429 6276
rect 24365 6216 24429 6220
rect 24445 6276 24509 6280
rect 24445 6220 24449 6276
rect 24449 6220 24505 6276
rect 24505 6220 24509 6276
rect 24445 6216 24509 6220
rect 24525 6276 24589 6280
rect 24525 6220 24529 6276
rect 24529 6220 24585 6276
rect 24585 6220 24589 6276
rect 24525 6216 24589 6220
rect 10285 5732 10349 5736
rect 10285 5676 10289 5732
rect 10289 5676 10345 5732
rect 10345 5676 10349 5732
rect 10285 5672 10349 5676
rect 10365 5732 10429 5736
rect 10365 5676 10369 5732
rect 10369 5676 10425 5732
rect 10425 5676 10429 5732
rect 10365 5672 10429 5676
rect 10445 5732 10509 5736
rect 10445 5676 10449 5732
rect 10449 5676 10505 5732
rect 10505 5676 10509 5732
rect 10445 5672 10509 5676
rect 10525 5732 10589 5736
rect 10525 5676 10529 5732
rect 10529 5676 10585 5732
rect 10585 5676 10589 5732
rect 10525 5672 10589 5676
rect 19618 5732 19682 5736
rect 19618 5676 19622 5732
rect 19622 5676 19678 5732
rect 19678 5676 19682 5732
rect 19618 5672 19682 5676
rect 19698 5732 19762 5736
rect 19698 5676 19702 5732
rect 19702 5676 19758 5732
rect 19758 5676 19762 5732
rect 19698 5672 19762 5676
rect 19778 5732 19842 5736
rect 19778 5676 19782 5732
rect 19782 5676 19838 5732
rect 19838 5676 19842 5732
rect 19778 5672 19842 5676
rect 19858 5732 19922 5736
rect 19858 5676 19862 5732
rect 19862 5676 19918 5732
rect 19918 5676 19922 5732
rect 19858 5672 19922 5676
rect 5618 5188 5682 5192
rect 5618 5132 5622 5188
rect 5622 5132 5678 5188
rect 5678 5132 5682 5188
rect 5618 5128 5682 5132
rect 5698 5188 5762 5192
rect 5698 5132 5702 5188
rect 5702 5132 5758 5188
rect 5758 5132 5762 5188
rect 5698 5128 5762 5132
rect 5778 5188 5842 5192
rect 5778 5132 5782 5188
rect 5782 5132 5838 5188
rect 5838 5132 5842 5188
rect 5778 5128 5842 5132
rect 5858 5188 5922 5192
rect 5858 5132 5862 5188
rect 5862 5132 5918 5188
rect 5918 5132 5922 5188
rect 5858 5128 5922 5132
rect 14952 5188 15016 5192
rect 14952 5132 14956 5188
rect 14956 5132 15012 5188
rect 15012 5132 15016 5188
rect 14952 5128 15016 5132
rect 15032 5188 15096 5192
rect 15032 5132 15036 5188
rect 15036 5132 15092 5188
rect 15092 5132 15096 5188
rect 15032 5128 15096 5132
rect 15112 5188 15176 5192
rect 15112 5132 15116 5188
rect 15116 5132 15172 5188
rect 15172 5132 15176 5188
rect 15112 5128 15176 5132
rect 15192 5188 15256 5192
rect 15192 5132 15196 5188
rect 15196 5132 15252 5188
rect 15252 5132 15256 5188
rect 15192 5128 15256 5132
rect 24285 5188 24349 5192
rect 24285 5132 24289 5188
rect 24289 5132 24345 5188
rect 24345 5132 24349 5188
rect 24285 5128 24349 5132
rect 24365 5188 24429 5192
rect 24365 5132 24369 5188
rect 24369 5132 24425 5188
rect 24425 5132 24429 5188
rect 24365 5128 24429 5132
rect 24445 5188 24509 5192
rect 24445 5132 24449 5188
rect 24449 5132 24505 5188
rect 24505 5132 24509 5188
rect 24445 5128 24509 5132
rect 24525 5188 24589 5192
rect 24525 5132 24529 5188
rect 24529 5132 24585 5188
rect 24585 5132 24589 5188
rect 24525 5128 24589 5132
rect 10285 4644 10349 4648
rect 10285 4588 10289 4644
rect 10289 4588 10345 4644
rect 10345 4588 10349 4644
rect 10285 4584 10349 4588
rect 10365 4644 10429 4648
rect 10365 4588 10369 4644
rect 10369 4588 10425 4644
rect 10425 4588 10429 4644
rect 10365 4584 10429 4588
rect 10445 4644 10509 4648
rect 10445 4588 10449 4644
rect 10449 4588 10505 4644
rect 10505 4588 10509 4644
rect 10445 4584 10509 4588
rect 10525 4644 10589 4648
rect 10525 4588 10529 4644
rect 10529 4588 10585 4644
rect 10585 4588 10589 4644
rect 10525 4584 10589 4588
rect 19618 4644 19682 4648
rect 19618 4588 19622 4644
rect 19622 4588 19678 4644
rect 19678 4588 19682 4644
rect 19618 4584 19682 4588
rect 19698 4644 19762 4648
rect 19698 4588 19702 4644
rect 19702 4588 19758 4644
rect 19758 4588 19762 4644
rect 19698 4584 19762 4588
rect 19778 4644 19842 4648
rect 19778 4588 19782 4644
rect 19782 4588 19838 4644
rect 19838 4588 19842 4644
rect 19778 4584 19842 4588
rect 19858 4644 19922 4648
rect 19858 4588 19862 4644
rect 19862 4588 19918 4644
rect 19918 4588 19922 4644
rect 19858 4584 19922 4588
rect 5618 4100 5682 4104
rect 5618 4044 5622 4100
rect 5622 4044 5678 4100
rect 5678 4044 5682 4100
rect 5618 4040 5682 4044
rect 5698 4100 5762 4104
rect 5698 4044 5702 4100
rect 5702 4044 5758 4100
rect 5758 4044 5762 4100
rect 5698 4040 5762 4044
rect 5778 4100 5842 4104
rect 5778 4044 5782 4100
rect 5782 4044 5838 4100
rect 5838 4044 5842 4100
rect 5778 4040 5842 4044
rect 5858 4100 5922 4104
rect 5858 4044 5862 4100
rect 5862 4044 5918 4100
rect 5918 4044 5922 4100
rect 5858 4040 5922 4044
rect 14952 4100 15016 4104
rect 14952 4044 14956 4100
rect 14956 4044 15012 4100
rect 15012 4044 15016 4100
rect 14952 4040 15016 4044
rect 15032 4100 15096 4104
rect 15032 4044 15036 4100
rect 15036 4044 15092 4100
rect 15092 4044 15096 4100
rect 15032 4040 15096 4044
rect 15112 4100 15176 4104
rect 15112 4044 15116 4100
rect 15116 4044 15172 4100
rect 15172 4044 15176 4100
rect 15112 4040 15176 4044
rect 15192 4100 15256 4104
rect 15192 4044 15196 4100
rect 15196 4044 15252 4100
rect 15252 4044 15256 4100
rect 15192 4040 15256 4044
rect 24285 4100 24349 4104
rect 24285 4044 24289 4100
rect 24289 4044 24345 4100
rect 24345 4044 24349 4100
rect 24285 4040 24349 4044
rect 24365 4100 24429 4104
rect 24365 4044 24369 4100
rect 24369 4044 24425 4100
rect 24425 4044 24429 4100
rect 24365 4040 24429 4044
rect 24445 4100 24509 4104
rect 24445 4044 24449 4100
rect 24449 4044 24505 4100
rect 24505 4044 24509 4100
rect 24445 4040 24509 4044
rect 24525 4100 24589 4104
rect 24525 4044 24529 4100
rect 24529 4044 24585 4100
rect 24585 4044 24589 4100
rect 24525 4040 24589 4044
rect 10285 3556 10349 3560
rect 10285 3500 10289 3556
rect 10289 3500 10345 3556
rect 10345 3500 10349 3556
rect 10285 3496 10349 3500
rect 10365 3556 10429 3560
rect 10365 3500 10369 3556
rect 10369 3500 10425 3556
rect 10425 3500 10429 3556
rect 10365 3496 10429 3500
rect 10445 3556 10509 3560
rect 10445 3500 10449 3556
rect 10449 3500 10505 3556
rect 10505 3500 10509 3556
rect 10445 3496 10509 3500
rect 10525 3556 10589 3560
rect 10525 3500 10529 3556
rect 10529 3500 10585 3556
rect 10585 3500 10589 3556
rect 10525 3496 10589 3500
rect 19618 3556 19682 3560
rect 19618 3500 19622 3556
rect 19622 3500 19678 3556
rect 19678 3500 19682 3556
rect 19618 3496 19682 3500
rect 19698 3556 19762 3560
rect 19698 3500 19702 3556
rect 19702 3500 19758 3556
rect 19758 3500 19762 3556
rect 19698 3496 19762 3500
rect 19778 3556 19842 3560
rect 19778 3500 19782 3556
rect 19782 3500 19838 3556
rect 19838 3500 19842 3556
rect 19778 3496 19842 3500
rect 19858 3556 19922 3560
rect 19858 3500 19862 3556
rect 19862 3500 19918 3556
rect 19918 3500 19922 3556
rect 19858 3496 19922 3500
rect 5618 3012 5682 3016
rect 5618 2956 5622 3012
rect 5622 2956 5678 3012
rect 5678 2956 5682 3012
rect 5618 2952 5682 2956
rect 5698 3012 5762 3016
rect 5698 2956 5702 3012
rect 5702 2956 5758 3012
rect 5758 2956 5762 3012
rect 5698 2952 5762 2956
rect 5778 3012 5842 3016
rect 5778 2956 5782 3012
rect 5782 2956 5838 3012
rect 5838 2956 5842 3012
rect 5778 2952 5842 2956
rect 5858 3012 5922 3016
rect 5858 2956 5862 3012
rect 5862 2956 5918 3012
rect 5918 2956 5922 3012
rect 5858 2952 5922 2956
rect 14952 3012 15016 3016
rect 14952 2956 14956 3012
rect 14956 2956 15012 3012
rect 15012 2956 15016 3012
rect 14952 2952 15016 2956
rect 15032 3012 15096 3016
rect 15032 2956 15036 3012
rect 15036 2956 15092 3012
rect 15092 2956 15096 3012
rect 15032 2952 15096 2956
rect 15112 3012 15176 3016
rect 15112 2956 15116 3012
rect 15116 2956 15172 3012
rect 15172 2956 15176 3012
rect 15112 2952 15176 2956
rect 15192 3012 15256 3016
rect 15192 2956 15196 3012
rect 15196 2956 15252 3012
rect 15252 2956 15256 3012
rect 15192 2952 15256 2956
rect 24285 3012 24349 3016
rect 24285 2956 24289 3012
rect 24289 2956 24345 3012
rect 24345 2956 24349 3012
rect 24285 2952 24349 2956
rect 24365 3012 24429 3016
rect 24365 2956 24369 3012
rect 24369 2956 24425 3012
rect 24425 2956 24429 3012
rect 24365 2952 24429 2956
rect 24445 3012 24509 3016
rect 24445 2956 24449 3012
rect 24449 2956 24505 3012
rect 24505 2956 24509 3012
rect 24445 2952 24509 2956
rect 24525 3012 24589 3016
rect 24525 2956 24529 3012
rect 24529 2956 24585 3012
rect 24585 2956 24589 3012
rect 24525 2952 24589 2956
rect 10285 2468 10349 2472
rect 10285 2412 10289 2468
rect 10289 2412 10345 2468
rect 10345 2412 10349 2468
rect 10285 2408 10349 2412
rect 10365 2468 10429 2472
rect 10365 2412 10369 2468
rect 10369 2412 10425 2468
rect 10425 2412 10429 2468
rect 10365 2408 10429 2412
rect 10445 2468 10509 2472
rect 10445 2412 10449 2468
rect 10449 2412 10505 2468
rect 10505 2412 10509 2468
rect 10445 2408 10509 2412
rect 10525 2468 10589 2472
rect 10525 2412 10529 2468
rect 10529 2412 10585 2468
rect 10585 2412 10589 2468
rect 10525 2408 10589 2412
rect 19618 2468 19682 2472
rect 19618 2412 19622 2468
rect 19622 2412 19678 2468
rect 19678 2412 19682 2468
rect 19618 2408 19682 2412
rect 19698 2468 19762 2472
rect 19698 2412 19702 2468
rect 19702 2412 19758 2468
rect 19758 2412 19762 2468
rect 19698 2408 19762 2412
rect 19778 2468 19842 2472
rect 19778 2412 19782 2468
rect 19782 2412 19838 2468
rect 19838 2412 19842 2468
rect 19778 2408 19842 2412
rect 19858 2468 19922 2472
rect 19858 2412 19862 2468
rect 19862 2412 19918 2468
rect 19918 2412 19922 2468
rect 19858 2408 19922 2412
rect 5618 1924 5682 1928
rect 5618 1868 5622 1924
rect 5622 1868 5678 1924
rect 5678 1868 5682 1924
rect 5618 1864 5682 1868
rect 5698 1924 5762 1928
rect 5698 1868 5702 1924
rect 5702 1868 5758 1924
rect 5758 1868 5762 1924
rect 5698 1864 5762 1868
rect 5778 1924 5842 1928
rect 5778 1868 5782 1924
rect 5782 1868 5838 1924
rect 5838 1868 5842 1924
rect 5778 1864 5842 1868
rect 5858 1924 5922 1928
rect 5858 1868 5862 1924
rect 5862 1868 5918 1924
rect 5918 1868 5922 1924
rect 5858 1864 5922 1868
rect 14952 1924 15016 1928
rect 14952 1868 14956 1924
rect 14956 1868 15012 1924
rect 15012 1868 15016 1924
rect 14952 1864 15016 1868
rect 15032 1924 15096 1928
rect 15032 1868 15036 1924
rect 15036 1868 15092 1924
rect 15092 1868 15096 1924
rect 15032 1864 15096 1868
rect 15112 1924 15176 1928
rect 15112 1868 15116 1924
rect 15116 1868 15172 1924
rect 15172 1868 15176 1924
rect 15112 1864 15176 1868
rect 15192 1924 15256 1928
rect 15192 1868 15196 1924
rect 15196 1868 15252 1924
rect 15252 1868 15256 1924
rect 15192 1864 15256 1868
rect 24285 1924 24349 1928
rect 24285 1868 24289 1924
rect 24289 1868 24345 1924
rect 24345 1868 24349 1924
rect 24285 1864 24349 1868
rect 24365 1924 24429 1928
rect 24365 1868 24369 1924
rect 24369 1868 24425 1924
rect 24425 1868 24429 1924
rect 24365 1864 24429 1868
rect 24445 1924 24509 1928
rect 24445 1868 24449 1924
rect 24449 1868 24505 1924
rect 24505 1868 24509 1924
rect 24445 1864 24509 1868
rect 24525 1924 24589 1928
rect 24525 1868 24529 1924
rect 24529 1868 24585 1924
rect 24585 1868 24589 1924
rect 24525 1864 24589 1868
<< metal4 >>
rect 5610 24776 5931 25336
rect 5610 24712 5618 24776
rect 5682 24712 5698 24776
rect 5762 24712 5778 24776
rect 5842 24712 5858 24776
rect 5922 24712 5931 24776
rect 5610 23688 5931 24712
rect 5610 23624 5618 23688
rect 5682 23624 5698 23688
rect 5762 23624 5778 23688
rect 5842 23624 5858 23688
rect 5922 23624 5931 23688
rect 5610 22600 5931 23624
rect 5610 22536 5618 22600
rect 5682 22536 5698 22600
rect 5762 22536 5778 22600
rect 5842 22536 5858 22600
rect 5922 22536 5931 22600
rect 5610 21512 5931 22536
rect 5610 21448 5618 21512
rect 5682 21448 5698 21512
rect 5762 21448 5778 21512
rect 5842 21448 5858 21512
rect 5922 21448 5931 21512
rect 5610 20424 5931 21448
rect 5610 20360 5618 20424
rect 5682 20360 5698 20424
rect 5762 20360 5778 20424
rect 5842 20360 5858 20424
rect 5922 20360 5931 20424
rect 5610 19336 5931 20360
rect 5610 19272 5618 19336
rect 5682 19272 5698 19336
rect 5762 19272 5778 19336
rect 5842 19272 5858 19336
rect 5922 19272 5931 19336
rect 5610 18248 5931 19272
rect 5610 18184 5618 18248
rect 5682 18184 5698 18248
rect 5762 18184 5778 18248
rect 5842 18184 5858 18248
rect 5922 18184 5931 18248
rect 5610 17160 5931 18184
rect 5610 17096 5618 17160
rect 5682 17096 5698 17160
rect 5762 17096 5778 17160
rect 5842 17096 5858 17160
rect 5922 17096 5931 17160
rect 5610 16072 5931 17096
rect 5610 16008 5618 16072
rect 5682 16008 5698 16072
rect 5762 16008 5778 16072
rect 5842 16008 5858 16072
rect 5922 16008 5931 16072
rect 5610 14984 5931 16008
rect 5610 14920 5618 14984
rect 5682 14920 5698 14984
rect 5762 14920 5778 14984
rect 5842 14920 5858 14984
rect 5922 14920 5931 14984
rect 5610 13896 5931 14920
rect 5610 13832 5618 13896
rect 5682 13832 5698 13896
rect 5762 13832 5778 13896
rect 5842 13832 5858 13896
rect 5922 13832 5931 13896
rect 5610 12808 5931 13832
rect 5610 12744 5618 12808
rect 5682 12744 5698 12808
rect 5762 12744 5778 12808
rect 5842 12744 5858 12808
rect 5922 12744 5931 12808
rect 5610 11720 5931 12744
rect 5610 11656 5618 11720
rect 5682 11656 5698 11720
rect 5762 11656 5778 11720
rect 5842 11656 5858 11720
rect 5922 11656 5931 11720
rect 5610 10632 5931 11656
rect 5610 10568 5618 10632
rect 5682 10568 5698 10632
rect 5762 10568 5778 10632
rect 5842 10568 5858 10632
rect 5922 10568 5931 10632
rect 5610 9544 5931 10568
rect 5610 9480 5618 9544
rect 5682 9480 5698 9544
rect 5762 9480 5778 9544
rect 5842 9480 5858 9544
rect 5922 9480 5931 9544
rect 5610 8456 5931 9480
rect 5610 8392 5618 8456
rect 5682 8392 5698 8456
rect 5762 8392 5778 8456
rect 5842 8392 5858 8456
rect 5922 8392 5931 8456
rect 5610 7368 5931 8392
rect 5610 7304 5618 7368
rect 5682 7304 5698 7368
rect 5762 7304 5778 7368
rect 5842 7304 5858 7368
rect 5922 7304 5931 7368
rect 5610 6280 5931 7304
rect 5610 6216 5618 6280
rect 5682 6216 5698 6280
rect 5762 6216 5778 6280
rect 5842 6216 5858 6280
rect 5922 6216 5931 6280
rect 5610 5192 5931 6216
rect 5610 5128 5618 5192
rect 5682 5128 5698 5192
rect 5762 5128 5778 5192
rect 5842 5128 5858 5192
rect 5922 5128 5931 5192
rect 5610 4104 5931 5128
rect 5610 4040 5618 4104
rect 5682 4040 5698 4104
rect 5762 4040 5778 4104
rect 5842 4040 5858 4104
rect 5922 4040 5931 4104
rect 5610 3016 5931 4040
rect 5610 2952 5618 3016
rect 5682 2952 5698 3016
rect 5762 2952 5778 3016
rect 5842 2952 5858 3016
rect 5922 2952 5931 3016
rect 5610 1928 5931 2952
rect 5610 1864 5618 1928
rect 5682 1864 5698 1928
rect 5762 1864 5778 1928
rect 5842 1864 5858 1928
rect 5922 1864 5931 1928
rect 5610 1848 5931 1864
rect 10277 25320 10597 25336
rect 10277 25256 10285 25320
rect 10349 25256 10365 25320
rect 10429 25256 10445 25320
rect 10509 25256 10525 25320
rect 10589 25256 10597 25320
rect 10277 24232 10597 25256
rect 10277 24168 10285 24232
rect 10349 24168 10365 24232
rect 10429 24168 10445 24232
rect 10509 24168 10525 24232
rect 10589 24168 10597 24232
rect 10277 23144 10597 24168
rect 10277 23080 10285 23144
rect 10349 23080 10365 23144
rect 10429 23080 10445 23144
rect 10509 23080 10525 23144
rect 10589 23080 10597 23144
rect 10277 22056 10597 23080
rect 10277 21992 10285 22056
rect 10349 21992 10365 22056
rect 10429 21992 10445 22056
rect 10509 21992 10525 22056
rect 10589 21992 10597 22056
rect 10277 20968 10597 21992
rect 10277 20904 10285 20968
rect 10349 20904 10365 20968
rect 10429 20904 10445 20968
rect 10509 20904 10525 20968
rect 10589 20904 10597 20968
rect 10277 19880 10597 20904
rect 10277 19816 10285 19880
rect 10349 19816 10365 19880
rect 10429 19816 10445 19880
rect 10509 19816 10525 19880
rect 10589 19816 10597 19880
rect 10277 18792 10597 19816
rect 10277 18728 10285 18792
rect 10349 18728 10365 18792
rect 10429 18728 10445 18792
rect 10509 18728 10525 18792
rect 10589 18728 10597 18792
rect 10277 17704 10597 18728
rect 10277 17640 10285 17704
rect 10349 17640 10365 17704
rect 10429 17640 10445 17704
rect 10509 17640 10525 17704
rect 10589 17640 10597 17704
rect 10277 16616 10597 17640
rect 10277 16552 10285 16616
rect 10349 16552 10365 16616
rect 10429 16552 10445 16616
rect 10509 16552 10525 16616
rect 10589 16552 10597 16616
rect 10277 15528 10597 16552
rect 10277 15464 10285 15528
rect 10349 15464 10365 15528
rect 10429 15464 10445 15528
rect 10509 15464 10525 15528
rect 10589 15464 10597 15528
rect 10277 14440 10597 15464
rect 10277 14376 10285 14440
rect 10349 14376 10365 14440
rect 10429 14376 10445 14440
rect 10509 14376 10525 14440
rect 10589 14376 10597 14440
rect 10277 13352 10597 14376
rect 10277 13288 10285 13352
rect 10349 13288 10365 13352
rect 10429 13288 10445 13352
rect 10509 13288 10525 13352
rect 10589 13288 10597 13352
rect 10277 12264 10597 13288
rect 10277 12200 10285 12264
rect 10349 12200 10365 12264
rect 10429 12200 10445 12264
rect 10509 12200 10525 12264
rect 10589 12200 10597 12264
rect 10277 11176 10597 12200
rect 10277 11112 10285 11176
rect 10349 11112 10365 11176
rect 10429 11112 10445 11176
rect 10509 11112 10525 11176
rect 10589 11112 10597 11176
rect 10277 10088 10597 11112
rect 10277 10024 10285 10088
rect 10349 10024 10365 10088
rect 10429 10024 10445 10088
rect 10509 10024 10525 10088
rect 10589 10024 10597 10088
rect 10277 9000 10597 10024
rect 10277 8936 10285 9000
rect 10349 8936 10365 9000
rect 10429 8936 10445 9000
rect 10509 8936 10525 9000
rect 10589 8936 10597 9000
rect 10277 7912 10597 8936
rect 10277 7848 10285 7912
rect 10349 7848 10365 7912
rect 10429 7848 10445 7912
rect 10509 7848 10525 7912
rect 10589 7848 10597 7912
rect 10277 6824 10597 7848
rect 10277 6760 10285 6824
rect 10349 6760 10365 6824
rect 10429 6760 10445 6824
rect 10509 6760 10525 6824
rect 10589 6760 10597 6824
rect 10277 5736 10597 6760
rect 10277 5672 10285 5736
rect 10349 5672 10365 5736
rect 10429 5672 10445 5736
rect 10509 5672 10525 5736
rect 10589 5672 10597 5736
rect 10277 4648 10597 5672
rect 10277 4584 10285 4648
rect 10349 4584 10365 4648
rect 10429 4584 10445 4648
rect 10509 4584 10525 4648
rect 10589 4584 10597 4648
rect 10277 3560 10597 4584
rect 10277 3496 10285 3560
rect 10349 3496 10365 3560
rect 10429 3496 10445 3560
rect 10509 3496 10525 3560
rect 10589 3496 10597 3560
rect 10277 2472 10597 3496
rect 10277 2408 10285 2472
rect 10349 2408 10365 2472
rect 10429 2408 10445 2472
rect 10509 2408 10525 2472
rect 10589 2408 10597 2472
rect 10277 1848 10597 2408
rect 14944 24776 15264 25336
rect 14944 24712 14952 24776
rect 15016 24712 15032 24776
rect 15096 24712 15112 24776
rect 15176 24712 15192 24776
rect 15256 24712 15264 24776
rect 14944 23688 15264 24712
rect 14944 23624 14952 23688
rect 15016 23624 15032 23688
rect 15096 23624 15112 23688
rect 15176 23624 15192 23688
rect 15256 23624 15264 23688
rect 14944 22600 15264 23624
rect 14944 22536 14952 22600
rect 15016 22536 15032 22600
rect 15096 22536 15112 22600
rect 15176 22536 15192 22600
rect 15256 22536 15264 22600
rect 14944 21512 15264 22536
rect 14944 21448 14952 21512
rect 15016 21448 15032 21512
rect 15096 21448 15112 21512
rect 15176 21448 15192 21512
rect 15256 21448 15264 21512
rect 14944 20424 15264 21448
rect 14944 20360 14952 20424
rect 15016 20360 15032 20424
rect 15096 20360 15112 20424
rect 15176 20360 15192 20424
rect 15256 20360 15264 20424
rect 14944 19336 15264 20360
rect 14944 19272 14952 19336
rect 15016 19272 15032 19336
rect 15096 19272 15112 19336
rect 15176 19272 15192 19336
rect 15256 19272 15264 19336
rect 14944 18248 15264 19272
rect 14944 18184 14952 18248
rect 15016 18184 15032 18248
rect 15096 18184 15112 18248
rect 15176 18184 15192 18248
rect 15256 18184 15264 18248
rect 14944 17160 15264 18184
rect 14944 17096 14952 17160
rect 15016 17096 15032 17160
rect 15096 17096 15112 17160
rect 15176 17096 15192 17160
rect 15256 17096 15264 17160
rect 14944 16072 15264 17096
rect 14944 16008 14952 16072
rect 15016 16008 15032 16072
rect 15096 16008 15112 16072
rect 15176 16008 15192 16072
rect 15256 16008 15264 16072
rect 14944 14984 15264 16008
rect 14944 14920 14952 14984
rect 15016 14920 15032 14984
rect 15096 14920 15112 14984
rect 15176 14920 15192 14984
rect 15256 14920 15264 14984
rect 14944 13896 15264 14920
rect 14944 13832 14952 13896
rect 15016 13832 15032 13896
rect 15096 13832 15112 13896
rect 15176 13832 15192 13896
rect 15256 13832 15264 13896
rect 14944 12808 15264 13832
rect 14944 12744 14952 12808
rect 15016 12744 15032 12808
rect 15096 12744 15112 12808
rect 15176 12744 15192 12808
rect 15256 12744 15264 12808
rect 14944 11720 15264 12744
rect 14944 11656 14952 11720
rect 15016 11656 15032 11720
rect 15096 11656 15112 11720
rect 15176 11656 15192 11720
rect 15256 11656 15264 11720
rect 14944 10632 15264 11656
rect 14944 10568 14952 10632
rect 15016 10568 15032 10632
rect 15096 10568 15112 10632
rect 15176 10568 15192 10632
rect 15256 10568 15264 10632
rect 14944 9544 15264 10568
rect 14944 9480 14952 9544
rect 15016 9480 15032 9544
rect 15096 9480 15112 9544
rect 15176 9480 15192 9544
rect 15256 9480 15264 9544
rect 14944 8456 15264 9480
rect 14944 8392 14952 8456
rect 15016 8392 15032 8456
rect 15096 8392 15112 8456
rect 15176 8392 15192 8456
rect 15256 8392 15264 8456
rect 14944 7368 15264 8392
rect 14944 7304 14952 7368
rect 15016 7304 15032 7368
rect 15096 7304 15112 7368
rect 15176 7304 15192 7368
rect 15256 7304 15264 7368
rect 14944 6280 15264 7304
rect 14944 6216 14952 6280
rect 15016 6216 15032 6280
rect 15096 6216 15112 6280
rect 15176 6216 15192 6280
rect 15256 6216 15264 6280
rect 14944 5192 15264 6216
rect 14944 5128 14952 5192
rect 15016 5128 15032 5192
rect 15096 5128 15112 5192
rect 15176 5128 15192 5192
rect 15256 5128 15264 5192
rect 14944 4104 15264 5128
rect 14944 4040 14952 4104
rect 15016 4040 15032 4104
rect 15096 4040 15112 4104
rect 15176 4040 15192 4104
rect 15256 4040 15264 4104
rect 14944 3016 15264 4040
rect 14944 2952 14952 3016
rect 15016 2952 15032 3016
rect 15096 2952 15112 3016
rect 15176 2952 15192 3016
rect 15256 2952 15264 3016
rect 14944 1928 15264 2952
rect 14944 1864 14952 1928
rect 15016 1864 15032 1928
rect 15096 1864 15112 1928
rect 15176 1864 15192 1928
rect 15256 1864 15264 1928
rect 14944 1848 15264 1864
rect 19610 25320 19930 25336
rect 19610 25256 19618 25320
rect 19682 25256 19698 25320
rect 19762 25256 19778 25320
rect 19842 25256 19858 25320
rect 19922 25256 19930 25320
rect 19610 24232 19930 25256
rect 19610 24168 19618 24232
rect 19682 24168 19698 24232
rect 19762 24168 19778 24232
rect 19842 24168 19858 24232
rect 19922 24168 19930 24232
rect 19610 23144 19930 24168
rect 19610 23080 19618 23144
rect 19682 23080 19698 23144
rect 19762 23080 19778 23144
rect 19842 23080 19858 23144
rect 19922 23080 19930 23144
rect 19610 22056 19930 23080
rect 19610 21992 19618 22056
rect 19682 21992 19698 22056
rect 19762 21992 19778 22056
rect 19842 21992 19858 22056
rect 19922 21992 19930 22056
rect 19610 20968 19930 21992
rect 19610 20904 19618 20968
rect 19682 20904 19698 20968
rect 19762 20904 19778 20968
rect 19842 20904 19858 20968
rect 19922 20904 19930 20968
rect 19610 19880 19930 20904
rect 19610 19816 19618 19880
rect 19682 19816 19698 19880
rect 19762 19816 19778 19880
rect 19842 19816 19858 19880
rect 19922 19816 19930 19880
rect 19610 18792 19930 19816
rect 19610 18728 19618 18792
rect 19682 18728 19698 18792
rect 19762 18728 19778 18792
rect 19842 18728 19858 18792
rect 19922 18728 19930 18792
rect 19610 17704 19930 18728
rect 19610 17640 19618 17704
rect 19682 17640 19698 17704
rect 19762 17640 19778 17704
rect 19842 17640 19858 17704
rect 19922 17640 19930 17704
rect 19610 16616 19930 17640
rect 19610 16552 19618 16616
rect 19682 16552 19698 16616
rect 19762 16552 19778 16616
rect 19842 16552 19858 16616
rect 19922 16552 19930 16616
rect 19610 15528 19930 16552
rect 19610 15464 19618 15528
rect 19682 15464 19698 15528
rect 19762 15464 19778 15528
rect 19842 15464 19858 15528
rect 19922 15464 19930 15528
rect 19610 14440 19930 15464
rect 19610 14376 19618 14440
rect 19682 14376 19698 14440
rect 19762 14376 19778 14440
rect 19842 14376 19858 14440
rect 19922 14376 19930 14440
rect 19610 13352 19930 14376
rect 19610 13288 19618 13352
rect 19682 13288 19698 13352
rect 19762 13288 19778 13352
rect 19842 13288 19858 13352
rect 19922 13288 19930 13352
rect 19610 12264 19930 13288
rect 19610 12200 19618 12264
rect 19682 12200 19698 12264
rect 19762 12200 19778 12264
rect 19842 12200 19858 12264
rect 19922 12200 19930 12264
rect 19610 11176 19930 12200
rect 19610 11112 19618 11176
rect 19682 11112 19698 11176
rect 19762 11112 19778 11176
rect 19842 11112 19858 11176
rect 19922 11112 19930 11176
rect 19610 10088 19930 11112
rect 19610 10024 19618 10088
rect 19682 10024 19698 10088
rect 19762 10024 19778 10088
rect 19842 10024 19858 10088
rect 19922 10024 19930 10088
rect 19610 9000 19930 10024
rect 19610 8936 19618 9000
rect 19682 8936 19698 9000
rect 19762 8936 19778 9000
rect 19842 8936 19858 9000
rect 19922 8936 19930 9000
rect 19610 7912 19930 8936
rect 19610 7848 19618 7912
rect 19682 7848 19698 7912
rect 19762 7848 19778 7912
rect 19842 7848 19858 7912
rect 19922 7848 19930 7912
rect 19610 6824 19930 7848
rect 19610 6760 19618 6824
rect 19682 6760 19698 6824
rect 19762 6760 19778 6824
rect 19842 6760 19858 6824
rect 19922 6760 19930 6824
rect 19610 5736 19930 6760
rect 19610 5672 19618 5736
rect 19682 5672 19698 5736
rect 19762 5672 19778 5736
rect 19842 5672 19858 5736
rect 19922 5672 19930 5736
rect 19610 4648 19930 5672
rect 19610 4584 19618 4648
rect 19682 4584 19698 4648
rect 19762 4584 19778 4648
rect 19842 4584 19858 4648
rect 19922 4584 19930 4648
rect 19610 3560 19930 4584
rect 19610 3496 19618 3560
rect 19682 3496 19698 3560
rect 19762 3496 19778 3560
rect 19842 3496 19858 3560
rect 19922 3496 19930 3560
rect 19610 2472 19930 3496
rect 19610 2408 19618 2472
rect 19682 2408 19698 2472
rect 19762 2408 19778 2472
rect 19842 2408 19858 2472
rect 19922 2408 19930 2472
rect 19610 1848 19930 2408
rect 24277 24776 24597 25336
rect 24277 24712 24285 24776
rect 24349 24712 24365 24776
rect 24429 24712 24445 24776
rect 24509 24712 24525 24776
rect 24589 24712 24597 24776
rect 24277 23688 24597 24712
rect 24277 23624 24285 23688
rect 24349 23624 24365 23688
rect 24429 23624 24445 23688
rect 24509 23624 24525 23688
rect 24589 23624 24597 23688
rect 24277 22600 24597 23624
rect 24277 22536 24285 22600
rect 24349 22536 24365 22600
rect 24429 22536 24445 22600
rect 24509 22536 24525 22600
rect 24589 22536 24597 22600
rect 24277 21512 24597 22536
rect 24277 21448 24285 21512
rect 24349 21448 24365 21512
rect 24429 21448 24445 21512
rect 24509 21448 24525 21512
rect 24589 21448 24597 21512
rect 24277 20424 24597 21448
rect 24277 20360 24285 20424
rect 24349 20360 24365 20424
rect 24429 20360 24445 20424
rect 24509 20360 24525 20424
rect 24589 20360 24597 20424
rect 24277 19336 24597 20360
rect 24277 19272 24285 19336
rect 24349 19272 24365 19336
rect 24429 19272 24445 19336
rect 24509 19272 24525 19336
rect 24589 19272 24597 19336
rect 24277 18248 24597 19272
rect 24277 18184 24285 18248
rect 24349 18184 24365 18248
rect 24429 18184 24445 18248
rect 24509 18184 24525 18248
rect 24589 18184 24597 18248
rect 24277 17160 24597 18184
rect 24277 17096 24285 17160
rect 24349 17096 24365 17160
rect 24429 17096 24445 17160
rect 24509 17096 24525 17160
rect 24589 17096 24597 17160
rect 24277 16072 24597 17096
rect 24277 16008 24285 16072
rect 24349 16008 24365 16072
rect 24429 16008 24445 16072
rect 24509 16008 24525 16072
rect 24589 16008 24597 16072
rect 24277 14984 24597 16008
rect 24277 14920 24285 14984
rect 24349 14920 24365 14984
rect 24429 14920 24445 14984
rect 24509 14920 24525 14984
rect 24589 14920 24597 14984
rect 24277 13896 24597 14920
rect 24277 13832 24285 13896
rect 24349 13832 24365 13896
rect 24429 13832 24445 13896
rect 24509 13832 24525 13896
rect 24589 13832 24597 13896
rect 24277 12808 24597 13832
rect 24277 12744 24285 12808
rect 24349 12744 24365 12808
rect 24429 12744 24445 12808
rect 24509 12744 24525 12808
rect 24589 12744 24597 12808
rect 24277 11720 24597 12744
rect 24277 11656 24285 11720
rect 24349 11656 24365 11720
rect 24429 11656 24445 11720
rect 24509 11656 24525 11720
rect 24589 11656 24597 11720
rect 24277 10632 24597 11656
rect 24277 10568 24285 10632
rect 24349 10568 24365 10632
rect 24429 10568 24445 10632
rect 24509 10568 24525 10632
rect 24589 10568 24597 10632
rect 24277 9544 24597 10568
rect 24277 9480 24285 9544
rect 24349 9480 24365 9544
rect 24429 9480 24445 9544
rect 24509 9480 24525 9544
rect 24589 9480 24597 9544
rect 24277 8456 24597 9480
rect 24277 8392 24285 8456
rect 24349 8392 24365 8456
rect 24429 8392 24445 8456
rect 24509 8392 24525 8456
rect 24589 8392 24597 8456
rect 24277 7368 24597 8392
rect 24277 7304 24285 7368
rect 24349 7304 24365 7368
rect 24429 7304 24445 7368
rect 24509 7304 24525 7368
rect 24589 7304 24597 7368
rect 24277 6280 24597 7304
rect 24277 6216 24285 6280
rect 24349 6216 24365 6280
rect 24429 6216 24445 6280
rect 24509 6216 24525 6280
rect 24589 6216 24597 6280
rect 24277 5192 24597 6216
rect 24277 5128 24285 5192
rect 24349 5128 24365 5192
rect 24429 5128 24445 5192
rect 24509 5128 24525 5192
rect 24589 5128 24597 5192
rect 24277 4104 24597 5128
rect 24277 4040 24285 4104
rect 24349 4040 24365 4104
rect 24429 4040 24445 4104
rect 24509 4040 24525 4104
rect 24589 4040 24597 4104
rect 24277 3016 24597 4040
rect 24277 2952 24285 3016
rect 24349 2952 24365 3016
rect 24429 2952 24445 3016
rect 24509 2952 24525 3016
rect 24589 2952 24597 3016
rect 24277 1928 24597 2952
rect 24277 1864 24285 1928
rect 24349 1864 24365 1928
rect 24429 1864 24445 1928
rect 24509 1864 24525 1928
rect 24589 1864 24597 1928
rect 24277 1848 24597 1864
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 -1 2440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604681595
transform 1 0 1104 0 1 2440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1604681595
transform 1 0 2484 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1604681595
transform 1 0 1380 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1604681595
transform 1 0 2484 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 3956 0 1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3588 0 -1 2440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1604681595
transform 1 0 4048 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1604681595
transform 1 0 3588 0 1 2440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_32
timestamp 1604681595
transform 1 0 4048 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1604681595
transform 1 0 5152 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6256 0 -1 2440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_44
timestamp 1604681595
transform 1 0 5152 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_56
timestamp 1604681595
transform 1 0 6256 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 6808 0 -1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1604681595
transform 1 0 6900 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1604681595
transform 1 0 8004 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_68
timestamp 1604681595
transform 1 0 7360 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 9660 0 -1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 9568 0 1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1604681595
transform 1 0 9108 0 -1 2440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_80
timestamp 1604681595
transform 1 0 8464 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_93
timestamp 1604681595
transform 1 0 9660 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1604681595
transform 1 0 10856 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1604681595
transform 1 0 11960 0 -1 2440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_105
timestamp 1604681595
transform 1 0 10764 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_117
timestamp 1604681595
transform 1 0 11868 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 12512 0 -1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1604681595
transform 1 0 12604 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1604681595
transform 1 0 13708 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_129
timestamp 1604681595
transform 1 0 12972 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 15364 0 -1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 15180 0 1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1604681595
transform 1 0 14812 0 -1 2440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1604681595
transform 1 0 15456 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_141
timestamp 1604681595
transform 1 0 14076 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_154
timestamp 1604681595
transform 1 0 15272 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1604681595
transform 1 0 16560 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_166
timestamp 1604681595
transform 1 0 16376 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_178
timestamp 1604681595
transform 1 0 17480 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 18216 0 -1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1604681595
transform 1 0 17664 0 -1 2440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1604681595
transform 1 0 18308 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_190
timestamp 1604681595
transform 1 0 18584 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 21068 0 -1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 20792 0 1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1604681595
transform 1 0 19412 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1604681595
transform 1 0 20516 0 -1 2440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1604681595
transform 1 0 21160 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_202
timestamp 1604681595
transform 1 0 19688 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_215
timestamp 1604681595
transform 1 0 20884 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_230
timestamp 1604681595
transform 1 0 22264 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_227
timestamp 1604681595
transform 1 0 21988 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23920 0 -1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_242
timestamp 1604681595
transform 1 0 23368 0 -1 2440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_249
timestamp 1604681595
transform 1 0 24012 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_239
timestamp 1604681595
transform 1 0 23092 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_251
timestamp 1604681595
transform 1 0 24196 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 26864 0 -1 2440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 26864 0 1 2440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 26404 0 1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_261
timestamp 1604681595
transform 1 0 25116 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_273
timestamp 1604681595
transform 1 0 26220 0 -1 2440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_263
timestamp 1604681595
transform 1 0 25300 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_276 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 26496 0 1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1604681595
transform 1 0 2484 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_39
timestamp 1604681595
transform 1 0 4692 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5796 0 -1 3528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6532 0 -1 3528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 6716 0 -1 3528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_62
timestamp 1604681595
transform 1 0 6808 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_74
timestamp 1604681595
transform 1 0 7912 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_86
timestamp 1604681595
transform 1 0 9016 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_98
timestamp 1604681595
transform 1 0 10120 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_110
timestamp 1604681595
transform 1 0 11224 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 12328 0 -1 3528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_123
timestamp 1604681595
transform 1 0 12420 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_135
timestamp 1604681595
transform 1 0 13524 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_147
timestamp 1604681595
transform 1 0 14628 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_159
timestamp 1604681595
transform 1 0 15732 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_171
timestamp 1604681595
transform 1 0 16836 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 17940 0 -1 3528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_184
timestamp 1604681595
transform 1 0 18032 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_196
timestamp 1604681595
transform 1 0 19136 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_208
timestamp 1604681595
transform 1 0 20240 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_220
timestamp 1604681595
transform 1 0 21344 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_232
timestamp 1604681595
transform 1 0 22448 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 23552 0 -1 3528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_245
timestamp 1604681595
transform 1 0 23644 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_257
timestamp 1604681595
transform 1 0 24748 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 26864 0 -1 3528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_269
timestamp 1604681595
transform 1 0 25852 0 -1 3528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1604681595
transform 1 0 2484 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 3956 0 1 3528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 1604681595
transform 1 0 3588 0 1 3528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_32
timestamp 1604681595
transform 1 0 4048 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_44
timestamp 1604681595
transform 1 0 5152 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_56
timestamp 1604681595
transform 1 0 6256 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_68
timestamp 1604681595
transform 1 0 7360 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 9568 0 1 3528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_80
timestamp 1604681595
transform 1 0 8464 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_93
timestamp 1604681595
transform 1 0 9660 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_105
timestamp 1604681595
transform 1 0 10764 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_117
timestamp 1604681595
transform 1 0 11868 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_129
timestamp 1604681595
transform 1 0 12972 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 15180 0 1 3528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_141
timestamp 1604681595
transform 1 0 14076 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_154
timestamp 1604681595
transform 1 0 15272 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_166
timestamp 1604681595
transform 1 0 16376 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_178
timestamp 1604681595
transform 1 0 17480 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_190
timestamp 1604681595
transform 1 0 18584 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 20792 0 1 3528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_202
timestamp 1604681595
transform 1 0 19688 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_215
timestamp 1604681595
transform 1 0 20884 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_227
timestamp 1604681595
transform 1 0 21988 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _60_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 24564 0 1 3528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_239
timestamp 1604681595
transform 1 0 23092 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_251
timestamp 1604681595
transform 1 0 24196 0 1 3528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 26864 0 1 3528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 26404 0 1 3528
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 25116 0 1 3528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_259
timestamp 1604681595
transform 1 0 24932 0 1 3528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_263
timestamp 1604681595
transform 1 0 25300 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_276
timestamp 1604681595
transform 1 0 26496 0 1 3528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1604681595
transform 1 0 2484 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_39
timestamp 1604681595
transform 1 0 4692 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_51
timestamp 1604681595
transform 1 0 5796 0 -1 4616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_59
timestamp 1604681595
transform 1 0 6532 0 -1 4616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 6716 0 -1 4616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_62
timestamp 1604681595
transform 1 0 6808 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_74
timestamp 1604681595
transform 1 0 7912 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_86
timestamp 1604681595
transform 1 0 9016 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_98
timestamp 1604681595
transform 1 0 10120 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_110
timestamp 1604681595
transform 1 0 11224 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 12328 0 -1 4616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_123
timestamp 1604681595
transform 1 0 12420 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_135
timestamp 1604681595
transform 1 0 13524 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_147
timestamp 1604681595
transform 1 0 14628 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_159
timestamp 1604681595
transform 1 0 15732 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_171
timestamp 1604681595
transform 1 0 16836 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 17940 0 -1 4616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_184
timestamp 1604681595
transform 1 0 18032 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_196
timestamp 1604681595
transform 1 0 19136 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_208
timestamp 1604681595
transform 1 0 20240 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_220
timestamp 1604681595
transform 1 0 21344 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_232
timestamp 1604681595
transform 1 0 22448 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 23552 0 -1 4616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_245
timestamp 1604681595
transform 1 0 23644 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_257
timestamp 1604681595
transform 1 0 24748 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 26864 0 -1 4616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_269
timestamp 1604681595
transform 1 0 25852 0 -1 4616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1604681595
transform 1 0 2484 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 3956 0 1 4616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_27
timestamp 1604681595
transform 1 0 3588 0 1 4616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_32
timestamp 1604681595
transform 1 0 4048 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_44
timestamp 1604681595
transform 1 0 5152 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_56
timestamp 1604681595
transform 1 0 6256 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_68
timestamp 1604681595
transform 1 0 7360 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 9568 0 1 4616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_80
timestamp 1604681595
transform 1 0 8464 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1604681595
transform 1 0 9660 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_105
timestamp 1604681595
transform 1 0 10764 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_117
timestamp 1604681595
transform 1 0 11868 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_129
timestamp 1604681595
transform 1 0 12972 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1604681595
transform 1 0 15272 0 1 4616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 15180 0 1 4616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_141
timestamp 1604681595
transform 1 0 14076 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_158
timestamp 1604681595
transform 1 0 15640 0 1 4616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1604681595
transform 1 0 15824 0 1 4616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_162
timestamp 1604681595
transform 1 0 16008 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_174
timestamp 1604681595
transform 1 0 17112 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_186
timestamp 1604681595
transform 1 0 18216 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_198
timestamp 1604681595
transform 1 0 19320 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 20792 0 1 4616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_210
timestamp 1604681595
transform 1 0 20424 0 1 4616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_215
timestamp 1604681595
transform 1 0 20884 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_227
timestamp 1604681595
transform 1 0 21988 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_239
timestamp 1604681595
transform 1 0 23092 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_251
timestamp 1604681595
transform 1 0 24196 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 26864 0 1 4616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 26404 0 1 4616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_263
timestamp 1604681595
transform 1 0 25300 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_276
timestamp 1604681595
transform 1 0 26496 0 1 4616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1604681595
transform 1 0 2484 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1604681595
transform 1 0 2484 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 3956 0 1 5704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_27
timestamp 1604681595
transform 1 0 3588 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_39
timestamp 1604681595
transform 1 0 4692 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1604681595
transform 1 0 3588 0 1 5704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_32
timestamp 1604681595
transform 1 0 4048 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_51
timestamp 1604681595
transform 1 0 5796 0 -1 5704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_59
timestamp 1604681595
transform 1 0 6532 0 -1 5704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_44
timestamp 1604681595
transform 1 0 5152 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_56
timestamp 1604681595
transform 1 0 6256 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 6716 0 -1 5704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_62
timestamp 1604681595
transform 1 0 6808 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_74
timestamp 1604681595
transform 1 0 7912 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_68
timestamp 1604681595
transform 1 0 7360 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 9568 0 1 5704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_86
timestamp 1604681595
transform 1 0 9016 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_98
timestamp 1604681595
transform 1 0 10120 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_80
timestamp 1604681595
transform 1 0 8464 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1604681595
transform 1 0 9660 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_110
timestamp 1604681595
transform 1 0 11224 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_105
timestamp 1604681595
transform 1 0 10764 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_117
timestamp 1604681595
transform 1 0 11868 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 12328 0 -1 5704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_123
timestamp 1604681595
transform 1 0 12420 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_135
timestamp 1604681595
transform 1 0 13524 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_129
timestamp 1604681595
transform 1 0 12972 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 15180 0 1 5704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_147
timestamp 1604681595
transform 1 0 14628 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_141
timestamp 1604681595
transform 1 0 14076 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_154
timestamp 1604681595
transform 1 0 15272 0 1 5704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1604681595
transform 1 0 16284 0 1 5704
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1604681595
transform 1 0 16836 0 1 5704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_159
timestamp 1604681595
transform 1 0 15732 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_171
timestamp 1604681595
transform 1 0 16836 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_162
timestamp 1604681595
transform 1 0 16008 0 1 5704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1604681595
transform 1 0 16652 0 1 5704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_173
timestamp 1604681595
transform 1 0 17020 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 17940 0 -1 5704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_184
timestamp 1604681595
transform 1 0 18032 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_196
timestamp 1604681595
transform 1 0 19136 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_185
timestamp 1604681595
transform 1 0 18124 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_197
timestamp 1604681595
transform 1 0 19228 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 20792 0 1 5704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_208
timestamp 1604681595
transform 1 0 20240 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_209
timestamp 1604681595
transform 1 0 20332 0 1 5704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_213
timestamp 1604681595
transform 1 0 20700 0 1 5704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_215
timestamp 1604681595
transform 1 0 20884 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_220
timestamp 1604681595
transform 1 0 21344 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_232
timestamp 1604681595
transform 1 0 22448 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_227
timestamp 1604681595
transform 1 0 21988 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 23552 0 -1 5704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_245
timestamp 1604681595
transform 1 0 23644 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_257
timestamp 1604681595
transform 1 0 24748 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_239
timestamp 1604681595
transform 1 0 23092 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_251
timestamp 1604681595
transform 1 0 24196 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 26864 0 -1 5704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 26864 0 1 5704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 26404 0 1 5704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_269
timestamp 1604681595
transform 1 0 25852 0 -1 5704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_263
timestamp 1604681595
transform 1 0 25300 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_276
timestamp 1604681595
transform 1 0 26496 0 1 5704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 6792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604681595
transform 1 0 2484 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_27
timestamp 1604681595
transform 1 0 3588 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_39
timestamp 1604681595
transform 1 0 4692 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_51
timestamp 1604681595
transform 1 0 5796 0 -1 6792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_59
timestamp 1604681595
transform 1 0 6532 0 -1 6792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 6716 0 -1 6792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_62
timestamp 1604681595
transform 1 0 6808 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_74
timestamp 1604681595
transform 1 0 7912 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_86
timestamp 1604681595
transform 1 0 9016 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_98
timestamp 1604681595
transform 1 0 10120 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_110
timestamp 1604681595
transform 1 0 11224 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 12328 0 -1 6792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_123
timestamp 1604681595
transform 1 0 12420 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_135
timestamp 1604681595
transform 1 0 13524 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_147
timestamp 1604681595
transform 1 0 14628 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_159
timestamp 1604681595
transform 1 0 15732 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_171
timestamp 1604681595
transform 1 0 16836 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 17940 0 -1 6792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_184
timestamp 1604681595
transform 1 0 18032 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_196
timestamp 1604681595
transform 1 0 19136 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_208
timestamp 1604681595
transform 1 0 20240 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_220
timestamp 1604681595
transform 1 0 21344 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_232
timestamp 1604681595
transform 1 0 22448 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 23552 0 -1 6792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_245
timestamp 1604681595
transform 1 0 23644 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_257
timestamp 1604681595
transform 1 0 24748 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 26864 0 -1 6792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_269
timestamp 1604681595
transform 1 0 25852 0 -1 6792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 6792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1604681595
transform 1 0 2484 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 3956 0 1 6792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_27
timestamp 1604681595
transform 1 0 3588 0 1 6792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_32
timestamp 1604681595
transform 1 0 4048 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_44
timestamp 1604681595
transform 1 0 5152 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_56
timestamp 1604681595
transform 1 0 6256 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_68
timestamp 1604681595
transform 1 0 7360 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 9568 0 1 6792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_80
timestamp 1604681595
transform 1 0 8464 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1604681595
transform 1 0 9660 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_105
timestamp 1604681595
transform 1 0 10764 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_117
timestamp 1604681595
transform 1 0 11868 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_129
timestamp 1604681595
transform 1 0 12972 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 15180 0 1 6792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_141
timestamp 1604681595
transform 1 0 14076 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_154
timestamp 1604681595
transform 1 0 15272 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_166
timestamp 1604681595
transform 1 0 16376 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_178
timestamp 1604681595
transform 1 0 17480 0 1 6792
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1604681595
transform 1 0 17572 0 1 6792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1604681595
transform 1 0 18124 0 1 6792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_183
timestamp 1604681595
transform 1 0 17940 0 1 6792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_187
timestamp 1604681595
transform 1 0 18308 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 20792 0 1 6792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_199
timestamp 1604681595
transform 1 0 19412 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_211
timestamp 1604681595
transform 1 0 20516 0 1 6792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_215
timestamp 1604681595
transform 1 0 20884 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_227
timestamp 1604681595
transform 1 0 21988 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1604681595
transform 1 0 24564 0 1 6792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_239
timestamp 1604681595
transform 1 0 23092 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_251
timestamp 1604681595
transform 1 0 24196 0 1 6792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_257
timestamp 1604681595
transform 1 0 24748 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 26864 0 1 6792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 26404 0 1 6792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_269
timestamp 1604681595
transform 1 0 25852 0 1 6792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_276
timestamp 1604681595
transform 1 0 26496 0 1 6792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 7880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1604681595
transform 1 0 2484 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_27
timestamp 1604681595
transform 1 0 3588 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_39
timestamp 1604681595
transform 1 0 4692 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_51
timestamp 1604681595
transform 1 0 5796 0 -1 7880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_59
timestamp 1604681595
transform 1 0 6532 0 -1 7880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 6716 0 -1 7880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_62
timestamp 1604681595
transform 1 0 6808 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_74
timestamp 1604681595
transform 1 0 7912 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_86
timestamp 1604681595
transform 1 0 9016 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_98
timestamp 1604681595
transform 1 0 10120 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_110
timestamp 1604681595
transform 1 0 11224 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 12328 0 -1 7880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_123
timestamp 1604681595
transform 1 0 12420 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_135
timestamp 1604681595
transform 1 0 13524 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_147
timestamp 1604681595
transform 1 0 14628 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_159
timestamp 1604681595
transform 1 0 15732 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_171
timestamp 1604681595
transform 1 0 16836 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 17940 0 -1 7880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_184
timestamp 1604681595
transform 1 0 18032 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_196
timestamp 1604681595
transform 1 0 19136 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_208
timestamp 1604681595
transform 1 0 20240 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_220
timestamp 1604681595
transform 1 0 21344 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_232
timestamp 1604681595
transform 1 0 22448 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1604681595
transform 1 0 24564 0 -1 7880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 23552 0 -1 7880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_245
timestamp 1604681595
transform 1 0 23644 0 -1 7880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1604681595
transform 1 0 24380 0 -1 7880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 26864 0 -1 7880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_259
timestamp 1604681595
transform 1 0 24932 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_271
timestamp 1604681595
transform 1 0 26036 0 -1 7880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 7880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1604681595
transform 1 0 2484 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 3956 0 1 7880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_27
timestamp 1604681595
transform 1 0 3588 0 1 7880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_32
timestamp 1604681595
transform 1 0 4048 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_44
timestamp 1604681595
transform 1 0 5152 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_56
timestamp 1604681595
transform 1 0 6256 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_68
timestamp 1604681595
transform 1 0 7360 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 9568 0 1 7880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_80
timestamp 1604681595
transform 1 0 8464 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1604681595
transform 1 0 9660 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_105
timestamp 1604681595
transform 1 0 10764 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_117
timestamp 1604681595
transform 1 0 11868 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_129
timestamp 1604681595
transform 1 0 12972 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 15180 0 1 7880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_141
timestamp 1604681595
transform 1 0 14076 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_154
timestamp 1604681595
transform 1 0 15272 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_166
timestamp 1604681595
transform 1 0 16376 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_178
timestamp 1604681595
transform 1 0 17480 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_190
timestamp 1604681595
transform 1 0 18584 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 20792 0 1 7880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_202
timestamp 1604681595
transform 1 0 19688 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_215
timestamp 1604681595
transform 1 0 20884 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_227
timestamp 1604681595
transform 1 0 21988 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1604681595
transform 1 0 24564 0 1 7880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_239
timestamp 1604681595
transform 1 0 23092 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_251
timestamp 1604681595
transform 1 0 24196 0 1 7880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_257
timestamp 1604681595
transform 1 0 24748 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 26864 0 1 7880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 26404 0 1 7880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_269
timestamp 1604681595
transform 1 0 25852 0 1 7880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_276
timestamp 1604681595
transform 1 0 26496 0 1 7880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 8968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1604681595
transform 1 0 2484 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_27
timestamp 1604681595
transform 1 0 3588 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_39
timestamp 1604681595
transform 1 0 4692 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_51
timestamp 1604681595
transform 1 0 5796 0 -1 8968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_59
timestamp 1604681595
transform 1 0 6532 0 -1 8968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 6716 0 -1 8968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_62
timestamp 1604681595
transform 1 0 6808 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_74
timestamp 1604681595
transform 1 0 7912 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_86
timestamp 1604681595
transform 1 0 9016 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_98
timestamp 1604681595
transform 1 0 10120 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_110
timestamp 1604681595
transform 1 0 11224 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 12328 0 -1 8968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_123
timestamp 1604681595
transform 1 0 12420 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_135
timestamp 1604681595
transform 1 0 13524 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_147
timestamp 1604681595
transform 1 0 14628 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_159
timestamp 1604681595
transform 1 0 15732 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_171
timestamp 1604681595
transform 1 0 16836 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 17940 0 -1 8968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_184
timestamp 1604681595
transform 1 0 18032 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_196
timestamp 1604681595
transform 1 0 19136 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_208
timestamp 1604681595
transform 1 0 20240 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_220
timestamp 1604681595
transform 1 0 21344 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_232
timestamp 1604681595
transform 1 0 22448 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1604681595
transform 1 0 24564 0 -1 8968
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 23552 0 -1 8968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_245
timestamp 1604681595
transform 1 0 23644 0 -1 8968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1604681595
transform 1 0 24380 0 -1 8968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 26864 0 -1 8968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_259
timestamp 1604681595
transform 1 0 24932 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_271
timestamp 1604681595
transform 1 0 26036 0 -1 8968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 8968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1604681595
transform 1 0 2484 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1604681595
transform 1 0 2484 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 3956 0 1 8968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_27
timestamp 1604681595
transform 1 0 3588 0 1 8968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_32
timestamp 1604681595
transform 1 0 4048 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_27
timestamp 1604681595
transform 1 0 3588 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_39
timestamp 1604681595
transform 1 0 4692 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_44
timestamp 1604681595
transform 1 0 5152 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_56
timestamp 1604681595
transform 1 0 6256 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_51
timestamp 1604681595
transform 1 0 5796 0 -1 10056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_59
timestamp 1604681595
transform 1 0 6532 0 -1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 6716 0 -1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_68
timestamp 1604681595
transform 1 0 7360 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_62
timestamp 1604681595
transform 1 0 6808 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_74
timestamp 1604681595
transform 1 0 7912 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 9568 0 1 8968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_80
timestamp 1604681595
transform 1 0 8464 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1604681595
transform 1 0 9660 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_86
timestamp 1604681595
transform 1 0 9016 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_98
timestamp 1604681595
transform 1 0 10120 0 -1 10056
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 10948 0 -1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_105
timestamp 1604681595
transform 1 0 10764 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_117
timestamp 1604681595
transform 1 0 11868 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_106
timestamp 1604681595
transform 1 0 10856 0 -1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1604681595
transform 1 0 11132 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 12328 0 -1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 -1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_129
timestamp 1604681595
transform 1 0 12972 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_121
timestamp 1604681595
transform 1 0 12236 0 -1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_123
timestamp 1604681595
transform 1 0 12420 0 -1 10056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_131
timestamp 1604681595
transform 1 0 13156 0 -1 10056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_136
timestamp 1604681595
transform 1 0 13616 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 15180 0 1 8968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_141
timestamp 1604681595
transform 1 0 14076 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_154
timestamp 1604681595
transform 1 0 15272 0 1 8968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_148
timestamp 1604681595
transform 1 0 14720 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_160
timestamp 1604681595
transform 1 0 15824 0 -1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_167
timestamp 1604681595
transform 1 0 16468 0 1 8968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_163
timestamp 1604681595
transform 1 0 16100 0 1 8968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_160
timestamp 1604681595
transform 1 0 15824 0 1 8968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 16284 0 1 8968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 15916 0 1 8968
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 15916 0 -1 10056
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16652 0 1 8968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_170
timestamp 1604681595
transform 1 0 16744 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_171
timestamp 1604681595
transform 1 0 16836 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_184
timestamp 1604681595
transform 1 0 18032 0 -1 10056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_182
timestamp 1604681595
transform 1 0 17848 0 -1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_183
timestamp 1604681595
transform 1 0 17940 0 1 8968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 17940 0 -1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_198
timestamp 1604681595
transform 1 0 19320 0 1 8968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_194
timestamp 1604681595
transform 1 0 18952 0 1 8968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_191
timestamp 1604681595
transform 1 0 18676 0 1 8968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19136 0 1 8968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18768 0 1 8968
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18768 0 -1 10056
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 20792 0 1 8968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19504 0 1 8968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_202
timestamp 1604681595
transform 1 0 19688 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_215
timestamp 1604681595
transform 1 0 20884 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_201
timestamp 1604681595
transform 1 0 19596 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_213
timestamp 1604681595
transform 1 0 20700 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_227
timestamp 1604681595
transform 1 0 21988 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_225
timestamp 1604681595
transform 1 0 21804 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_237
timestamp 1604681595
transform 1 0 22908 0 -1 10056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604681595
transform 1 0 24564 0 -1 10056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604681595
transform 1 0 24564 0 1 8968
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 23552 0 -1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1604681595
transform 1 0 24380 0 1 8968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_239
timestamp 1604681595
transform 1 0 23092 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_251
timestamp 1604681595
transform 1 0 24196 0 1 8968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_243
timestamp 1604681595
transform 1 0 23460 0 -1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_245
timestamp 1604681595
transform 1 0 23644 0 -1 10056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1604681595
transform 1 0 24380 0 -1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 26864 0 1 8968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 26864 0 -1 10056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 26404 0 1 8968
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1604681595
transform 1 0 25116 0 1 8968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_259
timestamp 1604681595
transform 1 0 24932 0 1 8968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_263
timestamp 1604681595
transform 1 0 25300 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_276
timestamp 1604681595
transform 1 0 26496 0 1 8968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_259
timestamp 1604681595
transform 1 0 24932 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_271
timestamp 1604681595
transform 1 0 26036 0 -1 10056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1604681595
transform 1 0 2484 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 3956 0 1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_27
timestamp 1604681595
transform 1 0 3588 0 1 10056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_32
timestamp 1604681595
transform 1 0 4048 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_44
timestamp 1604681595
transform 1 0 5152 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_56
timestamp 1604681595
transform 1 0 6256 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_68
timestamp 1604681595
transform 1 0 7360 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 9568 0 1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_80
timestamp 1604681595
transform 1 0 8464 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1604681595
transform 1 0 9660 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 10948 0 1 10056
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 10764 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13432 0 1 10056
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13248 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12880 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_126
timestamp 1604681595
transform 1 0 12696 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_130
timestamp 1604681595
transform 1 0 13064 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 15180 0 1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14444 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 14812 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_143
timestamp 1604681595
transform 1 0 14260 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_147
timestamp 1604681595
transform 1 0 14628 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_151
timestamp 1604681595
transform 1 0 14996 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_154
timestamp 1604681595
transform 1 0 15272 0 1 10056
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 16836 0 1 10056
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 16652 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 16284 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_162
timestamp 1604681595
transform 1 0 16008 0 1 10056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_167
timestamp 1604681595
transform 1 0 16468 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 18768 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 19136 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_190
timestamp 1604681595
transform 1 0 18584 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_194
timestamp 1604681595
transform 1 0 18952 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_198
timestamp 1604681595
transform 1 0 19320 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 20792 0 1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 21068 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_210
timestamp 1604681595
transform 1 0 20424 0 1 10056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_215
timestamp 1604681595
transform 1 0 20884 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 21436 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_219
timestamp 1604681595
transform 1 0 21252 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_223
timestamp 1604681595
transform 1 0 21620 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_235
timestamp 1604681595
transform 1 0 22724 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604681595
transform 1 0 24564 0 1 10056
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1604681595
transform 1 0 24380 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_247
timestamp 1604681595
transform 1 0 23828 0 1 10056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 26864 0 1 10056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 26404 0 1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1604681595
transform 1 0 25116 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_259
timestamp 1604681595
transform 1 0 24932 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_263
timestamp 1604681595
transform 1 0 25300 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_276
timestamp 1604681595
transform 1 0 26496 0 1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1604681595
transform 1 0 2484 0 -1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_27
timestamp 1604681595
transform 1 0 3588 0 -1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_39
timestamp 1604681595
transform 1 0 4692 0 -1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_51
timestamp 1604681595
transform 1 0 5796 0 -1 11144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_59
timestamp 1604681595
transform 1 0 6532 0 -1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 6716 0 -1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_62
timestamp 1604681595
transform 1 0 6808 0 -1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_74
timestamp 1604681595
transform 1 0 7912 0 -1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_86
timestamp 1604681595
transform 1 0 9016 0 -1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_98
timestamp 1604681595
transform 1 0 10120 0 -1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_110
timestamp 1604681595
transform 1 0 11224 0 -1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _23_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12696 0 -1 11144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 12328 0 -1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13156 0 -1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13524 0 -1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_123
timestamp 1604681595
transform 1 0 12420 0 -1 11144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_129
timestamp 1604681595
transform 1 0 12972 0 -1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_133
timestamp 1604681595
transform 1 0 13340 0 -1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_137
timestamp 1604681595
transform 1 0 13708 0 -1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 14076 0 -1 11144
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13892 0 -1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1604681595
transform 1 0 16560 0 -1 11144
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16008 0 -1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16376 0 -1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_160
timestamp 1604681595
transform 1 0 15824 0 -1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_164
timestamp 1604681595
transform 1 0 16192 0 -1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_171
timestamp 1604681595
transform 1 0 16836 0 -1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 18400 0 -1 11144
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 17940 0 -1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_184
timestamp 1604681595
transform 1 0 18032 0 -1 11144
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 20884 0 -1 11144
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20700 0 -1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_207
timestamp 1604681595
transform 1 0 20148 0 -1 11144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_234
timestamp 1604681595
transform 1 0 22632 0 -1 11144
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604681595
transform 1 0 24564 0 -1 11144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 23552 0 -1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_242
timestamp 1604681595
transform 1 0 23368 0 -1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_245
timestamp 1604681595
transform 1 0 23644 0 -1 11144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1604681595
transform 1 0 24380 0 -1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 26864 0 -1 11144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_259
timestamp 1604681595
transform 1 0 24932 0 -1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_271
timestamp 1604681595
transform 1 0 26036 0 -1 11144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1604681595
transform 1 0 2484 0 1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 3956 0 1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_27
timestamp 1604681595
transform 1 0 3588 0 1 11144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_32
timestamp 1604681595
transform 1 0 4048 0 1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_44
timestamp 1604681595
transform 1 0 5152 0 1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_56
timestamp 1604681595
transform 1 0 6256 0 1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_68
timestamp 1604681595
transform 1 0 7360 0 1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 9568 0 1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_80
timestamp 1604681595
transform 1 0 8464 0 1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1604681595
transform 1 0 9660 0 1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_105
timestamp 1604681595
transform 1 0 10764 0 1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_117
timestamp 1604681595
transform 1 0 11868 0 1 11144
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 12604 0 1 11144
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 12420 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15548 0 1 11144
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 15180 0 1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14996 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 14628 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_144
timestamp 1604681595
transform 1 0 14352 0 1 11144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_149
timestamp 1604681595
transform 1 0 14812 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_154
timestamp 1604681595
transform 1 0 15272 0 1 11144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_176
timestamp 1604681595
transform 1 0 17296 0 1 11144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18308 0 1 11144
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 18124 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17756 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_180
timestamp 1604681595
transform 1 0 17664 0 1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_183
timestamp 1604681595
transform 1 0 17940 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_196
timestamp 1604681595
transform 1 0 19136 0 1 11144
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20884 0 1 11144
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 20792 0 1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20240 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 19872 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_206
timestamp 1604681595
transform 1 0 20056 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_210
timestamp 1604681595
transform 1 0 20424 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21896 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 22264 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_224
timestamp 1604681595
transform 1 0 21712 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_228
timestamp 1604681595
transform 1 0 22080 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_232
timestamp 1604681595
transform 1 0 22448 0 1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1604681595
transform 1 0 24380 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_244
timestamp 1604681595
transform 1 0 23552 0 1 11144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_252
timestamp 1604681595
transform 1 0 24288 0 1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_255
timestamp 1604681595
transform 1 0 24564 0 1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 26864 0 1 11144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 26404 0 1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_267
timestamp 1604681595
transform 1 0 25668 0 1 11144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_276
timestamp 1604681595
transform 1 0 26496 0 1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1604681595
transform 1 0 2484 0 -1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_27
timestamp 1604681595
transform 1 0 3588 0 -1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_39
timestamp 1604681595
transform 1 0 4692 0 -1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_51
timestamp 1604681595
transform 1 0 5796 0 -1 12232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_59
timestamp 1604681595
transform 1 0 6532 0 -1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 6716 0 -1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_62
timestamp 1604681595
transform 1 0 6808 0 -1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_74
timestamp 1604681595
transform 1 0 7912 0 -1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_86
timestamp 1604681595
transform 1 0 9016 0 -1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_98
timestamp 1604681595
transform 1 0 10120 0 -1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_110
timestamp 1604681595
transform 1 0 11224 0 -1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13156 0 -1 12232
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 12328 0 -1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 12604 0 -1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_123
timestamp 1604681595
transform 1 0 12420 0 -1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_127
timestamp 1604681595
transform 1 0 12788 0 -1 12232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15640 0 -1 12232
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 15456 0 -1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_140
timestamp 1604681595
transform 1 0 13984 0 -1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_152
timestamp 1604681595
transform 1 0 15088 0 -1 12232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_167
timestamp 1604681595
transform 1 0 16468 0 -1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1604681595
transform 1 0 18308 0 -1 12232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 17940 0 -1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18768 0 -1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_179
timestamp 1604681595
transform 1 0 17572 0 -1 12232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_184
timestamp 1604681595
transform 1 0 18032 0 -1 12232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_190
timestamp 1604681595
transform 1 0 18584 0 -1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_194
timestamp 1604681595
transform 1 0 18952 0 -1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20792 0 -1 12232
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 20608 0 -1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_206
timestamp 1604681595
transform 1 0 20056 0 -1 12232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_223
timestamp 1604681595
transform 1 0 21620 0 -1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_235
timestamp 1604681595
transform 1 0 22724 0 -1 12232
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604681595
transform 1 0 24380 0 -1 12232
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 23552 0 -1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_243
timestamp 1604681595
transform 1 0 23460 0 -1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_245
timestamp 1604681595
transform 1 0 23644 0 -1 12232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_257
timestamp 1604681595
transform 1 0 24748 0 -1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 26864 0 -1 12232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_269
timestamp 1604681595
transform 1 0 25852 0 -1 12232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1604681595
transform 1 0 2484 0 1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1604681595
transform 1 0 2484 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 3956 0 1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_27
timestamp 1604681595
transform 1 0 3588 0 1 12232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_32
timestamp 1604681595
transform 1 0 4048 0 1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_27
timestamp 1604681595
transform 1 0 3588 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_39
timestamp 1604681595
transform 1 0 4692 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_44
timestamp 1604681595
transform 1 0 5152 0 1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_56
timestamp 1604681595
transform 1 0 6256 0 1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_51
timestamp 1604681595
transform 1 0 5796 0 -1 13320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_59
timestamp 1604681595
transform 1 0 6532 0 -1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 6716 0 -1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_68
timestamp 1604681595
transform 1 0 7360 0 1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_62
timestamp 1604681595
transform 1 0 6808 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_74
timestamp 1604681595
transform 1 0 7912 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 9568 0 1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_80
timestamp 1604681595
transform 1 0 8464 0 1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1604681595
transform 1 0 9660 0 1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_86
timestamp 1604681595
transform 1 0 9016 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_98
timestamp 1604681595
transform 1 0 10120 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_105
timestamp 1604681595
transform 1 0 10764 0 1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_117
timestamp 1604681595
transform 1 0 11868 0 1 12232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_110
timestamp 1604681595
transform 1 0 11224 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_123
timestamp 1604681595
transform 1 0 12420 0 -1 13320
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 12420 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 12328 0 -1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12604 0 1 12232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_20_131
timestamp 1604681595
transform 1 0 13156 0 -1 13320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_131
timestamp 1604681595
transform 1 0 13156 0 1 12232
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__79__A
timestamp 1604681595
transform 1 0 13432 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1604681595
transform 1 0 13432 0 -1 13320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_138
timestamp 1604681595
transform 1 0 13800 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_136
timestamp 1604681595
transform 1 0 13616 0 1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 1 12232
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 15180 0 1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_148
timestamp 1604681595
transform 1 0 14720 0 1 12232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_152
timestamp 1604681595
transform 1 0 15088 0 1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_150
timestamp 1604681595
transform 1 0 14904 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_162
timestamp 1604681595
transform 1 0 16008 0 -1 13320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_164
timestamp 1604681595
transform 1 0 16192 0 1 12232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_160
timestamp 1604681595
transform 1 0 15824 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16008 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_168
timestamp 1604681595
transform 1 0 16560 0 -1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_172
timestamp 1604681595
transform 1 0 16928 0 1 12232
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1604681595
transform 1 0 16744 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 16376 0 -1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1604681595
transform 1 0 16744 0 -1 13320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_178
timestamp 1604681595
transform 1 0 17480 0 -1 13320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_174
timestamp 1604681595
transform 1 0 17112 0 -1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_176
timestamp 1604681595
transform 1 0 17296 0 1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17296 0 -1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 17388 0 1 12232
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 17940 0 -1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 18124 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_183
timestamp 1604681595
transform 1 0 17940 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_187
timestamp 1604681595
transform 1 0 18308 0 1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_182
timestamp 1604681595
transform 1 0 17848 0 -1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_184
timestamp 1604681595
transform 1 0 18032 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_196
timestamp 1604681595
transform 1 0 19136 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_208
timestamp 1604681595
transform 1 0 20240 0 -1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_206
timestamp 1604681595
transform 1 0 20056 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_199
timestamp 1604681595
transform 1 0 19412 0 1 12232
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 20240 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1604681595
transform 1 0 19780 0 1 12232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_210
timestamp 1604681595
transform 1 0 20424 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 20424 0 -1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 20608 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 20792 0 1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 20884 0 1 12232
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 20608 0 -1 13320
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_19_234
timestamp 1604681595
transform 1 0 22632 0 1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_231
timestamp 1604681595
transform 1 0 22356 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_245
timestamp 1604681595
transform 1 0 23644 0 -1 13320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_243
timestamp 1604681595
transform 1 0 23460 0 -1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 23552 0 -1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604681595
transform 1 0 23736 0 1 12232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1604681595
transform 1 0 24380 0 -1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_254
timestamp 1604681595
transform 1 0 24472 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_250
timestamp 1604681595
transform 1 0 24104 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1604681595
transform 1 0 24288 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604681595
transform 1 0 24564 0 -1 13320
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1604681595
transform 1 0 24656 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_266
timestamp 1604681595
transform 1 0 25576 0 1 12232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_262
timestamp 1604681595
transform 1 0 25208 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1604681595
transform 1 0 25392 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1604681595
transform 1 0 24840 0 1 12232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_271
timestamp 1604681595
transform 1 0 26036 0 -1 13320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_276
timestamp 1604681595
transform 1 0 26496 0 1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_274
timestamp 1604681595
transform 1 0 26312 0 1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 26404 0 1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 26864 0 -1 13320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 26864 0 1 12232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_259
timestamp 1604681595
transform 1 0 24932 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1604681595
transform 1 0 2484 0 1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 3956 0 1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_27
timestamp 1604681595
transform 1 0 3588 0 1 13320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_32
timestamp 1604681595
transform 1 0 4048 0 1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_44
timestamp 1604681595
transform 1 0 5152 0 1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_56
timestamp 1604681595
transform 1 0 6256 0 1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_68
timestamp 1604681595
transform 1 0 7360 0 1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 9568 0 1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_80
timestamp 1604681595
transform 1 0 8464 0 1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1604681595
transform 1 0 9660 0 1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_105
timestamp 1604681595
transform 1 0 10764 0 1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_117
timestamp 1604681595
transform 1 0 11868 0 1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_129
timestamp 1604681595
transform 1 0 12972 0 1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1604681595
transform 1 0 15272 0 1 13320
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 15180 0 1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1604681595
transform 1 0 14996 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_141
timestamp 1604681595
transform 1 0 14076 0 1 13320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_149
timestamp 1604681595
transform 1 0 14812 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_158
timestamp 1604681595
transform 1 0 15640 0 1 13320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 17112 0 1 13320
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 16376 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16928 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 16008 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_164
timestamp 1604681595
transform 1 0 16192 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_168
timestamp 1604681595
transform 1 0 16560 0 1 13320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_183
timestamp 1604681595
transform 1 0 17940 0 1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_195
timestamp 1604681595
transform 1 0 19044 0 1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 21068 0 1 13320
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 20792 0 1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20608 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_207
timestamp 1604681595
transform 1 0 20148 0 1 13320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_211
timestamp 1604681595
transform 1 0 20516 0 1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_215
timestamp 1604681595
transform 1 0 20884 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1604681595
transform 1 0 21804 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_223
timestamp 1604681595
transform 1 0 21620 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_227
timestamp 1604681595
transform 1 0 21988 0 1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1604681595
transform 1 0 23460 0 1 13320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1604681595
transform 1 0 24564 0 1 13320
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1604681595
transform 1 0 24012 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24380 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_239
timestamp 1604681595
transform 1 0 23092 0 1 13320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_247
timestamp 1604681595
transform 1 0 23828 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_251
timestamp 1604681595
transform 1 0 24196 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 26864 0 1 13320
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 26404 0 1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1604681595
transform 1 0 25116 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1604681595
transform 1 0 25484 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_259
timestamp 1604681595
transform 1 0 24932 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_263
timestamp 1604681595
transform 1 0 25300 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_267
timestamp 1604681595
transform 1 0 25668 0 1 13320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_276
timestamp 1604681595
transform 1 0 26496 0 1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1604681595
transform 1 0 2484 0 -1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_27
timestamp 1604681595
transform 1 0 3588 0 -1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_39
timestamp 1604681595
transform 1 0 4692 0 -1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_51
timestamp 1604681595
transform 1 0 5796 0 -1 14408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_59
timestamp 1604681595
transform 1 0 6532 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 6716 0 -1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_62
timestamp 1604681595
transform 1 0 6808 0 -1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_74
timestamp 1604681595
transform 1 0 7912 0 -1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_86
timestamp 1604681595
transform 1 0 9016 0 -1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_98
timestamp 1604681595
transform 1 0 10120 0 -1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_110
timestamp 1604681595
transform 1 0 11224 0 -1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 12328 0 -1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_123
timestamp 1604681595
transform 1 0 12420 0 -1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_135
timestamp 1604681595
transform 1 0 13524 0 -1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_147
timestamp 1604681595
transform 1 0 14628 0 -1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 16376 0 -1 14408
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 15732 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17388 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 16192 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_161
timestamp 1604681595
transform 1 0 15916 0 -1 14408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_175
timestamp 1604681595
transform 1 0 17204 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1604681595
transform 1 0 18032 0 -1 14408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 17940 0 -1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 19136 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_179
timestamp 1604681595
transform 1 0 17572 0 -1 14408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_187
timestamp 1604681595
transform 1 0 18308 0 -1 14408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1604681595
transform 1 0 19044 0 -1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_198
timestamp 1604681595
transform 1 0 19320 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 19504 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 20976 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_202
timestamp 1604681595
transform 1 0 19688 0 -1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_214
timestamp 1604681595
transform 1 0 20792 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_218
timestamp 1604681595
transform 1 0 21160 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1604681595
transform 1 0 22448 0 -1 14408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1604681595
transform 1 0 21344 0 -1 14408
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21896 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 22264 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_224
timestamp 1604681595
transform 1 0 21712 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_228
timestamp 1604681595
transform 1 0 22080 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_235
timestamp 1604681595
transform 1 0 22724 0 -1 14408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24012 0 -1 14408
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 23552 0 -1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 23828 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_241
timestamp 1604681595
transform 1 0 23276 0 -1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_245
timestamp 1604681595
transform 1 0 23644 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_255
timestamp 1604681595
transform 1 0 24564 0 -1 14408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1604681595
transform 1 0 25300 0 -1 14408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 26864 0 -1 14408
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1604681595
transform 1 0 25024 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_259
timestamp 1604681595
transform 1 0 24932 0 -1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_262
timestamp 1604681595
transform 1 0 25208 0 -1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_267
timestamp 1604681595
transform 1 0 25668 0 -1 14408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_275
timestamp 1604681595
transform 1 0 26404 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1604681595
transform 1 0 2484 0 1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 3956 0 1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_27
timestamp 1604681595
transform 1 0 3588 0 1 14408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_32
timestamp 1604681595
transform 1 0 4048 0 1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_44
timestamp 1604681595
transform 1 0 5152 0 1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_56
timestamp 1604681595
transform 1 0 6256 0 1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_68
timestamp 1604681595
transform 1 0 7360 0 1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 9568 0 1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_80
timestamp 1604681595
transform 1 0 8464 0 1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1604681595
transform 1 0 9660 0 1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_105
timestamp 1604681595
transform 1 0 10764 0 1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_117
timestamp 1604681595
transform 1 0 11868 0 1 14408
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 12420 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12788 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_125
timestamp 1604681595
transform 1 0 12604 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_129
timestamp 1604681595
transform 1 0 12972 0 1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 15180 0 1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 15548 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_141
timestamp 1604681595
transform 1 0 14076 0 1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_154
timestamp 1604681595
transform 1 0 15272 0 1 14408
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 15732 0 1 14408
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_23_178
timestamp 1604681595
transform 1 0 17480 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 18216 0 1 14408
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 18032 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 17664 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_182
timestamp 1604681595
transform 1 0 17848 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 20976 0 1 14408
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 20792 0 1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 20608 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_205
timestamp 1604681595
transform 1 0 19964 0 1 14408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_211
timestamp 1604681595
transform 1 0 20516 0 1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_215
timestamp 1604681595
transform 1 0 20884 0 1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 22908 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_235
timestamp 1604681595
transform 1 0 22724 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 23460 0 1 14408
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 24472 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 23276 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_239
timestamp 1604681595
transform 1 0 23092 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_252
timestamp 1604681595
transform 1 0 24288 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_256
timestamp 1604681595
transform 1 0 24656 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1604681595
transform 1 0 25024 0 1 14408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 26864 0 1 14408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 26404 0 1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 24840 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25576 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_264
timestamp 1604681595
transform 1 0 25392 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_268
timestamp 1604681595
transform 1 0 25760 0 1 14408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_274
timestamp 1604681595
transform 1 0 26312 0 1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_276
timestamp 1604681595
transform 1 0 26496 0 1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1604681595
transform 1 0 2484 0 -1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_27
timestamp 1604681595
transform 1 0 3588 0 -1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_39
timestamp 1604681595
transform 1 0 4692 0 -1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_51
timestamp 1604681595
transform 1 0 5796 0 -1 15496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_59
timestamp 1604681595
transform 1 0 6532 0 -1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 6716 0 -1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_62
timestamp 1604681595
transform 1 0 6808 0 -1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_74
timestamp 1604681595
transform 1 0 7912 0 -1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_86
timestamp 1604681595
transform 1 0 9016 0 -1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_98
timestamp 1604681595
transform 1 0 10120 0 -1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_110
timestamp 1604681595
transform 1 0 11224 0 -1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12420 0 -1 15496
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 12328 0 -1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1604681595
transform 1 0 14904 0 -1 15496
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 15364 0 -1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 14352 0 -1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_142
timestamp 1604681595
transform 1 0 14168 0 -1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_146
timestamp 1604681595
transform 1 0 14536 0 -1 15496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_153
timestamp 1604681595
transform 1 0 15180 0 -1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_157
timestamp 1604681595
transform 1 0 15548 0 -1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16376 0 -1 15496
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 15732 0 -1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 16192 0 -1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_161
timestamp 1604681595
transform 1 0 15916 0 -1 15496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_175
timestamp 1604681595
transform 1 0 17204 0 -1 15496
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 19136 0 -1 15496
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 17940 0 -1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 18216 0 -1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_184
timestamp 1604681595
transform 1 0 18032 0 -1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_188
timestamp 1604681595
transform 1 0 18400 0 -1 15496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21620 0 -1 15496
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21436 0 -1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_232
timestamp 1604681595
transform 1 0 22448 0 -1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 23644 0 -1 15496
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 23552 0 -1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_254
timestamp 1604681595
transform 1 0 24472 0 -1 15496
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 -1 15496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 26864 0 -1 15496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_268
timestamp 1604681595
transform 1 0 25760 0 -1 15496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_276
timestamp 1604681595
transform 1 0 26496 0 -1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1604681595
transform 1 0 2484 0 1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 3956 0 1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_27
timestamp 1604681595
transform 1 0 3588 0 1 15496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_32
timestamp 1604681595
transform 1 0 4048 0 1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_44
timestamp 1604681595
transform 1 0 5152 0 1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_56
timestamp 1604681595
transform 1 0 6256 0 1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_68
timestamp 1604681595
transform 1 0 7360 0 1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 9568 0 1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_80
timestamp 1604681595
transform 1 0 8464 0 1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1604681595
transform 1 0 9660 0 1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11960 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_105
timestamp 1604681595
transform 1 0 10764 0 1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_117
timestamp 1604681595
transform 1 0 11868 0 1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 12512 0 1 15496
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 12328 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_120
timestamp 1604681595
transform 1 0 12144 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15272 0 1 15496
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 15180 0 1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 14444 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 14996 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_143
timestamp 1604681595
transform 1 0 14260 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_147
timestamp 1604681595
transform 1 0 14628 0 1 15496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 17296 0 1 15496
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17112 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16744 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_163
timestamp 1604681595
transform 1 0 16100 0 1 15496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_169
timestamp 1604681595
transform 1 0 16652 0 1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_172
timestamp 1604681595
transform 1 0 16928 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 18308 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 18676 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 19044 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_185
timestamp 1604681595
transform 1 0 18124 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_189
timestamp 1604681595
transform 1 0 18492 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_193
timestamp 1604681595
transform 1 0 18860 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_197
timestamp 1604681595
transform 1 0 19228 0 1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 20792 0 1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21068 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20608 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_209
timestamp 1604681595
transform 1 0 20332 0 1 15496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_215
timestamp 1604681595
transform 1 0 20884 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 21988 0 1 15496
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 21804 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21436 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_219
timestamp 1604681595
transform 1 0 21252 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_223
timestamp 1604681595
transform 1 0 21620 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24472 0 1 15496
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24288 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23920 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_246
timestamp 1604681595
transform 1 0 23736 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_250
timestamp 1604681595
transform 1 0 24104 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 26864 0 1 15496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 26404 0 1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1604681595
transform 1 0 25208 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_260
timestamp 1604681595
transform 1 0 25024 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_264
timestamp 1604681595
transform 1 0 25392 0 1 15496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_272
timestamp 1604681595
transform 1 0 26128 0 1 15496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_276
timestamp 1604681595
transform 1 0 26496 0 1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1604681595
transform 1 0 2484 0 -1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1604681595
transform 1 0 2484 0 1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 3956 0 1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_27
timestamp 1604681595
transform 1 0 3588 0 -1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_39
timestamp 1604681595
transform 1 0 4692 0 -1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_27
timestamp 1604681595
transform 1 0 3588 0 1 16584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_32
timestamp 1604681595
transform 1 0 4048 0 1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_51
timestamp 1604681595
transform 1 0 5796 0 -1 16584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_59
timestamp 1604681595
transform 1 0 6532 0 -1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_44
timestamp 1604681595
transform 1 0 5152 0 1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_56
timestamp 1604681595
transform 1 0 6256 0 1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 6716 0 -1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_62
timestamp 1604681595
transform 1 0 6808 0 -1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_74
timestamp 1604681595
transform 1 0 7912 0 -1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_68
timestamp 1604681595
transform 1 0 7360 0 1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 9568 0 1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_86
timestamp 1604681595
transform 1 0 9016 0 -1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_98
timestamp 1604681595
transform 1 0 10120 0 -1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_80
timestamp 1604681595
transform 1 0 8464 0 1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1604681595
transform 1 0 9660 0 1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12052 0 1 16584
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11868 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12052 0 -1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_110
timestamp 1604681595
transform 1 0 11224 0 -1 16584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_118
timestamp 1604681595
transform 1 0 11960 0 -1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_105
timestamp 1604681595
transform 1 0 10764 0 1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_128
timestamp 1604681595
transform 1 0 12880 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_121
timestamp 1604681595
transform 1 0 12236 0 -1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 12328 0 -1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_132
timestamp 1604681595
transform 1 0 13248 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 13524 0 -1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13064 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13432 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13616 0 1 16584
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_26_123
timestamp 1604681595
transform 1 0 12420 0 -1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 13708 0 -1 16584
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15272 0 1 16584
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 15180 0 1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14996 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 14628 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_156
timestamp 1604681595
transform 1 0 15456 0 -1 16584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_145
timestamp 1604681595
transform 1 0 14444 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_149
timestamp 1604681595
transform 1 0 14812 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_162
timestamp 1604681595
transform 1 0 16008 0 -1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16192 0 -1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15824 0 -1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_170
timestamp 1604681595
transform 1 0 16744 0 -1 16584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_166
timestamp 1604681595
transform 1 0 16376 0 -1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16560 0 -1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_177
timestamp 1604681595
transform 1 0 17388 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_173
timestamp 1604681595
transform 1 0 17020 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_178
timestamp 1604681595
transform 1 0 17480 0 -1 16584
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17204 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17296 0 -1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 17756 0 -1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 17572 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 17940 0 -1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18032 0 -1 16584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1604681595
transform 1 0 17756 0 1 16584
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_194
timestamp 1604681595
transform 1 0 18952 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_190
timestamp 1604681595
transform 1 0 18584 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19136 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 18768 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1604681595
transform 1 0 19320 0 1 16584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_193
timestamp 1604681595
transform 1 0 18860 0 -1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_201
timestamp 1604681595
transform 1 0 19596 0 1 16584
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 20148 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_213
timestamp 1604681595
transform 1 0 20700 0 1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_209
timestamp 1604681595
transform 1 0 20332 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_217
timestamp 1604681595
transform 1 0 21068 0 -1 16584
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 20516 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 20792 0 1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1604681595
transform 1 0 20884 0 1 16584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_218
timestamp 1604681595
transform 1 0 21160 0 1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_205
timestamp 1604681595
transform 1 0 19964 0 -1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1604681595
transform 1 0 23000 0 1 16584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21436 0 -1 16584
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 22448 0 -1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_230
timestamp 1604681595
transform 1 0 22264 0 -1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_234
timestamp 1604681595
transform 1 0 22632 0 -1 16584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_230
timestamp 1604681595
transform 1 0 22264 0 1 16584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_241
timestamp 1604681595
transform 1 0 23276 0 1 16584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_26_245
timestamp 1604681595
transform 1 0 23644 0 -1 16584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_242
timestamp 1604681595
transform 1 0 23368 0 -1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 23552 0 -1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_255
timestamp 1604681595
transform 1 0 24564 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_254
timestamp 1604681595
transform 1 0 24472 0 -1 16584
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23828 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24012 0 1 16584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23920 0 -1 16584
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24748 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_259
timestamp 1604681595
transform 1 0 24932 0 1 16584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_266
timestamp 1604681595
transform 1 0 25576 0 -1 16584
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1604681595
transform 1 0 25208 0 -1 16584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1604681595
transform 1 0 25300 0 1 16584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_271
timestamp 1604681595
transform 1 0 26036 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_267
timestamp 1604681595
transform 1 0 25668 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_274
timestamp 1604681595
transform 1 0 26312 0 -1 16584
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1604681595
transform 1 0 26220 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1604681595
transform 1 0 25852 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 26404 0 1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_276
timestamp 1604681595
transform 1 0 26496 0 1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 26864 0 1 16584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 26864 0 -1 16584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1604681595
transform 1 0 2484 0 -1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_27
timestamp 1604681595
transform 1 0 3588 0 -1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_39
timestamp 1604681595
transform 1 0 4692 0 -1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_51
timestamp 1604681595
transform 1 0 5796 0 -1 17672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_59
timestamp 1604681595
transform 1 0 6532 0 -1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 6716 0 -1 17672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_62
timestamp 1604681595
transform 1 0 6808 0 -1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_74
timestamp 1604681595
transform 1 0 7912 0 -1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_86
timestamp 1604681595
transform 1 0 9016 0 -1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_98
timestamp 1604681595
transform 1 0 10120 0 -1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12052 0 -1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_110
timestamp 1604681595
transform 1 0 11224 0 -1 17672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_118
timestamp 1604681595
transform 1 0 11960 0 -1 17672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 12328 0 -1 17672
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13616 0 -1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_121
timestamp 1604681595
transform 1 0 12236 0 -1 17672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_123
timestamp 1604681595
transform 1 0 12420 0 -1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_135
timestamp 1604681595
transform 1 0 13524 0 -1 17672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_138
timestamp 1604681595
transform 1 0 13800 0 -1 17672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 14076 0 -1 17672
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 15272 0 -1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_150
timestamp 1604681595
transform 1 0 14904 0 -1 17672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_156
timestamp 1604681595
transform 1 0 15456 0 -1 17672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15824 0 -1 17672
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_28_169
timestamp 1604681595
transform 1 0 16652 0 -1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 -1 17672
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 17940 0 -1 17672
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 19044 0 -1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17756 0 -1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_193
timestamp 1604681595
transform 1 0 18860 0 -1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_197
timestamp 1604681595
transform 1 0 19228 0 -1 17672
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 20148 0 -1 17672
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_28_205
timestamp 1604681595
transform 1 0 19964 0 -1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 23000 0 -1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_226
timestamp 1604681595
transform 1 0 21896 0 -1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24104 0 -1 17672
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 23552 0 -1 17672
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23828 0 -1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23368 0 -1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_240
timestamp 1604681595
transform 1 0 23184 0 -1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_245
timestamp 1604681595
transform 1 0 23644 0 -1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_249
timestamp 1604681595
transform 1 0 24012 0 -1 17672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_256
timestamp 1604681595
transform 1 0 24656 0 -1 17672
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1604681595
transform 1 0 25392 0 -1 17672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 26864 0 -1 17672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_268
timestamp 1604681595
transform 1 0 25760 0 -1 17672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1604681595
transform 1 0 26496 0 -1 17672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1604681595
transform 1 0 2484 0 1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 3956 0 1 17672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_27
timestamp 1604681595
transform 1 0 3588 0 1 17672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_32
timestamp 1604681595
transform 1 0 4048 0 1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_44
timestamp 1604681595
transform 1 0 5152 0 1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_56
timestamp 1604681595
transform 1 0 6256 0 1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_68
timestamp 1604681595
transform 1 0 7360 0 1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 9568 0 1 17672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_80
timestamp 1604681595
transform 1 0 8464 0 1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1604681595
transform 1 0 9660 0 1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_105
timestamp 1604681595
transform 1 0 10764 0 1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_117
timestamp 1604681595
transform 1 0 11868 0 1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 13432 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 13800 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_129
timestamp 1604681595
transform 1 0 12972 0 1 17672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_133
timestamp 1604681595
transform 1 0 13340 0 1 17672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_136
timestamp 1604681595
transform 1 0 13616 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 15180 0 1 17672
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 15640 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14168 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_140
timestamp 1604681595
transform 1 0 13984 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_144
timestamp 1604681595
transform 1 0 14352 0 1 17672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_152
timestamp 1604681595
transform 1 0 15088 0 1 17672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_154
timestamp 1604681595
transform 1 0 15272 0 1 17672
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15824 0 1 17672
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18308 0 1 17672
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 18124 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 17756 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_179
timestamp 1604681595
transform 1 0 17572 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_183
timestamp 1604681595
transform 1 0 17940 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20884 0 1 17672
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 20792 0 1 17672
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 20240 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_206
timestamp 1604681595
transform 1 0 20056 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_210
timestamp 1604681595
transform 1 0 20424 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23000 0 1 17672
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 22816 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 21896 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 22264 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_224
timestamp 1604681595
transform 1 0 21712 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_228
timestamp 1604681595
transform 1 0 22080 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_232
timestamp 1604681595
transform 1 0 22448 0 1 17672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_257
timestamp 1604681595
transform 1 0 24748 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 26864 0 1 17672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 26404 0 1 17672
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 24932 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1604681595
transform 1 0 25300 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_261
timestamp 1604681595
transform 1 0 25116 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_265
timestamp 1604681595
transform 1 0 25484 0 1 17672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_273
timestamp 1604681595
transform 1 0 26220 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_276
timestamp 1604681595
transform 1 0 26496 0 1 17672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 18760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1604681595
transform 1 0 2484 0 -1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_27
timestamp 1604681595
transform 1 0 3588 0 -1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_39
timestamp 1604681595
transform 1 0 4692 0 -1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_51
timestamp 1604681595
transform 1 0 5796 0 -1 18760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_59
timestamp 1604681595
transform 1 0 6532 0 -1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 6716 0 -1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_62
timestamp 1604681595
transform 1 0 6808 0 -1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_74
timestamp 1604681595
transform 1 0 7912 0 -1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_86
timestamp 1604681595
transform 1 0 9016 0 -1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_98
timestamp 1604681595
transform 1 0 10120 0 -1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12052 0 -1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_110
timestamp 1604681595
transform 1 0 11224 0 -1 18760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_118
timestamp 1604681595
transform 1 0 11960 0 -1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 13432 0 -1 18760
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 12328 0 -1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12880 0 -1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13248 0 -1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_121
timestamp 1604681595
transform 1 0 12236 0 -1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_123
timestamp 1604681595
transform 1 0 12420 0 -1 18760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_127
timestamp 1604681595
transform 1 0 12788 0 -1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_130
timestamp 1604681595
transform 1 0 13064 0 -1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_153
timestamp 1604681595
transform 1 0 15180 0 -1 18760
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 15824 0 -1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_159
timestamp 1604681595
transform 1 0 15732 0 -1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_162
timestamp 1604681595
transform 1 0 16008 0 -1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_174
timestamp 1604681595
transform 1 0 17112 0 -1 18760
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 18032 0 -1 18760
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 17940 0 -1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 17756 0 -1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_180
timestamp 1604681595
transform 1 0 17664 0 -1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 21068 0 -1 18760
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20884 0 -1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_203
timestamp 1604681595
transform 1 0 19780 0 -1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_236
timestamp 1604681595
transform 1 0 22816 0 -1 18760
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23644 0 -1 18760
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 23552 0 -1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_254
timestamp 1604681595
transform 1 0 24472 0 -1 18760
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1604681595
transform 1 0 25208 0 -1 18760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 26864 0 -1 18760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_266
timestamp 1604681595
transform 1 0 25576 0 -1 18760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_274
timestamp 1604681595
transform 1 0 26312 0 -1 18760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 18760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1604681595
transform 1 0 2484 0 1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 3956 0 1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_27
timestamp 1604681595
transform 1 0 3588 0 1 18760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_32
timestamp 1604681595
transform 1 0 4048 0 1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_44
timestamp 1604681595
transform 1 0 5152 0 1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_56
timestamp 1604681595
transform 1 0 6256 0 1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_68
timestamp 1604681595
transform 1 0 7360 0 1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 9568 0 1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_80
timestamp 1604681595
transform 1 0 8464 0 1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1604681595
transform 1 0 9660 0 1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12052 0 1 18760
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11868 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_105
timestamp 1604681595
transform 1 0 10764 0 1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_138
timestamp 1604681595
transform 1 0 13800 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 15180 0 1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14996 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 15456 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13984 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_142
timestamp 1604681595
transform 1 0 14168 0 1 18760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_150
timestamp 1604681595
transform 1 0 14904 0 1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_154
timestamp 1604681595
transform 1 0 15272 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_158
timestamp 1604681595
transform 1 0 15640 0 1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1604681595
transform 1 0 16836 0 1 18760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_170
timestamp 1604681595
transform 1 0 16744 0 1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_174
timestamp 1604681595
transform 1 0 17112 0 1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19228 0 1 18760
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19044 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18676 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_186
timestamp 1604681595
transform 1 0 18216 0 1 18760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_190
timestamp 1604681595
transform 1 0 18584 0 1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_193
timestamp 1604681595
transform 1 0 18860 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 20792 0 1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20240 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_206
timestamp 1604681595
transform 1 0 20056 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_210
timestamp 1604681595
transform 1 0 20424 0 1 18760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_215
timestamp 1604681595
transform 1 0 20884 0 1 18760
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1604681595
transform 1 0 22356 0 1 18760
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 22172 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21804 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21436 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_223
timestamp 1604681595
transform 1 0 21620 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_227
timestamp 1604681595
transform 1 0 21988 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1604681595
transform 1 0 24564 0 1 18760
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23828 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_240
timestamp 1604681595
transform 1 0 23184 0 1 18760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_246
timestamp 1604681595
transform 1 0 23736 0 1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_249
timestamp 1604681595
transform 1 0 24012 0 1 18760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 26864 0 1 18760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 26404 0 1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1604681595
transform 1 0 25116 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1604681595
transform 1 0 25484 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_259
timestamp 1604681595
transform 1 0 24932 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_263
timestamp 1604681595
transform 1 0 25300 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_267
timestamp 1604681595
transform 1 0 25668 0 1 18760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_276
timestamp 1604681595
transform 1 0 26496 0 1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 19848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1604681595
transform 1 0 2484 0 -1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_27
timestamp 1604681595
transform 1 0 3588 0 -1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_39
timestamp 1604681595
transform 1 0 4692 0 -1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_51
timestamp 1604681595
transform 1 0 5796 0 -1 19848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_59
timestamp 1604681595
transform 1 0 6532 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 6716 0 -1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_62
timestamp 1604681595
transform 1 0 6808 0 -1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_74
timestamp 1604681595
transform 1 0 7912 0 -1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_86
timestamp 1604681595
transform 1 0 9016 0 -1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_98
timestamp 1604681595
transform 1 0 10120 0 -1 19848
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11224 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10764 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11592 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_104
timestamp 1604681595
transform 1 0 10672 0 -1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_107
timestamp 1604681595
transform 1 0 10948 0 -1 19848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_112
timestamp 1604681595
transform 1 0 11408 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_116
timestamp 1604681595
transform 1 0 11776 0 -1 19848
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12880 0 -1 19848
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 12328 0 -1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12604 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_123
timestamp 1604681595
transform 1 0 12420 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_127
timestamp 1604681595
transform 1 0 12788 0 -1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_137
timestamp 1604681595
transform 1 0 13708 0 -1 19848
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 14996 0 -1 19848
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13984 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_142
timestamp 1604681595
transform 1 0 14168 0 -1 19848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_150
timestamp 1604681595
transform 1 0 14904 0 -1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16928 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_170
timestamp 1604681595
transform 1 0 16744 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_174
timestamp 1604681595
transform 1 0 17112 0 -1 19848
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1604681595
transform 1 0 18492 0 -1 19848
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 17940 0 -1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19228 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_182
timestamp 1604681595
transform 1 0 17848 0 -1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_184
timestamp 1604681595
transform 1 0 18032 0 -1 19848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_188
timestamp 1604681595
transform 1 0 18400 0 -1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1604681595
transform 1 0 18768 0 -1 19848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_196
timestamp 1604681595
transform 1 0 19136 0 -1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19504 0 -1 19848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_199
timestamp 1604681595
transform 1 0 19412 0 -1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_206
timestamp 1604681595
transform 1 0 20056 0 -1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_218
timestamp 1604681595
transform 1 0 21160 0 -1 19848
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1604681595
transform 1 0 22540 0 -1 19848
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 22356 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21988 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 23000 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_226
timestamp 1604681595
transform 1 0 21896 0 -1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_229
timestamp 1604681595
transform 1 0 22172 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_236
timestamp 1604681595
transform 1 0 22816 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23828 0 -1 19848
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 23552 0 -1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_240
timestamp 1604681595
transform 1 0 23184 0 -1 19848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_245
timestamp 1604681595
transform 1 0 23644 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_253
timestamp 1604681595
transform 1 0 24380 0 -1 19848
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1604681595
transform 1 0 25116 0 -1 19848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 26864 0 -1 19848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_265
timestamp 1604681595
transform 1 0 25484 0 -1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 19848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 20936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1604681595
transform 1 0 2484 0 1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1604681595
transform 1 0 2484 0 -1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 3956 0 1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_27
timestamp 1604681595
transform 1 0 3588 0 1 19848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_32
timestamp 1604681595
transform 1 0 4048 0 1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_27
timestamp 1604681595
transform 1 0 3588 0 -1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_39
timestamp 1604681595
transform 1 0 4692 0 -1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_44
timestamp 1604681595
transform 1 0 5152 0 1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_56
timestamp 1604681595
transform 1 0 6256 0 1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_51
timestamp 1604681595
transform 1 0 5796 0 -1 20936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_59
timestamp 1604681595
transform 1 0 6532 0 -1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 6716 0 -1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_68
timestamp 1604681595
transform 1 0 7360 0 1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_62
timestamp 1604681595
transform 1 0 6808 0 -1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_74
timestamp 1604681595
transform 1 0 7912 0 -1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 9568 0 1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_80
timestamp 1604681595
transform 1 0 8464 0 1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_93
timestamp 1604681595
transform 1 0 9660 0 1 19848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_86
timestamp 1604681595
transform 1 0 9016 0 -1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_98
timestamp 1604681595
transform 1 0 10120 0 -1 20936
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11224 0 1 19848
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10764 0 -1 20936
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10764 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10396 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 10396 0 -1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_103
timestamp 1604681595
transform 1 0 10580 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_107
timestamp 1604681595
transform 1 0 10948 0 1 19848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_103
timestamp 1604681595
transform 1 0 10580 0 -1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_114
timestamp 1604681595
transform 1 0 11592 0 -1 20936
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 12328 0 -1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 -1 20936
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_34_136
timestamp 1604681595
transform 1 0 13616 0 -1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_132
timestamp 1604681595
transform 1 0 13248 0 -1 20936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_133
timestamp 1604681595
transform 1 0 13340 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_129
timestamp 1604681595
transform 1 0 12972 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13708 0 -1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13524 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13156 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13708 0 1 19848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1604681595
transform 1 0 13892 0 -1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_147
timestamp 1604681595
transform 1 0 14628 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_143
timestamp 1604681595
transform 1 0 14260 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14444 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13984 0 -1 20936
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_33_157
timestamp 1604681595
transform 1 0 15548 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_151
timestamp 1604681595
transform 1 0 14996 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14812 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 15180 0 1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1604681595
transform 1 0 15272 0 1 19848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_149
timestamp 1604681595
transform 1 0 14812 0 -1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 16284 0 1 19848
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16100 0 -1 20936
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 16100 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 15732 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 15916 0 -1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 17112 0 -1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_161
timestamp 1604681595
transform 1 0 15916 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_172
timestamp 1604681595
transform 1 0 16928 0 -1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_176
timestamp 1604681595
transform 1 0 17296 0 -1 20936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_188
timestamp 1604681595
transform 1 0 18400 0 -1 20936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_184
timestamp 1604681595
transform 1 0 18032 0 -1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_182
timestamp 1604681595
transform 1 0 17848 0 -1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_184
timestamp 1604681595
transform 1 0 18032 0 1 19848
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 18216 0 -1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 18400 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 17940 0 -1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_190
timestamp 1604681595
transform 1 0 18584 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18768 0 -1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 18768 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18952 0 1 19848
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 18952 0 -1 20936
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_33_207
timestamp 1604681595
transform 1 0 20148 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_203
timestamp 1604681595
transform 1 0 19780 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19964 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_213
timestamp 1604681595
transform 1 0 20700 0 -1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_215
timestamp 1604681595
transform 1 0 20884 0 1 19848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_211
timestamp 1604681595
transform 1 0 20516 0 1 19848
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 20332 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 20884 0 -1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 20792 0 1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_217
timestamp 1604681595
transform 1 0 21068 0 -1 20936
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 22356 0 1 19848
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21988 0 -1 20936
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21988 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21620 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1604681595
transform 1 0 21804 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_229
timestamp 1604681595
transform 1 0 22172 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_225
timestamp 1604681595
transform 1 0 21804 0 -1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_236
timestamp 1604681595
transform 1 0 22816 0 -1 20936
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23644 0 -1 20936
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 23552 0 -1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 24288 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 24656 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23368 0 -1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_250
timestamp 1604681595
transform 1 0 24104 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_254
timestamp 1604681595
transform 1 0 24472 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_266
timestamp 1604681595
transform 1 0 25576 0 1 19848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_262
timestamp 1604681595
transform 1 0 25208 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1604681595
transform 1 0 25392 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1604681595
transform 1 0 24840 0 1 19848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_276
timestamp 1604681595
transform 1 0 26496 0 1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_274
timestamp 1604681595
transform 1 0 26312 0 1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 26404 0 1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 26864 0 -1 20936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 26864 0 1 19848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_264
timestamp 1604681595
transform 1 0 25392 0 -1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 20936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604681595
transform 1 0 2484 0 1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 3956 0 1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_27
timestamp 1604681595
transform 1 0 3588 0 1 20936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_32
timestamp 1604681595
transform 1 0 4048 0 1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_44
timestamp 1604681595
transform 1 0 5152 0 1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_56
timestamp 1604681595
transform 1 0 6256 0 1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_68
timestamp 1604681595
transform 1 0 7360 0 1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 9568 0 1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 10212 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_80
timestamp 1604681595
transform 1 0 8464 0 1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_93
timestamp 1604681595
transform 1 0 9660 0 1 20936
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10396 0 1 20936
box -38 -48 1786 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1604681595
transform 1 0 12880 0 1 20936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_120
timestamp 1604681595
transform 1 0 12144 0 1 20936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_131
timestamp 1604681595
transform 1 0 13156 0 1 20936
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13892 0 1 20936
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 15180 0 1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 15456 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 14996 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14628 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_145
timestamp 1604681595
transform 1 0 14444 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_149
timestamp 1604681595
transform 1 0 14812 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_154
timestamp 1604681595
transform 1 0 15272 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_158
timestamp 1604681595
transform 1 0 15640 0 1 20936
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16652 0 1 20936
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16468 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16100 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_162
timestamp 1604681595
transform 1 0 16008 0 1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_165
timestamp 1604681595
transform 1 0 16284 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_178
timestamp 1604681595
transform 1 0 17480 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18860 0 1 20936
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 18676 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18308 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17664 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_182
timestamp 1604681595
transform 1 0 17848 0 1 20936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_186
timestamp 1604681595
transform 1 0 18216 0 1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_189
timestamp 1604681595
transform 1 0 18492 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 20884 0 1 20936
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 20792 0 1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 20608 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_202
timestamp 1604681595
transform 1 0 19688 0 1 20936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_210
timestamp 1604681595
transform 1 0 20424 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_234
timestamp 1604681595
transform 1 0 22632 0 1 20936
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23368 0 1 20936
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1604681595
transform 1 0 24564 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23184 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_251
timestamp 1604681595
transform 1 0 24196 0 1 20936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_257
timestamp 1604681595
transform 1 0 24748 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1604681595
transform 1 0 24932 0 1 20936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 26864 0 1 20936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 26404 0 1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1604681595
transform 1 0 25484 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_263
timestamp 1604681595
transform 1 0 25300 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_267
timestamp 1604681595
transform 1 0 25668 0 1 20936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_276
timestamp 1604681595
transform 1 0 26496 0 1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 1104 0 -1 22024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1604681595
transform 1 0 1380 0 -1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1604681595
transform 1 0 2484 0 -1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_27
timestamp 1604681595
transform 1 0 3588 0 -1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_39
timestamp 1604681595
transform 1 0 4692 0 -1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_51
timestamp 1604681595
transform 1 0 5796 0 -1 22024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_59
timestamp 1604681595
transform 1 0 6532 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 6716 0 -1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_62
timestamp 1604681595
transform 1 0 6808 0 -1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_74
timestamp 1604681595
transform 1 0 7912 0 -1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_86
timestamp 1604681595
transform 1 0 9016 0 -1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_98
timestamp 1604681595
transform 1 0 10120 0 -1 22024
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 10764 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11132 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11500 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_104
timestamp 1604681595
transform 1 0 10672 0 -1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_107
timestamp 1604681595
transform 1 0 10948 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_111
timestamp 1604681595
transform 1 0 11316 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_115
timestamp 1604681595
transform 1 0 11684 0 -1 22024
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1604681595
transform 1 0 13524 0 -1 22024
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 12328 0 -1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 13340 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_121
timestamp 1604681595
transform 1 0 12236 0 -1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_123
timestamp 1604681595
transform 1 0 12420 0 -1 22024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_131
timestamp 1604681595
transform 1 0 13156 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1604681595
transform 1 0 13800 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15456 0 -1 22024
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13984 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 15272 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14352 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_142
timestamp 1604681595
transform 1 0 14168 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_146
timestamp 1604681595
transform 1 0 14536 0 -1 22024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_175
timestamp 1604681595
transform 1 0 17204 0 -1 22024
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18032 0 -1 22024
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 17940 0 -1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18768 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19136 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_190
timestamp 1604681595
transform 1 0 18584 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1604681595
transform 1 0 18952 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_198
timestamp 1604681595
transform 1 0 19320 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19504 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_202
timestamp 1604681595
transform 1 0 19688 0 -1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_214
timestamp 1604681595
transform 1 0 20792 0 -1 22024
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1604681595
transform 1 0 21896 0 -1 22024
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21712 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_222
timestamp 1604681595
transform 1 0 21528 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_229
timestamp 1604681595
transform 1 0 22172 0 -1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1604681595
transform 1 0 24564 0 -1 22024
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 23552 0 -1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23368 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_241
timestamp 1604681595
transform 1 0 23276 0 -1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_245
timestamp 1604681595
transform 1 0 23644 0 -1 22024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1604681595
transform 1 0 24380 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 26864 0 -1 22024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_259
timestamp 1604681595
transform 1 0 24932 0 -1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_271
timestamp 1604681595
transform 1 0 26036 0 -1 22024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 1104 0 1 22024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1604681595
transform 1 0 1380 0 1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1604681595
transform 1 0 2484 0 1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 3956 0 1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_27
timestamp 1604681595
transform 1 0 3588 0 1 22024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_32
timestamp 1604681595
transform 1 0 4048 0 1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_44
timestamp 1604681595
transform 1 0 5152 0 1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_56
timestamp 1604681595
transform 1 0 6256 0 1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_68
timestamp 1604681595
transform 1 0 7360 0 1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_80
timestamp 1604681595
transform 1 0 8464 0 1 22024
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8832 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_86
timestamp 1604681595
transform 1 0 9016 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9200 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_93
timestamp 1604681595
transform 1 0 9660 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_90
timestamp 1604681595
transform 1 0 9384 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 9568 0 1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_97
timestamp 1604681595
transform 1 0 10028 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9844 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10212 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10764 0 1 22024
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10580 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_101
timestamp 1604681595
transform 1 0 10396 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13524 0 1 22024
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 13340 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12972 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_124
timestamp 1604681595
transform 1 0 12512 0 1 22024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_128
timestamp 1604681595
transform 1 0 12880 0 1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_131
timestamp 1604681595
transform 1 0 13156 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15456 0 1 22024
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 15180 0 1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14628 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_144
timestamp 1604681595
transform 1 0 14352 0 1 22024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_149
timestamp 1604681595
transform 1 0 14812 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_154
timestamp 1604681595
transform 1 0 15272 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 17020 0 1 22024
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 16836 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16468 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_165
timestamp 1604681595
transform 1 0 16284 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1604681595
transform 1 0 16652 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 18952 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19320 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_192
timestamp 1604681595
transform 1 0 18768 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_196
timestamp 1604681595
transform 1 0 19136 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19504 0 1 22024
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 20792 0 1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 20516 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 21068 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_206
timestamp 1604681595
transform 1 0 20056 0 1 22024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_210
timestamp 1604681595
transform 1 0 20424 0 1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_213
timestamp 1604681595
transform 1 0 20700 0 1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_215
timestamp 1604681595
transform 1 0 20884 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21712 0 1 22024
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21528 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 22724 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_219
timestamp 1604681595
transform 1 0 21252 0 1 22024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_233
timestamp 1604681595
transform 1 0 22540 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_237
timestamp 1604681595
transform 1 0 22908 0 1 22024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1604681595
transform 1 0 23460 0 1 22024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1604681595
transform 1 0 24564 0 1 22024
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24012 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1604681595
transform 1 0 23276 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_247
timestamp 1604681595
transform 1 0 23828 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_251
timestamp 1604681595
transform 1 0 24196 0 1 22024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 26864 0 1 22024
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 26404 0 1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1604681595
transform 1 0 25116 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1604681595
transform 1 0 25484 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_259
timestamp 1604681595
transform 1 0 24932 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_263
timestamp 1604681595
transform 1 0 25300 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_267
timestamp 1604681595
transform 1 0 25668 0 1 22024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_276
timestamp 1604681595
transform 1 0 26496 0 1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 1104 0 -1 23112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1604681595
transform 1 0 1380 0 -1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1604681595
transform 1 0 2484 0 -1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_27
timestamp 1604681595
transform 1 0 3588 0 -1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_39
timestamp 1604681595
transform 1 0 4692 0 -1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_51
timestamp 1604681595
transform 1 0 5796 0 -1 23112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_59
timestamp 1604681595
transform 1 0 6532 0 -1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 6716 0 -1 23112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_62
timestamp 1604681595
transform 1 0 6808 0 -1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_74
timestamp 1604681595
transform 1 0 7912 0 -1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9200 0 -1 23112
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_38_86
timestamp 1604681595
transform 1 0 9016 0 -1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_97
timestamp 1604681595
transform 1 0 10028 0 -1 23112
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10764 0 -1 23112
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_38_114
timestamp 1604681595
transform 1 0 11592 0 -1 23112
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 13340 0 -1 23112
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 12328 0 -1 23112
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13156 0 -1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_123
timestamp 1604681595
transform 1 0 12420 0 -1 23112
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 15456 0 -1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_152
timestamp 1604681595
transform 1 0 15088 0 -1 23112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_158
timestamp 1604681595
transform 1 0 15640 0 -1 23112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16100 0 -1 23112
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15916 0 -1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 17112 0 -1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_172
timestamp 1604681595
transform 1 0 16928 0 -1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_176
timestamp 1604681595
transform 1 0 17296 0 -1 23112
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18032 0 -1 23112
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 17940 0 -1 23112
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 19044 0 -1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_182
timestamp 1604681595
transform 1 0 17848 0 -1 23112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_193
timestamp 1604681595
transform 1 0 18860 0 -1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1604681595
transform 1 0 19228 0 -1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 20516 0 -1 23112
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19412 0 -1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_201
timestamp 1604681595
transform 1 0 19596 0 -1 23112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_209
timestamp 1604681595
transform 1 0 20332 0 -1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_230
timestamp 1604681595
transform 1 0 22264 0 -1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23644 0 -1 23112
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604681595
transform 1 0 23552 0 -1 23112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_242
timestamp 1604681595
transform 1 0 23368 0 -1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_251
timestamp 1604681595
transform 1 0 24196 0 -1 23112
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1604681595
transform 1 0 24932 0 -1 23112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 26864 0 -1 23112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_263
timestamp 1604681595
transform 1 0 25300 0 -1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_275
timestamp 1604681595
transform 1 0 26404 0 -1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 1104 0 1 23112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 1104 0 -1 24200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1604681595
transform 1 0 1380 0 1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1604681595
transform 1 0 2484 0 1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1604681595
transform 1 0 1380 0 -1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1604681595
transform 1 0 2484 0 -1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604681595
transform 1 0 3956 0 1 23112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_27
timestamp 1604681595
transform 1 0 3588 0 1 23112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_32
timestamp 1604681595
transform 1 0 4048 0 1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_27
timestamp 1604681595
transform 1 0 3588 0 -1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_39
timestamp 1604681595
transform 1 0 4692 0 -1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_44
timestamp 1604681595
transform 1 0 5152 0 1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_56
timestamp 1604681595
transform 1 0 6256 0 1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_51
timestamp 1604681595
transform 1 0 5796 0 -1 24200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_59
timestamp 1604681595
transform 1 0 6532 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604681595
transform 1 0 6716 0 -1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_68
timestamp 1604681595
transform 1 0 7360 0 1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_62
timestamp 1604681595
transform 1 0 6808 0 -1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_74
timestamp 1604681595
transform 1 0 7912 0 -1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604681595
transform 1 0 9568 0 1 23112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_80
timestamp 1604681595
transform 1 0 8464 0 1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_93
timestamp 1604681595
transform 1 0 9660 0 1 23112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_86
timestamp 1604681595
transform 1 0 9016 0 -1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_98
timestamp 1604681595
transform 1 0 10120 0 -1 24200
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1604681595
transform 1 0 10948 0 -1 24200
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10764 0 1 23112
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 10580 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 10764 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_101
timestamp 1604681595
transform 1 0 10396 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_104
timestamp 1604681595
transform 1 0 10672 0 -1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_110
timestamp 1604681595
transform 1 0 11224 0 -1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_123
timestamp 1604681595
transform 1 0 12420 0 -1 24200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_128
timestamp 1604681595
transform 1 0 12880 0 1 23112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_124
timestamp 1604681595
transform 1 0 12512 0 1 23112
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604681595
transform 1 0 12328 0 -1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_131
timestamp 1604681595
transform 1 0 13156 0 -1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_131
timestamp 1604681595
transform 1 0 13156 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 12972 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13340 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13524 0 1 23112
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 13248 0 -1 24200
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604681595
transform 1 0 15180 0 1 23112
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 15640 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14536 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 14904 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_144
timestamp 1604681595
transform 1 0 14352 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_148
timestamp 1604681595
transform 1 0 14720 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_152
timestamp 1604681595
transform 1 0 15088 0 1 23112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_154
timestamp 1604681595
transform 1 0 15272 0 1 23112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_151
timestamp 1604681595
transform 1 0 14996 0 -1 24200
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1604681595
transform 1 0 16192 0 -1 24200
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15824 0 1 23112
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 15824 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_159
timestamp 1604681595
transform 1 0 15732 0 -1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_162
timestamp 1604681595
transform 1 0 16008 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_167
timestamp 1604681595
transform 1 0 16468 0 -1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_184
timestamp 1604681595
transform 1 0 18032 0 -1 24200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_179
timestamp 1604681595
transform 1 0 17572 0 -1 24200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_179
timestamp 1604681595
transform 1 0 17572 0 1 23112
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 18308 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 18124 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604681595
transform 1 0 17940 0 -1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_189
timestamp 1604681595
transform 1 0 18492 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18676 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18860 0 -1 24200
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 18308 0 1 23112
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_39_206
timestamp 1604681595
transform 1 0 20056 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20240 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_214
timestamp 1604681595
transform 1 0 20792 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_215
timestamp 1604681595
transform 1 0 20884 0 1 23112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_210
timestamp 1604681595
transform 1 0 20424 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 20976 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 20608 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21160 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604681595
transform 1 0 20792 0 1 23112
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21160 0 -1 24200
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_40_202
timestamp 1604681595
transform 1 0 19688 0 -1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 21528 0 1 23112
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 22172 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_220
timestamp 1604681595
transform 1 0 21344 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_227
timestamp 1604681595
transform 1 0 21988 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_231
timestamp 1604681595
transform 1 0 22356 0 -1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_243
timestamp 1604681595
transform 1 0 23460 0 -1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_245
timestamp 1604681595
transform 1 0 23644 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_241
timestamp 1604681595
transform 1 0 23276 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23460 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604681595
transform 1 0 23552 0 -1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23644 0 -1 24200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_251
timestamp 1604681595
transform 1 0 24196 0 -1 24200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_255
timestamp 1604681595
transform 1 0 24564 0 1 23112
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23828 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24012 0 1 23112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_267
timestamp 1604681595
transform 1 0 25668 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_261
timestamp 1604681595
transform 1 0 25116 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1604681595
transform 1 0 24932 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1604681595
transform 1 0 25300 0 1 23112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1604681595
transform 1 0 24932 0 -1 24200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_275
timestamp 1604681595
transform 1 0 26404 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_276
timestamp 1604681595
transform 1 0 26496 0 1 23112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_271
timestamp 1604681595
transform 1 0 26036 0 1 23112
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1604681595
transform 1 0 25852 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604681595
transform 1 0 26404 0 1 23112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 26864 0 -1 24200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 26864 0 1 23112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_263
timestamp 1604681595
transform 1 0 25300 0 -1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 1104 0 1 24200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1604681595
transform 1 0 1380 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1604681595
transform 1 0 2484 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604681595
transform 1 0 3956 0 1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_27
timestamp 1604681595
transform 1 0 3588 0 1 24200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_32
timestamp 1604681595
transform 1 0 4048 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_44
timestamp 1604681595
transform 1 0 5152 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_56
timestamp 1604681595
transform 1 0 6256 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_68
timestamp 1604681595
transform 1 0 7360 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604681595
transform 1 0 9568 0 1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_80
timestamp 1604681595
transform 1 0 8464 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1604681595
transform 1 0 9660 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_105
timestamp 1604681595
transform 1 0 10764 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_117
timestamp 1604681595
transform 1 0 11868 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_129
timestamp 1604681595
transform 1 0 12972 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604681595
transform 1 0 15180 0 1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_141
timestamp 1604681595
transform 1 0 14076 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_154
timestamp 1604681595
transform 1 0 15272 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_166
timestamp 1604681595
transform 1 0 16376 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_178
timestamp 1604681595
transform 1 0 17480 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1604681595
transform 1 0 19044 0 1 24200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_190
timestamp 1604681595
transform 1 0 18584 0 1 24200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_194
timestamp 1604681595
transform 1 0 18952 0 1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_198
timestamp 1604681595
transform 1 0 19320 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604681595
transform 1 0 20792 0 1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_210
timestamp 1604681595
transform 1 0 20424 0 1 24200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_215
timestamp 1604681595
transform 1 0 20884 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1604681595
transform 1 0 22540 0 1 24200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_227
timestamp 1604681595
transform 1 0 21988 0 1 24200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_237
timestamp 1604681595
transform 1 0 22908 0 1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23644 0 1 24200
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1604681595
transform 1 0 23092 0 1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1604681595
transform 1 0 23460 0 1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24380 0 1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1604681595
transform 1 0 24748 0 1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_241
timestamp 1604681595
transform 1 0 23276 0 1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_251
timestamp 1604681595
transform 1 0 24196 0 1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_255
timestamp 1604681595
transform 1 0 24564 0 1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1604681595
transform 1 0 24932 0 1 24200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 26864 0 1 24200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604681595
transform 1 0 26404 0 1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1604681595
transform 1 0 25484 0 1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_263
timestamp 1604681595
transform 1 0 25300 0 1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_267
timestamp 1604681595
transform 1 0 25668 0 1 24200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_276
timestamp 1604681595
transform 1 0 26496 0 1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 1104 0 -1 25288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1604681595
transform 1 0 1380 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1604681595
transform 1 0 2484 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604681595
transform 1 0 3956 0 -1 25288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1604681595
transform 1 0 3588 0 -1 25288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1604681595
transform 1 0 4048 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_44
timestamp 1604681595
transform 1 0 5152 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_56
timestamp 1604681595
transform 1 0 6256 0 -1 25288
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604681595
transform 1 0 6808 0 -1 25288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_63
timestamp 1604681595
transform 1 0 6900 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_75
timestamp 1604681595
transform 1 0 8004 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604681595
transform 1 0 9660 0 -1 25288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_87
timestamp 1604681595
transform 1 0 9108 0 -1 25288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_94
timestamp 1604681595
transform 1 0 9752 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_106
timestamp 1604681595
transform 1 0 10856 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_118
timestamp 1604681595
transform 1 0 11960 0 -1 25288
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604681595
transform 1 0 12512 0 -1 25288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_125
timestamp 1604681595
transform 1 0 12604 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_137
timestamp 1604681595
transform 1 0 13708 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604681595
transform 1 0 15364 0 -1 25288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_149
timestamp 1604681595
transform 1 0 14812 0 -1 25288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_156
timestamp 1604681595
transform 1 0 15456 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_168
timestamp 1604681595
transform 1 0 16560 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604681595
transform 1 0 18216 0 -1 25288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_180
timestamp 1604681595
transform 1 0 17664 0 -1 25288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_187
timestamp 1604681595
transform 1 0 18308 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604681595
transform 1 0 21068 0 -1 25288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_199
timestamp 1604681595
transform 1 0 19412 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_211
timestamp 1604681595
transform 1 0 20516 0 -1 25288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_218
timestamp 1604681595
transform 1 0 21160 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1604681595
transform 1 0 22816 0 -1 25288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_230
timestamp 1604681595
transform 1 0 22264 0 -1 25288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1604681595
transform 1 0 24564 0 -1 25288
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1604681595
transform 1 0 23920 0 -1 25288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_240
timestamp 1604681595
transform 1 0 23184 0 -1 25288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_42_249
timestamp 1604681595
transform 1 0 24012 0 -1 25288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 26864 0 -1 25288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_259
timestamp 1604681595
transform 1 0 24932 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_271
timestamp 1604681595
transform 1 0 26036 0 -1 25288
box -38 -48 590 592
<< labels >>
rlabel metal3 s 0 6664 480 6784 6 ccff_head
port 0 nsew default input
rlabel metal3 s 0 20672 480 20792 6 ccff_tail
port 1 nsew default tristate
rlabel metal3 s 27520 3536 28000 3656 6 chanx_right_in[0]
port 2 nsew default input
rlabel metal3 s 27520 9520 28000 9640 6 chanx_right_in[10]
port 3 nsew default input
rlabel metal3 s 27520 10064 28000 10184 6 chanx_right_in[11]
port 4 nsew default input
rlabel metal3 s 27520 10608 28000 10728 6 chanx_right_in[12]
port 5 nsew default input
rlabel metal3 s 27520 11288 28000 11408 6 chanx_right_in[13]
port 6 nsew default input
rlabel metal3 s 27520 11832 28000 11952 6 chanx_right_in[14]
port 7 nsew default input
rlabel metal3 s 27520 12512 28000 12632 6 chanx_right_in[15]
port 8 nsew default input
rlabel metal3 s 27520 13056 28000 13176 6 chanx_right_in[16]
port 9 nsew default input
rlabel metal3 s 27520 13600 28000 13720 6 chanx_right_in[17]
port 10 nsew default input
rlabel metal3 s 27520 14280 28000 14400 6 chanx_right_in[18]
port 11 nsew default input
rlabel metal3 s 27520 14824 28000 14944 6 chanx_right_in[19]
port 12 nsew default input
rlabel metal3 s 27520 4080 28000 4200 6 chanx_right_in[1]
port 13 nsew default input
rlabel metal3 s 27520 4760 28000 4880 6 chanx_right_in[2]
port 14 nsew default input
rlabel metal3 s 27520 5304 28000 5424 6 chanx_right_in[3]
port 15 nsew default input
rlabel metal3 s 27520 5848 28000 5968 6 chanx_right_in[4]
port 16 nsew default input
rlabel metal3 s 27520 6528 28000 6648 6 chanx_right_in[5]
port 17 nsew default input
rlabel metal3 s 27520 7072 28000 7192 6 chanx_right_in[6]
port 18 nsew default input
rlabel metal3 s 27520 7616 28000 7736 6 chanx_right_in[7]
port 19 nsew default input
rlabel metal3 s 27520 8296 28000 8416 6 chanx_right_in[8]
port 20 nsew default input
rlabel metal3 s 27520 8840 28000 8960 6 chanx_right_in[9]
port 21 nsew default input
rlabel metal3 s 27520 15368 28000 15488 6 chanx_right_out[0]
port 22 nsew default tristate
rlabel metal3 s 27520 21352 28000 21472 6 chanx_right_out[10]
port 23 nsew default tristate
rlabel metal3 s 27520 22032 28000 22152 6 chanx_right_out[11]
port 24 nsew default tristate
rlabel metal3 s 27520 22576 28000 22696 6 chanx_right_out[12]
port 25 nsew default tristate
rlabel metal3 s 27520 23120 28000 23240 6 chanx_right_out[13]
port 26 nsew default tristate
rlabel metal3 s 27520 23800 28000 23920 6 chanx_right_out[14]
port 27 nsew default tristate
rlabel metal3 s 27520 24344 28000 24464 6 chanx_right_out[15]
port 28 nsew default tristate
rlabel metal3 s 27520 25024 28000 25144 6 chanx_right_out[16]
port 29 nsew default tristate
rlabel metal3 s 27520 25568 28000 25688 6 chanx_right_out[17]
port 30 nsew default tristate
rlabel metal3 s 27520 26112 28000 26232 6 chanx_right_out[18]
port 31 nsew default tristate
rlabel metal3 s 27520 26792 28000 26912 6 chanx_right_out[19]
port 32 nsew default tristate
rlabel metal3 s 27520 16048 28000 16168 6 chanx_right_out[1]
port 33 nsew default tristate
rlabel metal3 s 27520 16592 28000 16712 6 chanx_right_out[2]
port 34 nsew default tristate
rlabel metal3 s 27520 17272 28000 17392 6 chanx_right_out[3]
port 35 nsew default tristate
rlabel metal3 s 27520 17816 28000 17936 6 chanx_right_out[4]
port 36 nsew default tristate
rlabel metal3 s 27520 18360 28000 18480 6 chanx_right_out[5]
port 37 nsew default tristate
rlabel metal3 s 27520 19040 28000 19160 6 chanx_right_out[6]
port 38 nsew default tristate
rlabel metal3 s 27520 19584 28000 19704 6 chanx_right_out[7]
port 39 nsew default tristate
rlabel metal3 s 27520 20264 28000 20384 6 chanx_right_out[8]
port 40 nsew default tristate
rlabel metal3 s 27520 20808 28000 20928 6 chanx_right_out[9]
port 41 nsew default tristate
rlabel metal2 s 938 27240 994 27720 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 7746 27240 7802 27720 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 8390 27240 8446 27720 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 9126 27240 9182 27720 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 9770 27240 9826 27720 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 10506 27240 10562 27720 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 11150 27240 11206 27720 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 11886 27240 11942 27720 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 12530 27240 12586 27720 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 13174 27240 13230 27720 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 13910 27240 13966 27720 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 1582 27240 1638 27720 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 2318 27240 2374 27720 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 2962 27240 3018 27720 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 3698 27240 3754 27720 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 4342 27240 4398 27720 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 4986 27240 5042 27720 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 5722 27240 5778 27720 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 6366 27240 6422 27720 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 7102 27240 7158 27720 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 14554 27240 14610 27720 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 21362 27240 21418 27720 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 22098 27240 22154 27720 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 22742 27240 22798 27720 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 23478 27240 23534 27720 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 24122 27240 24178 27720 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 24766 27240 24822 27720 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 25502 27240 25558 27720 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 26146 27240 26202 27720 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 26882 27240 26938 27720 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 27526 27240 27582 27720 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 15290 27240 15346 27720 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 15934 27240 15990 27720 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 16578 27240 16634 27720 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 17314 27240 17370 27720 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 17958 27240 18014 27720 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 18694 27240 18750 27720 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 19338 27240 19394 27720 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 20074 27240 20130 27720 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 20718 27240 20774 27720 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 27520 27336 28000 27456 6 prog_clk
port 82 nsew default input
rlabel metal3 s 27520 2856 28000 2976 6 right_bottom_grid_pin_11_
port 83 nsew default input
rlabel metal3 s 27520 0 28000 120 6 right_bottom_grid_pin_1_
port 84 nsew default input
rlabel metal3 s 27520 544 28000 664 6 right_bottom_grid_pin_3_
port 85 nsew default input
rlabel metal3 s 27520 1088 28000 1208 6 right_bottom_grid_pin_5_
port 86 nsew default input
rlabel metal3 s 27520 1768 28000 1888 6 right_bottom_grid_pin_7_
port 87 nsew default input
rlabel metal3 s 27520 2312 28000 2432 6 right_bottom_grid_pin_9_
port 88 nsew default input
rlabel metal2 s 294 27240 350 27720 6 top_left_grid_pin_1_
port 89 nsew default input
rlabel metal4 s 5611 1848 5931 25336 6 VPWR
port 90 nsew default input
rlabel metal4 s 10277 1848 10597 25336 6 VGND
port 91 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 27720
<< end >>
